// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
lwpbVUb1BtsqTTkDV0Xb+1CzCuYwocOQT6Yi+JdueKKlUgq7bPPPYZU5Usq51Ecl
gpmq0zJbl1Ztc2G32LO+3pimDCafrbVe+JdMrG9RA6lopDWAHzGi+Qc51Zwuzt9z
jL88WspjBcnfwZhHNb4TFNLTQW1E6bYVSEOcTlgMtAY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 46432 )
`pragma protect data_block
Dar5cFI58WH/ysRGa4gwz0utJd6t9ua0uxzQ3wO0yQRjRJDAvj7UEYq2ojbrePg6
Y48YdcO+L2HQViBIRM1ukqhi76gmiKB/Fdg4uj29eeavk45AaMUuBDK1EuFPLvl7
Hsr0WLTrQn6991IEuFLVx4kRTNexL+YypqHD3cZa3punBw0N3a/sovXD66eR5CkZ
MBvnqpmXz2QHur5rBmwzxx3nIEHc3sNob+YudXlFpRA9Fmbq9gArGjPa70SX7HkO
Me2rNLxtcgFbNZ3mpp1XECTtDj27nGakc4OKVUBuAmwXEmgmXCZOn2jateVmDwlf
+McDlhm/r4sqgrwKgu7V+5a067KxnLU8uE1MR1Tc33nijn5oYtOyFXtrAMiM1/j2
hNiJ9OPc3s1yZlkB7a/CpQ5aJhRsgMRxe//xhn/n/3ufMwhkgGztlg4iItl/3wgX
np2wDocB1JaN9a6xc6GVsjYblghZFE7teSNIDhYkFb6E7rncykcJLu1eRobq2sjr
MklidrKXOmKho6xGbLiONQ3BQ68OI5NPodsMaI4A06b9mfJzKEKXO85LlDylrBJb
1dc1EuVooha9gOtD84vIXcfvj+EctE96MzkLDmnWSrFG8AM5EXDnXM7MKDRdoRpH
OTPTFI08/RWA5cHZTVuJCwQTh5zc5X7kyjknCA1lbdfK1Bsrwn01tdLm5blvjc5b
Tcyr/msbRAL0fUtWNHLbAs6kfW/Wj8msDqqOQa8/Ypkc1KNsitcd+yUA8vTMfXpF
/EE/q0YObY6KpZsYynaND5EEzKjCijs18SooKK0vo0VPCC8F0NvGoaXYF4JuYoXN
QjYxwl1r5XENAFn73W8k1oELY4YAYObNBXd8TUaGEyUggDmLMCjG8jeCL0O7iGeI
sCkmpnD3h3EvRGucwCUk1Lq0ndTcFlvoNKDsDT0BXqdJPVNQcPDSqzvs2iTIdEcg
J87SE3Z0n5lxUEYD3golHE4ai4AnKorvZFmFp2BLA3jZpjvH23xRCWOnCQD6uh05
P6BJyIPOAbtH2jAoy7ykoC46zc+ckQNB6o+rJuyPcF10GYxWqJ5OwRDnXXDKP5zl
J2NT2RYxKtuYrvqSyWHDKHCWi0QW8RKXtNWx7m/HgXPkjaxlau5Zl7xvZQXPSzfh
0LX35pHEHYnLxXezwkpu+NZklNEn4v/lW1aMW0HK9hCJ3JZ//0Uu1/WF1e1yCtoi
mYz1RCK0hG4qjmb4bfZBGbQbo8hpe613+4n/53wkD0nJ/rMJN68KE74vZSdhbLU6
aGW4VviK8wJ5tV8GbEgGa731cUGNIAsKKIyHCdZ45fqzarftZ6NJ+cpKzt5CIJJn
WDLGhlp6cB/4mjPK+Om8CjPjQXgypHXwkI2JzJ1SWU5ACUsFsB3dyNm4fqoDbowa
sZUNqjHFXSYXbWz2UCdzS7i1uYJf0DlqOFvzNI+M83fjIeZQAGxEopeIMKCIyffV
7uEJsKtc78UwWlPT7S44z/sR7i4HfK7JfrkkFbxmfu1kAh1evKOoMdzJuk7QMTlu
ccZDS6MeUfF2dzQg8P2mFS8gu6SpWPRhl6FlF2nu95DmULiWntktiSclJjohzQsh
yfP6vC+0OeEVqFYo28eHhvWvRRBD5VVJfpCRy+SJp53k13cwOL9e7XwXULFkzmnX
xYpGxxRC+QFcLs9Yewc/oWr+PHFAs3xfzg15lLA9amGpeLRHhVycROEhl1x9DLWv
iOvc/XmrgTxCkIexUXEb+SU19tUrPjIcmN5k29L3E+DEV91RoMYgacZq2h3TLCO6
soqHZmV74J1rrE5KzUp0c/gb2Jf+BIMT/jNwXp8ixUExQ8JfIt/HjlyUPQrrfUIQ
TRViEMLe7tm855muQXO5Qf1P72cekHcdLCha2TaSj1H4CepG4KYKCmmqVHiIVX/a
dopn0gcVrtpKQyKIYOfYv7A4wfhzi0QWc8sLDKk62N6xB7CD6fQ84rtEY/d7odEE
Bw2PlODZATy9OhoW92EIUWkeDb2+xyArBQGc3bsuy8hXtPNYCo7gma/nspdR2Qx1
9xZBiVhs8rVphvjTha38DTDvo+XH+nmXFjtOq0eHaUPXpOSPSo2r2FBQXk1Auhpi
XkRlJMivnQiddFy/vClph5H9qt4uLC+a1w9nTYEkxz/elEvdIJNL3uLhptT0dlng
4liCgH8A0Z3rbaY3We9750x+6aKQlb0jwwF60qGjL5TkjJ67kdk5j4S/AIEF9o3f
o1X1B6Ci8ZcmmqNh/lhFNykjFC4DgktfOcRnFp1MidxCSG0nWcisXB19fRxYfx3l
1tFBg7cD8AuV4hYly5MOvdf286hH6JdKN+5a47m1nD7zWIyy3T3uKa7DQHi/Q0eg
/yUYZvrvi5SBPZ2jpapW8XQq47pgLbed6+ganjusJ8nVHLJvGmmcMRpJPlBkcArO
9OGIVMeM/uPX/IEfwbm4p3aAw1uGNXgHih119foPgatDsGEdjz9eNi2nAq71ymUN
9cm7SQ9JovpCIGcF6DBE37LsBybsSFmnL4Cv7I+3KlxRyvy/MJSEzYSlTeXe47WQ
YhQ5tuCx6IfYCGb7vXbfJRkBPqSM6wFgyc1YE1UL1ao5+D5Gdybo8ifBk/9fhVCg
+oLhNg1kfhL+n1UmSAllBohK5KIfeeLdulkCwXcknFONuqfvbF3b4RWLwGdlFQ85
IU+oWrI+ijofA1rP6WQqIQ6FBKJ8OtGymDr/GqS1IU7LVBE4noUkYl56bDyrum+1
fhN2+vwc8EphDoOogUQu2Me64K6xoyTzOqFPPMuWDK2WuntOwquWaX4Kg8KZuVsy
PjY7rzkzxvNbSmRA+yMhsiI3Xtj9cvl79xSE7hrnvahujh47/qBh3nML9Pm6z8IM
QNsKn0MpzNvmoEKRA5ZHwiPitt6KexCkMjUk8NRYXD4bLl0VKPq4q0n0VSHdXnxn
XASYLDJCs2pIOHrzwxQsS1jUlc30QgTFyGSooMxKiC/tS9yLmB/rH6n7/YKIjIb/
7vRwkK6SkFtBpNVnuxt1j9BxOtsAX6kU4NaA1lE8Ao95rzot2zMjuXR+NQ8+dEqc
a7NmmpgKeus+TNMyqfofUD/oNjJMjTVTjd5BxmBES6FP9HMdz/WGD2pMyklm25EC
5JRqJWoO5oobIqgOxpc5/id31M7Jmv0FdEd5+TpSDGNKkigZd2A6wmyPus2gaToJ
9Tu82vGsAKZihOD81yFoM9o+PEq4f21Z6PcPDJCXanCDRsrz8vMqyWd+nUOw+rzF
fHbt21cpj2ImWTMLblD2gpkm98+claKnKMA58kIDpPwxlyYklBNianZZBeztPKfH
rhiVSn+JTR52VamcmwgcnL1lea9crwu0IaYH4yg2WJRO1UJ+TW3K8ZLjKU0bZSDl
bO7Z3lbdArZZ5eZ+S5ltj7TLfd0Wy8Bx4q8+8O9ULbpNRij0Bq846QL3/LDNQfH8
3l2BBI3MT/xPfylZwE0KIaiOy1LgJZ20tIqmmQY4/7W7oIyACDtt9zz0r+Bb+aQG
8+a3c4VNvbLvXvnxhGdHY6cKuSBk9eStJzazZWUXxvwB0h0PhUB30mkxgLKv1lpo
+g+PgtyjlHE3+LsY7VX0wCgHtrfQ1Z5hGqJni+GFesZLzLWDUHpv4xjMc6m9s64G
m08mse/YnxroNBc5pA6zYRStKy0EumxgosLZzaw+ZIZd1aqDduRijin1QIRf8xYe
S6zYPgcyiZUdlFfQIEjx51Zubp2/asZfTFde4B5XwdRO25RwdnqmirTdDqtJPMyp
J9vucnV0L9UIYz2z0wsiwyiYuX8W4JmVAj+d9+fwhczhKPFMYOgQ8Ei45tLBoSkQ
V74syATRz1qvB0fdXlc/glWvIVAeZ0rO+1LM37JIpGUeWX+rvmASDTBFlv5lGULb
nUPa0dCuOdodHaa9hc9AJqFTG9VPw5SePI3fpcNqAmUPNUWV8r07wdqXC8EpkeNf
PR1pe2WwG2pTXJ/E6/LQxde0gVNwoAaVbEyGoQ9WWKGgt0nnsdFmLYD4R9Cq36zc
cf+Qj3ML2OuBPvQmzUuUy2b9VBJHcjXgNZNGKaE+UfmzQW75CMVLNGw53b/3DJqp
yH8HTT74LY7Ze/TMjG8KWZw+vHbGE1L9zaN2EG+0Rj3tq+aWVGqLf0MHeZicR1rI
+UFxAaZtxAL10htSA90CAMoryms846lb8aXviiDuIF73jhkeuLtshFJ4kY4H8Rmy
HUy/tbGqivY/JKhduxgRrcO1l9bpEL2u/hQ1TLxwHiq12h9fN+WJBR7EZD0uMBA9
Bxfg4TosENdoeHViB8dxruD+PRCm6RIDWUibqGxGWcM4Sfx4OBpOVJFVRtpyCKRi
ntaA2EwWPbxSjCYwuU4HYGPcGgu6K6NcjhwyMZQ7aVliRe+Ya/wZPtVubBt8zcTZ
7uOb2pjE7xnyeddEaKxE5c0YD08eeQhwx7cqXefc3wk2Apg318GU5OgixebTRQmY
4IEuBJajwiZ+whn4/d7JoLJu1qQ2zwPK3iPRSGxaVb3kcT1tmO3eKHJYXB92yh4b
7DKw/OnVZYS2j2fYsgURQVvxbue9hyYfZ/7KYH4IeVfzFPRaBQ4xUEAQ6+4Dcl36
+YWbYzTRIerkM7jrON+C9/qX99lbXE8xipuTotMfBOUlkUqWaAEmDZQhfku4iXnH
OR1s1ozmKi6wLlb+FVRFDDSfBuy02MNECMUIen8wIz1o01lbW4bDcRZbkugxU8LO
vz43zbKkNSv26fIm/nL849HpvgKaN9Hq5SsYxfHQiDr6AjBqT/feHrljov3l5zc9
w9ICXq/6goTpLazeLTNI6NY2ODIH8ksdJgw0ZorWvkFaxcWzq2MoFoGsizmauhVC
DtEY5v6bj2tgj6SM33eGSL5KVoz0XA2fFmeQtibYfa3nsfx9a2ZI6qgUufdqIrBj
qCzd7KmTnvXf5Ha4y7zfUjDcQjzaD36u4OjbwN+8jk7jwdMojthWMs8G1gZ4YwGE
0lLGL+nj/1lcr8Gezn4KnqxJvzKFhiI4hlASfPT+eWFtITZNJKrOQVSUkZi1Rb7f
U4VCiYP7w7uWK0kcO5aA6fuXiOPH8XE14T0vQjuTF3C3OM8B8TfDceilyC9oXqMC
EUsQ6Z5/vJIAovtF4NcBc8/OIZk0PYRIwlNyw0B8cTu2cF/RD6uLr9vFyRZd3z4N
wk0+1zrkSkkAxgQCbfQHFmah941OakbcWM1fMCUvXxpeVXr30xo4T1Rp/S/9S6g3
VbtBhezfJPfyUqpQKvTUthStRTQW3xFc2QkNsG7yJ7ttYplniKucOLsPwTL6210B
Yy9vCHa2l/cmHRJ+gJsiWRJM2hHO8Tma5CUMCPmqQBGWbYckLt2qdlLZEv7We5J7
n2Bs97ODe1QY/gH1cgky7wCmrdzV+VIauWvvjLaY7vCz0l0i+Y37W0jZcV4lJFA1
YmBoRoP8cfPuCJksEhHuSwZCczNR+R/135fd6IB3qbWmR4N0Yuiv/4UaeXk1nL1l
G3xGUTYUoLGj2By3H3hi0Rn47A6WMvmvF99w443j4DJTxHFybAJT+jq3qRfNI5+W
w7onI6tEm+WUppIC0kQQuQACDvB2RH28OISkkVAWg7j4k9AoKU1F0J72ywPb9BGo
rxa97A7DR3t4ho17dcj8OpP+Jv2zvWOJ9IKCxb5O9i22dHuwf52OJAIluoHnZWsQ
/aQ111qJwBPnJf7iFyRp5JwX7KofqAzd0SLPSTilEDBn1norZGNUKuqCLVzk1B47
KTo6bOQuzGQQt61TbKWpN924LuP67dfjYDbT+ufsaRYYJYzGZW7cDGFEAJiKfGiy
gqfvkds7XVnHYcHe6XPi/+KsYI6mICyJErBYJ6bSD92GNAE5kF1jpO6RFhM5PWsd
dqYIYjJKj+tOQ0kayaNIn3QK0SCTWOZcpktz+gptY2Yn9I1xAFrCGRxXwA3F//bc
vBK4XAZpZKdZLi73F8eR0mR7avfvQ7liY9YBHxZSNTZh+u2qQCvVUBLJVrnAJMnC
QD0uYIKWcPtt0NSG4JGv7oqnrFlW9FqqTY7GmEmYzSBzdSjdwJJOhI37j6HbSrc9
q3t8pTOlvYoYAMVyuWVqdMU8wo9YyPdfpGDoDzjJsD5ZgMKJnGdam1yLOxUtLQD1
KyjDueRwEY+RCJ4bmwsoySWd1yPkamJzENxTy+kzzZfNTA4l/C2d+HuJM3Ce9JOi
NxF2QkKLG8GdUb5PSEWYen7RlUsg87mCDLlkC14pYiCycE02tKmcoPouCkQXKv5l
OBjZ8PjY7M8FhxFkgg6WfgRmg2DCcjk8rL6ppvImFcMteC6MEX3A5NXJppn6Np+x
SrQVJILJvJwADt7v/hZv7G7y0UtULHXdy5u/8yYotmmEHWJqTL91pKf1KZsSZuBZ
iZEcoG82/c0GDZJlyNu2cLNXJbwm/2ZfYnXpo/X9EsbddXPxV12dx6QcDKj0z5Op
llpLtcABg9KhoiNpFNnb/eVnOiK95OfIELS9XALuoCg9QOoCXiGhqYDL1BISs3iz
aD7oYXNZCPSiyKKG7XFcH68gvsjbV8lm1xnP5qJxyIXEbbO3q6f2Ybcq6RfqqmzC
MxAaWyOaYd+/BDonSJ/dAn9XzVmJgSd8n2ZM8eJMv3TqQbsenXEL2ZWLAPTecQT7
vHYobzQD53BGJ3EVisJnqy9LZuuJ3yKzlW0E4XiS3LkoyL8G4nwY04k6EfNgtejW
ujqRICFp+s4+vimVMwvAesV5+ZqrB1zL26Mhu9qw1GhS0ih8pZ7eKR49U8c+vx2S
8T6StTuA6upIIHBMvAtJleALO24iS1daquYpeBtUElGZI29CaV17Esimde5MiDrR
/4RAeafy71SkS/UHND/tViy0PKM//NvMqsozhMbqNqtZuo5UbYTDz1W9gA8C2QdD
85p6T9BD6lGSgOdDSDUrzXF8rCeurBXHBiO6ADJWNN+6Ji751D5aacPW0I+JS7gL
uR4rQI46ZebC6XH/6s8rgPcae6sXCioAMUFldFUcoTJjSIzhC3DQQww7oYKNerTB
KI5+YUEqjq/+KmvXZj3ql7EEw0OPBV/1jP29nrpzLcEYTwCSO+AYyrSChpLl4ttE
oHYepP7JVxdS2WjZd72pqfeg65VwIc+HxGCYmca7SBQ33Erd1hoV/VZFtGa5KQYo
IoE7+AJOJ49BxIoX5CdaaYel6nDro4UIeCJm58ZVf00WSQeTufKV2d8nViJVcFbE
3Gapnt/iKZE3etCOpI3qfgZ5ej5yY2OMWBSiwNPpR6ZSVaVxT4Lj3N+2uNPng/uz
LAU00Zx8Am4l7qchNLEvL6XZ3qdV2RcD+B7Y5BmfxBirvxEYGRedJpoeD2WZoNzo
1KvVrkvr/L1hCrP+dhGfNme59XBwjZtAdlHQK4T6WWYR3cnIBpbM61pogxNtL+XL
NsUFLZP6Gn4pie3d9weOqSCVvqjEsqxRFLfi7TnqoXefA5+K5qtKF/2qgrVWgcZk
xxHNl13n34FejWAVcsjFJdqxaLRIEyGtR39chI0Coi5NEx7yu3LUQO70qauTF49O
Vm6ac22e5tQ2Uluyx+gR4OcY8WkBKSGX37tIh9iPMVdOxekuQeBxnvY2Wnc5uF3X
fl49IyWR744hruC1DEZpNlnZZR4tpTIlU3U8XlMG/TSYBfNDqURJlcyIH0krbVjm
LBx2tTABHxFPI1rOthICLQy73TRaXxKwMphUb4O53XFN0RXiT8FPVHa9Ok9acIHP
n7LSqjwt60p9YFWNatqm02lOU5OgjvNH5sZgXZLFKld3ihMQ3d/EUyLoMQ/YTYNb
3O9dkKa9ChxfZfXPoPomiAm+4DhEuFaLaCGFwXdRJAZ9MNl2TC/7ohGh0zG7jnCx
wQLKBXtsW98EH3ZfqfCPZ9q6lKuWyPAjPA4jOSwXMBkjj6i9V/BOVcMC6E9eT+DD
8n3EqRu+foq1Z+R/75/OEFmhkewI1QERxfzI5M3mhG77wIOv8ephabXVxkuy7+jD
dOUKpX6ufgW4SZqPyvouJqdJ7alXhqmPygoz7T1r6WuAzHXxpwKVmKUolfmGJibt
XqD7dkkBXP12nQ20WIhZYWFIflhOg0Zv/5c9W912XOcUs62zAFtlb7ju4x7OZW/D
vhx4bZYJBoIUE2nalj4EbDgvorvgU65HDHlUhURBdeRgtfpLiB/X1Xve0dLJmS+K
MRJTsXdYiDLFKeWtB+GjLDxahC0j8hrw0uY0NbdpPRm0POEYJjytzOaGmddDcSa7
gaqCOp/SYmNe0Mzj6zOb3/LGPWT1YEr7BiEwXFe6NRpU+0nGspwpnG0TGXC7ZOuE
/7McMUTKK9eL3FnBI9zH6lGYusUdcOcEIuZpfdhiZ8hBJVhqzot1tI5+ywFAN/yN
i3cPJLAR62v6MM7r5VQnRHKwr6qkHwONCMG2W26KekyFARGS0qrIOad7obFi32Ae
x/YP+zpfRMkZwTkksepXBvy2Z46I4Y4LHrBZHmDmiVU6Aa9lPAYopP+G+N879HBn
kkaNNunbThlLmMudOhjreLt1TIIOh6svpKI2CLI70F3Ff4nj9rhS0219W+Rra7NG
+IQU+BYn1lqM3zQeznLSUgrh8IFBTw3ejnmHvrSf/LujFwJ49CeFnpFlPXCWP8Lq
r/Kq7GjpFnShrz3MB9EfLblZDnNjf1q+BExXcAphKfqaORV3lwHvLrKpa1XUismz
nvOVjJTqfqw1aU1TBL4AVWn621h/UylralqWOg2SiBYq5pzDxvHi9bF3DmrjN2HG
bZ4rpqEtu8Xr83WXdOV2SdUZaApZ8R+zxHpWW0DUhJGUcQf1YtjWfgKIB8nN+07D
6xTxb6bWL1VPeeaf5Mhge+JrSSZsVOCRBaelN1+8wPiEFcVbrRwK46YXOPsQCuGH
WLb0rf49fkiFeDRMUZPuwKGJSdtD3BJOPqugI+IhLJlt76r2b0UXfhWvnKEOG8qQ
LDwMzCEwFDtMvK23WkdvxqPIlcYpE3fdWDck+wPplua0G4ZqPGWC7Rrfb+0xASxk
qN6WdVNAJEynodRBAj1ThvXQNSp4Ta0lB2sDP39M1F7iUbTO7qBOsR6tW7giHXpo
E/bUGJlbxWwZuiRm+EhPlNcus/i4HjXkKPFD+kzJis8Af/pUCnLcmpvSjvotmnuo
SSofPX9rW9/5l5K2ErOAH9Kq9M5K3XT0CieSFX+H22ah3fHp/Q9LSs4LbGnMWOU5
sUlSJ7ZHr+7kBIxdPwvLsNYLqBBtw5YsQE8OBnVZlqRRVrrHthwsj4NW3g1YM8kW
0OMTSw9Y0DtHKxmmY3GPFbUAgc34fjz4MfbJKPop9MN2xSZVraYytKE3woo4Ehx3
8BkAyhR4cwnxLzJ0+KXNuqirpicmAqk3k3Rq7GgEdwUOD/iRMRsCvtudU98oKmdT
popBghukNPT+8vJ0elfiZ+Rj0ESy8LNJbxYwwmN0HkINGptKo524LRzNutssTD41
B1ktoethD8Q01g0kRgMmeQ4/xbHgOjZiL+R6CS7uXiAiyNBWgtfVITTkTkS6qje0
RNWHcT8Jd/ICYfcZHjYI6TrC3lMz/VMJyX5rwPtJbsVIlLGwi5w3+tB+IeE6x+ZI
A3CTD0vUAReip48y/RVPzmiDy6Q89rEG1l3Jdwq+8PoWalTzHv48HApLAfOHoESX
jpZAOgdXlwlf0oym1PgtvZ9JFXmuyeiMpqJlyf+LS1GyxT4nUwuKNVm7ft73bw1j
Jv2qFLkiNf9VCuR2ikkqH3Xvq5d28t3wLqWDPRDDkHAWoVm6JhlhU3sKl0wZIbDX
0eI2kw/qKvofkIlULdELBHFIDgR9QmoEzYdFHFR+72TriwMa8FAXge0yrv4paRMG
TzUhjEnrZyp+avYGl/PkJogDj5Ttb9MvnFFYCoKYDu4IDmF5nuxKw87PMufi9dHe
8WVP3SPEYmzWZezQEtvIGOyB/70wKkggZMzsTnSiDod+EN6GVn6Eha7enTnksQoU
YfIsdB7SzdPUcaaaUyfSSXYakWLC8UGdEWC/L1hft8JTXzE9HF1ae0ZVPS4nr/hQ
Z/0HEjVnPwYT6EAJUcUbYmLE1mVUr1nnc3uD7yT13usdnOjpPitFh7DB4/Dw29Yl
Ay7dOOwzpOLhQupkCSHhQ6rq9oPHHUCbsUli5ZEhul2oqcDMzgozQZXFXxWrVv5M
KNxX7je7VQ9KHCkBK1J230m5g9VlcWNF+DMZ6DisARxRBH1oed74yI1Msts9V7eB
YJ7sL9EnakvsVC+0xBFFJhuPk9VEFq16P5XAsOnpvIhe/C85cklMsVf/H0yY6O5l
+OQwXkxRe6MsF9L+YxYS4pgb/9oufbMo1MCmXTCceXx4CmlKDhOwfhZrR8N3yDHu
eLdLE34Sj59IHUB3C2xLSZXLQuyfpFDRmErWEn8kJ1TVyeSOkI3RXUa1SaMMMoCR
QDjr+MVhg7sHovY5z0O5Z3nj72Xyg7od6MU8/tJrVAj53kHY7hv8KPX4myKP4w38
Dj7BgJ0p319PbYjV1JYAZyXHoAGXHWF1uuDnXTCVJWPmc5y62cAhVLCDa+LJziFh
w5SJ3OOXXOhjLY2QT4cnd/cqt1IVLHsqwx4LEMZXcwQWO9GxIZpGdBJHsZK9L1Bv
G35m6GoxAumGROw7BPiW+pAFgQeFw14i75YXE/WkAbzJq8pn8irdO8Px9wDM8YWC
JNmJG2kvJpUTkyahU38w5Oj+ToLn7eWQs+2/KZ1G2r93pmOsHskQ0EfwzlhJX4J+
HvAf1rJcIlLvhKt1pJ1JYTCMMywtmG5CDEADvsLyLDyeNi/CAy5kT0PJ+F3ywBDS
abrK6fiF3VtsPqTDHwF+u8vxWOBCbPex7KXTdVYpvgOiEdWnjcPgaQFzXKj/5ilw
/pV5LIRATCygP435rGmYjwfLacXlw1G0Ugrl/T02CNK8cCKD3obl34fDKAKhWTJi
QelwnThufKpWxQQtyEx9ESzJvnqGxQzrE/paPknNM86drbUsUiMYvrHO3Czyq7PC
9Q2tM6ojDZcO1HhNbPe50+AlblOKyzA2odVDU+OKgL2ap5oFkJDU7MCquyiTo2oD
4qOY4EDYLoiQKW1H/cVGfrM6rtDmI12hr8enjgc98Vuz7ktnsUcXdIxGjAuKg9YQ
+EOrIa+F1dmPQc4TrQdizU30Qq543sHFK5vg1L5DG3wq5zGfMlQzIuELra5q9NHF
L6/R6lDKTvOy8TELpIoT2Cqh0rZ0I1SN/58MMW1v/QJ0FJAiI67ZqGzvWDH8ICSv
120h3ESwLcofYN80QKOSw0R4RuEMM9C7UHRsQabut0nIbw90a3MdXUX7z1FTYonw
6twTA1w5xIlrthapStulF3pqTUM4LE737ZZvsc41jbVnq8+tlIx7BbtdWMQ0V274
11OHz7w8YKQI9KL/yQks6qZKquCGM/n3O9/9syDPOyMvWGyEgwWAEHltlXm06/bP
1f/q9KcFDZRO9q3i1MDgANCVQ6Siidmy3vZQu0c3hUDM+NIu7eYAFEahE84jCeDf
fPfZjBXG5459N0KztVyBUTpaB6CpUpNosFdd+cS3DMAQM36t7son1lSQAeo3zhiw
ogYsKm++JkeEY9H/sq46kb+9xPIxI6I8p6sSwSd2bIa/ZPt1TR0QrU3YtmkD+/yh
G8BQDo2mym/zKQLXFinr1O5nwKzVwJSVQ9DubHvL05ym1KBVm1NIO9HG6GbRi02y
3GXEOZ26GePnG1G2acBNV79y6HKbQz972L+/Ag2uLzy+DqGaVA5wFl6ceJhKjEcC
Y8ntWWVDcgjEsx3X86UGS7jgWstND+qP4tGRbZnHzVJKZjhqo4uee9NGGmHKrUXn
f42XaCespivFLAz11fN1cf9lnIdIUPqi2q+XzCgXOojs6gCgW+gAv4tBTQt2Qgte
yPFIHYFt6osb4kEn4vBl2dtOqGqlqq26Pgan7r7uDz/w9rx8S9duZgP7UUMXEZYT
z99dm7Etrz3xuoVChSNIIj6AYymGl34kw3Is+vuExSUwdD+/I+o8Tv3Z872eE4/S
5aTQkjJ4F6WaCi01dJAyQV6ByOccuF3stYcH3syt+cuJvk86adSLFenZf4UcaGmQ
4OUq1xPtKkN9YaYW7e/ifkKgXV0xINWH1vm3V1DLHu9d9OFPkwK7/EPcJWyrEzZG
U+QcFpy3GZVy9tw7+O1QRD4Dn7ExH/udb6qeSVCGyOsOn/JbswZtOXry+5P6Yqgq
zmdsEKI6YcsFb6WV9CePhgftTF1a212kzXBHJC/LGSkvtQthtqliRdvaQPqBgolf
jqaozdhRRaBR8A0XKrEuKAoxc8s6cUcs2G/BBjNyOqLNZcoWBjHbHtEfHtRr3O7T
EmjVlxIjb2Nqmt2d3B6Iz/u78BjgLu0ymCUq/BvWgv3XOfnKfmkXJobwVSDayifq
d5HkdsuolZqrzugaeQ9atwMWDxbS9eJ+N38zp7r+/CZVwOprVV5zrz1o+P5Nq7ui
C+9e0Ozv7vzLTMPGtdzOhZnfXw3yn6lYjez6qtC/IiGHaW7aJNjGbdMtwKLaSbYt
66aHehssEl7F0FVObjzk0nTt3YVR8Ov69Xa8ON+rXOW0kuIsP9YakaH1HM5tmtER
VSC7e4EJgxpmZVrO5dD2PxBZMIt4cSK7SS1SFIjzDH0bCLYwIOnIYzMkmw1bUHf3
QXVx5AveCepHJC5Lk/WiMJvgWD7abIznx2q/vZuK+F+Grqwx4QOpNqFZnTW+VU3R
7cbKloHK6Ci67/rSTmLz8CFszH6TTnsG4htV8KEnXbsbUOW55iHrv0Yk5uXkFyBz
VLU4jBJ9ATTPdMZOkBLy6CDRehcWFvEqpI+xA0QPDFoVGSMCr6Ndt5ALyHY6EtQ8
8MCqk0Vv0vZzGbYZkv+uIaNrMwDHNv8Ch4jiYZgmZ0mfKzEnQxj3A3RFwHdXUCvX
aiiZzhlhsGD3J3/X659Fki+pLqd1tXX/PEyYxFjoNmFPWCK6cejJCgHAlV+1IVqf
VAYRLhhKmWYNuAIUOXmCowmYNDVOFmv48QxmPNAW3DyzPdR1kaHcKPQqZFT/AVu4
agS7n8w7nj3C1FVvYTlsZLtSW22OM5QpeF9Wgg7gWBJ4lcXMjBiDpsVqyJ4DIBta
xHVUB4Xv8CnjwrPy2o0Qm1B2bR9etmHmqVMwYJ4ZvNJlRZoqk/z+Ww0Zh+iHR7xL
ac0xNwcmP0cPrXiksMS9nNouFfdvxkfNRaj0inMCVimqemV6cext5ZeNnv7rKWmo
tRdzOp58dvHCV68k4uoEhp9vtnvT/NQdSE5btBU2r+Qr8Ks0qrVfyt1dLYLzj2aE
a1esjDpKvgbcDJm3PxNYHhk8HaLp5f96XuHChCPpL7o5SiUP5eYfe2tus4tqsnPW
bsdOvaghVWjpsayEUO3XbTZC/Qj72T2Oev5Oadju6mYGNxbr9MpdL26xyDKIbV3A
wOoLMudtXMq5X5DF3QT/isXricn80ydlLTVYuHvRvJyG6wxiexHY/9XFbliqdzu5
FxwiWPyYoGLgGCwcC1+atX4Oewxii+sLW3hRuWxn8xRt4OVcDRkgPI1Oz294wA7o
hebwOypJ+4xUPsRd9I1XE73rgbBwvpR0K1Ks0QDenrQz0E5bukdA9m4/Rstd3Vm6
WE0LphF0u6dY9kVk3OUiSEQJswkFg0VVvkBq71c3pSRny8/Dcr7jHcPf0eqTDJhe
uTMQr6C9P1tAIXyqmPvHvJYxHlxfewlHUMTy7BBFGWIALAe8Vbf2vz7urKurv+PX
HerjuHtGIagjTUwYXEXp8UXvSwUIPzAUOTsfgsqOLMKZJea7Ac4ezwQMb2JcHWtR
l0hoXmk+jQ8u0wbirhrChXBCumYpi6Ez5jzDe/L3IzVP2JV96lylPQBL719jUYUj
L79GTQqVtrPnnRTP9/PWla0i/WjIhvXA8qlQkVlYA4hhU1wT8ILkBMZ2k9iZbvJd
CTl9id1mfUaHusAcj0quahhdDdO4eurAKZHQwh4hYfbG19Ed9RHAUIIVFAnbWEAd
2krUtRvmVAHYTNpzyrKNo7ABpUFIlBCIoT6BB+jHFkP5Ye5Fa9qke9Md+PhS5zov
a4r7IZ1gtw7GbKubiqEK4bj3MgkjLiThSgwlUkauPsYrmPqlQkNEPrTYCDcnUSJb
crSDUIYkFXs2aCIRjkr/0D93cQ0kWsqqUTrg2nLmvRubl3DvCJnfI2BfNemir/2u
o00w+Md4FTHmk4b8I0Oi1nRi+KwYnHOr9I6ZJIgqz6fso7BgzBMUIn4A5lu471Cc
Plq/oHIf9vc1JTMQo85C3mJeIPVbn3Jpd+Bp2AE17zoHn18mDPZhX4Ty9HUnK3AR
JbRIwP5P1wuRj+sO0SOu2Dfo+zyxp6fOG8rhl7rsUkjXbPoh8yfHihOkFBvQWLXt
p25nMkxxdce/c3bbIce/6sojqWUNFWzk0LfQO51AHyIhGyHZmeOecD0+FNDTa4Ld
VOi4G+kuJae3SqpyAqdQAlpYkY6/ecURrsgA5Sqe3fe+5jCGj4JRncfvr76KhRv0
ah7EmsrTc5IYfBxz0uOLJ1Vd290FK/rfDQUyNrkF26LcvoP1DnX/1BjYCIb/bfw/
OSMum4XX2iBL02ffzTvFmPBeve4RP+oVKxoHgxf4sOJHDTvKKmtBRsc7dR8Vl2Ep
QJUKb+31D6s8MsRM3bFZpNddPeKNak6W28zrMn+HRyL+Vird4Ov2fdQVFydvG18W
xX2YYhgegEgNlXXnwhyVSM5y490mZJjs7KIoAm+abI+T1H/5yNj4YoYIHN3iCR2u
xwV20nsM6Xi1nXPLiUgi/zKsLOvjshd3QUXxpSgoCiFUFgXkHztQCpjKJaIFpNmb
0HvFbUshhtxDtCIUY+i+r+mRBaNPe0WkHtp/qhbEyOEa8ZkH2VBy+TC1abSHd5kc
5odi5lLEAthWrnYZ7Jhmp5cd9C6KKXyHuXeoiOYX0nj9i/PBBAEPzBiX9AL5rFWB
IKEpVCMKHlJP/XqVc292Ung4VEW+SnqbCazvawshYDUDiKVHwprWNK2z/KVrnV2b
FBoOoObiE1fZxPWNPItCIcME3SW1fd72U191zgkW1KJCIf0Ct+lrtGxDro25kns6
a1j/LOx7EP2XZ371fjrcaexxXDiobn4OzAB+C0YhkBeV1dpB5DLvhIVd7T383dqn
t+twK6CljoTRzpSuQJjj7eRPUQCv8GtjMKdkLqDWQHNJRzLDBNeF85FTt+yQxi/c
eyju4rmXkVB09N5w21cHgTj5iSTWWt4FtcAw8kopREtmOX0k3sB5KvM1YNxWtpYT
uYJXKkITS66IM1P315x4qhS4J+LSpEzGTdfbnCK5oNGNIuQvu28LHgP6udNEng9S
A5iOHEwVUeISJ4OXaMbWRLj+HOaiHmJW0IIo8me6qqXyitfM3fz8xtYUS/KH+VBn
rXYxdZEDxRAxyedmN/ovzy1vNbemA+NEkXqZbYpYnmO19y6UpzjOM4mfd6V4NNrr
D64Z3DWZcPudOyccCGf1XPC/xRAV7LfCntsHJLhI2Nuq9UQ6k3m+5laeEqfc0o16
gf6uhuzMV8ZeNQitWQGzbaFWkH4nxS6y8U8VHmX8g293JB0bGAVPgpqGZImoDYgi
F3K9WDxXm/3+n+kMISJFU6i53YT6hlbL4sBetBkYx+WtX9Es16JWKGQPM5L0p6Jv
fj63lmE79cLNffW0/lifQ3lQ0lfVgPvjx+iBBBIHadv/hYxYXM1rxXMpHYaybsGH
5i/1BEgZobS4W4/Gww9CnliVG8SAEkgLTXspegqGaPpLrTzL+CQDGPj07nhpwrRP
lmFTWQl7SPSv8DhgfS6q6xQ0TcKU9BtyyRTwNjIAwVCLdoVaQcGDhwYmi0k4HXms
P4VCoeLEt4VGF8ycQbVeZmTBx1Kdk95Da/PUXLnqJViJVqYe8BWT3wgPbt8/qcdz
26XeVa6FNbAVAgGRBuAY5Ch91X9YuyWD/p6+xespr/wSPBAq4KOJz3oVDk1iPa6X
MHJWBqEPDMTPd28KRnpn9S94G17o/HB577eu4TAhjhJCJt8FbNByqBESO0f+X4VZ
yDvmXCibpOtvwl4f6kDTAHgtXrBKO76zZB2qUsnHVvfQybg7yTMJ/0lGNwXS8OBI
WZJLgXZy6Fpicc0GczBL6g+OtbtiYX0B7atY9pgJrrbkQRZlR3ZK6vPr5vHIaPQK
bp+whvhcA8UqDdQIwBFFklxwdPggUGC/26lgIhR4J4bYOosaqt/q/TXzmoJ6vrxf
snffPUwO+PX2Z8x+6b85sR5aNbv+Ar44zCb7N0jdhBPzuBKIa89pnnc0ODle7FXn
Q+DjXMaI4N+oLgoux0kk+q9QC7ObvE6DQap8Uvw6rjYo8suC9UcOoBmISh9tM/O/
wtCstXjnPkxz3GEMbhuCJivEbo7T6et4rVhCi7Vnyah6xBQsCB82hGDYQGpUBiPr
MeOIY+VJOJMNzaW+84+fmptPVWsZk05jdTYDbeF/jFGJFToUMgt/t++JQo4CCgwd
k0YXOThcV/olEMAb80b5Oj+EjEl90sBeRORHk2TfhLew64eyTGQkHUf/d3uijO24
1Z6JDM2ahKTnU9np/SV3r2BhPhB+CJW2O5JzbW2LSM8FFm8zL7GiG46G8TlgsqQ4
wU5/zVlowLRRQhSLtHWI3SyjI/30pJlVt5uwObb2TzTWBxcggcnPpWkA1dapy8rB
sCRMsd36R8jE/4ZIJ61JIaDiW1rqwgjhtW8t1qPQP/Fp1OyQjAmFUSuUnMjppLSO
2Mto+so9hhwP23qCDRGFpfC61RZd5IowT7hFIqIHBVwNZRq+gFWoTzyPt1tfClTI
UWq9zky3Ub1N8SvfwbDYV0Ha2f1aJmJG3nogYyAE4/fmu4VmgivPduhftbCIc9MO
1i94Zgu4SZ5kxJpA14hIsNeIhgbwrwBwk1C/cJuKMxCNzfw9qEpfO3xFpSP+OGBM
/kFcP2efM779djT0Ej22d/Q+FsN76ATmA2W9bahcTBbf9NGXG7Ppi3LoheAyVYfU
mwbK6euEy2xZcQ96xj3dQLBzs/HcQCgiJFZ6m8FuRhBQQe8m+qdWx0SUT1ytQGOH
ZtaDmwm5HGq4/pBwvYa9zEH/T462MpsM9AFCRZZVyDdVvtETKMXIQAie+gtm1laQ
heE0y4YnWy8eXy15G2UhdjMrk7caD55pjT004gvrFEHW6k8I09y9eKpI7VwGDvV7
ZLjMIo9cVET/a47/gOV+302WyDHaC0dIUjijSUhsx+jQ4xmJBPlKo+PmJSS8g81D
SaSK7h/JmrLJVkLY+jBGBcav7x+VprEqyLrv6RZ9+dNHG6aqkXPBfTfGjpK/bUGs
Pd4HNHuCLme6q3OTixcCpXFj8xha9lQ7SO0y/FWH98Zn06R2+/J9FyG8q/H3SUoM
7nk3lyPBdnwfvf9xuwIGzEjb8xdzocfiXn7g7Oh+s9QrzKYlsvYHN0o7KH8Rn5af
9J30W/AxX4WvsWI+8tJvXqux+U8dHohsiVK10MeGnnYWnmO2vMF+22XnVcIf1Gs5
NGYmaLeIf/5dZskvAoDbqVsSM+0r1bjEhiS4Mq3QO9cXRz/cvw5Vft7Z1RzylsLK
gus57b+uOO0bd4NhjF1KNk3xGBPnAdbeFEdad7j6jsnecZdNN5oA+xSFIDN/GdEv
xKdyoJnt63GUOjcpCwYk94wuQEYUjwVooZzfkWKT/UwQYiF4lHmFxUgBIYb/kH37
G7tPd8jp3NrTL0kk//1ek7yAkytL4eOwRbUE/SBnkN7p1yUGxE71zOaDs/IRuqGd
5C9xwZT4L2QOjX/2onU+Q2Tyjxif+E/HjCu5Dy4mpPPoe9e8W2J3DrFFZfwLKows
K/wF7XU/RHm9IcA6mQ0ZZVO9Q6v1t7NY476G+JkmvpUV73HpqvqauX4amilRL3LU
7dnktZFzuLTA7yvzA8rsDS2xFIsUayO5Z6SAXIdDe2QfEFsciNti52oBTdT7uljQ
m3+vMptzFbWoXoaWHd0yc19NgY/hdRn5V343lTCajbPaqSK9/jS/anUMXHT2O6PP
lUfQPlXiCTY5QOOG0SdfpIUnrrwMSAYRIHh3pETG/CYfhY6zLW5+uGhf/27Q3CoB
Fb5r1tJa7HwVchYIddAUmgv5HF5uZqhAMZcT9YXlZEhHy7sshLIxesh5mg2UNuMO
13u1D4D4VQYzT7/+BY5wQCMfy1ORN6lDO9f+eDUEGX2FMnGlyTOeM/1t4y8sGTLM
RZaLYOfAo4MWpd487PSkXH+unpc9493lVBTtG0uYiFsUz7imWQVq+jKuaiDok5Iy
cK/sfwNR9W17pLcbDnoXTq6rYYWAhMLEYa5IRjbg1H20vxNzn6jOLf41HhdNuBIS
AhwHIgE8AInQ8o2bMc7YOFWwgrGfemH4qDcyTIxLfwGHZdYhkHwCyitsZ46KGOGN
bIHdpstmzZAsVp9xb11cfvaxCpDNI9XpYGxaLsteupmXsp1l7hoMQaGSVDIcSwKY
XTAje1Rt7pVi/HUlKlzxtKqJU03xTquJ+FuFIKer6/fcEMaZ+ctkbBDqx+UTA3uS
ktTS0ZzmHmddjGIGidGXvFAmVWgT23yTgMrg5rGV7ghMzvleY5RrZzMXTeetr3+3
MDoM0Ba3/PtH9U2QmzGPCiSz+BuRjh0xUyWW/8tImBIM657BKJse/d0WjeQ8LtnA
DnxjWpiXifFqP0WAwh3vz19BI34i76xuercmLgGrb8WmfFIt1hb19aHDYVca2jd4
2Xy0E8qk86znEGJHF4NXzx+yMRZWsig57ZLwhghO9YuD5It0YegX1JlWGbsM1JHY
frIq0VIf2fmKMQEEfAoNyAB0OMAG2IqTRfvIz6051C30LAoOVYWcN3SZu7aDJ+PH
B0fWU/ct/B0SwEodi6rjK3yt4YfPz4yv/BdojxKpdEeMZp2xmZhjrjVrO/9xTySi
rX2C/uXA/VV20r9tND2jV7vcw0g5PtqsuvfUDkBucJ4/XbeTv+oTJUW1LojCWXQR
sZoSlg54ow0BzCGlg0Syp5gqT21wos28GqUeVLXyQUu/XBHKPhpJICwv/LxQheE4
kXQ1BN6lN+kfHq31IT57c2Na8PVTa6vx11AQJfPjonJkZ6L2pugapYG4YF+l2EKK
8l4Sd6dHOrQAa/0S/c7RyOksb880E0QFYH6MyNBuXvOswlXxojrG8WBE2FxvSnpc
Cdc6zRBSLs4PbVCGBBPwfv41NUeKnj2jUseiamEdlJZM18YmnuowYs3xxm7BZUdk
V3VCXpaYHhvEztw8uws1mDmawTqJnTf5c/8DlzvIEymndSQuA40JpY6PGZS1iS4r
+CURycrupPsy1C2Z3GtjbNBH8rXIH60vk9L1s2h0TX3cGbBqb4FUS0VOKR6eyPKX
i1CE9odzvYDsRRNxdItZLQqPg2tKTsOkSDWjg0VfKs+7y3YSBFjYG3D1rFgG8+nf
BDs9icz8eh+iAlb+W+2H6qrn5eBnt7rYKX0BEYS9edll0WQnOw5bI6mAb63rQEiP
mWGshu1o+NUsUYDgDWHZO10kf6xv8CRVE2DaNn0KitxwHEoc0gtYxFgurV1dZCZM
zmsHQsILxsL3JYBe36WeTBG82GdOUti5/+o/nHtYHM1QkmxkNE/BE7YX77t0eZjU
eoHMeDWJ3bTbtOp3RClpD+4IhpMTGk6u5TDiMeGbaO9gYHKtIVg3bPiMj/iy+dFz
WIC9+h5unA930whmERG4OAxAIUX1Nr/EQ1L3ojZXgsigfkoW82/bzM/oTpfhoyRB
gYtASDavUo/955jvqh0/QKpf+pmIsfs2pb62EtZeYGUYUGPOmLj2flcDHuR4BHBr
JOczhBp6MJZJizD8BGb4YSKYUSC3PtJeWw55BthSJ/uYusM1jD6Zb44ZEdsstQ1e
1Jp/hP2BLgvXCtjTAGhHMudz4Lbkyaw9INW4oAX/gsfDtAWUwnoL4LYtBTcPkTo0
QWEvWkGaRSF0f47E9Yy9UyymnLDa0eYVjcUxF+ORd5yrWRq8aIUayPVIHsARL+N0
8MahBTRonYFyOw9GGQKgDa9WTcmaYjQEaVqb2t7QakqspoAQRoE7gsjg0RVJvGOL
LG3uCLimP8BU+wobingJw4k3bO+dyjTZCOaVKRkMoaPg7xRllE3liYRklwUMwEzm
yLKoD1IyllGgeHc4yX7P4cVR3XeVUSylHXO33AsZ6ByDasOh67kGvmWGdvMufFK0
il2l1zcD2x9kkVIwTxv0UmQMqCttYWo7Hm4iN784UQ46Dcv1KI3PAgTdDKWfJq6r
TtIFBbmpF6cp5BYsm2EX3T9CZhzNfsEyeiYRScGTDn5jhMomZ4uU4MJqcDcpJcp1
+mBRyGzmezFBCOF0SpkPoR3o5GsMgveUkyL9dbvXAIA2A82GdDI8x+CsWSEhOBum
4ytYLQlj4tVVBi4aez40td4aZ9hMHc2Rieb31coaPvT3918Uezc94JlQAzRpSYpj
4THNRlpRg5JAiTBVkEtBnVQIkBUhKZzBauAUUiB7rwtYeifDKwWZEzCdHFQftQNL
TAY3t+pz7qx2tHs8DYA4i0amoJtqRmS96UynDzXe4Rm7gKkiukKE/jogRbdh4ubR
DtQMrr8VnhbIJNn8hBjuW9Uf7hrZBROO6IjrsAjNkOJgVYPWgy3BE3B9LigPpviU
Ym0zv2MfjkolgITD6loG8e70NwQMmZPg/0burAyPGxO5JfOMkYMcOEu56otqQINK
xKLgmlvwM7AuUCS0RaJ2pvC8tT4fVY5QJypn3W2IHVikL1X0YnFEx5mKrCoMAYrQ
9Pyu/01UX0R2zBF7clI8DPKGo6M+4a21yMPC2HShnd5Q6tTo44U52InqhNr63URU
VMLjyPcbfYq8oDp9df6MsKEVC0bLGJhG9NKSqxUeMFp1MlFdg4FMwRQ0XGtYz6gk
/YnuG+Wfsr/ONlE5dQ6RvyNajcGEmujSp1KW9/kfjijuQC4wDTqke16x2dlOlu+V
9YHX9jEFKafuF/2OfjpDfSd7qR6Bc2/IuKC+wgU+I991PbwtT8BvX7vkJwK0Y3xa
YfkY+KG1vsPkOc/Pi73MixDslHEgUu3DVzBU8p2Cbds/c7kdqCoxsF/3XknT5qwD
JHVTb7ZzVgfcaaJH/SroIm085wz2Q8ajC2XdY4ITVcMY1lA1jTBl2JXqE2C2F9KQ
rtMp/MX8vzYKRoosOYFYskvdQ+NW6q/2lQ9cvrPc171iaf6w59QJC+8RgEEvtaMx
3JjH8gBuq4lK1IEhq+QwY8IzB1Qg5Cas5/aJSgH9AC6+qjvNDfsaoYF0tb+I8Fxp
JGNjZzhAncePe82aZ/8XpsOEZgDRMqAiSxpjRxJLjBMbhBVNrAoapWzWstYnR8sZ
D7o8jOWcld4RsG/wuvAe/XGIxBNSnV6s08+dYz0F9ZNobUi1WaS7tbrgpvi78d9r
vJbG7EZI7GTKo+OMB7Zy0lh5PJAhfjm+r5y2pZNZvDtzASy3svuXcOSsaGV+R8/K
NiqiEfTNTVF6ydVnaEwnAafQ/xiPQGxfZ9dkGdPI/lXyCIsVLpWHZ0+DdjF5urnB
go+UecVzaTrVIRnutlF3KbJgJKr6YhCKGCfbt5+JqjAiXHHMdhJVeGsAFaG7Zucu
+rrfsTNFbBzKf4AHfHZXcs0dSiKAyxaFDThz4vxH7VC4SjIX+L7Du7/YfNm3z3AX
gqgz6cGNvnJr/PSwa5bNyiFgmRyaq+XhI6KUkrw2JdEMoxYxf9D6z3++dhaANb2f
yYvFTVFqqw0nw/hQNmdNF+YRUWO5iURLErsz2x6PPiW3qhiMOR7nsbeCKPd933Nw
QiVjrqGoSdYtCJYFRZg6ZGgrbOLdF+68Qbyukoqo4NkuA4fZmnc1TEOSa2k5o9xd
NuHmZl0uqc6YR8nDprFl1BQ8n09qL38CRfNvhL7SN59zBnYjvVABgd4Tbz8OXp7/
pdbhSK0VUF/VyrVhy64F/zQWV7S9YSmUS9y5/cf8b2ASujUqe5yioYOJvCD9O9jO
4nLpVCaYmJODqw0rOAjFL0BA2anhGJVBATElJY6FIfNAH+zsz9i79b7bdDBQI+4w
17AOH+5feNbUhFBRBFL18xp8oMMG901MZl017X7bPdEUWw5sGpuZk71X6PHRV68n
y0oDVxVs0vf78je70jOis/cauW37VQ8Jiq4T0q9+saMixmmm5aEGrMeW0UBxgG+P
2DpRXONCawdl6cxLuvh8PehZ/czwEdd1KSXP0mXBcDG1bMn+UR4YQLrXvjH6McE7
PE1i2lUcpZ9zHmG8U9muk8l0ftpay+2Mm8z+66EAfyZL7ySyBzL8FjVDwsQHmU1G
kcpT/05NLJsdYbLOZ22jRxoe0k5D+KlwXIN+xyPSoZWPHgD6aOYsNg0EcFS52tmg
/pNgxK1LlGDJlzzQJ0RXX0DUAWeYWdIDsAosSTRPStRngsgQhiZk7U3QvxKcLrRg
YbsAlQ+Jnhl9n9zF606AYxE7JDqzQ1UCSYGZ9JYhQbISMzOUMQaJMBA1mIS3ueXx
/5s3eX0hTSKGdsJBDCaq5wBriFvGLhfmueVObawgbUtd/AlvQOgxfsieQB6Ls+G6
//NsjHusTB5qd7lHDMA+97HdD+h2KzEFlgfU9MnbmqWkjQSZgUaZyxyoWc8uDYAF
crvJchc3nrmhg1yPEosKlxh4iqu/NlaMApnNzIDy6q6pOklrkhd+OCpTYfGosdMH
iESutCY0Zp41mY8ytTKA/gi3VE//dBztOfA63Tj5j1T6luZEkEsw8poN8Ry9/nmG
K0738kHdXrsulBcxfnNbiv/tCjiIbCcGjPw2aL5O50JFdQYPUvIJ+FuK1xmxE55l
+4m132d0q/eXHAEqB4Es+rW6nDFJyFkhxhmpLh3OPPRFlwm1x0GXqIZfdR/ZhwdC
qbJCZXzvSljg8V8ao5ax3bxkZZtv8IIsEh2RlECcsd+cTarAUAIWMSoKJ3CwVq//
rwGurPwmPqribZYBvAYNR5D+04gyF51o+pJXMvZouLpqt2gS8asmbBqVtgSxUxg6
VPWjj8jK4u5XxYByYnQgw67Gj3pisvRG0v5lFlbAt49ymL6NXAPz3SNagKUh0yKZ
SRvyHK6bUTemWUjLeNXNVVQGFgSICz+zWntbGVfK7CQVFaBxC277Cs7KyPgrXdh/
CM2kTWLUAklktV6cXSNy9TaAjQrdekfkD10VS5s4e1Ho6mVl0291S8RD/jNSz28W
T7dZkHM2e19tWwC5aZL8lMvqj3q6Ve0rHK689K1ofdEgEFECWpidNcJZ72C92S0K
XYECqptbGxNr22CHYgGFdvZYC0ki6eUIpZVe8EtTd3OtgAs7irlEaZC3PRuRlgGr
7f0B/kaU4JWy8mfQ2P5/PKxLKUHM/0gif+YoStznwsrDC5AtOF4NR4+OtGgu9Lwq
+r9ik4yUNcedKaxy2vzPqnvrs0AfdMGJDm90nI8H0jZdgr8WJAjr4Jcs6imL4+Bw
WJ9NPrkJ0RlpRb/jkwuCApiXwrw6CVnd2IdewDqZQVJ8dCd0DAPX0na/LifjiV57
VBrIqaXT0UtvUuLIejajtQLVK96kBJQrpc6M2PmfSaqKjHwMj8DxMdF2JrMMtIUO
MZgv+CLAE91UCDYDK4NT3m7EaXCpGdu7gN+XaHA6SPjBx2XdffgdQQn7vR9qSam8
f0TzTTTzgJvduY9b12UhompifI+RwTQX16V5v4XWt6Ls5IAHbZn2XouHrLBI459l
vTcEemHwdX+jLIxEYBQIsx1Bx1cvM9LX2em1JrKTuSbSVfJK0b/3mWnFeKokQbNg
ikFMsv5o/ChP7EckkayYTSJDiebZhyVspJG6kSL2nYNA9vR5YEU7nl0XgdBW7TP7
F363I7MQN7C1reOKaqR3zoiVbYsz60mfd0RwTi2yqiBzzJR/rS72FVHauzJrKdi/
6F6AGaHLlSjrITiSsq839oOqxQIiUsAd5WAaJbG3aRaj7+szzOgMf5pNjIVvkRe/
vNmAjpeSLOuqXRYzLXQfKnPWLWjfgK3K7bp68++22coAH0X1rhEbgM15IVJTJxbB
UdwraRWC2IS/K29fKE5lKJ/dppG2+HKJSm8FD2z4lsit/1QmlY9x+udXnflTvTqX
wtyFPcROljhwLLobbKunMV2kFITrEDyZSR/5Z+Oly9wXY4KADOhtpmkzVSetkaz9
V+k+UB/wYO+LvH07B/i/kl6FuTn/GS1Elw5Ron8Z2eg8QtDTwXzJfsNr+4GwkOS5
Py1ojpBUT4VraiOvkvba7TF8yD3wnjSRNSvvfaeP3OuNTwliAjcgn59pVG9PRFAX
dwDhsyKhGKVMdeCGRt9giOTgfwywb+L8K9LbhW4AK4xN+iVvMuUemqQsQBCNrZTi
L9KW1hSdb19aSHenyqUUm4vsqmicjkODA3ga+ho1yx4mQiQ+LoAR7o4KpNFKLAxg
S6ucjm5fNaa0+zo5W++D60qlEuIsNt5g88D98+31N74TgvhtZWEN8/+oMvXeC/Ha
s6lvDmVGqxb6LxHc/IG3JL6eZ/arNwza6Y0dgX0rp9UAGIAOCs2xtCtLWbmI8qn8
MMkiSTZGIIwbR++cvt6FR5XCIg/RhbV5nsOUOhfwyRIW7ih5P3/LpnvbidCI6m92
BbYyDRhpOr6zvctG9aBfMJtuxFbaTKhmCYYovDwXCblKU+qn4GympCY7PJyX3Rhj
kEEJ9nRs/4n2UlZgkk4Xkbuh8kKDCRGuqu2Hspoh6nvvLi2T3asiPSiap10+Wiox
HQFoOV89tD5+PfRSTDdmz2D1SyG0IGI5KdT6DItBcCv8x0Q3VPa9xTLn4oigbjnR
gp/jtUvF4vt2+PVVrgDhJGwH566hLMdSQwzzUvMDh0VcWOe0gPWF8JMyh8Iw6BoL
R4NpZXR9w3mVYp5tospOs9FvY3SGsupaZoAv4WsbczflXRjmtf4d3vdusF3LE+zw
V9RqipRzfTbBee1zu4tLhW7JHuHet6+HrLFHMliQFYgXMjtFSD4vecs0nFgNT5Lz
LhGXnedBySxHhrU7fJoVBvjEEZntDkijcdKnHqLCrqKJ3/lMIQBlOKiTVAe17scw
1xCoR39mz/3wfXDBTyooAiVbal96ZdoN8TVAaTidgibxXAZd5scd+koXgesd5Dmk
R/jpMDV1cxpyf4p9bHhdJav1mo9Wgq0jG4K7GLYMModUptptNRTVn0+hYkmfG3Ds
Yupfg1CzNw50eMCRhRdpsnDjiHYFGSaalKjGmh+OYrTbGUcI3FqLqsVyG8urwb6O
zVu1o5eRi6zFkjnawKHiBI6MoCpWt8g1f9ecF6avrJguaA1Gau2HJwBf1Cm/lI2O
vZU+O8rzqFHBA7JL4SZukBLLvXnU3EWZuDRwHye3zdTPjfYA+uDc2HGN+kTqG+in
H9sjHO8eeg63WatgozJKmP/NE21t4mo6/kTpUGNEUUkT+4RkYl3/jfHIBdyr87xu
cnlu5evJOUMSh4wJY5uC0lmg/wOwqM3PxagO098MW6DRcw0ZlDJI9kVCBpuequqe
hSbxPeAeOhiybsnsfuAmELjLPlHUeIm/jbg+8YB2QR6uw4ea6bFPX3N7PkLRINgL
2W8SCsliAOlgZtN9UP7Er+ohtjBe79wUE2BKWpFWp16fXXnNL+TkFsHBfbz1BUGm
EFceGLqwiwNSK4FApxB+yJWchszmep6i4rVBCZvba0bGTYF0UfA4ZYxmunr0Z2Qo
ONc6+a7lLWh3pcxhZLxqrX7NsvR45riURlOHSojMh4nkQhjFCFKYsoSnUU/JFpf1
GlutVkZIE0PB7ZfA0uMKUxe9RGrUbq65LB2GoWu18v/3sJvzWUQtP5jxKe9NMgX7
/QNfcccGMW6OnqoQHLjhhoCJE/fzA4PpT+y1DkoZoDwQeOdnBTDTXbjLhP1ABgbe
zoRE2kF0QVjZSOAJgWY624X2FLW0fsWNVBnipT5z+qcdG5LSuaAetinemeIlXlg2
H0L4vVWokuRezyFrpxWFYCvDkB9PflXZXxsbKLLW5y/Kkpri7B2UZg/Ry24/lIJG
8LDajWZen18fj84InUqC9tZ55DXJoh5YwfT1a9IfRi9u07AfR/b+x/APjd69H5mD
eGhxCYcV2aXHQ5og9u/caASM9I3a9W+uknNWvGz236iaLqvAc1xVNF4zqTAWHraB
/UmvnEmKdTvKmL73XCo/UM7ljB46CAaLRUCMhS+FX1lCuGnHPGF1uISutaKutmwL
tZm73KW+QDO9GvVD2pAshfp+TGKo5xPcYSF55KhZiLUXONJgh9u7Hb3K/obBRuu/
Nrv2qfIfBBwOgNBMcbocdIhCJdvve97Vh67k9Ukx4q61rc/ZB2YXXatb0/3xYOCJ
YLlYR0HVGJ9kRxUMlibE4gDeVwiVwbvhz5KOTySvf+k8XIr2FmBeCkcyoalniBzj
oC4jd/L+p1D7XM5nVe62ig9gHOzwJVpsQqx7rsYIXCEVirthdC2XMxcSM0615TRz
LoEv51ZNapCcKCHp2Pa/rwQs7Z8AghaQqaZ34wSz+PtdSSShVMbvc6RNFyPF8SXk
zl82PfqF4UpXOim5z0o0Pr1lDS5OkQSoZ0Ak30puCcel3GEGNguzhCNntxHrk6Mv
08m6zgB4XIRHLQDhrJObiR90l/3fwIbYOOEdLstSf/DCC1quHgt61y8r00Gw3akp
55GB1yj/Mvcz2d2KezczIMoN+2c/OxcO2nUVMLIOKfJhu3D3GHf1bTSbRUCYHWIJ
EYt4647owAlP+ZQ3OFeFbAuhASQhzHN1YqMl+D5CTQr3Vrk+yn66Gs4vaK+DfdHO
Q0an/1sB5pDFzKsKPRNoiSzj4QZVKjqnpAjdApEshQYXohsJURpKP0bYa+d2x+WX
eyUlI0rFKbNvNi70V84/71NBC3+qpknlKsi2ryG8iIEmseouuTw1G4JEJsOnf8PV
///q2uAj1kJLfwjbtkVzqiKQLd9IIgDccdLI9+s/QkFwY1oB7erhTHhrpzlPB0Le
PV1dwCWlGtq9eXdAdx9VyBvnpYBBqSXrMbcIom+Y+DMFdpiJYgjVT2PxCWXFkXSy
g/YINx86/CCKbH3TbG2wUA+PbpVbktFv9ZEjtefy83cTbKmsJ1peoBXWIO7reudP
4VvkVcL7hjmvSz5OcN5sJhFBrg1g/w51zz3TKj2xfC3Gwv7nX0rYnKViURA5mbca
lWOr3UJM8Usfexkrpt37FbGenAnV4aqgynFksG3x84HzN/oDrE6kZx5MCT4yeAXs
u+34RxTsapGb9/AZ1bDFDSNZ0oNG6oaLIt4VsPe0P7puO2ewJ0pE7WBXAKNRIU1J
j0NP9DDFNgaIoaVjwpmszfnQjgGOcJJF7js1JcYJuGbtF2OW4r36pPJb4xLSfxbe
H6OxExqM6hJ5kSml49uBFK8e0G8XN7iJmq5PhvL5Jt18bRPaDcBIsh7a9L/ofH1l
YK8yy7eWNsyGDGl9br9V4W+huGa9lWHIzit827Hq5KqCnOSnarVJzVsYSWnpTibG
/hLv2dXYEqzlQ5ZwYMbpkEBLTRWfmHcO3lAs525L4wI7FNYDumxvQZ5IAN3h/ipB
xw9yauZsvQHqQ4WySO6XuKD7Moppp3yN6pO7PrQFREF210YSI7bbjuKQJXJz5w2c
rdXHMjdqFAJU/erBaSr9j1G/JbnZZAkfD8U53mWOAHQ8oHGDRG3orVQW5I4WPuVJ
mEcYDjbLXoW3OnH7g/mMPp/i+Eb3vm2Pu3PvnZyuznrqHcrh+3+fyAcCqaw7/Q/m
Mgts+RbEO8xIab3543dMIGkbodshwPApRSBDH8PLcLlpkxxzIU6QhYjJm133SVeR
lHNI8XtSMvV9ksZktT/h3W5Eo/xSR7p9YRJsVhQcMACLW7yidqnpb+ZNwaUAsCIy
yQczCVvUIQuWFxg9F8RIBfIOV/B/zvkcmOtOak8iNHTJfh2kS6Fy/iWyTOVthjQH
lzd66AuTXuY2hdKxGySg1GEKP7C58tOGHp+EAxm5fCdua6sAB4yp5KdcAIeENVbc
uOKsN7oJCkJdkvHO6IIL+jJpn0wThfUp9ahhhtwpA4S9aEiSsV4FsuLZJPcrnbap
02/kiGRgH5l94B5Z0+nwYrHgervaAbQg4NBdoFOBRrvBi+gkQQH5acKCHnKMURSR
g+YQsyb1Xfd3CGTI6cc6Xu/q4rlNxulLajNXm4NlMygliZOy4BoMTt8p7fXssByd
aVYE7qrZmhtRu+RFtd82RnzeR0Wg89B3f0oT4TJnTXDj6S+8w9hqMZClxlIj7piS
4spce6Oyvq5IXz8csSx0Rn1WDQ5A8T/TpPBZ0LcJIWYi8b9AKrffSNx92bxBg0/t
dNuqOh5tQcFZxGHi8/vUgQaNUtsOqvmM/z3F0S2DhHvTvEfD9d9v+4e8K1NgV/lR
LYYx8NoejSp8uWp7qYhGl8CLRAAEDSEVS5SC6aywbQ4w5NPWZKcSFgzPTR8sasLJ
Lt0il5bXJ55IQt+DjcCYnp2kI0y0pm94138oHothLUHoHza0fRVHnVyFIo1oQLZD
Wkn14Oao5Zl6cLsk+AGdmwNyYyMSsfoOYN3Vwy/2FUjp8WWn10knzZ2H6JXcCZnG
UmaBo+LVqyl9b7foKftr1Z7lIJwJmDFnJU+8WnxzRI5pjFEn+kQVep9IDTlOuwBG
3AnrMFuYVK2ZFoeO+B6fDMCN2OkVifdkBTOkzeDFgsO0BUA92M792IgMzmYWHACt
wQtpslG5yq3BOeMWqlyFu0mhgKL+G8FRRrta+KaYVzwwu5gp//hcn6q9WYnKVIiT
KYYwu7KdBIg1bS2IkzQp3DO7fT6Q0y+0G9j3IwIJPdrHLeL0eNdchTlc0bizU6wK
g3En2AoyVcuU4myY68OQU+wPiRE+uhiIA6x4GOdJvMuAI5MOv3PKgYSj8XWQ3Wus
Zxy8WqtyyOAZjVSqcFdXGQekLBk8j6mxz8yiOiIyUbm7lTJYzqyBXhiMMxrX0ZOn
3jo1xWNNBauwqPJrJWJKyvqNMUdNNhMoEWuK5WxNFefSepx3CuPh6SKAgHsZiDhZ
wzlONakl9+himftVQ3x9TRT+ubQcRjJyIRD6ZqJcHO29aP4GYEcbnJ+Vb98mm+Mg
+LdNYF4P+npx0OulAb4OFK4i2xKPdJN86iwc2/VwoRUPh7Jx46xJ+zOZP/CvpuzE
7PyGucjXL093JW8Ih2BWYQD1fQMuHVHmOLAReC2iUWPX2veU3VmknHq2VF3tg5fN
UDxMzTrQGfwU9x3MIfDBUL2qp4mssDuf2W9xHni3oQtdnJiUHndytXSSwVtnmMlA
N6gfu6Fd5kb0TWjKdJf2c2avq1wYGFQBQYtCthnW7SHzeO3TDCdfRl6RaxpXUoQS
KbOyHXW1G1oTxJh45yNB9idc1B+bt0fxAjVNEfr3M0IeerrnFSSh/6QayOZ6/LIg
kjcAqpZUSyaY/qKCukTym2X/+slemdqL4ckWKDtKgHsfVjI6FUHW7vaJSTJk9ff0
9poOcRbi/2ckU99TsiXj6dL6y+XHt/R76Sy9qkMMee8xFl7hrsAMOefbmOEE0fIQ
jkOtYUqxH+qTiVozNl3OiksTI+TUDAuctXs9/TkUQvh+CinN8EoR+4sD0/1LqRxp
mwiB+pq6qIJpVfjMqclmIkVuC4MpMqs73O7NABUYUduIo7leRg4fJpM4Utfkfava
1qJDncljPbJXscOkheECXfnIuH1x3pzInTnD4UeLBWyy849KTOAFGy6VmTJDDJjy
eD83YDxmqTgX26LVx1IaZagPyw8kiSbElrg451Op/2L0b03t2UeOBpvjjmCP3L36
na/D9a/n7l91kwgRvE9b7PnHrIUrGvLpClUxnk9uEaDCA7rmRLRfZh4ia8W4EsGf
XNUsggunyqaLoj8sWZjRsGdDRBTp+dy7yD6TYa7fGZOWzXCKNZsx2PJIXIEau6nG
Mdb1nupaIHvhat5yp3XRX+z6uocNlyaHaJafYCNSwl58HP9GBL13nZ9gB5URyQeA
Mki/FVawFElprH55TCLncgrPLNRWHEpKEeIx/KcOsU6GxjsIVq0aaw/t6PRimjsx
uZ95p2cizjEpA/QEcEnldHY1PR1hIO8T/ejIYeVf/7+sgv/QDyDCdZ3L0FJtiZkm
BPJHWTVe6/dyWtA4/XmbEcR8KFiw+uy5vhDBOf92gl7qnF3lt7QCxVp8nKShbGKQ
IvDOlO+SnArFZW6BG/PXYVHCUvqzFheth3UsdIegXMTKEts+2tbgEn/YXn1065Eu
rOB9b5ahuV/E5cukYrd0iPVYlbA5Qo7/9fisThNigPH+oRRCSbRYWBewZbpD8YP/
7kfhsabvLgASAmndYGow00JD/qP8PvC9ESaGEf8Zzx2R/BohamJjXuyBIKDm9j/p
VDO4OVpmI+IpYdDmbyUQ/QAwQNZP9v07jo/tzq951ECek5gCe9bcspOg5N5OGuYD
tIWP2JpXOCsqOj42Nmzc0P7K72coDbOnqm+lUttJXIn8LpU0ORVKqauTC7Ewgqz3
W6PUrtD37Lu8FdGDZzHrzpgyv08Wbgn4QUMG6EzF4DAj+9ame9GsO/b1+ro9XKuU
utAUUzL/Y18BWG4dul2TX8s6Dmb5eT6Ypn96x/Qd6qsy1+0YC1CKsJgIfA44tj8j
n9kOJ3z4Y+W5Uw31lEh9rnvq6q/bcFN07o4gepJ+KxA5Q3AuNZsW3xCi+JXbWQC3
OSCgbu6h46vGuqln539E4Y3HVi0uUoSw+obvitVc4yPlVgxtxFIJymKbOrqrDuBj
DmypfX/vdGsrD+6NWngrYSb1inNz/GAHBv1LZpAIygNeVtSDuSo2v+5UAk2kFFDb
VZ47jJcZhP3AtSqr88Db7DUv5Q4Ay5Ezjr52GIHwks4mh7V9siJ1zRx1b1s7IC6B
KibGrtsG+GES1qfg+gP/jimumpGHfkGneSCVLIQflQLAtaYMuJCXaEyFe3NrV7CP
K+akS5ni0CfJq2MmkpkzaACNdCgEymdWxkAUrofYUKupejPQl/j2RYJRiVe3f+GL
TRU7N+0XaS11WDn++YGWPYnjGrlfDLvBeQLmMDRUSxiQLTCacmxEps+0jDPcUndX
epgn5Rg4WYZCdTAN/W1cV4E9b7DetQu1gqc6XxDyw4djTFjNo7/Uxh7FwnBrTaEj
k7e0wi/jQo8SPG74ZerGi/J5sFuOHSeMEPMWS1v4GGbUUhFlQ+ig8KOT7rZu/gLl
N4OTRivRTHHJ9i0FambmvV/DU8W4olSZwZRTp4CfIOot1dsNLIJYAnENRLXBApXt
FeVicPWb3LPpnIAEuiuQ4a0FICeVJ/jzv/W7JbVOFHqBRMEwWSN3f/xIsRsh6oO7
ZukQOVKMKw2SD3q9h38q9kHy8lpe/Z7ndipXJspzLMoRuPmC3vQ0/xWgGv/6wj5Q
sVPpBAhw6vp+TQM2tjxcYbTDeXzFE2J0LQPhNB5Kvstne4dyJeXdQmDWAIViQzWO
oynVGxxWT+0xpFUaCEJIJLYcbUCFm7kF6FF/s7TGVHSJFFga0ZNXx/2IfYlqsyYH
j2VP2YjXnG3k4MCJjd4RG2n8X07UX32cM1bloNthgTtEqVp87t6UpqxQULxIsMVg
RcoHZWfBADKXYb5SS2RrvZqb1Ld3kVrTwA8YUwxljl8dbz1msbgTT3BvFtrduAuS
UH5mlP14Sv4fxJhjwFxJjvUzSKxkVJY0TowNXGav7qlY120aw+gjBvsgIgL34wfK
V6WNgLsBD/o1vN1nJjBAEU9D6Fe+gkNvT5KTRGsZNQw6gtBtA4/02xBmn21bwqwZ
wOIDRC/VfBKdRnckEtYWf+Tqo9IgUb+2zP1gwrWmywnkFvwtihBeCyT0sDGFtys9
vzpJPmlesJW7AYqvCDHEQs4aaZ8EoQBQYUqTa3Ix1uZRiT22kGkeXckvWS6FUdgY
h4fVjw1riyCnm26MB8bJdaUYPfkTc256uVh9yFs3fHNxDaGGoOPyqbKL0h4T375d
Mc4ZPrdVtKRNR2Ggu2jCIEKjDxORD72YYSB2gA9o0uMeOyvXmRhjGKs8558XWgVp
1QvIy2N/hl1APhOA3W9pHXZehQokjcscwlK8GpDfmYe2yalY4j8HvhAi1tOZZTUt
f4Ysj4uBrueKGgK5ZLl6omYt38vfrGS4cEDsZZTaBYk8wRYWQkkH53xtY3cKFNxl
/6R+q6biDp0FM0aqCn0OEAB/lGMPorP1cjY0RM0Lq/qekH0YYc+LipufplTwnlKv
DhQA6ul94kGf/P8s8jdLxLiL6aSOjGP7DhaaGN73OUiWcE+txop9Quzrxz2wlTrb
UdkkeYNTkn2ToQy1Ud8LbVt50QrN6s1gINaUkExg8kBHErN/LABqR1skIvKvJ+/K
OH5O8ln3dLMSViU5UWSaZ4ExhkzIWltJSF9MTIt5KxXZmm1q0WzbBt7gOF3CQjuB
eROpHMYJ9P4gteW/gkaJGapEwmVikM/l+2URtfj02K5+AuYVHjCcxUIoWIO0qv4d
xFLjlhZ3denz1D6ebQLkwkzit+WmG47NHGhhYNjfVnAoAExabntR8e0NlpvrhZyH
qhg2OIO9C5L4Sdorj2u+xEcXZJotQhcsdgxfyKbHUzFYag9JPgva1EXU7v/PvepI
RgrNiq1UgXuAjyp3eVXoeqLp8oJhq6eF+OzQbQD0O4PmecX8u3M222RvT4MoK7/g
k7rmaJV5tFpYtkLqoMMAnfSry2nC+PaYSQkucAR+q3o+0xTvdALStD98DcYBSblM
OHEigI5r9+mWUctt+Lv5zvmdheF+bgMLoXflAJVXt+PfspJGIvYmG8V2gvHBrlQH
Ad5iAODIOnyNtNlkelVc3adbE0ZZfPXRwvyqjiLk+OcPtA9foqxpnTYUL9XyQUKt
FOLT3EOtqQgew44q8b7B+xN8BHHFE7/ftbgkyXogkfd0Z2cq8JxYQmEEcTHIxZCD
0JUwx33XqiFslGroVNEqJxRytz1IxCX/kwT5wgpdqBDfKUmaJrHL5aHhHEyIuidd
xDEQBXlHLWHCtq6sS++uiKECPFWu9jyMdO+2K4H8mPiAayrMnLVRCqGNk6eBvyei
kw+iDUt28/86sQRuHUnA6maiuLzZnBY5da4yUa3p54EcbLlVipTgcgQ2WDZ0PtYt
rb03ArFEV/e/BWtElkoaW5kwHhOrhpT7091Mwreh3yu45n88j9hWZzKXrqU+LNs7
0PpV4+LZ0pUFQ0T7fvraOKnGRyVEuhXZqUBGb52oG0lqN7rycFXxTa+/vCB8mrAP
EBbil8UkCtUrd4GbFQBGb/lT+WbfIIeMdlICQF7ZR0JUG/Q8tgrtmW2Fdjxt0vzz
BUEsdv7dhwLuKE7pDFh/lg5ZCLpJZMMmjVbXSpWnCDVHOP1Nb6EzzVtmLxk8yTag
E1Te67k2vzi8LtayzhZ0YrWXK16A5Hcx5cNuk2fqn7mTpqY5pZuXubaLAUS3x3l9
DO1N2oxmJptLyCIFTE3bP9MoXZSilsiQat6X2s3yr+vsVIKKg/lPhTDFO6xA1++n
yvrevppLswNmK3EXHkp83rpYkAIslxfk55jnP7IbARmuMgfq4LwE8kPL5+YkewGu
as2/hTXtXXgT7VwJvi7n8aAiS6AIadC70IhbRipvhCQ2KrWCSaXjcqa7nopOQ3qT
pnI+PlJUIcLh0kPz7BXxVJc5nligNSqugfioWmMBJIQkHe2kez7yemrJqIAPDrpt
pl3cpZ1wOvdyJUUdaXSk1ScELsYwYjsmf8g9B31GiY2kdqL4+AGOl+I58QMeMCeW
KXLHRQK0B3LsW5olJ5kZLh9JpyicpP93Ne6v8nb86pC0m8i7jqyAUP/h6olv1J/+
VBToDql2NCFAQP1JI7lHS1bJ9nS30e94fCJOohfBL6AZH5boF60t1yBOyX5nTVl/
Uz/ygJ9D6fZyTeROX+7S+gH5gR1MvduN6oeygid07D1qFgv5tD4JYKCmr+L+UrkC
uAuF+/C8XDD6rEio41RwFI3g/cPqwhLdYij3hOfwGyrWwExn2B+ScnXkV6tx1Yj4
oBfp3rRhS6aSWX9A57ceHyq1dkMziBj+a8p2p9xBFq+gAvGV2q/EQs3F7wYddDRL
SatKIgfNuVwZk9Pa+Amk30LTaCZKfw4Kquzh8Y+YpONDasJwqeEuewT8DJueUqSW
OsXPxNRATysniguQyp5qzjAAAM4A1WuTZCWnx6w75KOP6tccA99bMPHsSIJVo+9n
cab7r0wHfCg/0W4my1gadAy7QnlKHE5KRubl9UtJ7yQb3EeHmmxAbMtC1qNBmMDr
wsgczkeCHjb7wvZGhBwGk9QGU3lztR9LN3NaMaO41s86lGlkFkfnYGWEHaFRm8QQ
Lf6eNyV/bb6zHVwYxjMKImuOMyZZkaUmP29vfVh7JJeugbC2G45P/qZO+cxwGbs+
ODTgEIAuLKIBbfIQZWFKpeSLkXbl29cyMPzHS3BwQFmL54ouhWc6VxQWyX5DqnuL
/hxzhdKQEqXA9d/WIQT+153Lct9AU6jMG/1LBeu3sEsZ93BwVT2IHFRqfh2igvWf
28LUF/Wrf/nY4mXx/Oj2dLKf650+gWoQcXA3n3kPt1XLwI/EHcV6Fdcm46KQ2I6O
mP3h/6Lwi2kDsbe8kfJ5Iafg/FG3Dhiq+EwbyQwPt/QBVTY3dowhcU1HWrjJEg/T
QLEB8tFAYt8sVhGeciWAhQs3MksZlCJnMJKuNmWqgYGTkWLYNbat2ebiJz1WW5Jz
JaecWPc31u9UsImyS1IY1Uf2cU2sCWQeycc6N5Li+S3ZIc8XHGolx0DTN2jen8KB
2kQbK0pq9YfPufcDtbXtIW8o294HGjP2EfRiljTjYvX7qO9h+rhfrU7KAdvOl5bA
yaX24xeDzlquLg87f2JjCE0HtcaRk5gtosAayWiOOsORDxznuHCng8WMz0g1bkvL
T6kBXpuFYx7V01gX4EDavSvGTcN8UNmmp0tXYvN62Lc23wwFJ6DKekkJX7eprj8C
xmb0VOSTyYhphYL9mccJ2iDYQsXui4at3q5FjNN7jGcI9oiQoeRh2Pcg78TFj0T4
vrvhjKswAWT2lFBloiYvppt6Q1NKnDd/j3pZUavQK5MP7KDeFj/kHos8MQVB+LdV
u1v4f5OeoKovlu60MJ95cY4HKU079STiv8UeBdaXJdkRilZniaxAGh9kKmn5CVUl
cI+FdZ6Nw4souq2d9SWCt6hX5mFsSCJ3O5HdPVNGW1/gUr25ah7zPgYZH8WPUpV8
P6NmdTEZ0nmRUVcCrqRUkbophVNs03jlnN3VVLCZwjxZhAy5hHSSsZhRC3Fdlncq
kCDXgvoCN9g9KbNpw6KwDwlObw3KafPYAnoJ6frq5dqgAeWzHlJGT9l6Gp0JnZJQ
3VBt7l8FUl7qAfMZ9B+7dH1xwH7N3qWcRta2BPxd54pmwfQGEQ1/bYJ108NyziaK
nK6CSDB+xqQN4Xw61hSLNCeX3bTSYz79hRxQG7pTwJlwy6/fytVqo/lN0Dy9KJcC
Wb6/P191EeU7onHOR7WXK7GPLEHMqS6NKSxYtp8dGIeMBQpRpvmmKvIieXuC0PHX
1TTyYBcyBeB124491NYdhXHhnbdgw19jQRYpwWV5QWeQpR/+y9VS9QxZ949GgEBH
H0lBWFvq0BUdPYpyVe4Uq8JgsUBm3+5A28CbCtgdrj4sKzzd0Nh4W/iibQg36JRL
mfZsQ8YErkwO3iJePi6PWYX2bL5VG+BHEHAW7AcBYMTiOhFdi70lycqvOUp2wvcr
uNgJUhrKECWHKRLmApVcRHVU3EQGY021bU/CyjbIeMeBmbB0TtJ95lE7kpblzvO7
EPC19Qd8+B0UurtjSoWmhJ6fU5epBrJXBJ7TtrYNkYMPT3xf2zjePuqzaWDD18C8
Qjce1gccntv41879m9gOrAvphG7Y0/QQ4gj3DBCYXLLd/1tqfxrvCzJ0KN87hnxI
S/anVe61WsNn7pVXm/8gVCNjUxgmrdChMNWR34KX+jR9WTW3kOLRcRw4U/F7bV79
0/Rv5+DHAT0c2UdNlstDRRQCQuRQfPcUxF0VL1aPdS/JC3sSitFv2SFSFcYxBLtf
K4dP1xta6NOuzieMrKNE9Sc29RJaiWUL8ex8vWluyKxp/E959JzRcLuHM+Fj/lnR
JoJVvxz5Bx28+WSUnrcbfhfro4A+pJONytYvvN6X9dQseNwr1Op9NPQx2z7o50Gn
86R+slYRXOWuSRyIAj3BbJT7gFQHFpR0b7zCVqXTr1t+u/yoWL994TaN+6gnR7mr
/L5S0a+n/voZStDecVKFXFL82z3xYG4eFIdmEKHY4JsK2o1sMoC1jdTAYtw6qKN6
bxkhOcNYb0Iar4ckqi81/9C0v9eji6vgHWS9WBGfDILhLcu2y/1SJ9Il1Jw71Xjs
wMORsKU38DPOqoxESGhJntO9XmeK2AbqFY0nZAsKo8JYWy6yuiOn35ri7qwTwxIY
Lm68nQONgtRdVmTtNXQ7mZ4RjoY8XflVkapUpy7IAImvn/7y9agUDDx00QYHp6P/
ZUEEGnA+SmBcT4/ogFwY0vDoybt97GXiwsz75HXWBV99R7Vgf64TEdi/bt00Frhw
SiPDOKpvtQywdywHOACHvrvigKfCp5bgVrtFNn+4Q2B2UFj7SSLT9NtwUMLCi+kT
jZnNsz/t6sVPL+OcqrZ0MSl6W8c/JhgM1I6RItNYf3X5fg6TWSo8gJa/vMokcW5q
ez+lHdpuLd9acGDPmYFaqSdHvToh6ZCmmLS6WQDlNV7fIf7HrA6peeDfMpExNgCj
mg0Cy6ITLjNP5s0NodmLG00wTz1tmXWBn79Z+3NfS3suwX794khFS7dm4Bjgi1bK
439rNPPNi3BzLF8hPdKQ+Tb6EKmeajtpSGAKXeezuZDwj3eeYJquTDaOsXK3LJSt
5ZBG48BlingYuGjwLlnDzIMbEqb2vv3lmfbv+EzcxWmOigXEWo/hU1+bEop/lwWm
IRFP+u/MdKNwDNxDfgOKXs82KwwBKSsUUq7AhimbebXd+F8T/yWRhuTXKvoP9yMt
YYSQ6ddGjtfuPKrMX7j8SskDSwPQ4KdwA9r4AnoDCRK0q4y4E00pPcROCBylUHC6
6CDhgy6Q27e4VvljbRqgVmZQgVnMxIf0btPQVAAqgmA85qWtKtmGpUQoeKFFVWAN
Ag9XhvP/F4NXdqYWpOjqn0DwxAz9Plb7FUnXu9/VT+5EwmPD1xdXzNQ5C3/6I+I/
arydIPzC8y9p04LYj6SM531uzjCoVSr8Ni8iSzmJm6hxxzfJ1ZgUedQ6FvL9/1MP
OZetB1W9p1cKfgEzP8mX0TJ2V5uv3Pd6inBL/ZKN5V8ENtJhCbTAjgsu/qtBprYe
GiPznQhHrjMvNlqcTX2ErY7pb2LKuYzLLtBDDQfSci+5CU4eYpMTMyX0gJ4D2ust
ZxBmS71yEQosxS1FAJcR3x9lFLCqD1xv1boMEgGV8aHy8CDuxJ/cw7lCCwjLZJzG
J3RdfuXXNGByTWA0H5640bRivwPiTS3uZTtNv8whtWOpZij6y+v1GI7m1s4Bd/Fk
I8N746HvJQep8Z28y/T3sMMaKIrCBzfGyZwQNWBEc+3DVgdsSVNprXuWwj1sViAc
2KD7JP2RaJT6E80rFe7OL8gmb4UP0CTzpu5ctLIE2Rc58nyDBAaVtcy+hg81gB7O
NuL/E+AAgdo5C0bA6WD8HdBoL5WchcUCK3o6yhOAI2U2/0Yws1mFIxqD5euffpJF
Lrvq6g74XUzOx5tOB9yI+Fqpc7bXMFoUIig9jshpgmevP2jF5ccKzJJVm7xtiRMh
Gn6MI6vodm/BoGHQ00KnP9rcPae4/PqtzPTQpMg4MRB7jinL/OpauvKrH3Ii30Gd
DAd2NKTAbtXhbf/UxuvTSgr3zJERgEubmrNDyLuT0cXIxCfB/SqSf//ImgES5aln
aZI1/pBXa5vmMXZD91HsOlaQg10+zBkdmhB+9WjoDYuIM/B+z3Jtqqh9wfLhZcVj
oALc6VHDB+HQIQxFsyojMxMuSG1bAex/+mZGQ/74KuAl5LFASaYAxnbS6D2bJM3b
0IiWOyZCkuEJzYkyzGqR5QotR8wylGgkBo8I526+QcKYgmUCaRXl7D3CfhqheuDI
4HdX25v87trCHOnro2X6yya6v15Y1H4oHEKeoqb/H13QMwfl6E0nw8XJcANQ3Fa+
LlrLedL8yJAYrCDHvtnMmKCSRgj0GNijBOMXg4y+bKceBwrq+g3NV88THvmVClJs
g3Ncm9ymX00+8nk1uPAft1ybQ1/KzNOhtxOOPkXsfhPe+5d0F1T+jF7qA3si2Z65
9l1MwPuIu7M9K61YmY6wbQhOV4vJV+Zo6iBPRz2IM00n3tyNbeu8AQx02praFgEn
xP2Z1YPkDyt791hF1tkDdQ0Q5HcePmufNBn3uBzxyZ+FKSykPwUihQUS93ObJktJ
rfKqfNZQOOwlWiOE3rZvR88xzfaza/bZQce3iCPiJHr30b3+3xjq0h+Rv8gC07Ix
eS0fNTapBggHAbRF2NlwC0sFj0yAYrD2ggZDNlBLBTZ1g3i+9xitnQ9PJMf1eii1
IJ8A1mdIlP+MjChLcyyeCGVMx24k4B5PPxRd7nOT7/6jxPUARih44E6LThJlrXuX
RX37PLgu6Z8tUK6bepWTqXMbcWaSayTZkbGekDkFwoLGLEvMAyKeLWWsUlo6MlZ2
tv1UKGQtVaEl8ez+ldziIov+/4Vodc0jo6KLzzHhtLp5YdW2BIjNPnbjm97Bk5hY
R/suR6TZ3UQABnIPRbyPZ1l1Ffbl3MED26593hFkqjPdOmsY86U1kw/BmAAt38tE
9MinqlCxdkUkF34M1ty5WixdPJG8FEbm3PwO7OenpO0qq9vheNs0Ktfl7tI+af+a
5OM8k9lwOSOHYS2PnxMpRSmHZZSH3tf57ux6gSt6eCVMfi58UFRrNu0vF0MEEvKe
Tdwc6GGH6wpmY1HuWhNaS/T1p5Knqkag1GhrydehCg9JIjikhkaRAowylCa/7QSr
YAislQnqa+e1TUMrtURKMw5LKcV31r/ITcyPt95hJv4Y3qijvW3xXuguMaaPmESp
T7DRBS4hZCeByTuROPEjpTLTzeZOT1dLIemkpcCg6XjCjcvfGA/MVtEwdkFtTx/O
rCOGhTN9pZXaegKjZS6m2UdabHNPbKTUVossIOkofXrnOm+HEYZ1dAMqX3gHMSxv
SSwvd2OmZkZD//v/2pULBPRyPpLyktpsWaxa2OfkNlnwC6XipEYtwBZuTyqAkUvI
8VYCg6cZ3Cw+IQ7JsPpB80XJe06KzCjverm5du3NXwM0EDnYwyDHvufCaHQs+KDn
DdZKXQYMqiQBIhGc5ErDW3xnSOJvERioBp44VdW7t7nyvOqLn0aPRP/LIKIfK3Y1
3MpImPBgrGCwQ4g71mnR+O1cVs7fkAnXO4nx549vu0xlpIBcvTfUP7UU8vipX5Jx
+ShA1Ait3QKnTBF7Fnz0vIcMOALoMVYoe6xs/LMxQbmDeQN0Yd05M33OF1oZrTNf
1dpBXTuhbricKOW4h0y4lEazzcK4H8oE8yH1YKJj8BtUyZKF+RLsbq6Y7WFMDDwo
t+hDvrsGFM7QCYp0wIGOx9LzjJnil3CbnM+lZX8QPnQxJr6TojMK8UVz4sdfXjJe
sFKytQ1usML2bfegAnMnYueCXTXc4pG5Zgzsujh2dW/czvNWQAypeMBFg72Wx02c
G15FXy6E1uJIkBLx+rZ+4EGc1ujnJe4QIjw5ArwuDzmWZbhL3GsFbCe5VkREmEyo
tyixxunPtEcrvqV0y+Bmi14mm7grxx7BQBBRb2riiQXY0pkiR29FMnOfFnJ6tm9D
lyYGTrCg9SVZHF9g/0Jk6Jc8m31L8jD1qVlZ/WsJMDiD0C7erqVYw+/0xN5VgnBR
kC9CVVEdmgRHR8ui61p+GbGocghMp2j/ONwtETZvfPMbj8fYou7MKk+sq0MgRpkr
wcUfPwHLqEwXO56D2zLqQILTX073JNfYzRNNLN/Fl8vNYB78RmmGB4CxRJo9Ev9M
62nG9+MiHMLNkj7W2FP6fON2XIGyRZqZKV9jWavset2dXYRFwdSOPkq4tCPA98lV
RWBnGMXx0pnPydb45OcPMeLn/r5V0PobRGZi2b6fHxKyg0ay6w+GxLd9ZQRlt+T5
uXzznQNHUE8Yu8KjbK+t3WIloFIQ0BuM4IFnKnLQhVrwrWjR4gkA4UZIIjaFKmJj
WQqW16x4IMImpBJ6HdR6DCFfAZ9ueGMhlJf0NqAD7yobBUpQPhYz7SOR9t7jf2MZ
BATBFk9eudV20LU4cmT7dvyQ1kDPW+q+iGBc/PWHvJg24gril7E7LoA6ZxK/A6SW
QdIYD/u/z3Yg4LTQs0C99qy+nDFpRj3YdPlMmso1ByXOUTtRf09zCIZ5WATG6oLM
YnPwc6BfvZa9eFwbuQ1TRdGwWAXlF+FWqxUrKUyVhln9dtVXIlPKN6p384NeEhZF
yD1CwwQf5Z3clxGshCF6flAIJT6rQZ2I3FDF78P3qc1qSOOHsNHhhD4xCL8x7bOJ
T0sOpcOH0J1zGi1mSueBdQ8Bf+QAyZZq9eED5UlpK6sdJ45uNjKeIStEqtYCOuxr
+8CRJ/PiwI7I0Dt5VL/sqYtCg1Bh73gPQCcMfcuKwji4izmZZUzzFH2FqL75HUmW
irZ2j8aZ8l6FkXLDXEzsApL+EyPfKXvN1rjfwfAH7NgQAOo5h75qO9gTmR8rZqoH
kRPkO25gHYzCRmALZBhsMkYQTCuAoWf7PeAvu71cibZvpS7TSbkL4JLcuu7tOqyp
peTe5eh6TVRlLLviaL33KcnutofXPJiAHXr9ioUfH41QGVFgsb4IpyyQLpsx3NEv
yhKast1o1+Mdlb/UYxPtZ+m9KdgIHIFd+S1AaWhc8zWz2OwDZIVUAz/RHA+H/xPt
xghBTkDH3KnAEaGfblAZHygKH34UJGQmGmbjY//QeRN9bsglS3UY5IaTebFmLzYj
ekaE6ekCpvPDCOZHDrsmIPwrkRREA2uSodSScxnq729Eh3ixH28vtl8jJjL3f7aG
f2DLCtyyBagxkk1d+s6uxIOjU0vKmAPb4hQsc+XCZjnjcndJvHd5mIKWEAMS1NyS
9rakYkbBBvXqQYVJwgGM9yOAZyana70RvWPRQiJQFOepCZn7XZ5Bkl7UyFv1zZec
MZm2PfL36a2IGrgl6q0dONvDa7SJgv8a3yGbrUYMblDTjDzvl7HOOvj2HWTwXETG
ymILc5j6XvTZnlt0L7hsCONo9saEZi0kXpXtIJFq5ymgkcAxHtnMwAxIscEbsjYT
aIRzsPtvo5LeyTghepf4yy75FvQcBfiDudbXaVauHA5rekskdDqQLldZ9eemmO1s
2PIjJPKecO4cK+7XUGj/C+ZwJMOh1nuapn7Yyc0fjP7vvAilaRxWeDlIA53OS+0s
e5DqmtwRnVxUXMhfbMV9rTzltsjKBJ0ZIpkZfCXOm5+6whoSETpesc9jKW4wJknx
GZNB2YrQai0vR1jOVVoCGqdBTZERCrX7nEPoJlX6Y2+WKjvJfUoIobObX9oE317U
ugMO/q8RVSt4jHu1IkOMTNPZulfBPf0ePIi+FoL0L1GVHytsZxH3e9nm64Qp1BMD
GV7DMZam2zGf59UlxH9gkoXre4m0jf+NA03mtpyF6Eyi5646xJcdT3hpLGlJGbIc
Vk8FUnCHf2L+W1K/s3fVs/QBS3n8Sp3u20TXYgwPFLvJ7hOVcqQRzzZyHNlVvrnr
ZyGjUzZgvybB/pQhi47+DkwPVlWXrUWEWexNVmSPt23yvi4n/JTVStK1VF39gsHs
MUeAbjMnnV8OVRyXUXChc1yV/M20Zt4keE1+dL9nzYtqNbpbJlPe01HGaL8YTNRJ
JLZF2YQg48qJIPvpMvhFq7bzWzgRolm1+wUnlxNdyOUNpXE2Fhm+QZIfE10Ria3v
LcXhCY2fB6BrdDtqBiSwe1DXRf9jmy2JLd9HqFoKKkq/XXi+2qcNr9X1QH+I+rPK
UkfQBBD6GxSW4KExLCYm0rW6e8DwX1MzF8LzWsCJHbTHdH/tFyXQPdK4moYLrkJl
FuscdkZao4WPsAcaEjAqmnV1AgX71uD1T20VYTLJFNpO5sUTTkeMRIzcthJpdzUR
8Hx9gzsrCXL8Uzte5W7R+nALdRnB0bbas58t0pL6p8Oh2asP8QUIUvxTdnPDTNqk
NUPtTMvCyZ7+NHfnxbKCMjeWnvcPBPUoUNTrE+9KV5EALOhwYQrHS/Tkd64AYC1a
3mcv2ZntaUXJ8eML54r2sY0V9pknLF5ahjGOt2cIDOj3NelhjFNAyAKH5tsi5Hhm
1rGDtEK9UStKgLkAzhMhM7t5dXNjijnt66iYejDuD7NkAGFp9EMrXPK25ogQrqxR
dTVsQG85WyWyKkXx6eXQyEwa4+f/BWjFhvF2nUvYKjsP1JaPVtl6l0oL2Pzicjrj
dc7McaG3RYzX6VVhSAzez1ahoJD29eylfCnfgD9x2jfkDUKVM90roGI5OkT6tq7J
fMu/tIws7a16qKH+ZjSik/s0ya3bgkBuuckogygkIR6oshPnikHdDqUnrvi/ymR+
hwGpDt1rzzFk54NVCLMnc3UlKx+PHel6iClZVcKh+DXYQc3jeOh/y/eY7wLkcP0O
TcOWi6dm4JA/rpyRjqU1QRjJUZgdV9vRf7SHlRipHovatozLS0+CZvJtqZh8vpwR
BFrXpsMMliH5IJkn/MKvKeKktu8R57nMzqxiGpMmQgoelVvWpKKFqBYT/DnqKQye
4NLTVsKpG9dfftSTluIE3w9iQeJPiRZI4pSVaAtScoS9+ONuKl96NDiu/840B1HV
A8MsPpzBlbNKn5uWIJhlKComGFgrq4SSh8mqw9GaPOVT4fLXGGDzjlAs+VuGglOB
ad4eh0ehgHFnOtxA8Q/sE6vkznbhiWpeDxu3HHjma+L+4OQg6PTkCNZS+whxSQt3
olcjE8VRYQzu1T2jNx1rFfNXp8uHSIZU+rXB35+2+p+w96RBtOsSgGguB+h/FeEj
UD0MCR64DaatdTW6O06Kova/yvhLhIO7WZNT2EI0xo8EdWD9+8lshkaVNQy9JJm0
PhdTY9KpPiiVBBJ07lFuIQMWlXemkOCiqx7SRnEpZup8ciTy5VZh7w07cpvBTXAL
Gg/fXBHYXWEPVSQMu2dMTs3RVUSBXIQXf4tTRdq7+Juv77J65kiCWrsI83Bu8r5Z
WauRYvFHCDwjHV0wGKNZdv4+bh+My1ZObxu1RRupiyOJAJf6u36Mk+z91qWF1B5V
lvJFARWiyDgSTz9CjC5rZPIWme8v+dsJO7NARlGT2t3lQjkd8oelIYmc3DZtQ7N3
FjWHk0GQB/ttlaqE1w/QxiI8s1lv75ulQEBM38gw9pYIAIqXXGLDCkNv7oQuSZUc
Fhh4iEYnSEtUtEQZhNNJ3x3Bch4uM/RYeEE+ZtREfeDOdIwKy/dYVER6v62sX4vw
nMK+aZOH91oL4tGicY8X6XkMIT/AD6ZE31TOPWBGM3W2OA5lgtoUruV+KeNJY/6O
S3Wg7jlSnVMp+HRy+o6q65vZoDpBpEcz30ImwGAyvGwK3lvcuodLeMWBghV5hd2q
80yuZBnOj6eD/pvhBBgDeFAnKGQDAI8v+5UOryIsfS9ldOV892h65RO7IJDF5er1
IHu365zUrGbObH4Ju9oc84nUzyWI7krSum7sXgX/td73l3WpkxBuFCUZQaRjOiTH
QW0wfXkwEAcUM8u8/9efP6alIE884ZbmoYcgGt/nb4okTK0o3h+nBHs+/x29C5lj
3LFDZVlLsEuWprx4OHlqmtSNXjrezHR9/GOWeJRzARYYFGiRVLsMytDiVVA3fQ7D
dyZdXeS/lr+buVuQMiDqog8Cm+VBewumYkPMvafL2TaKhzX1ZBSllfqmJbttshTc
fQAYznA318CkhU5QVmS8mgY+3GiOfC8grPu8SLIjED9W6d10XPA5m+FpXmAjAlOL
5/iuL3W8+kMDSetdENgTlRabQZJdKRWKscKCw14WVTudvfZ7oZ+Bt+iE1yssRoJ+
xe/peT+rcQ7lNAH9gkWql7V5ObaNtF9YWP5+YTfLLLz8DSvET5Q57spZy2cqVuov
/ZLwsQtj/i2TNG7TEVQQz2nJ/aJ3kcb4ZUdZYlQMsqZa2VoJdbIp97wmQZbh69B7
488NVAOaQnZsEZH1OHNBPVwiq3NfUn+XxD1AstpDfUu6PpcqNY76rkDAZZxs+ot2
dtPwQBGa8y7T63taup6erjIQPq0KMDPfozISZIkN7UA2/oHt+O0P32dAnhXhtQiW
DKtEWCIs52+WvdDpLwU3RaHKXwEbZhwAL7NAdhymHvkP1Pg4G4nivvo0VKZOc1hw
UfciG49QGN/j9HrtqH57m1kCpsrcivdeSdgxgu2vLZ+5lHazAJtuj3+TKg8Pc5nr
GfC3tGMo8toj/gnUt40i+rGqXbnFrLBa3OhHDGeB6k4UxepWkHydDE30EP15ECGL
G33/Cn4+vc06VY0Jbw+BCOOs/eksSayquuLGTeOkQwpv3Lv/Z0GO01WUciNlwW+y
KEvE8j7HdgyvMSJ8ZGBU3+UWND634haY/h9seGXOu+z/16qRf16mGO3OeqARHW7F
aAGDYFsjpxS4tExdMJ+B65r9LUiSLuLnOZFY5NHNpONMIDIqvR19BYrh4LVr7LSJ
rgLDimvoKY/M7g0SA2rRjnbv1CvKq+AmvwWKHfmqSS2DPzdiWmsXTau4t2M1fxAL
e636a6oVj0H/cXSmV3G+0lL6l4xwFJwIeePHXS+p0WuPgF7KIpowh4UzgT7Kd/hV
AirtPXdhDrhD73Cnn2fYKuYqGboG9zUcft/C3CORSrJBfqIao5kN7dKiP6Jo3dH5
J82TOdi5b71esCKI69BmZHUvgqLU+n2SpW0rTGbb+LtR4wSqRhOvWStm0RNumF74
SHvcO13+j0IBFom7jm2yIn/MBriY4lXkv7z72wxrG/yqlph4s1VqBxewG+Zi6QVO
OT0ssZfxRYUB3QpV+0jFvM1DMnMAgNpaB/Q751gaV7Df85wrMpGhWsuAHk0xGPLJ
ZZiP0hFQw8VyzGfSiWy3hPW3GZ/cZDqJxJuiuhGhIVfJpnS5BnzJj7Z7FDuz9rNF
3ojbrSHBajjCtJ2A1eAEq3K2gNB7WTY3FyW9/J07du7Owq88kO2JwlKKh6IvlLog
rcBk+ZbgfheJwEDtDGqkZwFn/CLcVl6UwVUxavm5r9uBz838AaxynQ6+Pc8qYNZH
7oFgRwnRjoG0uqMrPQPG4HdMOg8FCBbsz6zr5KXnppub3H96/4pOnLw6Gp/dPsiF
FCd09nhPhmWZ+CLCo6dtsHbxyqHHasqg7mE/9U+2/I47pVWu2jKeCbtskOF0rXU8
OwmU47QNwXnnAVGMVm4shBM7BvkBG0KXVXIr0n1S9RjT1fgdBk56sQe1lymrFEao
fopOoTtnZYET5RjbgyJgkYFwi9ktMQdFBxgOg+yMAGsBvLi54u6BFRWgXcQivanY
YVHhEg+Bi2HJxU7/E7a9mBk74kyY5YnsJZnpZTA2yAPJpjUrYR16VAorGrkHFunH
Ojb9l97S4uEoBgGlN9tbVZpK6Gb2qYMUhZ0x1xmJCxMlaSKtCVLDS+VqwnQLhOsM
nRfbg/xYhwd4XxCGeB0NBIV766nKNppD2ThXArtY7VJd99czp1FHop8V4mlplFJQ
i8jHlddTknQrBKNhEIZgIxvN9plEpDa3sg1eWC+Urslwj7yQM8StS7gPedume6x8
cKdvU93sCnUNWKeHXIDirbL8B+7UQclpAXsIcGunB/0GzFwdTi2ZZi+DYt3ECwbb
p0OBMMJM5Mvl15OyNMt/YT3tZRwJp1+RdUWYhWKus1qfqyslTG94uOegZrKxOmYy
EaV11CUdjLfWIqOX2kXddMszczzOVt/ia7v+0zwxBsD1iJfydk1Fjr6lqSVUgp0D
n/iIuBu//aBMZPDOkruZuwUpqbUGnkrUs8KpgDVDnmgygIqjwMEe7nGks1Ch9pIB
ABEgjyIchIrBEO6Odgwj5P1lsnpa347NapMNN5yuvMjdJ+tc9sIxFI+brN9EqrjL
uK9a/+IfI84oCuM1DWHT6rOBv8dmjKcZbDerSC8pn2vJZcXko45ZeanJD+H4DwaR
Ndn5bZUVFtegnYhpiEQSwTt2BMJZ7ukQfcr2N1pQF7vhftm25TR1M1Lzmy43hE94
l43UUexBF6FrIPYHDyQpYy9JD1YT+rvZoT4MYscq+GYJfIVfqHnp4lebYwt0M+mh
UMhLl7wl/Bn8AUN5tgJquhkbrE0m6bw95C/ek1V1szyfrzYd/oCM4+hkgYNoZXy7
4WA4PHd0AFD8Wg8KY1nVJlp8JZA2O14USmCdlAny0M4GVgt+CJPMYt5DmP5cbb0E
sVZpxsSm3Z3J/rlji9PBqSOmHVtU1lBGfiU4B9IbZtdKX6PD9zun1ApsTE6U/QXn
B5AY7vTkOA3DKaTXnIpVV4k+AWHygZmOtGT7ir/JpHcMwkZxWtrWSO0q9SSYK8me
MIO9T4qnwoTl0/tzOf7s9VVT4yCeP0sDnMhFHJHS1mbmUStGEUigRR58ARnQxPPy
aUd0z8/6TJC7vY8W+FVyMIsGXzSK/A3j5Jec6xTfV32ae4OqdxiRr/kWRXvS+wyq
9LHGKkSJb+taOJa471tLKjdOqLw/M0rovHQcJZtbsWow82wpOW0XyuX9zHwybqXU
LXqO086oHGbg2GPfzDXKoXnkZojZ0fEfZKABwcZ6L/2nqPPqmLGRLw8m5Q3RhGtI
Q41OlgLC7kJuqVNCrN34Y/0+OXOTYm0frexJFQ8G3Nx6iAqeNFrx7Lwughrr41vi
6FrmM37Ym3XspiRGlpYjQH38udKrXGvGdWRuFtWPas8EZ84UB/u3ajkXWyXJHSBs
U8daWzkRzN+qxobOWR/Vqx9nMloHOZ9l0PtnuOVG7K9OJRyrDuR5XfK6W3Ykj3gC
I26ONVi7oYTt+gnvA2XhVnwcuGcQNhoHsACxH6flCmvlS2jIJ83NDQAgTYR9dYI9
ytBYcv+R0lc+6KAxDJAQ+OZF1LMvo6ouVu3VrbvDnQEjVDd+Lr0Hv7ELxfkOYQzU
Xhj8jwEAqvOhZfMRBLMZTihkYgWvITNqZiJapFUIP7kAl+slHCzkZsxmPbmSYwGk
t1tGj1sLBzdJB6RGP9LtUikgHfn/T3SxLLU8GRwX29/CPkus/oMIQ/WafekgqZl9
R9g5+tO3Okxmy0jOtDmOfZTu3H7KdtNkE85XEPv8/OpzGA7EgIfU+QC9xCX9Jb1V
r9qo6FxqSegF2T8wk2Jz0jaCTpMbjXbFF+hDI47ZM8P4VpI4FBZV85MJ7Qns+0+8
RqR+tvr7XP8iaopdboPUHA/lsNRqY78CQ445W8/+Xc8hNoYwpzpkITe0n7OWxglz
b5HB27vRxuqd49tRv2RMiTkYXnbd7CYeHprpI8r4FWTiSbLaRm2FeJR1LAII01Q8
R6GpipOK8wnlfYMEnElVSNxgsbxMPeWHNLbkaBKDZOqZu8fznSwfUJtLjahElwOV
+bL+qBYCobVKGyB8pTOUtLexopj5w/nDs3jOcPXbifhtLezqV+gFMC2k2pAbTJBX
F2WznfX9ThAhpERr0y4waEx0v14KeLru3hgYLInXjZV5eTsuxqMFS8EgGD7OsJ44
glm3vqvYF4qyzp8D0/i45qeO23QQ2L5o08IWwwzOQaKYmd6Tg3wp9uhSLHVK/7hN
/HRZlxZmt++uugaP0W8yGLP4q/NjOKHal6X4sb00czXnagLQdUfnL1Wyb1xWTnFo
s1lx1ebs7OYEskmB5HWhgtKKWpGoTHExv3x33zLbKGYlu5e6s95v6lGjEGOFOwdb
2cJ10b5ZFfMl0L0c4xUZJYXJC07N3Z8MypbYo1fpoJiLyR5DlK0oIPSocPdQh5LM
7yL78LvXO0oRoklE9LyuDJYna+3O3rKld5qoPo1SrKDKnktXfdi50QET4zaRSMNl
M4O6liG970dlrPVh45cDY4JSTnp0V44fJgokP3H50PAbMZRfai/jL/gDgfPu8Ot4
G4NSi6dscxYsT/lxJ2UECX9+h/LNzoKlVFylRbUln0+l5BVFZsl554uDdFUA1Abf
Iq9a+9U3Cpnd3Sw5266bSQ5TwK5sPXhahQzPOucxi7w60/dgsuRzwOJDtJAnTqW5
WRXIXJe0XlA/IYMD2/AiLZEh31tg8xSeW7+P+Bb0OJ4YIw5K2Br+QDK1hUq0mHsC
J7FNeYd1HPq571AtrAOjHeRKMFLonRy/oI02DVVkIdC6MhH2Baoyoovz8fa6CQ8b
d/vFkgVmt/roZJFEtb4xeLmVRAK4wU3YqewKo2o0IgZaDODUuAe5wkN6AEuA72vt
fifYC1ECz/1lMPU/+TsLi9SCl7xw5QFap+VqdDzJZ+5rE3OkWwjlia0ufsrCBH84
+YKF8eiZTjx69uOwVqswJBT5nBUi4D0DbgIOMIlnT7eImMJedMURcx+mkr62yPzo
+xI54LWk4tcyOFkKtNs9CT9/WR6atfPk1ydxIf+EM55G60LHBz7Ok8foANHr/nrw
LBdqm9qc575RKY+Om2MGGIPNFYNQO6FgVCR7bG+n2dVgyaTMunF7uqg5dz7myT7I
wQwtmkMLGbFlcASQ0lPThitNfGx60xgNyNMWFyGVPo103wjpA8B21qXTISukgq6n
ziCtB5vmq4cZEpIKW/oezge8ErzKSeyM17IhU11/kZSuyWbsW7E1ItR7Y/m9RYwr
tbMe/rHXCDF/Q1BWbDQAw2jMldQNdLtDg540VxJOVNk96/hNSOgh/R4R8FpVhQZJ
CrS90FZlb1YCG0gcXiwiE8CJRXLWz+9vp+HDib+OEduCQ2osl3cXESAhHVs2I/Rs
IrUCt0dImPDVd7qz0e/QAvZxPRVhTRedDxq72T2MEUoKpcdPnkzsN6Tn1O/VkrD4
OZ5bFIaiuhBQDWugmsaNGJzfbE8EP35G7BKmfqCXyuYeeCGey0/U8bCJKcWE77Er
l0Cpg5NIB1WAW5E2UYYlBE3mfc8BIVFOToO0oK7KSfRIquvY4chzZQzOHTnrNSTv
/haAK6Ru9AGQLj1jDL/v5db4PdnQ4IVIvTMto2TQFgRxhvykvHoubWKqGceFuUa5
HWUJ/d+a3WRmaTjxPlD3MmzOmqfanZWiivabBECZEP79+B7A6VLH1nL12Y810OGV
OSiw9PxYV/6gE+MDJRfMeHqz/IMClJD89Hj5igCR6sLtTo3ncBZPJMJcRNEAzyva
YlFj52xYaAD+KmpQeKtxvXkrPgo2jOiDb/EpzS+SPwvXHj5lFRURXinYyQva1rZj
D15bz+fz1aTaiTvMK8M0AFAF2dpbX6IpyveMDz7YdhwSRz3GXWVl7p34fH95VIpz
6+VsZ1HQYeUXZ21DvnHPvEyLJBbRsJ3a4oRarUxW2enGrSbzdaE+rH0zorJCzY3t
aDZsS5joAC6LPvVkCj0OuFukb7+oLMfGk8dE2LDSVO1d+hi8Iat7AZvaSzQcMIAu
Eso0Fmbm1lSpt3BBUySeJdUBAavTyxYOfIHN5j9tJi+1ZseIN4LwvvMsUx5fk0eO
4nitsbUtyJK2/k4Iounxn1yIPedS4TeB1KXiiwFIR8UCMMu/9DFsDraeDcB6vLAS
CopVndTRdgtw4W0lQFEu169f0YQCb9qHWhm+aiWla5sDO2mXeT/vwkcU0XNH5FXL
osC5FnxBuhTd5AEeeYL7GYKvGpKIGP2uKAiZWm5WUDToYH/c67lE3UKMQVAbnouE
6RRXUUrNE0yUBWbYvwFtdw4U/hVMSaw171P7HdYnwti6FLlel6GWhRhDiE1bJSZb
x+Xgpe4Z4lM1AmXdX3MrUV1EdqHAlLIfIiH2vU59TEyZ0KfhlavulKRMsDQTk83a
FRIzVCbIo5Y/7mGtRCXUuto6QdWKOEJgmRDJEpwQL8RXFzLeVp4lf8LKrf7BnSZ0
LW+Q1qFqSRcjroI8f610Kmt7hg8x1+AUaNtYMLPuElqFowo6KFDgQZvpH9dldqbe
vJMuN7arsNoooCtoJCZ6zEY7eHsPEjWqul50jnlEW1iN1LKCJ+12jOzAzI4vuMTt
+BO7fURpwe9wElpUvb5GP5fpLVBIj5yj4JBm6OXGavlfJv+8lyZWB/gfaI0bcDa1
irc149FoHHv9KqQ7VNQ3bGkoEHihwAytijA4l2d1hCK5ZTF4+INjs/gJ611Uqhqk
GM3XvpsCNp5owbCNhJXRvhgnKBfvFe3DaUFFlvO5pmM9D7ILZw6JbKmrAxV8GChs
WLMs06Po0X+0xQqpi4KzC3gsyUDzRvL6yH8Frc+ttua5YqBgamnoMEBJqXGqnCUW
cxBJZxpi7+q+KL9ehN8/8txCsa8XQGI9uFI3KpBS3sSoMycf11xMotTXEpnqi5DZ
b0NymEJgYXUw3+kZFGEZZ1rIrRUWtABmrgPrYnklMwafejJM0FgZt+Vp2fewAbPA
AceznRFdxjBfjdIR42BIlSQfYgB2Xwj7qE6xoCvn0pClHrUAcGhtC0XCFxvTy6Ot
0ATp1SNv8RdNcDCwanrJeY/FjKKW9EMLcPx+BOSOp0nj8mmaufPMGqPg4YJ3ISFz
ebwdKt1JhOD0QHDWiOcBYOLQEhwIKWm7RB2oZukrRWjaX4PwJLsQgbQsg6UAdj1I
kPiMubH43psaRkJNrWfTYnaiGWRuOD0xGuApP9wJ8tEcYw6VRTSL7SVZQCkhTJas
TZbSM2Kq55DI7yUR2E6hOcrpftdYyM2MqxGEpnQu7eJcKJxdvFhRxE2FXGfxMI81
LHFeUzYi+FLBa56VnrEYShxjG7/x05VYVpZacmastVPOwR8XUxycDUSo0M5aWYNb
dkGRdasQuTJFsrXI1SgJjfgAJImCBCSzmVhTGyRpMBvxy94x8zZMNZYEk3xraqe3
mmsumdLgCxNORmIYV+w+dtmEqpv57q/9sKbk0K5GEGlYcIdM2ze38jvcj31A7l4w
xAtVNn250mfTfS0zUG+b5mZ5ft6HYg/1mgSNRRbz7nEC08+8AaPRGQv1uknRulPo
9CIkpMWmhij8ziHzN0aTcG7z9F/uUK8OctIwXDIXydLt3W8SVpLXFGnIHh0mvOTG
i8MM9PbOcbuKt7y10zfiQGpMtDkkifAuylrjqvMjTenr8YD562MQy/RFLgcdyLEL
hmV2qDzpKwbgj84EMQ+nK37DwRlMP/onWjI2R/2EOAIgzBZXfmL2UVfz8r4HCFfL
0s2kKjkY0942rkwJ/XnFCNs3cv4M0yeoIxg2yDYJbi+SR+Sgk5b+bJtB8YcfA1GM
MW2R0n9qmuywWpiq7daX01Q0lvMxyB4wGYTwFy8PKvqw5ZiDL3AoSdOqU2e1vqCg
baFyomubpHoKaYjL3TUH2uHnQkIDvTVo3IWhaskMmmVFcQ1w8gIkgWS/YltCDVso
9CwEQbqMMnmE+wkqD4PCboBH27taQigyU9BpAPS6BbH5QjsJSkYFkhOWpvxlWXiw
T+7/bENCaTxyVwfYUY3kbTx3RiUL2sWNEKXwKYQEgVzujJom1fCfJ34ocL/4NGcT
LXDPXQII2eMK8hI/+V2rsPswOUaaDXZhtkkZ7j1PFwp+CASvJB73JmB3YkZKvpVr
bFDqpgPGKmqAbZubJTdMKaPTbMNVVhFatuNDtd7K1XyY96bs2neo33B5MVc2jgWu
MGY//tEvrKjDbPodt3rWf8xnrP6klY5SNrfkAHo4PB2LnH4idBADLbLHnksWj0e/
WSsdpSoWFGK/CGz8WGvcjIbho7NJQqXiS/xT++Prsldf76dtJKocjfmJjoFE9tc0
/ducImL8M6muIUD9tEtjKVDHa/wW+FU7Ct1cu6i2iJOlncAK0mMZk6BEcFRMomCP
ENjmzfZ+6EyUCtZ5WRr0zdoaY5XeZ45YpH6vWPqTXKOOjijTCG/7CHAQpvpSwwct
YTy4+aIyBvLaJiZvKCfDzGyPBAHw9W6a6vCgKKhj68+gLHbhhgpSAVdEdAXdywHz
Ny7d79+OADURscMCDmVQ8r7uJy8uLbrp1qq/Q6qIfq/LUlDhgDMe0Ka6i6FxzdaW
sh9CZ7SS0ZOAJvjgW5GcBJf8XG0ZEH+j2G48WDeAyKi56PDssnoai7/uo9LRQnLX
lV8fgVGUl+Ivnq71lErrmLeRvSJ+nJNI4oGJ7Z4pI7J/orsIIWYKB/dlpv0IgUsQ
bWseYZ1BdkAGKxnPujvoyCuFfY9HfWt+CGv+hUkLBQFNdHiM1tRxAa6QCnBml48l
qCmA9DgymHNkgu6LNJS+GZLq+ZQLN0biVqRf+7WVfztJxyDq38Xfva7bb7BlTcdJ
TzCkfOmDUnqmJfoZ1D/n6ZShSrpZO4eEVPnVMc5CjtRlCc67SuO0HmpAKEhcNp/d
JIz/7oKTXlroYsz2lIOW/vzc0e+iLidji7kFJ5zRB8VXm2p7PedDqvi9JKP068oA
0nmQY1SqR2wdy0k3/SsJangXdEiorvdpuBGdlXsoxX7kc//AjkKse6aPEw1ra8i+
CHuG0wSQNEq7M+tE3uXoHBsKdHpP78lfg9C+rm5VWwDKpBYUWjI7fj6RZvB1ZBYi
OGsAx/gvaKp5QSl5LUm81HHQjqdPd4S3FQnpM7D1JTRddoQFBe0L+YgFuXBSdVeL
rNrHB1pjxumwIYScFGEShYgO+RNqG1/MLQUFuuxXW+BfO+tHKR3xVTtp+ZYGRv0H
RQk8Q8wQy0d3PvGCv9Xv4VxQp/lc5atbfvFs9Xw9vX0hjXT7iFzDzamDq8xUkRP/
0b3UzusDcL0fQ/k0PQJJRiZFNIRh0YEZrqFmfsDY/0NLueoQArfY5E3IMHjF2ubh
qtstG/kR0hw9GimuMKH344rza++MCAfCCR07k0Ss+OR/7t92HvOjT9AXo1SqL0Lm
0mLwDQ3lP+7BVz6W6B5uNLn9EQxpD9mC254+8N8ho/6UD+oXJ7gfD6fJJZNqGLf2
b4HA8SgxLTcmQSTE+IjPX+qvFgoYWZHOI9NOoQVQNKaYNH7V643XiihH3nbaTKXz
BLKD8Je6WBCZCQDBZxZZuFQC39JkDgxWPnvalmPUQvI1V8ZlEMyhILUNF1uNnSyK
VtzQV/KxKheG6BydK4GkaZZikIc+lV4GbitiLwevGosUhz/5voB+Bl1wqHVLvNWo
dXgI+mJ+xdoVSQ3qzQoCx+Sjz02sC90SyIFY1FtwaW/VVPYfjuYIPJpxCKOJVbkS
RvVb1dGdjdTtbEB/gcEH6MHO/lnM3+RkMXhl/9uVlcoKCxlWDhxhbjKqzP+CAZ1i
9HEVtDVMetnLGy4ybybP9I3jQhlIwSpjaUnJtZd8aFFeODpJAxNLZHD2wftz0QLH
BXPbMK9sGAklEmGvr/RDmbM3nWcyqB7Repv3P6iBs4ybsZANFV9affWDbc6kKrbi
AZdqB8JFMy4cm/V6SY6wAg7b4JTemWmBhVxa9XJUQNZbDyDEP5uMdJvv7ITDjjTi
amb4CaGY9nTaJrhcHMIjOje9NK6Nq4v3Oy8yLUnCfp//rgXHXe3nfg76vSIbBGjY
HxBTAHL3P7R7QtrVOu0WtUwjUxUTMGW625oop3nFsV4PjHQWC5IoMsij4/FP0LYL
FAXnb3EORyqsq/u72A1UVN7NnYwaWD/esDCNRnNXRwZdC8+H68k4HL2PUPgdRHhs
H3igmLKd374o4y/YQHJXUzutIcjkF70zUlMU+50w6d7R0RkOSi5X8aDo8s9rP/PJ
fepeQ2yLVriWy2NV3i1aZyFemKDYKW0YrYhw8VzGHNU5yK219blt5AGCF1BMcHos
6lHjOpyjeNInet+Ub60C8A4p/5UcmfL4dKad2YlNj7qgV64WOa87NwmiwkD53lj5
YcAUY0Oa0lI8A98gr+Rb9aMyiWFJd6+WzmrVETdrctiBd11hYYzhXKh+4mfDgOzs
QBzsfPGONsBnIaiRuRAaFCdxNeCqe7Q2HDuYD8wohoSD2NVBYvqdspLCmsXNdw0n
Oz0s1Ja/LXGIwJlSPMq2eavqFSYxWWNcUTTE23l6dRK7Tdcfb9wBTE32B0s75+u/
eUSsiA6HOpiMvYEf0v514XrpjaIp9WgJU5c5WM7znoI/PwUqaMcsLaIK0kYQhDCD
B9sbi4/hhQ4iVm3BX25FWgU1MQ7shHmNirAD6fsaF9aqrVPMXYEkTBDIVN1O83gg
tXWENgvLdyAqa4CBTNO/mHzVjeTvTOelxyh6rdQh5w+mt64T1gmA21F0ExqG2CpU
pKpChEHVfYSn0vAPTpEFEA/D3pg+WEcarGGuTe6YRoOh3ZtjawVkOEjd43IfIcBI
br9pwxd+ZFvbjj7pe96NCml1EhTmXEM3mcvgnHpxuV67qK0FGxuc+SfPH8HO6NBt
Tssc28IKvGlnDSRWQU/lcluFJhX0sXOixibMsMuq38I21g+4jb2/oFz2vM8Ycq5O
tAxPDH1tjVU5gmvYkjBFyzdVhw2OBRx8E1cpuqPaqoOOm2Oko1U8pPg93OFtv7uH
cGhQEq4Tq8Linsx4jd36oKnQ0FK2MiW3bvV0zj5KVM8HdB4dwIl2tjxvRxPobjSZ
eV07MyH39PjsB1LHfYvMQ8J5LukSCwWcNMWFQGj2edH4wfCFfhbjFQBzYBWiF8Cc
3feDtd1wYoiWLwqQ8grOw8UyJMMWm0xmijUDUbJCD8cgEpDIcTblucUwh8JypYkW
vUVU8yF1S2kh3+mhIn+Mx3i42Ou6uIOac7ws1WfTVoBY4bn+5y89CP1Ep9B+Kq1E
ylZ0mnkRof74MV4qd6kaul4exUm+AuiPqvAOWCY1dXaen3QFb5NqqgdO46jCFKBI
laRPhrSc092E2zTZKta2kyk2tX+c8iJLzQASaptWjuBEwPnVKde5V+Be2o/weG/d
cBMi5xNxyxdY7GuUs9g76DXCmsEFovKjcmoURsDCY+FJzXJ8+rLrfyFBytspPJVA
E1UL2yFpJo/GBWnhxg/9+0K6Z0vlmc+RK18Qvx+o7S2lK5RSC34o7+L6gGFdXzuS
AoZ5BUDKEfQqjJmWEflitEFyLiHonhcrgr1CnzTVZYqOV/98G21+IwQsTeS8tAqG
ky0y2+7oCzo4mdcbqqMCTqzPpuznupOJeWieTN8Gz+XDvcAb6eMjnvr0Vs1wWMe0
A6fkxsK5nXLemTOcKD8b2RcxBDyvxtAJwabc1979pIWi3bU3KePEyedlx0H3+htp
RJDRUH8wtO/5Wzv1waE923z77Cwo6R315OvTB/NUDy5srgUbuR6dz8AqTmsrLMCl
UHg+StSeYyL5f6gEUC1KKWPOm6rrGm2bA9VUt8MNaBnKZ47ApxLVV2/3UYFc0eT+
3LPW7KYsYOvLrlEo8yfIQT5JDOQKz930na0M22CpOizBUq/g6531VO52WcgxPtIy
CANvwDu1h55+p3IE8CaA7OwSGKnHfbf0wY00NHdmHzUOcyVz6x6qcWbXcUy8MaCA
8hqNv93VE1SQCBSbAL7SITg3e1gJUotRRufgrrQf2YybXIitPDJtwyRhP8IwGzCB
Cmmx/SfKZFOJ1DoVXshCwM1EJWeMEyWsGFZpAhMyoTvQqpzo+/anac8TrJxru8o7
959Ow+6cvmofTREJ5bZemWKp5sEHSN+z/PUvch09+5RDjVWb1GwpDnNEc21mZokb
YdZ43e/RxHfPfywqQmzfdZCP9BUk5O+OnoB0HKQQM5MGX1CvM12vtUxRBKmSCeDx
Xref4K7Z2n0GdsLRcZdvln/u3vz2F69mPKltjJwgJddLzWigS3hWRS3xRyNkHSuO
MwSLqaQQBO28A+1nM6vf02Cy6ywuiw8HGpPEHjT821q7pv/7vyLJ/Vh/ZxqUI+ar
RrLvDOflESIXFvt4SmpXlNGZxos03g1e4kSBZmFcEhMUY15FVQswdl0iRXsvTxji
iOhw5neUeDhoaG0lIBJEy/UnN+IcM3WV9LG6okWm1nv4gNKoj9k8R8lJSg8tomwg
L2PZJV5qtAMsYNPzgyvhzOP1hmK5VtkXtcDJzOddBMeuLZGX+/fTSJXuwiRoUPT6
oBuuDBGro2pGBxeM811lD0z09T7MCQeAb20W1B0uyBOY2UDQuvGBfkaX1Ii5x8RZ
daY6uH3158L016Borb8btuAa5vKRdakO+40Vc22n+dfKEAOqYAw5lcKropNQ/wNK
WiLRDT5l+4P1DzGjjRhkIi+jgWeMuGC7p4ua8gvTo2S01RI8dzTL5suI+1THomtU
2Gx2o+6t3o3ldmPh+fwYTeeUSIjSoK9qEeoJgBtfT4bIrhrMJYzR+gngB3wAfCzu
WXVl7kFaDKe+8tqFsraEvrux2LmMaynKBKVSv48Zd/35nzYfpFab5OdK2zwXnec3
1NqrbRHy5mrr7u9Hn8lzuSYVV/T5yKxWTx3d+Q9PnSrnvdS171P25v97r04dc0j5
OI9AJKmgz3MlgQl6bOL25+MqAcODyrYmW30L55zOCL0azfgEVl/KYR9/npRSsd9E
JpMEmxpq0eYKD7UQFg1NgysSXPB4k/AzrrGScSLCmWt8ZH65Yu8jm+KWOW0gpQmT
dsoVioq4jv0BVnes72S0jdydAtDR6UWl157eCIvJwAEdpA016wrgOSBVvGF/T6cv
aJQ79OySLIyirtxsKMcCPlI/s/SXNwtfB97Hhqu+YhEPYrY5M46bPUW3CjX/ypCP
UEcZFNB2UntGj2lniOHpZX35Rql7fahvX2Ed0BL8/w/L7wFgQfzPP35ApcVv4dlY
Aa03V0uiUhmADI80WxBByZ6C6Lw73FFUTaRL11Y7ELyslDsqw9aAYZ9V0lMPynFB
hVoHhKWtnkzMuPHj/pqQq3NnRdQ6dPjTfiIb+s/tKvIEIAgf+5ZKRI1LZHNe8Lxs
9WMgK3wv6uqM6Y6wKK2xlC8SBvYt5+jze93ntWrV47jBeuu21XlactZjU43ctj9R
4Fi4J3ZFkxHbxd2W2MBSTC1XDr1cmIBPxNyo4z09dCvzm8dBJSTNQjy2AR+nSmWH
v5RgS8+/XkiQI2sR+/OVTl+rKatxfgaBmyAQ5CF3oIjQfCmc927YBXytcaqwln1T
CjNlzCA9hJRtyvksQF1Rhtefc5GG4CK9WEcdwvnzc4Ywl/ZHy/oaGxFjpXyWd8T4
5NnZJdyETXzvRoR53XClWLNxbGnN9fIkPEzIGWFQQ2iSEBdWLFVLgjaZf5Ch8beM
8OG/a+LTL7QAGKHNGJ/d/Hzsip5ByFNy4xW76Hica5Pgi2Bc1puS6wzw9POBJ7IE
NBzZZod4Jr8qnW8BDoilC6BUruOYN1+nKMpAtpiX56zswJyAesDoYENjwbt9N5bI
PA2eeBITZmgznhC1rNUKcvSW1hr02BQPK3MXl+9xpDMhqYL0451ifyUehQhLh4Ex
cDcvA85wy3smNTwl5iK7GK2a/YAF7G9QdOVmhGX6uzFA5k4Y7Jmw3DRV+CNOZP+U
03mQXWgBLW3pbATYjPuYFdvlQsYVHbkPPUA7xIpfqlgajzpy62ue3e5/+ZIGVr80
rxYoGN77JD49evdwoxwBv2eeYYcbDIeHTqR9+k4hoW0qTBoP56JN2BeOHo1LMDVl
4CSvSjc/Fl72OuUNh81XzF7E4362qSzpRYItyZzSMTBhla4dSnq5BzSBxUsitmhv
J7tvzMlH8hI2BPajAi+oL6GI+yjEbzoMrJLqUAd8huECEhr7tZDxrSZLXpAydK01
4sWRlmwmVE702U50mtopqZi6gqIxmUM6+6pMX9M9X/YHngM7tteC5K9ZLvOMVzRh
HBIva5JQitV6svkBZRLKxYiXr41KrAfc7y5wc78oQxDiJQXTfqUaAhZvmx+UD/dQ
LtugPs35pKnauPmMBZwl1YWuqULiuj/7sNHvy4kePNhl2tZ8IFtXz8OOYgDfr/O/
E4X+ItbXVQUxUnr/G8eoF6xu5J+Rq/j3a+GCWZ4sRFe2vJ4CXqWZHKsbLW/DKVCn
xkYblFDPXS2mnKzW2LAJz5SGSnEiT9BD4IFrPiKwrE/+pqYgo7iTgoE8SoTqqm/e
vkI+l8RFFf6Dl4ZIhlChiOpA0r+y8R4ONcvkYaZG9LHFKdTUzSomwQJnS23Zn+ec
1e9+4lP05Sk6W66CQCtm8MJo5ViL/slV++y0XTfPvJIsRhGFNL7c6r5dPKzby57E
qMq6kAJCqYtWyLVoino2p9XbmE3bWf7RK+8+eqc6f2H3N8VacLAVi27dr70N7CBU
eynFAYt+HzZBt/IxfjIIjG5I4FOgfLT9aLN47h7Jgzp256e/3PqDqQKK09/Yqte6
w2xpSCz66rbWgbbYZBGLZs6i6e7JNFA3xp509nZL59qKJPjJLBWuBW8+esIai0Cm
nJrB7b+vYtbjtYuO8pwPonHe1HgUwqYLybIroyFIgKV8cATXG9xv039TONrIZHIH
iwyIkrMEW1b1D8DEZ+UTFVtCHVDrgutEXBT8t6bFeNgS+4cdJW5Go88IwEuXWj+C
fPAgLJzIjU0JpoKx5g5XpT4ji+RvknIvk7NxKYgiWxhvH8zZrAYGp91L9Xe2mW/q
NtCy4kwklUEA/79nPFVJXwq6tvzTXRhZmHPZeyq5SqEUORUcy8Al5kTIXLmov+M5
Bj3KOQ2SERezW+D6pX/11AJezJqWkpDusmhz6kjksAjdHbBKG5lvDfXxI8U7SIBg
wDMOpYfA3MLI49gwpddv2deMiXuqBCbr128QTQLQrA2runHcrBOONFeuXT2ar7TZ
lvXHgqAiigYfz+0FOMkdpGPUCYovtyWWZuzVG+UDVXUBMbTvKFhO8nVVAOTwUMss
MSwkTtH3RpIOzu5qP0aJCfOzwgeZ2pNsw8NMOAIWRfIbsHbJYSfSpSfy37zKUt+C
NV3vHotuX8PW4BpCaJwK8iNKJOSZuThco0wtt5Xl1p6RRTJhSnOowL/n/CmOkHfT
Jbsazw0XE6tJyQKJkc3R4khyz0JhzU5a/oF3FTzJM/CXKsemk3GtxmqUxvNZ76p3
ScYr5+SEaOY+F7PUWrtFQlHFqF6toVydMaW0hfK3e25GrxpAiTWTmwvtBU/EkSZL
k/RBdSj0RhShFoy/6UKK3wTiJKqIPu3CUzSGHQe1Vss8dYsvZK6qfK7qRe/HNxwx
gZV72O9NSATeTAlAM8h41oza4PbDEmJ2guPhnR27cBpeRWMQZwAI2kPPOcmb8y+l
bzHOajQ7K6Z1/pBhKoYIS7gqx5ZEGnh97H6Iw/9+JJcV0m7p8aBfEt4FWzJPScs1
Cu9x7768lh6V7SWpIlZtgmGyg7W2B7lZjsyAgHf7PIVcW2Dn2MRRVLYGQuwhEt3d
eQbBIvxKkSRkzAwoIDvWwiTVf587rbOA1KfRmufsDKyYqD/i4qOMU6AKleflMToH
qziSgO420776JLHGgLcgq17lXiftrQenK9CmoM6cJ9MhM9FopgvtV0uMOcCTip6X
fcPEvhFVjrQ8sEAU0+YURpfiGPWRNL4HGFF6++oNTSkvdCeMU93OSlOCdxqPVnSK
+YdHXWeeij7q8OCf8EBkRvUH2TvV7i5m1KL+csSkKdunVgs0UUFNCxGjby1PeUJL
NhQFAimP9gCHIw9rRrPmlEjTbiuUFYL0Hn53oDIvDV5WHGg+6jER3IR6LEfCiZQ3
hXd3DIv1kH0aTJmW4DkmrCkcd93sWj2Oy1B0dq0XO+NaIPH9mSGM+9IW17wbQPJq
CsgXxDu7MaHeaaEOFwW2QKCBBdme9JQ6erZYRfZtLen2wiR65bbWKqqmGZMXDqa/
d/qnL8AsEfX2smVSvYGDcCqoSz98RWUiXGH64jBpNXDwyBthqAYDfoy7nfzOkfgj
V1MnSD6UOJjWMlyh8tG/bi27KnGzi50dJI84tcSRQLPoRlsCzX2xRgtXHZkine5H
L+mHiQjFfh4QVdHQZSzKt7DmiSXFnXEkvsS9K0vqYAXHiiGtR9TDXAIW6MMXuZe0
yL7dnSufRkIALkB+a7ntIZiXkSMFFU+pyN9xQ+RbIX2tgMIyV8LGEFF2wWZ5Dr5+
pXx5k7HFEQpW2p0zeMTSLUZFkPKtnfWlo5ciiTBa+ayvWje1xQ0uzedkLWgpdgV6
m4zvn+nq7wHXM8Lv1XG+i4A9CrRP6SD/R1Maff+BhM4UWHb/ywOS/zo6IJaBo1iU
v7KJhzjCQuzzycpkXhkXnSASkBn1kAltBecO4t/9WnIVKwtWBTNx35YEYmvUbzml
yjMcFl59j2kNwTMaT9kRGdREl/HUQRo3A2+zpZ7a1THhED0wo4HI3Ux3dKvISWA6
U3R5WJxgGnRTfB2RzrvVd5WXT07iCAUEWCD8sX/A0ciFrqyuFYjJH0U8BoKG0rmn
tvOcB2jJoUPE03u3QduOhCM/1tXAlo7yxxL5ROe1F17mMHeIZOlQnq+fpMwRpZ6k
QIopcyhWQwiSta1d5cFlkDYzlVtHXWVNXRthVaSgFWfOaGOqbKT9LEHicAgFX+BU
IfobAaOynyuhVEr6J7VK5UmaoJSuHcFsXOFTHSD6A8SmckO9KwvSa6o1UhrCUb03
vfo+npqf7sM3veviQ9G1/fD+tVZ6QQHPbfQKDhBY3P+tsDgQDMy3pnuJapq/D4AV
kH3rpbco2xP5FBMDxmwiyul0lPDypgwRipI3yzaYldkGQ+ntIxKVp5FRxRsbGlr+
pF14o/XIGLFfyI7upyM8o7XdENJveppbAe5DHbRTXUIcIe1x0490FgkZVDpCwbqK
7ywLyDWyMyYAs4hgia5VK/6jXbsjto8nL+PDW8pel63Qr9lP5iUKf4Pbswsn34u8
skd3Q6QLsAAaNeI7KMlPXSUt+atTKuxn4u8J2QaDnzh8TfW8BrcN7OoQTMsLuYRp
VAuvlUDUQLZfYY+ZXNV2DEwANAunjU1OryJolcJ+GprFyqkJ1KMonkfNdgUY3nUp
fBouCXsNXWjgygGdoMhelfp4gXTzaYnjRb9utXSwOxVQo7dFKw7wYEtWY2E6GI+L
LnuGGzI0vnzVLTVMlP0UWL7HZwrwu5mkxLp847U26B9KtSKWmErFCdo8voUXkNhF
1tVMxUnze5KNm1ygYk7THQL8fNxShaZQKWDYFkJ8SUXzszpK0qJtGznYgVBeH5R8
TVDoxOHg2gtgNc5Nd1n7pPeedM0XGU/pf8K1BFFNg4BivNZy9ABbwIhd3Fe37ead
YNA2bS91VzTd/j2OtfvcKKV34Sbjdmsw8H0AicYiAjdmaKwpjXYQYS5QgpeiMXSl
C4I0D2+5Df62r3denQIsowVKi8emPxWDKN7GEBl+RLJEdojEBqIKbrsJx3QllasE
ZgZfqKWVulcBz/ZVssL9mpvYgxF3jyDHPaSApvKgZhuMVWjO7H5fK1/XsZ0uErHS
aWFoAAGX/jRlUAbHTlHOW8IPzXCDRDDmpXeZITTtfLSGyT8T2Xri/BENN/Xyn7PL
y8DuRK045CtiJ3SYUbxWPdGSMDwGNoe1hT84JT+NLo61GavQRAfIq8OQ1vh2QoEd
2B1UW/XsXh2OvNZ7nbKBX7GQXOv4LyWa0XwSg+x/KIGtZhKA2+7t4rv5KTENJiaW
qIe3CFNn5wGDbmMDM3gHQNRd5Pzue6Qi8Ip48NpG5B7gnh57u6LAJ6bBddmegkZP
rOyp+zCiqiym6D0qLDpk1X8asCgb70vADbf5d1HEqnEJSAS5XkFn8D3bT6vLiAXe
VWx5YTzsgfQErKPtuy2iOK99figZ0fwsqOi1jSTVLK2nQYfo4WtKDk5HMaqgwqyJ
rPjK/N+WIurnOHdmeyU9NH1uKGx9+yHvLQ5Gbd6aeB3xUV0nTcNQnQ/zc9b/7FO7
B0Rwel/J7dPIkHeFEx7w2Q==

`pragma protect end_protected
