// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
sYBANmYFMhoSJavDZMSjL/bcIUM7kswi5wFAWagM3pon/iL1zTJpxVSqPlbHHX8h
5v+Y1GjX18QTn77NJpskG3Q+vlEyJRCaXsF1hBU9C4/f55sJoDeLRfVS05HCMgi5
QxtAm0CbYzlRUhEiudbWlo3j/xzw5y3irDHmDnn1OWg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 23568 )
`pragma protect data_block
zSapKTT0ivlWNa488s18hoAg+uVn+mvRKXCeUcpVzO4LwA3vAywz43cTOLBoDxMq
dfWOM7ILJW/FVsJPomNBbSYRef58fDgXJ+5dNf3NWZ8CnjAcnWe50iGQNYrsWUN4
5Vy25B7PaLQTVz7voijDzQjlVnlVEkhudCLw/ujLlPBv9iLfgDaa0TZnwdWQHCVZ
vMwrbqKIdGqea2qKwjrV8p399PAGiH/W/25DJtt5vp6CYyDI0jfadRYSHq6iGFEm
51Egxu1v2LsaeWmixu53N09FzWnoz+ztoHlMprMYXT+D86EEB26oOZO00MV+7i3T
dfkm2RpSaupUYN8ScJ9Jgqo9g1CVTlqmy2fAXOyvwexTs40rFFPhmn62U20DtLe3
xx4V1a/QE5xkjxOJsOX33LZI0BQN/jbcIUTt+z53LI5BrpC20cG39Ho0PVHzRqeT
FSXFxEwNxP2EEF3XnaQIRduECFd+7XMSVKGM71fY0dgsryoJOTwUK/4mkxiPiK8u
PPczWdtTXdyMwBSOotl3ZwdpPzsa34uprEwp689Gk12bpuZm0dVE37ChMznwIhmf
KECcZr+ELFSROn9OH/IByYOehPedbAn+gYehF1jNM+Z9SgNs6jxVsoJv3YgGxG+G
ZsbO/t8kOQtag0/jBjuOtZeczEttDzNKQttHCSguBmdRAJd4UkCVjLT/NkSfxOLr
ImCzI8wY++bUcEQ/ocqg0heSWYrmgY5U2JDmDJCYfzz+IhZpjhi8A0pVlp4gX5Lc
c/B1NXT6vZ7G4sK3MmxV5SFYxbI7QpQUHvTnDU2Df7KGnG92b+/ZMmVp7v17yt/h
U5Ab/2XGM0NLE3PYvRXpMOrtoL1CzhrkAzdr8HL+3VdsmmUpK1PbmuJ/nu1/Say2
CEt88hc+BiYIYWn/uMrPELrWqIJWRsfYx2pDnngn0DdEvEv9n596BMAxxaoyqdZ3
nwsYmkjqrgEVNLIChiZKVtYV7Bsc7Q92kFQHATC4hzdF3ayYvLOor134iZTD8zmO
mfrUrsEXZn/UWzM2qIG8OgyL+bl9EprQDhHOsHzOQ+0iKlJaYGZfkt0km3rG+g3W
efokSesyzLBfJEY4pflRrCLyAp3kQbQoJKKs5u+2+s3Zt095kcYTnxMGJ7pNa54l
7dIUSKcV9MbG/gTZTkFqBKK5wIkpMK47QxLBlUAxJhxMuYXlVJgbyl0sp2Iwd8Fk
b49pHS16ZEfADMwWYZ9IGABoQDlwNbbvB+YE3nNrPPMXcqmybiMBPe1SZAVJV8ad
5Je9rOsuLdAOLGcgtz8ATIc5JIrlimOgkwDTRaVXVShr8Rp1QWb9CdCcHTVFjmNd
R7gbGKjFQeoSaJi/3gXt0PyM4zelF8NZRobS3yCp7RPMRY4JQ0yJfmUYeolkgQrQ
oR6to6KdsclkDCBApNkJ4GCVRs6fF5a7aA+dqOq9M8P2XcMsTpYh2Kr9WwigB+9K
3RfV0kQ85p5LSh+DzQr3PJ77IeScOB9USPnuTGHQoPFI2ZigFAvx/E0nJgTtseU7
1Sy0oaymeuxKJYNO+sPz+kumZUpgAuWBW3F1j4k+XeyTogjUE1a+pdPgrkkj88v/
7nW9bDFHsmdEL7HranyQ8Uiu27Dy4FpI9WKK0kUgCYyUB8ISYRBbLyXFrv3IGRn6
XFNtQBOydRlpiFm6OotoiP0BiM+bIzHV8s/NM8oeFrxahbH4ZFvCXhANZIyFVxf+
0A1m/OW81tzTFGydZQgr3fJ/2r71GRzLcbLPBZVOAXzHdmDp87SexDRf1m5FurfO
VsubCknYqlOpm/4ITSLJaPT9KKz73C7RbNfNJhe2jpn8V67HUSOQiKgJRrD1kEpB
QR/S08IGDiVpTlMLLaRiJEs4YxS+yvxEsBE7pD1XmnlZ0Csat4nAAENjak1YKJUc
WOgiZM5vnN7+GwRpHrXyfPd0DuhKfKxdn5pvNjq6nSmKRQgKigcNV+f244ORD+QY
AC6LQDR+bVDOvWRm7uAQkFVIYrYT8v0hMqc/YRz+SuXXiWyNgJXuhLSDv/JGJKNz
PCoNFmGVwudQS3t+m3b4EdO13QLAzDowqpZkPRuoKYuKFd3jUaNCzsUqc7SpVLs/
CuHLq9/mQ6GAEVSYiYwMU2s621vz8tZ2AJEYAjyjI8XHvZX96+TKbFE6el7JVof4
EDOOSYFsAOmh1k1aJeemv1RpjT1Rh2+eFHr98S9RFOMZ8PU22EPWazSS0yyHgy5X
P9rr74GBeoaWP3f6vdSftHxARE41W34bNLU1UgioqyAQ2HcDd4isLW5UsT4JGCfk
ed4ZAt/io4cSUm1smq4FXjZE//wt4kiT7P6oKLRpKNjwHuzaAcvf+C0nk0I6xQlm
xM7+lJBH7+T59BTICLr/0UVV+SHxSpw9OiuLUpPgt1rOA+6e6bVcA2oBrWzpDfoG
KiKPXX9CY42cLtqb87pEZC9uclYIEsqGvWCqleGXMMMQL8EQlRHIS0x0cKrk+qwF
DCCDr/Znw28p/a+lDCVECyKYj5A86VsZ4TX6AoLYN3R6TtxrXKekNowMzClFFjIu
aik/kTLuwKlPfgg3ioC0u+U65alKvmRlP2GTqKeWhyHzgzLbydrOGgh/jDo4XCTd
FCXfGhBcqbKVSanxrplyCJydwWGV6w1GKIx0Zr61wBacl9PonXiiD97QmDcUJwIf
ArA5YdNzeAK124GG9RTvkgKUIE7azieH8FMnP5uKV3GCFb5FqWKRdNrcdSE6FZuT
ThQW1s8zBnynjus/01nhUQFjYocT2hrVVY+zR9bWHdtSjxbG5NaEwkOxIQ6Cu0Ak
WNIySyi9iAq0Az1ITQ8bODStrZ6gqpDCOaM0pCedYHJzoDqnDs/ks5X44xeH2HvI
0m+Ob8bFoCQCjcoeTcQokS7bJt/KXned5bmBL5nr/g9EiO1DH79dv8a2NQOZg6OJ
Rwpr6tF6ubAztVmrGByilgLIKkanfv175kx7zHwTmLF4+TF7lBcqzpSVU1l3Kvb9
pRotcwJBFPXoeD2opf4842p2TH9/QL7Y/UGwb6rLihLyjno7oRInLiQJQ7Zun10R
eX3hOccMjyOOLxIPuGXG133goF6e1P1lgKS28UQSTvO8gKRT1nfDQxqQkK7mjVt/
oZ+kYnOEcwF/HZpFgJIq3yJM4sNdfq6GvJv1oozrx9HdfNepBpmL9onfdVsaFqVE
MRXlpq95HaUeXW9OCGdafkOMb8sDaHd4pySFIqwQskjA4yy4boVJFC0cCZimUpIG
nhWLObH+1gJEnAZjXV/8xzC6YzKPlR7caG9mDSXHa9Y6a+BJ7666H2BxUdztOm95
i7GtbH09rMPlXAbJSpqWWiTdPcSAWEp33LDNDDYHtGpjkXkDEb6KA3qJktiNNAXu
y0qLZwhmrZHAnydOFx5hLAhNO47wPgsAfn4XMFtwf1R1ZgY/Ru3v/LFHorkUDWT5
vHWxpUc/BvD7RQDiAoyilopxCN8hk+29g7LbZSsuaNkxsfZkw1N8QcK0x+AqgObQ
QuQeDZ0V7Gxtjhion2h/suXWQlPYgmVhgmEnDpEYcy9wEIEBDYkACyOlD+fSmcSt
8H+uNyX0w3tJ2M3IeyKOENfBOF+r96nsX2IIhY73NbMS+XQRtPCcvLPJ8i4Op2cO
9VSzZNiWo+r6S3/oGwsY19hfufuB3aVVM/N7m5c3xqK9JCN3LdDzq0evMih1gIOA
/+CzlFT05Q60IjPGirXs7oAt05dybTaZzvGUhAqjHxOooBx5HPNDAFJuLS4DtceO
b7NJnaV7JrbjqbAM0V5wsqOImFsZcXSHMsBQlwsU7py4bjDNF4WI/x54zh4yDHxw
8UbdciNSAV14/tl8FDHyTVgJrymm+iUxWUStWGRVq4gn0MP2ttM48mHCIhww0rXK
DzcqEa4O30PqBm7aX0jUKGfhWiSEG1mCcNv8YR7yrf2STmzCFj1p0+EP2Y3ZTAx4
Ui38hEMpzMud476sTOgmMTrRNM769zaYPy03MNnv3kGvq6AsyKHKUP3ctA4S3KzG
v0vNcYaBghhnGdhXXt/jAb1H5JO5URe5vhYcWjgQjP6eBRe6Mrdu2tthA+LjRZ3g
l8M9va8YAwI2bTZ/rEa626q7d59jF96uf2LoiSuT3DAjh0Yps7DLkUAHeWeWPUk2
nKoHqG9/Hu9+f2GhjBjLZ1VWbsvQUZwy15kZX9+6Bz0JGVJO7PJF0LwUwJnH+xH9
W7XV1+GtbTRya5ln4FeKwf77UoaLP2iIMhgu5h590I2YTaRicjbQaeOR/8tWcNaO
o6TQyvqTjDH5c1etZ3tapcIzFoljkRfWlbDv766CzHexrSo+V8ZhREHG2A+NahJw
3mSlFEcxwarrQoULuQxsUb5IcuuQxNQPBBTOKM9KdNQjKwGrVkpbQxedXI37KGIU
NBr+sZb7mRVI2+K0wU1LCtvP4Y/W0LntBIuZzBcl9Sf3DYU+OzYBMffBfPdpha3Q
CvhkB4TNyVZbgsxOYtVB0u7IUqJ5rllFyepZLew7hhr0mfg6Ra3U9eXiphEJWAgu
CuyJtsCYPRxhOR63c9bXPwgX7d1Xw01RF35yvCLbqSI+q5MCLQ6vM8wAO9K2yopN
MsZ8EJc63mNWzzBPFrgN6+KfD2HDehYuCT38zr/aKZ6xcT6r+AI6TlBKzws5/IYk
WVMxE55NkX9og591pnLKgkJSfNjfF7vOziCnAibU9vA7+v4qpdX2LJiiCvw3rg5v
z/6r/SKX6K5+ys0ry1GsTWPC2lrf936q+9RFQKiPfvzCdM9h5Kxh1NwxvDcHON4y
VxfZXwDhMrJHZB7vkVW6DLN/DiS4Q6F3VGgvDQf+2KMgCNSck247LSG7KAX+Lt5U
Jygs4NTPB4uxNSKBk79zHB2UO0VP/9WtSWLVZ4Akj8AGu89QcTmNPAkH3fbceMxW
Z34txVK5iPT8tSOvJVh8guyqOStND96YUOf3ahRvT+O6hdATiiTNeDCF6ivEzGrW
+d+3bSBOcjNNGoX7H4h26DX5cYedatnTViBq87B+37bXhPjOComCcDSRW/3I6NPn
sDW/KHfFGuBU3cTCllqxHXtuQQZHqDV7nblyfjBpN9/wNVsO7Fu1bAnrujY7ISXZ
SxF2cq/bAIcH6uT4B9OQqkA8BDhl6rYXU98QwpLQWS0NjHOhJ4K/R7sxypQ+bZg/
Vb8fEF5zmpHWiXvv0EeQ+ryMaxbdf3V/jv2C5fLvuq5dm+ZAK2bJ18LCyryapyrQ
Y6amPzG1DZs7p+5XHhlcwYGlPqbNtU29M2joyy3S/zTP0e6kTwG9CzZOkzVKEO5M
qTbQkIcdoABFaq4MFUCFthh5cbzq55eRqSkTwuXGzgmrCBIu9LQRdgMN427R0ENP
57GTGnVVnnznDKK2Y2XnjQPm1l4UZ9+J4pDWAVABSH9Ky+Smtzty9OXoGE3X4Dif
0iRltsaSrlc3oGosJo4we3jfCYIkav/EOPyHCuhO0Z95SPBqtiTq31YGRoDUq/9V
TIgYwkhjCJlPYu8Svzl9kZHuPSb7PsaooTB2Lp/D7XIdskrb/wG88RsR8NaFDPcZ
m+5AqcaBJFaW/rTkSG2urpflio4BD+FIcrM1fGlFG0fQc7YotCBuSNFpB/Uzv12/
zbDRHCChxPjdsN6KoySm/mjDzMGboQrHRv+dQf8yNllbABzEAmqXGaxWpTnNAzoT
Otea+VK5Jp5vFPCIxs8/YUtjt3Lzb4WEhSzRbguyEyWpMJsmNMDBQy/DUaz5ETbm
pJQ2a5vHvRqR3qgMYz6x7Xj2YF/s+TLrEK8YubVGdF8C/Z9RSDr2XZVEjbRm+hK4
h2EehXFJpFXvgXJPZp8kxPiAlecXVxkfvysVr+MOSvq61Cq9PVLzLbWQ6fUtOiT7
VaRUcCmyhw9lt+wanBka265Dzc93X7tq2N4MGykGCFc1Z6t+BO7c5vaQBxRNrKd0
645N8VDeQJ41czJlyRT/ZifHhI/bUsf1F/OTF34Pi7a/91AELJzMPZN5CSDM9Jqt
cgjpeNXNg9mYz3rPCpZmjrBSVQCYwOsHOrVfshpNckB3Oi8X0QbFZyDmkKyEBAfo
0IJ55OoidU+midsZbVXCYUuKQ585d6JTnrSQXIaQFcw9BxzDDP9v+H1p0GmryymQ
71Z8zlZEyUWLoJWQ3VQEAPsfw8UnonvoHaCdg0wHFQBHFsF+sQqxH/NXMWr+H0NN
N4/7vPBuEnyyxpZnKIu/lMDA4UuknmFGaI9eUVQwbuiSYJjIuwN3oq3Ix/6djMq8
SnYmnY4mTlRw/mpNXJ3ZKtqyrZYkv6BgVp0e7TNLlaEnUI2qC1/0M4S7z9bnW70N
Ym/q8T8zFNcmGzaUfLe/XgqF7d5O7/AvZtKIheYWev8TEShcmDZg2r5nFCBxXHrU
TRcCHbCaJVG+UPu49xcZa6zlfkR7Hz1XJ14ra480sAzcaqCDEzPnqXcHVU16CYvQ
gXKGTcYoewT1CjOi2yc+l4fTwzWv+wYidEOt9iWGFmoWLPwzfxF2ABJt7elK/9AT
jiSn7ZyNSzDRDUjLg4+kfT64PnwaIu+K8fcIzUYs/Wc/TXK3Cr3x302ZtULLvZi5
83JnOpf2f4sKe9+ehd9hkgkZIMPeT+GtVkMxm8uAcX1yYyga2gSECPYk13Lmas4r
acXc4qFcBJW6Dc6YvjEwxMEipII0PcMw+UA/CmKxcIWu1SPzTc+tRWpZ/gfkeItk
cP/yiX/9gvC103XIZ/AlSweTt1xAOKCgYYhiWpNsHxuqPzE6E2KuxgclOlFqwn0b
1PiqHqTVVo7HCEwW2IUqczPf4MgrMr1A9T/xCONE6a2OjKQr9RQdNNBKFXB2zIqa
u1U919KDj+HtEROs7aG8CKiGd8wdyPBdmbY13dj2nFqwI3EoMWjpoY64REULuGhI
JrZs1wu1Nt5mTuLFi19qqUB7vQLtyqrKbAAubirbFokswXiAhZrvC3fs3axVTSuy
dWSlw/AwK8OkPVj2RB3K5bR5nePnkdDFRl3DuC6OVOOJ/SiuzpSV3JNejd5LClAx
5SBaPvLGx7Wo7kvOh9x415xvbpWh00Eihf9jezlw1CPt9Ck9Tn4CLD2p1Qoa/KLa
Q/2hg0ebW5SFetDRarnWsCnN+jD81LyWlAcZOd0oiM7VTa4sevzBhQBmqAvFlBpQ
+zmVf1J13p5opMj7+eslBtrLu4h7McsCkSpQkPBWWnKZCACsqx9ohM9Dsd6XSMAX
sqkGa5Om8VMoUwPuqzhq8nmSfn3GihGlbbYiblDCN3DhPAAOVFTpH8ecvSuXc7i+
4xVRCDIwVt2ORNGo8UeV30uZ0h+V2otpL0CPCnxrW5CuuvGnOqEyeQ73ALqkFo9X
00Uw3B4amhyheW4IcBDE8lwIWe8+2H6LzPDOpCW6uLx4B3lpjIDi0BUm29HUZpg2
sphuo8H3HwkdXH5EaFXw6Bi7i+4i538OiqpPtMMx+r9eBsqmDwgIMEAhVmG7kTvi
ARGNYyHjl5zOsZIo1QkJ6REc/zir0y8tzChes8n35YOctFtFZXrkeaaZ9Wu8l8YU
wZWRl72bG/gaj6tbyAEdZYbvnGLK2N/Q/F/4FRQrL3x3GZbW5ESGc04vI6imZH4z
Dw9dO9O8YiPy578mpc5lG74mL3qVPv2hEgB2JpQKEk2+qvAcVYgWtfo1xcLFF9F8
wdU5IJ/BCA2dpGaXYrEjBCzGkJIcdkKbRukSoPPT49Z2bSNPgC4OybRB0+KUNn0V
t2EGN68+GbmDflcCJ3PhZgrD1YsKUE5rOwosFoDXezl9V754uP4wLPibIkTzpIQI
Ndeq15lTqS+yl6Ey8Jt7BAu/cMT/UGeoQE/2MgwASkmmxPw72uGFrWB9KAc4Fevg
fvtGONgfFNyU+h71MuAaCEgcijRrLWYakbXNKZ/cy4YyPlJ8dEIvjKN2wPTEdumV
GDAazt+PPvI41qB/tva5Ot9Id0+nqjOvLELdB2LS3jhNV8ubnPkNGNya8+8AHfKd
M+8/f6siwMGiPPv62LbSbzWqQUEj/wn4St9O7WMpZV6mfLDINXzfOeLMiI5nDHYR
Ra8LH9BYvx3O0i60ztDd/anZ2d0kHKS7dcCl7VrJgzhDijwuKUlp3qf2LVRsA04b
6EiBZACSPvqkH7smsJMjB2IKxPY4HmS32FQw3h21uf7/yMG1ezIasriR/7+/SReh
ehuvTFK9tTMzOOt8TpX05c1IKGK8VP3KydIs/WB0zGOwot/8gnBKsItJCxV8qmRG
Us/trL4MSdBUDMP2XEaOlIKbjCivdeFG1piIe9SKw2M4XUAW143+zW30UqfGTac5
U3PXhoKVTpKH3m3uJsJQMwCYVk7hfxNKx4Rn+gDvcICtduAgyev3txivgyiRfqHD
I1KB/y/7imBuPmddS+lh8i5s6LqnDZM79550LXgZJUhBVhW1uBt/O58io83Qg0hY
uE2Dyl9/ImA33+8MqqdO+BWDJ3/de56msVVfvgcprb/x9UwaxRhuXk5aHOOuffhS
xLt5L1feGhrIDuWJoYyiHy5ZLOwsd78J8tPGyh9pLkPYsiOVyD9waTPT1Z0JKSFE
+Ej+tIm66K8q+TfTOih4QiOyqdN8AcHbBo/D82dhlAF9AXHBk94uRuguxSCC/LGA
bg3rEDpW7H7ZtyuIWuTZMYav5KcWoesgwxcYC7XW1zBad6+8DUGh3Vr7Jn9uAfYD
bh/ALzdYk4HuqAfLML2CENgBZ5k2dVCopFqadFg+uxuPdJ4B83YqHfYhVrNY9Yx+
+uwVHfRD8ziaQVINpETFZhxV3QgnTqJG8unnswERclOQ1NmJipLHd0YCNIKi81mM
7jUWBlyXQljabue9i3wYzgAggta0yfsILqNt4v+PZE9gbeCldEFcs3U0fEb4Ik3K
Y1gYeYW3ROAAqsq7WDfTJjBeibRqFU2Xa6DkTO03mhXMOGp/ioYrwMtfwU1R7FeI
PZl7smTL/LPQ7vQjqIPE+0ei0k6OVhukvDddBquVz0eMZElwTeqSDkBxjzJtDFPK
uTxwZXCddQjF23yaVvgREgMbMY+HwY0k0+4SWIiSy9KMDCu3uQwlxrioLMpqlGfC
mzP2wQvllJ4WD8C6bx545AMtYG9ADt0Ajz56RSsogpG8L1Dv7olIRrx8knmC+hMX
VeLXmNL8F546Viunnc1EP3pDvwPDA1fBSYedlvj4zdf32eymhkTXPT46Rvt1dFfz
s22ugmj75RC14c04xjJ05ohNx3DATsEMkb7uGSp6qo9EaCoZSiTzohSlrZQlvHux
wFtLVVEJLs7OMibFv59tMKcUsvQSZbxBpftyoyHyil0YnfK5pEVGyF7bsaIF0Mq8
Ho5fsWuwjvrxe95pv4nVSRaJz7plmKsbuXtbJEgz+/+cOu1xQiBrEyhNEdZ2julG
zuXqHk+mHphN5o/44CROUWot2LfzhEXPRm0994Lyv/yGi1HoOanc3to946pgDXRU
/Cgd2XftMNSMupJmN+1MXa0cbZDs8Kylx1VnPJ21QcX3fvjB4gzt+8P2tze5kwqT
RFjhLLzfELRmR//as16twlu7tvJs5KeVPsenCNmVEPDxwjRQ0kwwDDT7GGYQkdxY
nv+vb/PqrqL8IERR+tjga/KxPRi3K9rqnliR7woA6qMHOKqVeS4XjqxPquvIS9da
Wc3BFXzIGrflGCvrkQIZTJv23LVJ0DmWegEZ6VOODmAQ+aiUmIxXQpmfDXa5z5bp
p26aAAc73VOjHy+ZsL69cDjfdmL3+KNh5+K8eJu0beUoQuNbxmHgqP0a1WQir1N3
lhpPwz133TOYxLAhJKZoEeFhDlxctjP5pmL62GexOBODE7/qWJfp20Q//e48Pz7r
Z/dgrhbjkm3xSYvXDPwKv/RipyfCBKydmr/vJPFW2nuOgzjQNRsSnK5ch+vzEN9K
zlALZWRdSyo23Qtg/tCloCEW6RCWFwMY/t4m3kStYbftCrrSP/5hz83mU8pWy1Kg
zysA9drHE2AOiXUH3lVyrHmDhVFbjZRRMDTm8kzj7FIDI4y8OOacDapXqIyWGZpA
Tz5b5wfxOJQ5hvlMxg4R5O5B1qKefeW8OrxlTZuLVYDtna4GYFw3zUGDwRq4Tp3H
q7LUNZ7sMqKISYZQNqTwK1Lt+Fm7OpRvI6hUEs0l+YWmls1TRB81i66JbZ279u8T
Nsqpxm6Zu1c0Z8yAE/BJ+ec39MbGHsVQSBKF5RvfurNuSWIyn6xtz6BUoiZO4iL2
EfERjVO/1MaKed7mDnptzeYrl+vAvmQMhkQSzGqkV7dVyE6/y7R02QfVbRUldEQf
9z7x521QvYT1q1PEpGBq1kAxSDlFjAdW0W5/pmJtZTVgZMiaikhqOkti61Ioyhvd
bBRcmexMcCLuHo60VR7+Wpn59FLs62eRAkJy1i8yRnSEDNkaBrLy/4BEz2S8oTSL
zy5bn42wgiTQoXIi8tIHWmzsxIdiAV/Xqj2Vxbg3C991+vgux/6OPeVo7Vndb1TU
MysqpfbXKQTu0FubyddpcYIRcEZM2jN87rsLEuqtTu3JR7W5FByf4JsXwTW7Wh8D
sY8zadqJZ77jAPQ9ClulqiE35F9t2NutSRpSXpsA6wSlwcLBx1l52it5y7nwpU0B
ZcFezf7t7r2fjZbYDBOUFAf6v1vZMpGmXyxO8ZSAI7JxslMvkLX9Sv92wc3epv3h
RMwRtmpbAnBIDZci7ZVstdAnVq4D0dF9BUmjveYARYK+B1gl7mltjEoHrySSGzr2
3fB5wREKEC7cMWzslQJYYkQCptgQq/dSlGlmE+jLgVd5cKOVcQyWLce6z2yi0uEx
ii4kXlTParNL1IQiiZbumnH3N6vHShzF+qTFy+Mi1zgTmZDTyYxk1v7ZkiGXbYCu
MUl5ikPbGy8TED3xRWUW/sbXe/ZYCCppxPMlkazbCBLHRzKTHOq2kr1iwSw56nhr
F9Yz2VtMPaxKagloztamn97Aql56YcoRIrXZw/fXrs4oeRwDx/rtCStVNHZGyP0L
iCwyXYekczlx0ULGvln/V8lhMD42+KfPjF06zcOhj1HpX/i+Y6QBJ8SkOGb+iVfH
toNjoGYqItxHQjsfL2ofwyEP57mnthZcJ1fbnES+L2+McOyIA1fHdu8bnndh8aZe
eoJt7WYTu1NkdCx16ktTrjWStrAQDiIZe7l7/CE0WvWmmnmR5K5sVNvR1YfVWfd9
yYs8Cs5p5NXar8e23ylnBJR6iK9OSzm00MciXrrDgoZ+EhBaDwb9z7e20G6nyhl8
T+D/c1h4EEFGBBJ3sLCQxL6foIFETX3g84HPpNWHoB6Z949Y4zvsG2haZ4+nLLBD
sPAHX5GsCRjqXBkUpefJnKBOrlWSXN8BjiJLRS/uiMBojxbYskI7wn+BaAdu7kVh
+uQpKG1dPELtXpnXPoUKh78qfbcthS5003Qgc8qKvSEHI1d/Y6i5YL5PWomooG3Z
4ic8dJfzyyEral5lHfPnZ+rH8dCNl4zjNUhFcTn9xCaLPwjhbd64Hmm4/ePpnIZD
jvDzA2q57OEU4GfwdCA509gKXerciMhrEJy7rTsOiUIr3PuT0VgsTV06gsJQB2qp
6panjop/mJ7oHUs/yhHlcVZLMAUGQUpeOtbrIvEMQVpWe00HGHEdNF63qeC2sCIt
BIYYkRZAzAmwIofXlwnowOndXMt0IoR/j3AHNC0hrhoGslwdLzLXWKk+woSlPUKa
96vGdAYt5Bcj7eYEHH4O/Gh66QTqMK6rq1cZnOsYLvTvDUiGawFLlYFBEQTxAkGm
XIJvYniPAHOPHqPJUoD2dTe97JfVBI771DeHGqI/ANuUlpYGgw6kD4eF8W5CiVNp
LB6yrIxseMbtAW1mwjXZjm+r1ku/NdsawteVXFwha5aMFpTGxeT3mw+baHWr2Tk0
5fvpsDSk7womJh2dpBbZs48rK/HEmbBp8leUVQNsePIUOT7zrODOaCQSMzx7FtjT
LSrihH4Ij5ceawmx6HUSUCzhXxlvuwm6WuGcSXbObWc0ppe24S1yEkCoRbVzmB9k
Z5COhoGuWXlQjPv5CzuwxkTdpJEv3fPvEyeP/wlsbwD93M/0pjOe0/7z8g4wOFTl
eKggHX+3ixvaEkrps3svAc9QZKjhgbUN+I2fqh411ISLY0g4Ze0C6jsuSwPfAKQJ
7XVtbYNcp+9tSz41KZOQTzP7Q9s3/w96eOkS9ryRKh5JbvIw8fRioq4oWIGxWcAD
+XFFtbbtWVJgNGMR361HcCGW859cxE64vL11AxpYJpKvMYppUITWHUisz3RAYEvI
CynrWysDuc+jTAZ7vN8m4NzI5yDMCAFiH7EqTBslV+w4FgizCoutG38QqGXwQike
sSqx4qw8+om3k4GCBjxsSyrYqdU25DCrIK/uUVjU4V+UxhPh3XphewMYbpAKYXIM
ovVlHpgcH8dpcWdOMkDIvEXodfq7nO8nDN7b704+HahGrcCBqo+hP0OzqWQnX3e3
84QC54l3T/skk8zE66prCOv++sOePWkeQkp53l3qZHuTRME/NjjyjTBT5iTX1+fZ
EDFfNapmWRUwfkAdAhlhg5s9gX+3vWJh7HdRCLtVsS7Btz5CMzc2T/f/LxdCeRDj
/WmglUZYJXcs1VTWSlPgzpTcotPR0Aiqhze3vSudbHIskZkpaTC/DHdtiDi4Sa/C
1XIV/DHOLyiK8n/XkVJM05u416MpR4drnSfD2HOo4n28uxVFMAXq5qaekMwotBPU
4LUb+zBAJqMLj1wpZ+5O3GffXUOGJRQq1J4eQbvNsIBFRrEOsq2kJb5bS6SxKS7F
JEp85diP73pvKWek4Waieanuoq4hY6yDZ64BzpVrhycDQx0ENCoBV8DmmdX6HHty
B7UEQCjvxxGQwaioW/BCYpBOuYSWLlDh+kCGtNlffmVZkmkRzmsA1ps8jkD4uhKd
8frYaehFYJefFxJh63D5POoioU+Pkagx1+Vte5agGXxLzRpWzhuVsPqm3DpdQS+e
hmD9xGwOvrXJ5r7qVQrohq8ynd2WlpWv0DVCobeW54Xl2liy4rMHl6pC3XXcbt2x
SHNi9XUksCrFjCI09h1Dfi5vCeGJ8c2h5Ojz0rZ/g+LT6FxnVywfu96D1NOwAo6q
YMIg3hzJhcYUKYWWlpL8mI1V/0KpsM2pDH1Tsvga2ezacWuc07GaQK1eOiGeUyp0
QMKrUfQwhhL1k+pdPWtMy9X9AJT25Fx6jPfjiVkUoibuXXzgDWO2afPIWRVDS+AF
Fu51uG8Ry9wCIz8CjR6o4vL4PCm6r3tyQlPpSZrd3FAzZrGE5TDMTyLsXl6EEzbk
DtgntEfgRF/jHsyItXeyZA2rulrqBdE9Pcat5kXMGmhfxiVpw15FYFDwquLcKXrp
vfJ2VSieunaf1Z/DsSfa8B8xmBVRuCQbeBLBZ4iFk0dc9OBftPXO5koF51wWxcN1
QtkACaRfXSQ1aaOxifQPy5cdepIi5Rx5c+v66QAMs8HSQv3b201sexqvnEfJHAJ9
q+WvSysSPO7QWN+HBZzwX19mH1DRCLsTm2xWhPfQfbgED6jvt9VZQqIu/TTB5eZb
GjzDU49kDHvP+0aD15AIvqGuFzu020OdZpwLguT5S5AWtDaizZBPwX7N/8Ej8koZ
PsIKSuzQVCNDiOlFEAh8+VN4Aj+MFrb9Th82O3tsPhFb3Ddjv6qWX8RWeFTsriOX
g8eL+aiJj0MqGZWWfKZeSclUZaYsRcnluBWzL/cQVL6fMshhMjkguDbPunDyYmv6
w/s2fW67qoU/pFadPhA+NIYLE4FybPnUjaXcVydKgKVjQpqKxIvCN21veMam1afv
WMcAgESYJKAITcoYfh95EqYABa7ystVnlz3//r4T2oWW+F4X/0VfaHWiyyoWIy1a
BnQRyW57rMbWkXMwSeN/15MsEEEIcglO6ZywpmtLNLYC12Ba0SXaqejIG7RXbkFB
eyZqVZuCqxgi6QVHSeI/4/7AF7XVR3YXYz+BJWmT7Zfl+PnJpegQJCKlWZTGZZ8w
HDLonHEBMTQlMWj6cW3aoFqcXRxs9CF9D7tMyar4WvtkhhpfeOlopBfktAkQMIUt
LOPsCsbYVauRfG9xGsL2RaGD1kGE12dP83jwvDgD6ZOAOnaE9FO/fEbjOLONk3ex
1mrApCnqJZtBXS0ezBoTXXVA65AmSwh1KrrbszZI0oPUiXnry1Z3rxsOf4PmRDrF
/O15wKY4G4YIWc3+okjm5lQP0n/JF/7k3tXwei7kOyT35ZKlkAuRZluHMuJhHcG1
/X5krldSUKshc02PlCd1NCQdCCS5+90//UfU1LYJgMG/UaMloCzH98C54jVZiA8N
PnmCk0wqem/AC7VkJ9jEwIo5KVa2wlya9wfMyaBBmaKXnuWz87o9B0RDnBlPVknA
QwcUpsmjxYiWYwkpjpaVHkp5t5gkSc6o89Fgdt40dyeh3VM/t6TgbHifDPArnT5D
b+UBZ8x5o6BpgcXpxTg6Ux2FTgCT1FubfKgtEsIZQr2YUrQvwWH1oZwGxQx6I1Dz
OHlFV6mYBDN/jLEHRbTPJCrmUIlD3qxmt7cbgb1kSPQ3n9eXuyKUn0EzkCJtSMO7
J1a/z+COWhOGFmk8HgJsRIuOxz8tuNeOZgQMQgmnGdlC+DNTy5gePFvEZmQAMVlu
JziL+R43G7jmvoB7438681Pg0TNhxFWb9xosNSSllY/+VUHm8poueHVR6jo1xJhX
fmUNSl2TOCnLkRyjFFB08tHcNJhEy308aNZgby4ZsSdDr9lD3cSt17DPJ8zfQtxl
0K3hcyhALiGx/VvlV7o/zCkd3VxwI3vIchrcCkVfPp2RcgVNSP/+/xA7fFKFe/xO
eQGlBfCoxKGSLO0CRUd13Ge+reITLlffPos32sMTWV1jgOuaoMwzG8g4k3jCaBFj
JTTwylDbQp2XOutmYFTHBpNRHeO82CFHzVC5tcW2O/lzn5Quhn83B6IsZfusUHHq
CsrIGYvudb+6M3c9cQF9xNnVUAYDibhUhb6ZSIQVUxh1hl3Nu6vKiQEYdiC9J2yM
ma6OlxFlDF4EiUi+oYgSfy0JzTh5uKbDtjFd/qaqS9wt+qukRMSOgKXz11iAuH84
N/CYBtFsqC/t74Mx8muezsk9y7nxIwYe5N5PD9Ruta2gKcbpr+piJEzMSasYUQAU
ripzyVvU87NqiroSnAYWHua4Bx6dMaWvMs0ClpJVexoYTchktIYdcaq9Ye8fd6Ke
JaY9Q0dkisq2v5QrbrHRM5E4LsuWU+QT6tPgwtA78/PrWA5NaSPiH1ycuALCx9/3
h9qR/C7bR4oN7T+WbS35gBuoL50dwuhVc+njXS91IY0Bo/0skBuykYF2huYMiVN7
teUz2B5thuMqhNwGxCy5MhMqL+spTztfEGdLvzbBGfULSpidEssVeH0d5IqUT76W
ZsUpYAfPNYXHe/CJFrEsyRgRuvmN1/8wJ7ScTKntk1k9atlHdum81gFklP+/sD+k
DKD9AxTW85LvCdhjxNlytSqb7SD7CwKpiyv5/3ODC8xASVPnVGHim5TwgDjPFH19
2lh16b51UzrbInxbDgDl2LHmp3U6eAKpUliMRCd0axYEU8DpeS8j+D7Im8Kv405y
koXtjSNxUJJWSBur9sXO7+dxiWaJYwjzA0WAgxadMtPqEMkW+aecwkSIbeGFGDQf
gdiqzH6fGin2qTXdbZ/zkNiHUq0BPBR1Vo4o8sdKuEas0IHK/T7mEOm+uhycs306
k4AoiNdZk3n/CUKPHbRra29HerY8zJ/OVxY/6VBAVms9mr4VKgnzK1ealIpAVLzV
IAcjlV0EZn83qVvyp8N5v/DoB7HV4h/3hhys/5TWi7PPLvjXMuC7HnoqozbtHnHC
EX5Rz/zeRRjUuw6pVb77MRibhRyQViBLyrLlhLng9b56hKvu7gY8NDQ3uZEGvkyE
5T7MvBlT1k6aiPGCqA/IGIkqVj9Msw3K/DOwz7ML4Ev/bgR4GcfJjOvPro5UJNQu
tRBzYoln57tGgPuFJVeuzNYb/YnH71SUTYyLonS7E/WUqhVW3k3GoBJeLfrUpg65
XcXqJV6aUHgjrA3nLLFqhLJgiSc7iwtM+jbNh6Rf52BB49gs8Gy7Avd25gzT5vPX
gY0+F96tK0+migMdqMQiODTQbruoNtXyYXpTV/LDvuh6Zt34FDD+wR5OF0fGIZXM
kevvg27MuqnwEWXKcufOXo4au1zJczLK5m1abjM1LJMWNWU7pQABpPIsfEq3TWYD
IccYzSfrfiabgaa6AtfpU79Rdqwjxq2eZao2yUq1KoHHdUIquPtc3SXRgEwKArjI
w5xt90FRd1AlhmqaAwv/dDbXnclIvgGze3A2RdEwWdnEE0Tq5NfLNVAQ/yaO4v8Q
idUIAZfmLviagvzngFTk/OSX5OpCVM+76FF9WnKmH1khldJj3fNDk3zM+u9irq/c
1Vbg33foSfH8kMGu2uDLQgeL86U2na9+41FNFP1RaRLzW8e/dQX43Ex82oVVK0tg
AaoRr73jxlzdQrrpzrtdo67bxmIppU7/A9Z6MAVAUMlrhXdOJ3WgmoCVlnIvgQGW
bVfkAr2FpbB/q1jpEV3hGaXLJ+cUTtAVlRhlzlHB0Sw3ueMx9IcS8aqeWgbMpyFh
iKeUF0M8/S45fRPlseb5Z9LtlvRdLG+nf03wPDmLVegD8Qgggdo5sQZMeD49l7n0
JyxXHbCYwVTbveE6EZifOqK4uJzqDyig0wYEtQC3mHsZp8XzxCkvFQQdqwMRWTyU
1snDB8fXlSxKFclu3o2FeOQ6Ov3Z8obcZgMdWCdgt7P10rJ2mc7nYbrE+cehEvr0
a39kwJrP1K7+UYQ6p337rjQ4jpP8nJEcj+GEAwRyPG+mhWDbs6TjH+80HbxbgGda
tT34daHOeAm8jXMblnYEoE+v+sV7QgDbt93PYDPPJJJUEDwbr0mXKmzEc44U+sr/
K2Dj7hWRtPj2qiD8LgfizSMJG9j5HGZsFTF9Bz+me1kjsd5CAXfbmHfY/SE1pKQS
V54ELzw1lDCvzaxF1mKJ5gPas+yCHca4pemH7xyQ5fuIlMWctMbYMeUD+d1Dpx7/
OAS9UMSWqsi0qrcZw94n7Zd32LC5wH8k50DG6AR6MLsLFiv2f8qlNQGd9Ew2OHxj
lvJVabG9EZeFyPyk2AlwlgGnbLhP29k/oL7Tst+QKpdm3rC9TwppBvoRnEa9WQLH
I9JRPPMOigXGfdeGM/RdL49HtHaMNCwZ68TcnKlWvDSf9L/4iaeWGAYzdnFom7VZ
vrsynelHO0N+6gJcD14UG+Qjp5DVvqbGgKwUSToGqFhCHr3at1ehkm3HEsrh3MTO
aW86YT4rh+wjHESVjt2lknBPV+YHYZdMiTh5z3BwpxxhebQxuidK5ro7b9fuWPdW
xLKPjIsSWFpnM0IJqg89sE0FVo9YwF89O6uQSrxwgHw0agTmin2/3HXyy8kBHSbN
HHrzF9VTt6yyqU2nsn+QFPMkowB0FCiiTbiwYDy1eQTJn6+qcY9TXHS0KP4U2IWe
0eq8Ut36GBsS7IE/85Jqqr5eO5l4ot9PKQ56O7IOtU1+5GHl37OSz5LimW2md2B1
4i6j7V+uYymBkPZ/4a6bROWEPBYCb7o8OSpd5NBSKMJYkVTPUMTbqtC3idSzrCyK
/qRL+4b3lo7qFGiyviZYbHNDDkXpW5Rsi+mpPk2gyoC9hF6theWhr56F2UftJ7Ac
qiLViJFazSAsgtNoDBVwSrwXyqQEtnn3UfFR0E4I12BZyB/Py8ZvB2bXtKx42Rxg
qT0nJCsq4xqxEyq/kzMng/d1qU+RJw2aWQVrncpK1tHBkLNpe5MI1loL5f9FQKep
leGXP+uDe6cSo/a3hiuFiuFLL4KaexgzT8WPqgRQpsyKsGe54EFJKbCxIWQ4OeVj
zK/NUq542ysfk1SR7zKZxgfTU8aOJKY+X7tXZp1IDrAtoVBBUR2zQAcD1lkooMZa
gY/quyw+xEF4Ohk+TYPOVjIczUvNEPDEZx3663DBl4gMv2bIY6chAOiNifjnfcPA
P/1UWrWnyWuw8JjWspBjUyliB7soN7FjGKC99B115/dMW5LNcz9PW6e/DvUAtXsa
VY9svkXUq70/Le3xqFgK1BJjhqpZ69QjnpgSGblt/gusf45Jq/t+B/Kt9MWC/rWQ
mff+aFeRsNww/PKay7493jPjGXO6V2IzKbSRhP868P2GXPyNQvIy8a3sYEhminE2
DsvWNn/MK0+Y3V6fSCE+W0AYJ8bVCq7393eKBbHeh7bukgMBcsHuGSoUwFlzy07J
orxzQJ0GAIZKpJ4HCe905yzP8jG0uF3lw30uTsaKCxoJwzqg/uW06DnXqvsRZkKf
wFB8/PrPp+Bef2RWEddbjgPvkx17A2Or1Lg+dYnbOOV84Z/vLadRJwRR36at8lsR
3cpqge/sS3PZUCOUoI0IbAHqbUMXk32SKEmSfxY7nVQy9WmoUVeg7t/6vG9Yvg6k
DFAln8FlJ3VoMpax1a9M11nheujYvyirrBQ5Cxh6maE6gSzbP/POIl4AicG+SW0J
lSx9BBiUijHa2FUtRrOKG9EBSe+4bz6SvlrQUX3YqovK0pEAqdlR4zwR39QNteIO
JbcgWFQ3b2YorXX/+9hZ7bCgkvqJq5m3pihTqvi1CDfwVeZ6NzrSpzhIRIuVt9zE
9MrI/UAmT08RbKapH7szyGAgl78gnpyTGGISeeIq5m3SlZ2nXsvlcXHYnPLkY4lW
doAHlCwCPqiRPNeVKO7L2KqzMnhwuZGakW8MTBgnSFR+C98zzMOQBQvZLVLknCDf
RFdMj0zKeK8xhCUPzleZOmQH9i1Ilv/p/zoYquhT4ziJSz/xGsHKTAmuxOTT5evy
lmodeJpOE/Yz5KFo4fCxJPbRlG7bA0M6WP5TBKKlIBLNlpYIor7xnJwc2L2zA4Ty
FE1I3bmv8QRphBwpmb+b6TpCFSluxP6Skdg0uTq4ZWiMldovo4ts0aPDPvBUQ+5B
tzT2IbjdVC0BUUWjk9D0zrmepJKbf/ia7sN43Vv6BSBWhKgZjGp9IhGPdHmju0aO
rEBskOEpvrxtNgT2CzRoHpY0Mvmb/bzjUuF7OYSjZUmR+EDUZTrN2sb/w/0Pmq0u
wYfrWUALxi0cjRph7uDmItJlFLGlAHG/j21M1SsVxfExqU45OFx/5ArXjKLNwjHy
m/dim7ZqTLgWyPYNfWKfwWgTMxVpzEBy0om23JTokaYW5YzF3iDjootXwaRFRfOM
VRqxBQdTI33DcZxGEmsUKxiv1uNwBBED2+Qfb4SVCGFLzuUkJbt5Lc+ZAbj9pAbs
AKvPiRCtZtprTrc8KTcGQMrbyKzFomZPlD10dDQ/Dd4oUfXlNyP8l2ftksDlLCmJ
n2zTLQZat/iIzYFEMNPGTZ64u0FTUkR1Xm6MFKomFLDAJfzKaRhvj+zfFIWnZBUx
12yv6eim+U+rnqTkSHusKZ1ONItCXTLChddzl0mQKetGyXR53k4SlI79VXmoj7hQ
0nglCaO/T8C+JTz5uXnmj6fPJWviwihfR7rz9joOgDejFsZK1VHtUFY7tse5VoD+
kq98cdDoFrUrESTHo9WLEr01PRJvUg2+IuV6YXhnzslGCdVNTUfXtQWxNrBCwIzY
zZd4WGSKVR+Fh2RdogXKK6JJNWWevhkvc4ttU/ahxEV+FWGxg13HyQSNXr+7WoT+
HkPZI3J8NCMY0LuW1CdM7Y8L1rZPE093Vjyo1fia/dR3oDVDOHHq5oPrVW6k6cnP
cKGCSaUbZ1kJ5TW6zvWmlGbZ46xViii0aFY2BiAuJqF3stvMYNwqSGXd1AZsIwFK
t4Z6MK8i07+mpVLlCRM/Lzq1DV6Q9AlRXi/OBf8JEVDyY3EG7BplqY+5UzJUyY/T
SUY149CBWZj/dRjbLKjWdEQl/Unvi+iBQrh47aP2vA3sam7o0DD/2arE1zpDPa8S
pMCricKXw6xzGK1yEcLpuzXAWvo8rC0B8tWkeahtDzuHLIPUTqZ31XtbycDkrk6l
BtUtvUgtdFSmB+fwjuUoyMPws91Ax3mXylX6/GaYT+vqhDEGs9vk6rWk/BDFw0g0
cTBC+6nqli0hBv0q5vePrU7to36RT1O0X8/R6BhcW85radwnN+bJAol4jYvnH14t
aPZRmyzadzBoWRw/A03TY5KQP1YGN94UQG6Jdhjshm36brdot2FkftwMMmBriBSk
R08O58EnP+5K2JdbJs6rGWUXcvMFPcKf/R+CNy58Y6X7iaBinp2P/qF/Cp0MghkI
MQBRfBbSOQZKVNzviVK1zHtKSNhM/YXIBXsWKOhnjX6Vlp7mDlx7WxD+fpZXHUIo
2ksGBZu7UpZ0RQmadMGVfghF9m/lOurnF+Wu5cDwybYn0krAjQz0qZx0NiY6WHNr
hFfBuBKQkJeYhxfnqAQn7h3KxJ8RBcXOhMCIiwthgxtoRbbDn23cdnr/UEcq27MS
ZteDdQp3lmCAC+6y9XuXm8V0pWCFIq/VieO9JoaKgHBmTLlbT6W64AXWEFzEvjYP
732xm28pwBCJNq88/e0nbAFEFbgiptnWdmZ93aYCzZQDaLJCyfp+1JKwb0IlyLfr
CF34Jh7oUGaJ++WxK9cll6WxGR9cfrTf+arVfeqdM/lGK05TDFRbpM7rwIMneDta
ct8VSKsBI4kHhmQ+T7CMopd8e4JGY15oEVKuwMdimA7XKF5InTTOGpVngtcwvgtK
vVuK+RTVQzvbKslYvqr4cRG55qqviwevKGJONLqlK7bMUrMERAYfpWK2s8vGtkH2
tO/4t5b/NvgvQDVkqXxfW0vl0C0zAC5mr0ul3pYGuL/rhZ8gWYgoWPTQbzgaWYKu
eIScdYlMckobpWLo1w2sh4sDV3G6s0E9gLTziwu96/Eb0+BQpqoVA1lUoA+MlH8U
ezdMx3Pyo1oCGiv59lZvxhHvaby6FzX60M7YE1aByFVWpgA9aUKy8Pht1BJQZO0u
irdm+chQ2iKHmCdENKdXNjU9Yq4XCGZwuTWcrfzTPimcmFUwZ6XruJ50LSGeND0v
jiBNhNtjULOXiGUi+Iwupp/4/pLsYZmWK8w+sWX1KYqwsaKeGpZw4YIkKCSEibeC
xzs1BTcy+2wizhgZZjLWVaQjZsDNb4b7nC+aBNMV0WA9TJw+eNR9ufgZTXd/7LNp
RD/KEXFaI2BVK1SrJSmv/NWywGjwbhbMRmutJDzXFe1YT3sWAabzXDs19k1tUKwy
LR/TcWNRIKP/hIpmFB59eVPdSHFIz3YK2FHravySwVrn0omO6Y95s6QRMrS4E/nb
y4dodUAH/BlKbiUhjJSAr72D1YQ88CBRDSMnuXGZ/kAOYXKnOwGGLxseK/k4DHMF
hldLAeCGiBwYfef8F7uG9NJ4z3GLjbMikZB4fKx//2+MxxD5ALYsvyA1M8Incq36
VSNel/ofnRn3ZqFSccQPCmF0TLRJX4Wbyj67jMzoLnbJrOKqF6w7QnOkr0w0vfIg
671Jp6WizqJx691dXPrrydzzvOnJ5jtAVrw4FixNyBZwB1bSFHgJ28wPRFjjAXDj
kVllJB/WynyHxbVJbRGxwlQFdkp5kC7h0TWstQZQjpISV4hkt48yHNjPs4wZ+fYk
yalJWXRiKBaU6f2HNZCqElScDR8iBQdINtNK+ua+mT8eDja3Ew8kuR7JnK7nPiMm
NufEU9Nr1swNCdlELw7rogjQtz8ARe6LBVmtvcnrirpsJjUtCONqzvAQeiKMQDVh
2VNt74hWyBRPMk8GHOk/HekM6ZW1yunfebMcwH5ebYePF28aaIrh73aZD1dlTIH9
rEFdJaO8d8rOFtvGCZMV5Dzlwz/8Y0NI1i0HK4g8WxJagHaRISbxVc4IIje2jCym
h5BgXeE6Pz5Gu9mpXauHi1iV0AzZhQ2gYwNmmYkKqpXITb/zUaCdcOa2uwIykDPd
0EVx9Ax9jgBTgViMqpzKy47k2gsn1bNOvbG15pECrwHwl2Hm5vDC3hkS0StDpHbC
mvcch3qEHM97vcpcjDV8DQmO/AempnInPllTaI+2YKmtl5QurD80Y3FXUKSRaLgl
mherqK3J06PuZi40Ycqe+R2+uXmclOyx/shNKQ32vEvxpipGeVCo8KyJiJZpi7sr
5mR0GiYLMa+fn8wfYVYGos/LtPGLdMIXjbP4xsyYejXREaGkeMfAPBemWUaY5gW9
LOg1QHoG8qiDzYYfmqj1iKIMCTJmHBIisReZyfjCU4RQkNhRPYl19I5UXKFVlxCG
eo2IbVdN8YrPijDxuE+jeEO8c2UGUoluXdDAr2gfBUv2zvGPvt8bpiSGqhgEvpYs
iqEe/aXyFwcNphLLlk3N63z9LKOGLsqGUwbeE9cns1J0oW3DmVfdyvxuNS9tILSj
K0D4fGjG4H7XnlYUYtYX1W+/gShvi3CrA1+H6uLhnsprxAjRMsfvqew4QKhUoCeU
NKP//cQw8MWXlSxstM3ffvcNRs4QDsQzv2X+a/DfvZTMH/kPxea8NOlLna6hgo1L
23J41JF6T1nMYZNp0XGVqGB41lIRU+iGMLFiPazIrHMNwzk6/ImBmz31iPk+Nzl8
aKknUJqC7IvIC68n5bcaVg+iG1guDfG35LVGAdtmwDDrOEgBpjjxJ+G6NjGvj4cB
6vandvlOR0IkUfO9VwmyskMIDLsk+T/EzNj4NAV10hxWDO2hpy3JDY95aap9GvJe
IpEKIrs8uKhH2XVBbnQO+rnWPKqPCm8B0PiTVU/ltoxooSUjPPrinN+I/JTLUrnH
Hao2/OEGMZa8KzxPIX8zz46v1j4HJq8Yhpctgu8YfK0ssyX+H9MIedq84vrCjqvu
wa7cLm5qcXJ2A0WIZZcv1UCyncWlE7k791tbmWhwQb6XG9C1K1yEqAmP8P2IIry2
k1xhAChT5rKrHJN/2vG5/xSXETDNW+3CHtd3R4X5WYZn6Jb3iTQxvM5zLM+SVlCc
6HAXEFuDS7cajAXBjMpg+I7dDLijhD20O/CwJFSQKFV9ftvo5dCcNSch5Z2XoEF2
8TW0ReDM69cCQy+LkUaUYDJ0+hGPAlvDAhH7Z+QVkGc+azdjWiLXKKZt+LxSMfgN
AMHx5UJtpLCoT6KIGCpfTv2PpzBwDd7tqakSEs6BpsXAda9nVVOzRE+hYa/nbv7I
n9TUBrightn2L1mKrMdLLM6boL1ABPChtBJkB4SivWF+WaZ8rcXomIYWPRBsbILo
KwrUVU041g5cerQLGHm0nRTQkz8R/RsoLFW882HqLRxLH/S0rrWbUyuhK80v46UD
scdu8neEYf4VFcN8PinZbJShriRi1k2qHZREBFIEgsxzOn5xGDaea8KU8TxVEnYy
IpgZUYwMQM0rB76sYxDrhyk+d03rLa4FCzZgGYKCY3WFbcysXo5z28WXV9VhFXr4
VzVUfbUINBGRUwDXbkWe/KYCu/ysd0UUkj0KJKoVP6RTRqgD4X896k23IdHkb7zy
gSwS44ET8jC+Nz90TJwGwBih+Uggkir/89w5Cyet7INDbEbPzvqbyr/XlSZmpyij
ErnWzQh8rG2ZrSmi7OW+LXkVGqllnUqprFwwl9uoIpxHVeNRpo593xFeO8IqYwSm
t2aLko9e03xmFS6F9gucURWT20Lcti2S44k5LdtSsimUT7mDrWvn+zeRy94MV5k4
Bpu8I3os0glIe9fzKoSOw5QPvbOFc2sUxv2LeHWMV9uozzfGXjRJYIRv3PgHUlFn
HQvPhvoCwwW+09qEzH7l1LVBELxFKRYcrWZNef6hQ2hW0ZbfU2afTqMi/Pabd/Na
FOx/4z3qvsNDAfp7Di+XteO/XT8i/2k1XY7w/wc2KIAxQYDl99QGF/OxXU2dYJDu
mTM/tg2uaRyqqM7yRNrZvvmxUlNaFJh1N/zs63ttTIVU9HSLzEW1BRLni73naglI
hBg3uavYFaNsx4Ypk16HB5ZHx3yBU7feXgPluTorT7Y8hcixqZX2PQNW5F9NtDaB
8HZ8Xrtz7DwQFnvlm/9xRlHl0ZeCC1dGEvhkaO4rliw/5ataa+ohlp2QJMzr6pw2
Dx7TOp7qCgAMrB17f6Lv6Gik6p88k0JpRaeEGnkbKpks9S0KilqF3RmTjzE6aIRS
R/plhpMD2vlCFKlw/nxWAgzJYAq6nvPUj0olajZRr3P0nshvr1LV4ViSY124xlKC
GkUeo1zBpdmscF0O60ytFYRyT2cr9EEkhG3eH2c+rpfqyZd7ot3rZYZsKh8te8h0
vJNGQPpQHbi21txZypz+6WP0k0UgxadLiB9MBG6yJuCFKmKsX91nv42Tvwvi9Z4j
OBe0iZq665bUAsGeQIeCIeVilrFwIPODcRprc+DJuEfKhkgYGi7/ZHK2hDB9RBjP
rorv7oXREOvBSm4vjv0SehLlVBqoTcFRWcg9CxipFTme5afWMb4KtO8j8jBUY98d
G67o+8jowWBhA5TpqK2ckSXvY7gFn9lrXgqZaMLAzQETLMkZx2IWJKW1zGYmbU6s
Zb4Md2VbYwmJ6SzwIchmqSfv79QqbI08vt//NF19zUvpIC7HPHLKnvkEY0KjR/hZ
fBOsB8ZPZeaLrTbxTf5PreCYvymxLSlPrJFHY6T0fpDgG2tlO+YHarSk5VZmQ4y6
x+uQ6jvBHF5fOAeI9I0eWbFbpTAh3J5sRbGBFDA4WyKAKBVoab9v1B5fvehuCoOB
CvDWXt7krrwlcG9NbYACcYsj5TlLjfs4quODJxVhsmlr42gtpJoIwlyrJ1QOYoO0
oXjn2hNILHCTaZ6pRROvkXVscYYDB5BCp1O5uU2PDa74bobMvbUjTjW+rZuwxLcp
yNP5c8aW47FDHTZBZFEP+gkp/d7GnLVvu87/iDjCzql1G2E896HGAwhW5nHHWRrF
kH+F4g2L1Y6JW55ZIpos4TW1tnGADzlK4Qb1Q2rcHPHkCZzGXON8npODfmuml0S0
BifhU4Se9EuNdacr8NyV2q0lIYaGgTo8719v4bDMezK3QlciPv184Lww+xRtxbv/
kzvkWXYbp/gB3G5B8/B0au7o837PfOMo6hlO7zxL9TNzzuJ7MDf8dVt9yO66XlWU
fYKEePnbPYtfoLQSZq5XjeG+yhhwfbtgsQCBPBpEQrieVDvwVEuQJvZZ2HC9AphH
MhJVBfvIZTZvBBYBnJ8bs0gx52xKdKdDRoXEIYrp/wFAqGO42lZjVtUsOUHE8m2N
eTDcU3E7EDt7XJevh19rx1hJh0zZXrVeT+rD/RaibHOdNtHz/UGizZu5B13Zr9rD
/ph7WTMIt3Cqz4eNV5wGQkq5WZhVgbs8+F5QCTSHeVC1QOVuKpIDVERNDli5C5yD
c15+W6o5DQ76MVFpU4WcE22jO+UKEQ11x3lISb5JNhRXhIvvPIvXj1tvcfB+Y70d
cVMZ4lH7RG5ZfPLqSqNYSqDkaKf+k1YptBAUVhmrOw/oZ+YN7VD7XCV1ZKZJ+BuO
7HIu1SK/HKb93pJ19Uf1g/6hpnEGpQHS3SxxNNhppa0QQRAKzqBnVIXD2z6cSODQ
Jy/Q9E7BSTEa4Kfb7sI9lpPxKoZsvl7pS7IZJ6ZibFXZWKGJR8iJh1TZoppgTqFV
0ywdvWEgvxIpUns7dqNqzOgLxV0LFBnstb0UJqjLMwZdI5Zvp3ffNIk2GqBwpUPR
3hqrwLE6ie+nOmRJ2Jg96HcbxtFRv2cLavoeRNXML5yrI/j/p2cYFer8qdqucYtH
v/lcbUMGr7u7rs0crbz4jbz9Xhzm0LIw7U/l7SUM0/zTg/8vIEf/dft1NolXbegK
7c676BNLwNKENByN9ZwpLlOfKn2FM6fOuCKZOcD7uomQqbWloj4Eep67/wAa0Wix
JS3DyxfmWGLYC564Z2Qk9op8WUV0sV0J0nqReRe01bi7jX9pv8vki39uSg0D4dXu
8ix3Z3+/wYGdsDFO4coW3eOyB1wj0WlCp5Z9LKGxbcRZDBK18mlfyI9EKvQvpSy/
2ByLzE/ZG1l3kbxQ7D+Wb5HQVWhOomsgw9QF1bu2xLBZeXhjDz57YP2JBm9+pEaY
bd62i1xJMjfIvg33razCYIDeqCA5z4/9RbvB+jhkj5Sk65Nse9QeLMCUVGEC4dTu
wjL+cHqGnwIYiYRyiizXDV98qiMCbUu8faAtVYORBQiLsiWhc0mifqIZkZ6gA8R4
bwFef0MwuN5KkPnkS883CR/3xrLWdbGqlvSAIsB6KiNC7YYrh5BkCPw9JxY+9cVI
/5SLTP1kXvY466UVswRK8XECZth8cKv6meRbJTql7+HBVBa5uSYAXjVKmtmt3w6j
gsz5HQl8r9J5J+hYTfn0bn5mN0zgjreOGTsrOInIiU2dCPsulVIPk23fQKsXdYru
+yzTyfFJCDWmt0VSx2BjqHxqPn+anNkdpBiskzMLN4E2SZWBDNYp69fjG8mYL9rB
TgzWGNACuQlf4IBK51ohNjvKJv0bB/Tqw/EjZufmSexrj26yPLB6Q8VfT2dYHw4x
5FlDIALv9XfXJk1Aik7UoQA3MPxj0h9/E7MSdLim+WTRQGV1DZb7cGkgKVFaoWhx
JmrsyKxvILj/eY8VQ8UgdXpNqFSYmMSIoFHenlEdYvioGAxi4GkJzVD/vLd+ftdI
j7maShLgzN69EZoGqi8aqIxr8t0gL6TmQdQlWSzLi3bbDQGTcUMkPKXQsFO0Ew6x
7Yb6JPoucHT0wrVmifmVXIzW4OORvYTZZEXocnrbb2J9tuHOwreciaOTyXJonHR7
c6sILnQKKR8WvMdxn7wXVRQX1aas0Jv1KaOkzlRR0mXOmQh1bVfCW4JYokvdEL3v
2wvhWuKvoCCXtVr5Gcl1yZCajJgNEl6PgI47A96AyR+NERRuEDTreD3dortMOznJ
W2ytLB8u7xhyyyhmmpe+Ygnim76wAqkXjqLet0MDqh36n/g0UjfV1TlpD1HuQAQn
pPllZYgblXXOlRY4TyLv7WdYaVUOMCqFhxMSgjdpMyq/zwZiTt911GpOuy7zZxOm
OyCUpPuRCR9FJ9tzCeOPJvUk5exUYqYpVpSWkrv1ACOHa9vW3QClUWQwI9JFXqbm
1wLKFSbCpbwqCrMhU3et4GQHgTasObbFTj+rpgxhmzAzu25zY2Ft8XN6guR6sPij
+y1LuHuUEzodJuFrJS+ph9oPbcJ5v3HpTH97ONCCkG8YISVoRFdkihBM5BYRhKjl
dbov5zLZ7prj1uqiQmu9p2tX7dmBm94ZugK1gIra4bajlS9LAsZzU1WbxsMsdjHa
VBwqULTbk5Ylh8oDZSEB/6t0AA7nHSgLOWNFsKPy2lL1K3qydVkCL0c0TaUDvHG9
SGhd3cxahOWlm1XNPwEroLph4L2BRupkgbxWoZcOvfpUmC03HilmOtCVYhbo5r45
bcqJ1fUN40jVTy9KQykQ3fXfY5CEs0xK4vHAwuIG/KUFxi30x+3TFD+A7Zz8naJR
FJIzRNVxCyL6cNpWWAflwQ3MV60U2wPpeMDd+OdiXb9iGjZGmcnEFAfMwiCnFY28
l0XBWTRGAwepqiVAuau2Mgi+yApxcMLRBmalOkUTzWhrPISvRCBjP1H/Y4+nYP7x
qIwQf6DaHbwX8yYvVLAMODoNadr4+RvCMu6w9J3OgNOeN6iRusp3AUo2axUXOCUa
Zlh8CTr1TQMd7VJjD0dT44N/P+4TuyIK1TNRFKOtyyVgWIYhXvOxXwdojfhD5lad
bG/p28AY8mC06CBwHhYKAXlMQkNWR72wRiG1jKzwbLJCyQnOv4BvjtiMz+tFWG3c
+uwl2+8mxovBDTNYvPhCjIqBElQl+NTieejtjeQjlFjltD+7Sq0cWyUTVyEgetaw
eIAO2/vSX0OrFO1cPXAoImjlA9E89UJljYIwp+b9Cs2hF+Y13AADXWZkpNpY1/dH
XGTBrVdXhLmmDT++q7g9r/5ftoSPhilGWcuPKDRqne4J9CaGqXM6cikZV28jXsRh
cr5+ycjjlZ+IlsXJcrW8xlYnbjzDvM7s7MO6xuNiJWheMxK5uZUEnHguroIaSwAw
Xse3jqRQ36+gdvQgSrV1BXnLkBGxIpnS2e3osxz09rn0l/C7ESdU02h8d05iumMU
LgV/s16RYHCMoo7WdqZLjc1t/4vO9e3dPmmLzb+dQrN6ay4UYj4/5nRvoqPZDdO4
i6P+m8TSdo3Uq0l628JbEnDu7rWpZ1x9DMfeQVyYbSy5dVTGXF91S5bsfNv8KLEd
H9B9xCUk5iJuth9prgvEi2BT2EtaNBZUvkJ5W45kvMO2j8zsyhCKgbTQQmebzlp/
bLIGX5lyKWxfHHA52KHNX+AQcg2ww94hEFErNYUuvCIvLR+ymzfBu6KkDo9FRtlc
OGSDqBm0vLtns+Uza5ZzPqBFelo1bXUrJF8WPwNFgpHB4vVVnav3aAKVecJKxehh
hk+pxXzlfYyMzJ16uzsRKcklRnyVVhXZjJCKcGxNm5tEVwDqxBqcSi0TXZQs4NwN
0C2qUFWmTSOHj0WzHu1o4CVssrt5Pdk+LEjDjPeXS2dkmD1Y0eE9rj+nBZQWpKMV
5NMxuEEh8rHtIK+mrdVQ8LMtCXFmPXgtQcQsO9CBHOCn/raFYeyh5s2x7PrcEuUG
oAPxv/dBfGv7cf8YMT8PkUUydA7dvYsxuoHEJeoLk18VcWaEjfGeY5Q5YEb5CTW3
co81RjTPZXR4CE8nLP2KUSljoPNnHGGrtWgvy18SK1nPQxgZjj9PjAPBVEiBz6fI
Cppgbe+QB7nEO2CRY/S6rQa8o9LZOrvoTUA8NoEIuAPOSnycAzx2uI+kzR+9XEcB
djh6wKh/n9XmDp8hAoZ/NcI/qBIGi5KfZCY7eAQmNKF5zJMbAwPCDb5PqNSALhe9
5b0ppR/4RZjaz2h9vQcZz5zd6sJLjP/9lNrM93wYhnuQ+ta/9D13L0KLDlrIshcZ
YH9DrrJ5SPvBI0fmbVCkIQcGpzme3Pm2VyIXgj3qPW82GUG5A4nLMG/fpJbtG95+
5VbIB1k2QJnVtX0kAODGujXU44ps8mW6ME8vN23MAsPDmndPOV3b+lY63J5vuDWs
6YCYX6zAQrbk8ExsrRgUnmS3/tnJmduTUOdBQNaeEIO4TaINrpF0eRQQ99cYSofm
cV6Fb4VGi8EI6e3Fg+pWkuW/OHt/juv+JI3qRMqEXf5ds0Brfma22pqTF5rBVZo2
Vn5SeThRnxHJooU/ocD0Xy4QAXDHfIn1y9qLeb7dxvQlCv8gejU6tdr3HLTLyU5A
dC6OPRS4Y2Y2BITFpI0OB41pScBn/SbmyKX/1X4CDGh1+Isv9LI8jBxDJdx22WQf
4N+iHLL9xwnpBY4Z10jpIePze0hlc+k8fQ35Lm2Do1PZoxoLi2mxqmeDc16hhvFd
PoLvHkNaxhKrI59Ruv2rMmypEaA6jec8Llgv3YIcJksGTtBWpJzNpUwRxTYU5o67
gkHta7MBzWrpLywmnaX0O2t25a3VHTaVc0Xema6ZGMm1pf/+GqaMXnxO3GOKm+4S
zjrRAeMA2A5JsBBNIptp0pN6W4FV/lN/VPXyMhKFYkMCu7JTaxAyiVF+OVbLCkvT
TeEYEfhsEMdTgCatyRY4VcLuCgxIj201PmvbTJGFVdudRhJQC95j3Le3ZlODDplm
aoGkQYED6H0twycoximBMT8jUmYM4YzeGya0XS6xCcqWxCjk10nwLZUJMZqh7dI1
xiqF8eJEGtt3iPpWn9uq5fz/rtOOX1Fghj+RLL4zeL5VdpJx6Ho08IgAfLbzomph
pEHqX0YJtCEXtCdpV9xe6iWt1lwdqRKXJi8yRG2Zt5ZeGuUAG2qy1S4jSlOqcmoZ
9myI5ZD105pOXfxHfRp1I8obr+4A7CkK0ZDTqIUFwIET1sqpb+SQocSwHvD3bcXt
yZSb4jjBm1S6DLz6LCNxb3bK4UObbZisYTcSWcTgZltrxnF8Zcsc35gAmFdDgubg
2waDkSwCUofXAyoFF62i4YM0bgqqIZAKUfnz0I809AdpzkfA4l713Y510fS7hKLb
raEi0Sp7YDaf+IHGOFh7MUfJ1tRba9gOYhICB/43i8KM9aAsV03Mgze2zS9Xvs6V
22I6RBSvj2i+Krr7pgx0HThxyPuSYvXgiy5pa8n5SRVSTH6akt045Tn6dMBx4bva
BT1Agh9yl0zIV3dgXhDhFNam7Hvd+0Fku7bGgi3nWOAhBRfwzTXs3RbvdLkm5ZEK
jJYiI6X34ZukbNW30hyo/rRRj/MbaJ3IiFcgW8dMMRFh7MtQ29LqNRMYSq5tHsgD
h+f5HgIoDy9cGIvryff/bUCYpZXIjVyf5xs4RjcgGTnSP8tTtulQ+ntCkJcGMFnI
ZPRyd0qKTObep33x6NMnUgjrU6jQIKmoh5MJBUfYMcTmB8VNygv0V2XWBO1wR400
CuzzAc49tzziZua7sTImbuDRra/14K/hcanigd5ftND7zEv9BJvMOkaqbso3g6Sg
yz2DCIup6df+sFajbQb0myD/5sRKDKWsZ7EuyGBCEcCBWF5GEao8W0tY63dugrjL
jONDR8Yw3+Mh18ZrTrhVL5W2/D9gP9P092D43/I+i5OJz8HnIYWv5cCUyBjJ713J
eKcpcW5s/d0etZLqTqxdO/oLwIjGgNOP68yIVYfeA8U/ZINQwxRgTMgk1DjaFUhw
V4+hArVNY6YIAPkLBiPrEP5Wn0QRfBPReNKitC8LU0yGikRG7fnvRjXGylBGQFru
i4tcfiGcCt0G/47Pa9zKMv5T7i0mNCsO0XXR1BHhlvirtMKyP3qZuEAxAlmTbdqA
CQUHYG6/2JAngU37GEUQljLswdUIxekqf4HE9DrYcWXkgUAN50hv8WT4JQtJ94ol
EDh0sZb1OE8IcznhhJVTZnxDMioikcpIPvHa52gEv6Wkdx4yBwHsEprrbmzqCm9B
3EuWAfk/Qfq1biLsysATi9ojxfB1VzuuEbDtbFDLJSLf2hxH9i+Ci5YlFd0pT3mv
ts6u/gliTVt0iKJ/oeGtMa6F82U19tvfGQUYv2ZTvvPhNa1QJuv6zQHV1sG5TvMT
gtjn4NqIj1CgDHaOQlQnJiIYl/T6t+u3WpbL9nJwkEFOEItKTIN7vRTOC2snWXvf
Uz4NTWUac1lWBuSZk0tLD6OGUyt5gh4ANQWTB2ZjA6lcDR8e150M/vu8cYe15GCz
b++IxgHDoCuiZr8ps0jNpx2SyFrUBI2mr/bgdc8WjAIGYeLDFVbMOxA1NTP3jY+w
noElQ5NZ/DeuA2+LRmyylAJwwL03gWEnu4nCTJxz8pf9jpgsF5qTTtrGSDwX5yIY
8Rj5iuao6S3SPyMjtt/WEAcKG8tkJk8qVoAXcq3waMgckU2p9ipDH49fX55TnhJt
LL2RrVuKbgAnNrJR9M2CscwBxez7ZAoOvIUSS6K3pYMlZvI9ACYidsg/TrILwxM0

`pragma protect end_protected
