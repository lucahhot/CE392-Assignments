`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KVzxb+MdnUSl1UgTPCA44VrkL72OVfMETu4upSOzw192I0WXjwGf/JuM7ezszrc1
8xLcL5BqRl6yjfw/nbIC17rQ6A6jbXGptFoE0lyWfTHQJ8xIWGPqMHIhiQN687mM
1H+noVBXiYUadOYmxQMN+yXJYplqZnZkQhudrNAVfe0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14688)
4GjU+IX7Y8VqnL4eRxlJMyggubNYnlEiok0i2MB6RmifK6cR/1/KNV159SF5AQCq
Zn47JhleJVWSWKOqMU7wgVByQnRmZ0NQQN4T0XbOx10qgbHcX3JT4F35erEdUno5
Zr6d4JNzhExn7o4Y8d8xWaD/oGNtW07v5dGsUWkWZEfEN9gYKYTvi664zE3x0OZf
0QElvex66VDsUMbiIHjpdrZEeL1J9Sw2WIzRiAEGTam5f7SJlfgA444bZvm1sQsU
CBZFRZHFgGeqPW/iV8rpT+epoaPLDvmW336cflbq+Her1JuWaqaWUeUH/wnyUFaS
PQeU0Q/V2wufqWeijjGgwQC5jzW+hm2TUitZiuhkHwjQJ196r/BVbibI2bYLOf9C
A5Bmc69nxO55K6/m+dDmiH5C4GguCBEwD+lfUwdYVm6YYCPG1Wl3n5cMPFsvJ6r3
f60aKWsJdiGxbxv3DG+/Z5YYl5u4N762+6KydpzridL2u5f8ULcxIaFrWem03ary
IJ7KykCcBDrZFrE0i11wnAKwzzguQbYryOOxIgS7v99YxN41+Km5POriPd66JwGt
WUAXdIPMr8aMz3RvkFIkLzwdHfMUXpv73lzlhD3PsnwEUE0ONUssauxCMBMY/aNQ
PhQk2uAzg1Q5eNpJx2bQhLiYX/gaYqejFcZqIskKhdfGE0LMxFwPUjVOVjhGAF0g
IwR+n2tlPKr+sjHQSZg5Kwkui7DZYwCQ9Gmkx29opKz1RzWtCeE6PP2U3uDC+aZz
cCY2pmMNfWsurnX/3MpW807wS62yP4qgpFls7cNTrxQSlvUvcVdp5W5KSkgLFuMv
3uijgG6hskepjT5UipBTiBRhSbhxbJHFwz1XlKXI0T2+l+16jxVpVtuA5CVsAwWp
fCcKJjg742HrAZFqWJIs0oqk7EYiRQ7pSYc+X+NG1l7toFQ8mjKtpLS4Pf1P4Kdh
O/FkzLmBSB1aFvCxeim0Odetmz+JdLs0j0V/j8U0UZMWwrRYdQOk520fkeCzE78a
AttOqqzJXsN/K+U8uIZuBfrGAnfHfhc8EwX4j7EkFuhIKJBoLsmpLyWoQLZnB3oP
tLIPkEYRXHBmNl3AnIXJ5qO7Z2s5yPn4wN4wIWdtu/l5rncRJspC/qDCIG1hRYn9
48ihtW3JYW+L2lqkjuy8tG9jUS/m1iAciHSQGDXUV+3qARmg7giRJLRp2R3ubpKL
FqMhvG6MKW67PTmmXoundCKRceTaOdwSMCnSxahoslebM4Xwtl1scdqEbCHlF8lO
AE0s48Ix1ondsiqKXsHfBcNX1yan2Z4qAcTa27QSZrmdw0bui3HP28xYaJTJqT4d
mQQYtS/u44+IdA0Yknp5y8XKD5AeknOeB97nJls7XjlkqzYOszv2j8q5EnIL2nRn
kINhiGBjn3DwJFhKH/DvTS85WTGJU/iO5OBbSed2gO5ceQQg0Ub16gufvgEyxixY
miyyfE6hsIhNFOr9NMI1ZrKqNds3BVR93b1MgUlwWSYW8Vm5bXOtYva5TdvNhWB7
mGMPfwK/yb6++xcIR/lwR0aDnNIGyeYGTn6+A1+8iOTzfDJpuQTnpRA5D1VIsb30
WwMf5nWtda2r+c8uA9+UuJX/uHGcr9G3teZ8adC6V+NBZDRsibMVWEiJiTssukRa
eb2nntfENQpjBQrWRhh3ToPMtsat0LffvK0MN9ywoxFQpVr+jMi15Qf8TRIH/x0V
vHOBY8QZ11V0PNfWkwHufbirPUECus516CxBT9HgprXb6d1qR2k3v73CFrzQY6Km
LZo6TFW0ldhA0EQrXxOOwc9niUbF0THHStNHLYc3JPgWp+cbOId3CkEjTg298flQ
csiMAyhTW+krr9bm/ngrTuwpk5/YErmRQqQAaPZJ+ZGr/WhepSZOl/NDny9gmlMl
qZKMr7KCOXEdluM6Lj2xdraJze7kn/IIqu4uDwI27XKiSCiNq3+iGD7PCn4gaxmN
cJFYjO3K1zuA9NS7wIUUj6j0rNhUcEga8CNtUQR907Wqsf6W6yjy2fzkOT0DSo4p
/tGgO/UzBJSC8+cX0valLPobFhH4AAq+F8WbvGEIXWDCKHoGHoFLYsqVBXxMSFRm
nvs1/c5mTyNwlmhirrxTfjlin7CrpexgiBUuzTxtafR9qYLJ61KMjydEebxmQjNZ
Qv8yVMvzPzQ5LiD0vtyr6v9Zp9d1EyScDLPvveVM5gRqZZt3PC93c3TGMZBfNdxv
m5aLUESuPZXiCLMu/MudwG1KuZvX+biDlmaRbWvAcJk/unL0invCc36umrXvjnpV
yP7Qeki/lBRh67qcXJxuzI3GCO+Ki5ERfJ7hPaKfHPKx16ZUJOccy7CSUgGHk0mF
yKwfitWvfc77kDsl6uj4tGAYr45PG2ZQ8Tg+8UnFC3PNqdNy/DRpMRU4ILDoIaWO
cbs1LEXlCgrNbWthYnY/ETieypMDNLSeAxtILXZA2vG8LttyhPkXxsgzaDeRx8oc
8MxEoQHltgagtX2jRgguC9mdREnxMoT/kqgm771+lbTMfweJczsYJYgX+3nfLTKR
Fh/SK/wRZ0FAb3BpKGoaqIL6bOY/Or8Cev97enITkUQGT8gMjoRoe1ZbeCnm0dTe
PPzuICbKaI9XKsTfPiPlQ3wF17+04QFnOauxOk8zhsFzW9VCrPD/fCyXHNo0H2wI
sWtM+2bAqK9RXgyrf4NY+fB1DOPQBHKlq/wemqOZ5HfrP2wrnGD9Z9wZzCNsU1+j
pVS3qlsqWSQWoxN1n65q4wlhxc73XsF3SmHxOcb+6I8qRG6Q4HRA1gdCUFqfwS2o
QMFRsbZeDECeaXNoXfht9NV0dgkgkvQBj+HogCrTrgzd7vsioR8l46LGF/hV2D/s
mVLRSECkE/j0qhTlm3PwjtS1OU6rw64HbZKbX+NI9rGv6RmbVssds/H79SPGz2uL
/LwDjsoBZ2G9gcjN6SLcPIUb/Mt1/MnCyyk/LyhLU8pjJT67zILxfbMa9ZXX4CPa
nHp3xDgQ4pfSa9QE/K4yXwWyYuJmdkRPCFgiTafEzZ4wKxFF7IAOcoGWnOfM0WZc
4wVYLrSIpu3X0AY1SGTcmwkW7esiw+fSnl5sLBs1QrdFnoHyy4isqy/cUhVFdf5s
TH+SkAlqC/GDLRiX67s5JS6ZJAidfjjSrVLQynwBf01rTadCZEfynCnSg9OtZC90
ixtyQ1ykATZQNesHJSvp4z3UHQcr0bjOpzfXS5TFpXRVlhTFxZXTBgfS71ot/COK
BsMOIWifPu3DX7yyFwaEALL6bnRoexqDAW+E6hES0ihBhEdw8NBtOCGNsgwqSe/q
0bOnPWFvfuMnew5w/ZJ8s8mJn7jpJjCGZxUeatYlif7UO3Enj1PmiRtqlC2q8LA5
aUsZ1Y/e4sFYprYKcIRwhVvtTcb0SZeOD4IoOp4tF+JEue5kX8Uyyzb7tF5Q72TC
F64xV3yN7GlUObs/ALQE4k1z8990hWyg14lemhknbYs7gRrysV8myvMjduVDJQwz
SNEhsNFHIgNR9E9/4Wf60qaAvOSi/VbZSNoR1yZXj6rRtxpO/SeS+9Gld+3u8Ziu
3YJWDHQH4G5ywso7PBWPufZzenXw4RUR8FwFDCiAMa0Ppwft/m5cHI9s7G7ms4bh
U+8t9SILCwijULctcApOq4bXWoXyqC/YwiYPfuzc+462w9ZFeu82ZPw19RhuodQv
tiJC01tedi15RhQwSh6lnaXBHw9fboQ5T5D+0399Wzz7vCjAVARNX75IGtrPI/ef
cROIwozy8jDQRLNPP5Vb208nXYzrhyd7AF1F1G9WOFpRIq1/WMb8Q0DmDInbTF45
3XfA0xAm/6uIIgIhSDPcvdrVkB1JYJi8gn4WF7RcCZwjq227AiR8JLMOuahHiXRd
od5LO+Oxp5cKESOL8bQNrxbw1+Gvm7du22N6JP6+IBIF2th9VZR6mciBmhcWq/ye
oi0kWq6B9fF7iOKS+WTJXILM+SDivVdLYolNpFmk77DlIUCZf8ygHjLyF3CEophd
HAWFmrixYxj8MJUNffeXvH1yPeA9BJqabGzk3HseTZYr/GjXiTKTINZg2/n1rflx
mgtXcNPqZNmw5aMWc3ltYmJpjdnyZZ5er1fGy47vm2FoeR8/ppn3RCZ0m6SEIek+
OEq/nB6rg3AlsZn4jTSI6NO7F8q1d6gfQjvXvHF90RzTN0+Pcny9NDicJszX8vXo
UOLedR0pr3NDHO9PJ6ZdmclBiMStlquYO07iRtgHMwKHnyN7MnWTlyzxAbgn1OTD
oIku3pN5K9Qv/s4ztpi+wUFYxENcCEMHqSrOEBUfEZrZXsZukBaEMivqeNMqsOE5
MKWorenHwJur2+tsTJtb/bCp/5BPUL0TyZZu3SfjGrlRfHvzBre5wJueCFSfOSCD
Pe6qo3vJ9Vg+oo2I+Tb9fGYiKopRG2S7VODhFBeJ++87ecbxE+5E6e1l0huDgpDc
WcugFvlkhUHMesKMkSSarIuQZR11Xu3sKyfkCfBXUSl75s/2kmXE94xLNGJLDA4F
76SN07+xYbk6CL1PQg37ON0EuI0s/DDhcV98VxFpegdL2ld2H/shuScaCTpxhJQ8
DNmbodcyIjl2qh4gw2oO6HPvZyKv6RduGM/mM10kEkZXXjoEqQadMO7u7TU4Qpn0
q9iMD0gY+RTreBurjCS/MuuPbhTYxFkGawdJC9JyBfSv6Rnb5fv8Y5D0xZjheo1Q
JZCEY6VGi25D1iT22LXVll88XMbKEuKsNRLF2oSJBHQ+h9GS64FLebxAXPGcQz/I
M4oS9SlEoFdow+OebDErE1/pOSZzTIxiIgLgxkp+6VjjJdvuuBPiV/yoqYrJb3Pj
UW764rnsRa/zvQs7ROfTCwcMfvUew1AOMBhtbfbuivkONuH1DYi1fUKh/wA93W5P
1/Xq01WnVhkvtZQCbsjdI6qJPa5N5ganiZiQ+fzWJo2OOko7jpH9AlT8b5anqyrF
/UGww14h8GwYDIVBNWXlnFMkjtrnv2CjZof7kUFN6O5I6rN+WuXr0OKkPyXEV5aV
zkj3UELUSQY0mDs94itdYkVK8tOR66+20lJcwpKp1ZduhGbu0/vs2KlfFwtgqUYB
iFyNJYX4bbLtHLgxZp8M1BnseUJPGnGdq29IsKtqE68aoP2qNaWRSQIseSC/IJJ2
EFT8FfxGDgJHicNfW7kQ3bWd8C7B3r3f6hHxPubytS5SNgaYebLpJgpW4SuQREVE
uiTc5/D5lZbklYska04DP2UkrkyDLvWODrBB71sOc+wLKVXpACFej6FvnDhF8VwO
Ln9zjsgjqSD+/CKwv48frHm5r/N/GmuiDNpj5rGQxni4FGZzrquT0QwYVjQZSoHy
fvkTIYlTy3/pG8X9zYfeIP+t2HdcVpXiK0jqenQXycHu7t7g59IRGleNz5NxdLC7
KGd9muldXeE9k+OQXPlmd97as2/3ghhq7CIJmV6z6+rOQahVESpC6i+1Sksx8J5p
KhbErJRXdSuH969wEHGuMq1Xhn/ilj4Whkbh3FcUywanavVX2bax9D+5dvOcEBfd
vG15x6MEqLVaUQspyNjCbUgMreIcvoc0yUnjp/N30S9quplrwdomMltA2lHbz0x2
2F0k/afwnF0ebft5R94Bkq/QEfqktYXs3P7AwEj61wtF73hwg2atV4yQPIq2oA54
rM2FvYj/6ubES8H/Y4grs01yXuSRrRk7bkSfgoODZfROlhUwurrvq2iKpb2E7beV
i0OBDdTNzVJKAtyXnC9cUOK2z6WUfrcrbmiCI49gJFXaY1cUTJFQYGELTQ7puJI8
d2hNeGVkkPOfkZxvo16jn709LT+6bUF7gGkrasAlIkUcHV/Be1m7CO52yLvzv3L+
xEMuyXtYyyBFySE0ExYvfTHcx7IBG825nFbW/+4s4Gre6gf2xk+NqS/oelHkEIbx
+Qra0QdZRh538Qobe4XUgiv22dOhs9Y639dRTfgOtGBHB28bLqjP0yfBB3bwD8yw
NWyglUoIf2ov0p/K2QOUwaZf79kdlr4PIb+nUsav3s6y9ViFsZU8kYUw+477cS90
mpKQ1aZdiUwkYed0/NEM4FUR4MEypmoHKMujVCrOYEf7jcqyPJXDTjOhbya0N9no
0MZJFFjw72EOIc+aZYH/xFM+6fBvRdPCBI0c92rYNypcJMHB6ie7y5pR3jA0u/qD
onFegMAFW58J0VGj8UnUptMnYV/NlshiDBSLhCpae39p7w45pEUF1RhlL1ZNJrZg
4KwFLTr6fEQK8KmKzYeEH2gUGU+GWHwXhkL7VO0YLjJ9O9CqVbD298yLK993fmfG
jYKx2eVNX0kYOlOiupdxWcA9wvlwwUSwDUACSj8loq+H/WKTWfwa4jCJYgaLFr0R
tRLBQ3MklvUv+qDd1qXD08K8MPOtUO3zgRH1mYasD4lNtGo0cMScLrra/G2iH5GT
uZeL/wvVucJMPOB7dIca/3fzI+pGWNUDJMTEIB7TwtRQL3QrYZhBeOMbDC0M6329
HocloLGit3gMhBIOeM6GD7faQ459nxvue6DB2q9QllM6aiMw2MMjjOqJSVvHO9ew
Y8iOwxuHl+uxaATh0w0eSM2EgcTzu4cOs6u5OptmjyrypMhLEhxKjNYY45bAqKOD
L8klGb/LXwM4WFxdM98Xlhz9nuesG7ifnhOYlzlafap8gNJAx89iQxmCg8fy/rNi
4py1DGjske8O7V8RMAihILRLJ5we3ZQVUi5uL8PKQZDuLSV57QriYALe3RguCygY
nJbY/kZm6Mszoe0sb4EIAKH1wWUTaVGo6kpCsC0LTuoYijp23TCFAbrFd9gAwzpm
PtARlzJu1BTss/zbC21UEWMTokNfdLj/Kf/ISNyofpzc8fWte/G9KKHV88jPEsIL
FGUHLXbZsklcHr+ZTsgPftfUkzXxXzLiFq2JZo6vXWQJcUH9ECKjkplW/oAQokAo
ckZVzHtx+NudZGHNRj95VaAUbVvF3QeLSNSW4ExdPUv2sOn8ZiR8AeXDQce5FgZ1
rUyFgemp+JpJLEL5lhW049bkeIwJSWv+dpfzyCyOse7lLyJVVliseFRLJbdsnmsn
4wzQ1eQF/ZxHFBKnS4t9A0XF4lnXUZP6UTrk8hb5/1tvup7dOF+HqNBIG7nzZ42t
BXsHMYCZhkPTyA9ZXcGVb6e80N6WwCh27N5qe+geF1hwEdcrPLD1ygCL0c94J14W
JDc2ayjwk+2kEgETPPjU/aMmrX8hBgCbPFcksEGf/XE3X97mnIlsTX8hame1Sumq
NzAb77CINLlaqAJtpeKpxGki0tbSU1uFiZZg76xyQXkYpR4esrFwiKtL253gpiA0
ibk1XwAPoDgfcOYGLE/5u5DzjymXc3MLX5aR/3JFuHuseTvzpnGwa44y6qWM+d7U
Q4BHT1aUc7nk/cZlGZabduo78Q86ce+UiR7UzfccClzDBqRmk5yRQ4a0m4uoTSTZ
yiEruabk6RUJJ5X3AeAo7ssBYzTzoqHV7I3Vi3OptnzQecRX6qj354lBaSDyL7lO
T9Du++3R1n3OKr06q9tQqn/lHM5l/gnJViIxcOUDI8dvNwYAJUJc0ENL0OctG2ii
mcXePQqM9S2SxBnylHhpjH/uVS7M+PsuLS4O/afvqjiGQ4lI6Hc36EGRGGozjQq9
3BaUZK3mWtwvZCME/J+y3+oAnQ32B7lMbA0IrMEd7N3iPdPZqtn0dpFdH33GMlQQ
15OfHTz7uPn/Bk0kdvNyIwcC9H19ZVklp1stBSmXqYURUH3hfjKAwMgLu7ydDqsS
qUm4t33HtGBr/t0tb3DBwaQagYV5tlJRDTnDp8TEKESnHuorAZ5q4IodpxWr6xQx
mhcNSeg1x2CYx6gkvo3BiGj79kEX6C1WIP1K95J6Tgf10nY444tKdfZ8tI8jKhX7
cKUWvWKG2XyfiPxkV4rLS+sm74ZJAsNTrhFbON9INaobsd0zNi63CMUyMWguRW5Y
Ivc5ZXkMYTB7ykyxzs7wGQGSikI5tlzKnRbk2KRCHRrD4MblnHzfHGDJbnewt+oS
zYgneYLoTgbFRk47+zpgOGucgXw4NGFxrnWkBQxBGBQSGoujnsJc70WTNI2RdJkM
l2Vwii9qRFmKg9RnTB5A0qAzf48VN4yA7ZgVWUq4m9U91OBkhWC1H8i6sfY/TW9r
a5jg26fm7fHCA3tZ9PlkAwNYtDFqHKi3dTxKa/QmjPH9ET/+O0lusxW+d26zUabO
BYJsjbJQw2F+djOdQhEgB56eVdG5sw9NDj46nPBQcgXiuwT3dOWvA71k+T2NfREx
BFvHBQRZ70wBof41aTLqqNRfWZKfxL7W5zXPBGn1ky7HoWIZ/Wf475qLzRXwY4lS
4lLdmMT6AHuRjWIfyHpw4T/zqzjiX9HtZyTWA7GZ+YE5dP6NbJqw9agjmIKQFEqX
dgqCmbwcXLyiI/Y8MgeVEamMLTWM57ThrPp+hTHYhcnX6OXN1mIodMppM4FHabJA
lQZua71mZoGNcOutZq2Bdf+JFGa/yaVC6XwgxECUrNDtwYupkTdH4wGxFioCTiqW
VEa5NO0l9txpaQFExT8OmhBAx0N7FS+wkRR6loO9r/e1KQYn/2SYHzolf/WdOx8A
eIQJlbrYRYw+vr+nTv8g68MZK6pXE3lnHFf9neGMtFUT0q2tGXoHUUH7eli3qcSe
klHEvDJ4BDrge6mKP5S9SuoFp6+McxE3q4LwI9YtybLatskhDKl91X7uqkSXfOdo
IYfaNHAy7xu5K2k4JALvaGP0c0Hp+IiKQpdWJnnySmyZOa6toXfWakyn7wFyWMci
MeSSKiA9+hAmy1fzYQr9Oh2Mpn13yh9DbiMN352qAC0Qy0CKPYP8sIJG3F8zOoWP
SjXBPPPEctJSeZcx5yRuWUq2MvJLJkjaIZ4Lkk3cpryp5Uwj5Iz1lut0Ap38Tt3l
WORm6pOU8j710bcv3BLtwPAVpzXe7CbOnOY+4mKdXKmSeH9Etv9BSjFlE2Odjolw
cbceVupuoQ14eKgwJ4VTIHIAt8Xtbpww/ayHY1zGRkYxhItJIk/4HOA0S/0rhEoV
qx9C4nb0e2m/7Rbq4XE7X0zeQnn+TqBwyORU7wVaOIYfxTexYmHtD3/+r+UrbZ9m
6z0wsjp4MuhT9hcq5UtwhZkkIhewNzc4zMyZaSzJ07R/AXaQcJ+OOzLpaqpB/pXc
HYV14UT26c7tjCDAXOB3yJCrR0BxpMYURb/voYYBxnm/u05QSrXI7cItRZ2w70R5
Yc4H/cOMVw/H+uKKAd3EdA58d+mhH1pdDMWFlBq6c22cUrBX5wxiVzn2CVXrMJzw
yF/0TJsDRd74a17TKfd/yX/Z5OQI4meSKOnoPPJEMrwRCjTx/Oud/6vyzhTbjJe3
Yx4eRNYuu6iBYmwFUnxETdOPrHvegngKHbn7ESQbH4AHcLEKHGmu7cIV0Fpxb1TR
Oqw92GdtX5XbP7ufcQJimOd0FRrLEwSRt0OtF/yaLYNGMXZIPr8wSdOtduSt5T7R
QukrAB7iquZyKlEsddvo27E0CegMfCxuTrr8srSNA4Ui8xCQxDmv9WBOHWr1zawP
6k18nVZYXqGzXdpn7JkCMbHCo+M12UIwlntPE4KJ5fm6H4OriYyRGzMk5Wcgzvri
t1aGfuEB0XtmVwzBK4n3lS9CPWj5HRAIl/wp7nJLLJrF6YKIoxsqgEdQrHwDNseM
5wtCPwxrH2hGvkD/RW3/r2DtiLbWC34MNn+OiyhmIF0bzm2Wi0uMVEf5zjVhBtiz
W8vA8Imk6H7d9Hciu3P+9czF87JgAAWSpCnc7+83HeNnNcx2QcLbdvVO4rY117rg
PU6n7lLeMV8F14qKQkFfDcwrg9/FwkgDOE2V5JBqrn0msCrXEXmNRq6BKgWJBof2
V2lVaAhznu6Q8xk2fXLRKOzkLfOxGo9saGCg+O9nIizZMiW+H1mAfG3M7wT9W59c
EJBZAKQl63PwaJZIQpaoU5WO3FshPZLNJ9Z5MQt3etFOaWLyH5+cunwX55TuN0SV
hSu5G/0CjgHuveRt0dc7Vg6t8uyzZIZh2M96FAMrURA+8ZEM5Bm6y02G+tRZJ3Uq
+Tr4UYlUhkVQVZg/8NIR39GWe9fYWqVTzOHCrj3j51YFS8MrKblo0KuGst1BHUTM
OVDw2wGAv8I+PYeeYddXpAOMm3CGolWzA+CAueTAKSDcWDUFhYqyRtJETLKJlHlS
l48eXq6raW9qQqAfw+M8N5U+kQ6sppUIb2vUEHm/ALmiRF2IPjiQ2cVTXHl8hf6j
W21D2t/OOlUJsalgxm5pwVigaF3TjAAZo0RHjCb6bNmJnUmtYM1j1Yx/m1HkTNTe
MS6yID/dt76FCmJ515yQN9IaJFdDsAScUiwo89oKq44JOWZLTlFlRQuAunUWjM6l
3OhR7NwT4bYTwcuFafGQOOZ2vuC7PiJm3DDh8HSEPjaDXSu6YDWgaucW5/026r/u
iYDV7Jn4v2vNAYfNB00T4I5lYSEQkHuqYH3wCmkMIeJ98DCGFi9i0itHGZissy9s
OuHgXYtFJwqgkgdiD/ssClpAgLItM97qt16r/dXvOBJYQnyiEH81urPTFaYOKFtT
e/FxOo/9KFTHsAMMU2jb7Yqa7CVV3vz1Wk5Cu70lVDKxAJp0nsJ96m2cMNI3mrvM
me5ASojrMBjs2upitXgql5vz8yn67nETt83ofEbYiL+McmEj5CgyqfDPIvSnwZns
EqltdpHsQ0tkuzLiIOEFZUa0eD2eInHhqeX79IM2srSzuHLvYJituSneow2VUjJj
/B6lu74D385KTfG50H6HgGIbgMIcWYE9AeiZPQoNLDC94vSS2rk4E0fzXVZtOOAo
sCGcQBDSSf14tljjExBDPgNH2G7Rl1OnoZ8UPkaiwYG6trIBejhZiYqTgW91wrn4
+9fAQY6R4rFB+tGdThtC0/xlWOETxvpbWGSc8WznelKGfFtk9FCuD96TchoIM31F
S0kWTSiirS7fH33LaAtTNpt/MJsBzHOHHnZl2LYjFLp149hPADRGmGbbHkRM+MNl
ecLdNpLNErjtBAPLGlYr4ML0/X2MDKiOt8lakNA+cH9Vyvyk09PlCgqDxlGjbgtZ
qZiFeQFVeKf6t9AupeQrqf0UYqofc28zNGn4Gr1UnFBFpPDZekIPPLIYd2d47LvW
EZraN84L3TyaUKF2ray2brhGKn//s6TsjFkSRAohF02ZEvpc5dYzmePn40aEgstH
I5f3m5eVVzznN69oXAihCxbkxkFzPq4Z5fCyU5JdKTVTIKB3KWvvWlSpw+kVrIiL
yZ92RIMg64dtUSgxLxokqHXct+Nh9TfvLGUOBeiZcy0iiIMLesWrkl4ycuZc4675
E+Dy48jiXhfHblSy5ukilmpRyvB4rEAtc1aagUQf8vKoGAixT88IRyFytljIEMKN
D4RRo6nAQHkcLSwNgsxWsqi15XkKZmEhVShQg92e9XcmRcVYS1DehZwz36SDnCty
HGQdrdcZMQF08arx415dLtGK8P6iZ40zNuJaFHKBQbY1Fzn6cM1U4jvAZzvn2BvF
3wZ+5ATWiBX1tO8dUOMNHT77SLj6T6JC7Cd6eLCtFHqGmrmD+noVXiBWjtn1aapw
c5YyfLcbsvtTmj8SGSpiT3FVfYV0l9DlRsI2D3Vsy2p68NFVMbx1zY5pSP3AyeJh
jg9dSYZaocxl1T9DUkuAAHIlH9P5JJBDCU7p+nXDVqPPXdOfEzfWsZoLPkPQFTzj
qANHlsYStAN6oCdbPsxNeFienH00vv6ocdwtQ3vf3G+jkAzTJz2XDbJc3pX9hXm2
rxGemFtRxc42pZAlR+A2VM85VXAvNScG7IctMeFBinz8ywdLHeDgtLdeXg5P059m
RUbNsoNGQJE6T8dR8Jvi9y16fyTzXh4FFSJ4ycwk/Je3G3jlm/v/n5g+zIz3zaJj
1nfZ9EYBYoMRbkzSO4HAftF5qS4WUVB/EnXiupL93cpsxZCz+yhkC/yJSNtr4rVw
/2n5iWjtJo2SHRXSq4criBDVY2zvHOKqdT/kH8YZYm7ERtfF08PmKOxKZvgN5Tw5
HHQQU8iwkghmM1kJK+ID/dnRrhN8VU7tegH7FYTNQtdq3ZXLg+0J0fo0KJ7TmXKL
zdUixEtOZm1P9X3ryP1y7wpTo4NkvzhIwPZeMGbegyydyi7HV7P+2gMnj4K95ddB
qxKZHvqzj+ua9jNxxJEGpm5+Xoey2BaL2T1y9mcUbGP79Dp55JV4/p7KYiItK90i
MRfAHr4a8bN2tpaPy08APKmTofq7qyrlgXPpK5Np6Rin9u190da/VSl5BuG4kBQc
Xbh6M/9JMwnAnJtNmdw1vRArZUGbLfqs7DmZK7VNpSWhgISHB+36dlpeYJqMvy1b
pMB7vsXseQbOD0XUiSdEgwhrSKEAESeJ0AaoC8WZf9GWFCgrmfbsoXC8RZ6xGbGB
3xaNsx6deL1udeuhxY4sVKD279XqNq28Q8Pp7B+A9vhPYlgaEaVvwor9EeJxjpoU
LFXhFkl6Jhnwz1uVeGDkGMTWPbR+6I5BM2KlAClf4iI6VdGXVFPlH3wpfsINWd71
7SDfqaadVYe+h86y7N4MIcFvRv54T+5hyibHDxg3a9aRJEHtsiuH21Mk9JmRxwLC
FmPQxmosC/DtMQTVtA1aRfWy1Esdy63sOzAw9Goz/R7DP1r1oQEvTRVNLOXbLO3D
sqPcwCpk4bKSjHSxW2QWjjDc7mPcvaMmkFKKZdPHhgl+Z18bBYR7cHgWWHQSzxti
eUe+H2Axi/y5FFQvgx3h3kLWUBUU2wgtl3+wr0Ibtotp9y9b5ZhGdXbTrZ0k6qNo
+CZKma3x0wfcCZx5mXc0i4gJ/Xl6dMDFByb3pOd83tkussrBnCGjt7k6KN2kyLIV
qWn8M6dDP0+dEQpR4n1VnaVKuqnGSz+TaBmBQ0UQbmAjUHYNe2v0KaTrd5Vy5Ks9
Q/3AeJHRMobfkWu9iRuyYvps/OnjlKs2TxUbPOGqLPgvaAeSlXXXyv4KDJeqke8t
sYZIfuy2XCB4/92JOCcmvH8BhSA1gwgHv6uuk38mVASfFC3Ppb3CtWw7FgnNShC3
JALAuRfX6/Xwh5x/K1StCg+Qh1nUW8RyKwxPYI46P5xxfm6RbfZ05vOF3oAd99nF
JCZFN6XXeFOJQOXj8C5FTqMitiQluosYGUtcGVelRvGHaBHO25Hm3SFy/1j7mxuZ
wgUCWYGJyUK/PuGDEiFx613oYhHmaK2XxaJv/9JcGWuTpZblL8k2wl7E0GbQ4pVu
nApw9+HS1fl2y9nu6rxdoqXnC21nq6/zRWnYQ+wMJ8NvCyjt2hoVn9i6HlpJhWBD
jDD/BbfSfCL/rlILN69isgb/HL3sqhn5yVl1Jx0n/d2eCr2qNSz6M6smshQ4Nh2c
WA4hrEqwcWrrNiUOIcsSXLiy8M7oNuSgiDiZbmlf+Zx0x+tl4glFaU1mXESNMFcl
ccE9EDY9lwsoowqYMgwuskvuvO/kxr2T8iD2+M12Q+0rS+l2uz99P+SgdY/d7Jvg
u2gEpmx7M2XzL6cSJNFR/cVLfHzbbI3cxJ+RdtEpY4pYczr5guXZVkp6RlizC3GI
PtmZVc5k8nfpJqOIcN6CyJYx5IFkYB0hlb3UXVnEam+Rpos/amNDPuh+Hl1a8G1d
OCEBySH4pBPwkV0l0bNQNI9WdvYsaOa+xP8+4Tsqek2aGilMArI+ZQQrSojVzZ+F
rI1VTeQQxRpbC3OcpxdbN/zW7l1uRDsWHd6+OHGeUJECrQmoE3zyhbhrruHpTPpm
QF0qKlgczEgsk4oAAL8ICY5h61tsw4d2cVj2wiV02lO06tSbfbijAwjjqnFThAUC
V1k/shq8I1Xpi2p2B4hpENWS845rAMpYlt+ofhD4NvpqmEe8BRVwden5WqRBDJVu
GUAbNEWNUdxAdL5KXF6zgHWSQhtFzR4djvaJOuDPKag4kX2jx4CkiQ3p0RpCNohI
w7I6YZf0wnCHb9giHZY+jBakephjUR/kPaBpPj2jBqR4A9P1j7y3nzgU3RaH4DNN
DYi8zTkCwtKSl5ee80sfC7l05JCOkH8HvevQbK6oE+7fNNrYM/vcABAh6NRtRGIP
VGf7dfHJ8NeCTOa/Q8BCskxXvs7B6TA0xzDLH6Bq7rzkvaUcrp+UOoX8PKoOlvYR
Taaks3mfieZu99cRa6fxCqmdpInbBD75Jab2tgf0Iyw1CzCuhkm9h6h/m54oKYPx
XbnieSNn/ezvi+zbx83pMrMh7gmsU21I3OAU48JRKEYpuFQw4Ds+wCf+fVyPV3si
RseEKVyf/EQ6nWD+S/34rCvL6oFAR8GG1YrCVKY8kQ/TIkKqjI53jqDH78871NAk
S3QsqiIoyBHTrR7QEu9Jy7aSXFBHVrDpN3BgYucEag9i/sk5pgIXaky8OM9FDkqA
K1V2biv7ZTYGnP2y+hQtpMp0wNmycUr2o7R/rrPvYCllnRyK959g/HkNVItZep8w
bIJyFgzRlJfOnMXUfduJUEyuXrSx8m7HTHlzpoAAfIuGR3Za4/Eae00UBG3WWvTv
49uQnf/NRqBqz5EZqwPp+lLY6lOnr1ezIrwzWYsLNMMHUZcS2Hi9qsYLlaLtL751
ykRUE0DOLakhBlJXnboQsd2bRnPOPOiQ1+9xhZPHDDhgx1faaEkBam8Hh5PLVYTP
5oHWgox3aYtefTht+iWCK2vESHna4WULriCAlqZtE5Ix7Fup6EKV6Zg+vUgu7h/T
rHRGHL/EgMetJizMf6ndfAx6K+/E+ZI2k9lA81Rld4Ko3I/08WYGb/Y8cH6KWh99
uJZyKfod5zFZS0+frbWEK88yOKnbCWjLfuzq2X4EMO1DVu6xTmOd/UrYghKP+rDT
x8ZeaFxnw1b7x7ODS1QITVXD1Kas6Dl0uho53uNt54kS9BEpeq5ega3OpUhAy/16
0udIQn73G0t1nLwkS07H9eyb+gvuEV/Gd/H3vnpC1DldurTFNfigeHiaWoaT3gJR
RaFFZ2qddZ4ydravIoIVVHi8cmY2J29IQOgdfcbn6KOzOeBClAI3u4HgpSjcBSTb
ifZFpBD/nR/fUAx+/nzF2gX8m1eSPjShAveEaBKzDlPNVCeVIvmvTap+tHuqcH7l
qylnW5MGIu/EmQiUEFiucLCradYEhMVknMSOMbuOi1wKrwbwslQ50j155CVvAIJ4
MrWRREbHWyfkJgVUsTpd4i5j0/ehaKqU6pbdbRZRX8zI7Fc/sWFObNVMALPAeWMz
IvefV3E7eJt1zmukFbO9wR2uBi1TiY+XIBLvjaRXAfeBLuQmKHbxx8UmJw0svdN6
qDNdoIspVVPHK9oyct3unNlBxXPNGqrT0NbaPiuK0YxVQ1SUZqg1Pq6XfsEKLeIh
ePPsMaC1lPptWEnFRTbm99R0N+wRMb/R9E6u55ALCb7Y/hwdcneTZxWdRIr4f077
+OCI/g56NMd+wrn4DCBwDqCwA5Ro+MdwvyWtM2DPj+uwTIU+lxIdadUj2YAopy94
NEo7kbMwAKcy62qOBH/YtxxM0LwyMsiV5EmPKhO95zRT1QXDqEvScz2KBKfEcHa3
WCVjznB4Tp+bWgJfRadQvE8+oh3CseU1ZqtHdtBumYrDb9odSKnqqNjwEieyfdBp
iXVlpTxFjx7sS0z2NVHA1T3atcuAJU5Isscls0bM1+MWHbQVcFZxFmHe80qJ28QA
qFIop60L+ruNr8yGmZ3nSV2XiADzBKT2/CtMRlFkdP4Ewu2dZCvx9jnYzuuXIYWF
QBadxkefKzWKPsT19AWdvTtDtTxY9acEB1wukMZUpoRBiP4Xtr2fzOHyEk3y2QBx
j604MXxDYlDI7S6i/cf5jDYjb/n6l7cywwgx8iqZ0255xKBKw4xi9puV1mXYzFxK
QrOQ7mHP6kpk6aGOVXKvCsHHjHOQClVqY0nQPWKA9+LEm7lhmuBTNkb8mjtfMEgj
N24fK1B3SNvEPIZzzccVciqRO2mMdMTf4FDXjZTNO0U4BvtfHXqFjH/wWk6KjGg8
wKy5/Qd4WdSPTK3PKSXDn1tSi9Dj/381MmIwjZYA3ksGQ5YBvAhWYJj9GWOgUjfu
p/3crUTy4SEIuDdLbGXgckonlhkP0u5wDZGtSuJnIaj8qExzF4Hg0SjSkeR3d/b2
W4cq0mjxHCbdwy6S9WKmA4GVHN4xFUvtjMHngF8gC0jpgPkD0oZsS1Plz+iFzuQJ
I0PPFz+8HRinwDhOa4KAjPSUrDXncumlQHalePrmnAGHmGnZPzoMi991Xtc5XvJi
35T4PdwEJSnxi4CE/t76BAl4atYxUspuykj60M5dSfxIzkm+OBdEi26kT2NBs617
rn+6bEPK9CXrD2SxAe5SeCpQcPWganpEIcdLnF43jUuKGxZ0PnDO/lLhEJsOAdBj
rXdqrBYl1k1R4IlKBwskfFrXnRii64qnnTf4RYRQNH86KEvrMz76zF8oVAad21Rs
juhAfmGOxIqlzYcavTShLa2g3n93TzSjTS5kvWtvRZXJL+NfI7ybXZYuDrw46Yfc
NnxVPYgp674CSntEBANOEZjHZw8llaGIdD0VNVJtiOSg+318nFQOyQf9N7iz+bHh
KosKFGmYbUgzHstwKPtDcxTP5RpsETvR/AMTemDWsqdyfCqCNzldcWF/cACn+paD
3PDX4FoV6H9v7PQtePce/eqghqTVfZtGrVEngBVCAGk6+fgcYPimPMxU7yPMb8GO
BvDbnRgRg3QT6IlSL68QVeWWg9acZRJiGkrzUZQz/s5u9JF7Fb9Y8vw1y5XMFoZG
oqZ5jDv70q30cXI/mK9KFI+xw8fcuPxG8PRkwPY9UInnL/qWTlJXmlMJXWXFQq5/
ifUtlGnOUw1q1nBOqPnk0WeJ4ZfzGnQZKVw9/rGrCiroeZuf0EhL8hinplq1KBAu
xw7WOBsJaKnuX1tHx09QVD5e6RvzznjTUhYXV7a1FHyaYQ89Z/39D13GEurG/DoU
QUWAMz8XpuQQdZ2JsHEUbdTm44fVQBJCFzTZz+2nh10DooUMvsTGoqTDzQ75/QoZ
y334lNWQiMee6jslV0up8nwlMFsCAFxfFgVUASRKVJCSrQ642R12XFEArcwUpUk7
et6uzmBrXvGMS2pu87KkXFOz3tDAPyUcS8I5RGxYaWcTfSNCeEEcHmtkYZNZCbGE
s0lJ0rQ4WtXrNrZpYaeqD1sZWZReNqWWKY9Can8HUZvP8FoZEJpzOMAl/pOwWcSP
uCWec8+c1r7fkIscziWrtnxNMrnWVrPo/NQKjjiAoZCPDo/0Dk5QHiUqZ257ybDL
1vhuecsN2Dpc22mF1clBZ8uTJ6Tme7k5RD1foNE93Rh2O1QvObfhuUO/v1M0gT4z
8HUPFCwYBP/MQGqBiJWZdZOM7vWmTKlmM4ByOZrjYyZCrCB2r9/zyKp/19uz9kon
nR5uo3fVsze++g9VoWFV26X/V542w3EYxOlCyyorJUQxwsyqXAgKOfo8p0PWNpCk
MNybU2Pf3Z9kHQlQpyuArdVEP22tQ0YWayzDs+dIS2Fo6w/93IYOlL1i/MI9GxII
ht8wCelLFiBuPFfTlGoIGSkHGa/o+yCSXYvwRcEn1kwYdrBYFpNCvQl3+7qcMuBO
+2RFlYULlSDKmTrKy6x/C6fFxHwVY+yxAtBPqSgBGwrdEvWHVgpKiCO58Z1Yjwot
m28RnMgnfY9aEXufc9D/qRWsH/A+WoVbEF8bg/kxOOkUftrwaBcEbk0gnzJnb9pp
536O7TK8YtrI2l1rr+lQaoMraa7z3LJR7VE1RU0cuogBmwB4u75r7+CyKLXuTRSY
XjkIF3/PsGWVKLb+lyJXaAuJA/63VbKuZODR0hvRDFqHu5QJ1WkbT6QWm1NeD2W7
kdpHkaGGcrUBQIfRG/aQ9+yeoWrS4T5z6UicnLDUYYKyiMxUvalfSg2JPe8pHdqH
CJe2KPsJDLWv713Ol1kRF0Sbx7lA57NqlwJrxq4BAvRhW5QQBSqXAQbTpoy3XnjE
2X0BL9w9xCmgMGhRj+BovmRAJdLplGvijLQeCqvm2d9GDFYjM31QV7Rm37A101rL
tPLDA4+L6d9fGX6SSy+JKJMLCBWThptZGM97MB55qpxXn7XjbELTK75Dpd2Ybn01
Fpoe0VupXColqckD9NcR71+2Joywiy9pllNIXPgsU+H4xDrWG1FfThv4GqT/gE2T
7onvGDw7b8DM2pNXiG2jcnMMrbdhZkgVDVbDx/GzzoTGwwe2KpEnjepeX1Uf9Mes
ZD37o6+yK2wJa7p6j9msTdfBfQyz62jzQTz9qjybQYPNflARyfQAzQafIUzEJ70B
EroEHNRnjTiLvVJaXffNQF/7rIIzkLiSs3ojWBeEFZPiAqvrcD6EgUzRbP7nwOXk
DxqpF/t7IicXwhY1Kv0hnr/cUlZaCgxyhlGe5gNu5dZpok8zIxEv6Dk0844rq90O
P1q2Uj7HrqrNki3JIcShbcqYbmIH0+3xfpZYvn+Y9/o2fMgWsL/h/CMVgKXGNJUd
Wdj5N3rOtYIwVvO0tr87mkicgoP4j4+UyAZ/mm11gZ26w+8qdo6j5Ud8IT27O7xt
awlWJTSqlyzHG49Wj/PIupTivO1Nk4bTuP15m6AJVmpceQstgMIshr95+wJVJjSx
yCPLEInpmDrvOJO+EhKB5kydIU7uvrtVboaggGcdzsZdahOgxKoWWsI/9GqEihEZ
+ZCcN7PNpET1a/vAhYDSnbs2jqZ+a/Ra723jxQRwse1IQhKQau7ABL3aP5Z5uTZD
LCpNs3vLlPbU0xMGO1UfiJ7drsVzoMlJfc+m/ZG6BxMhT9zJgD9N2kg4Dqy7Cy43
Lnij4TzdsVDVClCrYbwBi5AkIQZcBu4RBLLpxRyMHqyfHtIuIorEayFvBekjZC3G
ZrR2n/UaouM0/dRJALXpP6n03ZBPfHre148niovubh6SegiE1nbY315BfOJEkaAC
IfOmBiAOHcaHY/uuvjZAEIlxahcR357XpnPqmw9aVFKCWF83x4no38c/f7ddNkxe
c5gefbgIMkMYuoEhIjbgr0IKr/528rKHz5WesRlfdw8+VFdxECZHAZ94CqToPgxb
moBWk+MLhIHVeVVTzshB/JQV1CvbpUL7Flc1P6/JluNL5O2kRSdVMKoe3mqJCHJc
cg9z9yldSP55xhclxXs9bcPdFMUXmwJ6Xy0g4ll9VPXnT3zMj7/e2sR4fUfR4wFA
8pwKiPHkQJGRc5w2fGu4nBK6x+/PoWWgBjo2JBtz9T/1aMb4ySHhLsPNpIt2PBZS
CxiBZ4sqHsEMXbd0c1hLppz/LDQh121IxWQeI8abk0wMKmYXucbiGUlV/WSFA88L
yJxibGSOcwcaQVAiot0cKcP2FIv4/D7Ix7IAALAlGkdnkjIpphCf5AHmvx/UnH06
SqaNibNjY481I1KhmE8KDpYMFeSZA+UlVdzqnZPChK17n9dVfqgpKXevRNiUvYXf
dm7x+NWnzhZibYrl/29g2DyQAte7LLiK3Pua3DmVOvO3GajS0qTzDJn5t/UPiZMs
`pragma protect end_protected
