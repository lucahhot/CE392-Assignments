// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8BcKMuBSYfF76JleiQh4t+VwD6UcbsVISLb1hukiM45CcrvRCAg720v9XqikIC7N
vZF28k4KxHeEoaEm/ma+EgIk0eX5V3jiPhw79+3tWaX5rOXFSB/LLcttpVuJZ9hj
+ghyHz6fBKIloGG2NWYPMKu4zfofxes52rFzMMgWoX8SvxwGUpNkQQ==
//pragma protect end_key_block
//pragma protect digest_block
tkcdwGZ7EpU6+Unybvf8MVzmzc0=
//pragma protect end_digest_block
//pragma protect data_block
784NL5kFpJzYTofMypOs4Rc79SD3/Vvugo8LK8cBnZi1dB90edoUJGkr6rBpnnG7
3phoVG3ezF6quP2U0CGDrYEz/0a15mDB6pE5aojFwqB2gcjkCsY6hKTuKlPsnKyZ
mQLtT43y+5NK6wMVgY21y7Sw6JmYQzRLl8dB4WKSr8Dh5HSxrBJK6Bz8GwHJL42O
nSu9Kp1JrpQnL+xYUr8pfvAA6A/FZLeT31hd5S7rvKxq/lvaAlis8fEE2MMLopqY
yowAV9oq5lruwZcoHczJj+joq3Kja373tzTK4PYbXSdYS+uZJwwzpexYdy5gSNwj
aNA2+FFjd6Bc+tw7TUxrjvDGV8ZAvzfyqrUJ3kuD3djHP7rrCO4hbxUQkSaN6XGX
xf6zFA+o+2X61aUo6fLyKq/gGTzQ5hvAXNFUG/FHxh5KgPP+x0mr4KBMKfhpGNog
URszOcFtPfxSNenYX86SVfhwHm/OWfnjz1SYtdwauQffgHzCYvXwQCExfoEpkFv9
FFCqTczbcU6lK1UKB3EucTyxMaxS9LolkLlc2VsvX8otXalGWpgB99gLVYh7Tx5S
0N3Ry2wuNbXg/X6j7o0V5iywgZgk86UtSEq5C10umJzZN/I0hbQzLa6TD7ShZ+ah
qNFNVf9nonqCZfc+YNj4F3wW9SYv/zeQ2YFxaR77SizwXkINlotnQsOxOzEbk3K4
7vnVrBJrhfc3HLl+o8wsXypohV0QjfHFfp525hHyeroJJx1H0tTkrLAV2msVHW1h
CpG9dLXePU49w1fUej0J+iDP2zWqUN7/kAsG/AMzb8f4TXU/iQQXuojjEfWpJb/w
KZP3peoIk8yHLtabeelzbw+zc4clJ8IjG7iQMd7bH8LHL5t+csRMUsEx1xkJCJRT
cCLNVyxtehWKom2AYsQDeEwLDUl35p19XykMGu5FVaPQw8/Ii99ydJ1Uk6+yDI0s
W4nCJv0cwgGt7okp1rWKELU6YsQzjvXgYoCYCVDy4yG+xksE+k8pVg2VQODF2kj6
uFZeG1stqQL08Ac07jmnOXSEmup0QX0BnBYtd1Xi5j3q2Q0G8morGG4rR1BXj87w
bZOowUxQy9nuUT9fz9OGU2ZYe9OcnU6lVV7gF0F05lVbYZAB2NMEAhKW97vTI/21
drvTaAmEINMbGoH/X3uXgwjkuAuYzHk01T0na1rb2NW+i6E4XiJWDfGiZ7DUbYBS
zW5+DEnnuxP6Zw0VoZBN8/0hWNocd3FUFGvQmlf22dPhM+RbyNEJCxSQP5m43CWC
98UAm10f4/N4hFl1LESI+f6sUmnZ8AliqYMFwRPgX6y78f4aRAdv39ULtGth+T1L
hmC2vzNfuHnYqFua3cokFrra7o3adlOLwDButkA/6E78IBYUXZHLrZPAx7HvxfCT
qjJphjHAKy04zJw28sgzr1aOI427lCg7Aip9/fHhcZhYMxTckfpzZ9UExqLr9T+t
oTMOjrIBZzm4ER1buEL9nxnvjAMy5AgN68e6SRwDB9BSN4/ZzqMFCr/uvNQqFBCg
h0f9/ZUVDbGkrSJDroy6PTlJ81OXH9l75qY5neepsYDW/6/CrHkgxaeJT186wsSF
JLNIw/+9wNvb1uY7HdOb/Gzl+3c4hB19Lxse2V413zbybrP9c3eypSZMTOcGDkkU
UIZ8z1VVRReG6d5G5MBln/sYbPZ07HOzIbfoh79UvhvQUeo1SrdDUVluN/wyAjTF
uVmP5okBrW8Azr30FpnqK30hugpSus0y/t8Bl9qTYBz62cnVTdz2zfLB/H/h5SYo
CPLXZmZOL0MLmClfaqWnmV1JLgVh9za5DjWojRa5qdbXyZdiAweKk3tsnB89pk7q
6jjPqhqe1qSJcGMQOj/bG5/a3Sr7Ie+WDvQfFdCQ7oXfWTNDOJ4uPIlgidH+GJYP
yxW1gtvB8tH6t4ZO3cyHRzg9x9wHcUAB+KII78Xpcyg00vp/zD4KA3sociMN1d/1
r+lZHxS2/qGXYnEXibEJexMSJzkzFdaWdxuPABzdaMihy2Y8hw3ub/ewYr0h/YhP
eldzzMJQUkMx/Mbg0I1qboyd9+/tdt2kyL3eLI06gEm9oIYFTBQAUXijnGWiVj13
pz/dyEtNvXfCQx9fNvcqyWw0/4mVN76ikBTIfyVSDh14SKARDf3ngaN8hGC4U0gp
9X1FcSou8NtSsLrmSOkGnAFiCygkih6qH4QXNXyl/aVW2QGWORu3jRja8iDPTV9J
yZkXBPoWbQ+/nOmpr2RTzRXqEryKrY7jMJx4TtXLYR+gp++sQLPow+XhKElOh0wz
120NMhlO6ABL9SXY6P9Cy1uh3qQOtzlpYZ5XVEMeDzavYd7YC9AUs/KefI6YtjiZ
Yi2kOAkJ0Zkz9K0SqQH1VdQATDstk4QS+u9hLi9i6UppqD6cbmmWzdctCSXYwKH3
Jin/qoF7J6Gtepy4WUECMCGfpoC/DXr9Zwofsg9SEwAKsWlSQVVUQb2x6RnYcjbN
7tCrk022Y6b8g2/PZefz4QftkPilWlDJTylrZq+kj0EKzYpYveWxjHzsiXdNKyk5
0lhdh4hQAc9S2Wcw5zTWrpeIO7JP8Mct9jWiD76IhexfOXO6DezJfUsxZKim+c8K
P+EY/O3stXluzD5yb+UqFHsdJVaXB/pux5Gjmw9XuTR1vRsQmL6i5LmHPbwB+4L6
we8+ruIUGpo9Nehw9XW9ITCxRAkqsWjza1K9k4oWE5tvIjtD6pOxIpTmNKM574On
izLSML8tvFy7kEzOeIj1FrfjU6Z0U1Wjr1siC/R3lyeoAA4wlXViKNvxpSInTfgN
uqTX3iVwDIjOdPqN2MiZu8tfcOOCJoZtQdZivAANAl71zf1fmYhwikzIGfiuBQ1S
Y4Fo3WvjVP9bD/GoU2ma7+6HEdx2OmBgUQLf3ucKB6tTEDzxveVgmxc1eWkJVqKF
9OKcx64PVvATFD9U8CyAXxzlp7rkaB4xSffBxZQAeJxqBBa16vCVRiFJOiJqeqZl
vFKsgi3FziJweLvC+6UUJHHyZpaq82wNgPFpe+STdIrX4xBnISDI1RDmZbKhMVZP
4mBXkuHKu+MKULmJivi98BKTWB9kqL9jLl8JspWpKK8c9Xvma42ZLxUx9sXeCw6n
QEpOqs8rx7N5JHP2Du42AiIsAxk/wrt28tMM3gKjC1p1K/enEMdpzGdeB3WxoMbz
QpkWVGZHRb8BH64Y7zYs9F//+9fP4ocw7wrQQu2i6cMzgqYjPQi75WELAwmkS3Ar
4cYI6gcelgfR+K/HMqgui+7iKUeUYb2IyStny65XL1vC7lIjXLyCY4Y4sHIQHkt5
3xqMJ1AAgisebVr6vYFgoDZSm4nRBvj/UPB7sQff12DLesAuKdS1fH4e7ViNQbdw
rN2JbUWzPYmLcQeFHmO46uRTzphy7U6Z9Fm8jDFkEbIptbktJy/A93BA2pSOzNJZ
ZA9HCICyc/t4smmAH0sAEUEde/jLikhwaP8P6W4N23cX1N9ZC5KpC7nxxvVwOtwa
ZgHhy/frGCXP8vUPwmML0x389nkFA6X26tm0//ANsND0rwFJwW2QouxIw4F9IOU9
Xm91Ek9zuvoth5M4gGMFEosBbqF++axP1HOO8d0FOOwp60eoen0IKo0sPTIIWnou
Jz5BVh6+zxA5GzDOO4U0h+BGaBm3Ei5CcvVdngcmsFHdZKeCEYOBTiRvfMOC8pm3
LsPNwkWcbX/3aZU91+Py8sUwmH4T8xfYZPOUo1v9j44c4nxMkP3W6DOPCxEFRWO2
mPdywU37btqxSJoQ+atEScQ3h/mHnZd147Xp7Tdlf+pVsNtNGWvpc0iLlKQx8pYU
WUMl77NIBIHO6Cu6HpvsYklW0HyVpFO7NAkWXsW9rcH4UaIN6AxPlkrYrWu4TAQQ
pdLXuBaRlmw8p+Z98+ghMSvM1PE9yAHuRzm0shB+aHJAOwpi+YXcrZ0NVMY+mTcU
ROr0+aJ2zGgU0IhpxRNBcumbDbldWmJ40aty4NS7rgIT9xs6+0n3HClnHUoEx9BJ
kd0fNXggA5O6RSqSpnFtrFJJ43rfSehFJzqwEI4UvJfs8LM4cUrcFBzNg2ncFnP5
U2OQ5aIOAGcqz34LwzqMwX4eSsqfvmQPmgtYSxqb3Pk+faI2T+DkKlA67owmZ/dO
1g5ikhZJDM2mb01sarQZ4ANbfT8+/iu122JJPbhZVO+bCfMXYD0GoAmmth/KMiy5
fVOrnmVzk6cXVPG2Vw1fsvboUUV0FrGG/5Ji6rcopyR64HTUfZY5LGreC7KJfu2N
qzNIbAKGUtRSBJONjQEkDH/0xB0kIY6fUZvDywSBy/kEGmXCMFBllcmcCeT/MqBH
T7AMRrYVcPympP9cHGREOyAvD+1Jd+WeDvKEq0+N1hzrxs8GXDE+zCDGMu/CHsj4
DD5PcyXJasJLUNZknuTkj6UfksILD3VUq3kfXXEYhJMwfGFdUv1SfFPT/ar8O0Bj
pRO4B4QjDBe0nzwY7DhXHvqPn5V/svMMabcFp4rkrLdACtCkTgEwvaPgcrc6qDHi
crWFl8r5T/uxF8APOfTnSJ8XJTEd88L9mQv8M2XklZeolbPIMn166tFXlYo1tyBG
oqjV1tPSHUlvxEUPP1EMaMcU3WuQmZZ6FEM/X6XXMr2Siy/kXjpysgH+25v6bdgv
J8gQIa5gVjqhfkc+jNkcAZ1VfQmtz/VQEMQVc4PPp60ch3F+Uc0v7EtVoi2wDnNd
FwMohwPINt4/wth81xxNWTMfdT5h1iZz5TnthIrjhze5/91Lfj08SzztGev4jqJK
1nzZsYROM4DyOaLfHvvWCW1aaZDCefPyezwSMhwrG08TT2HJDJ9Jc1OjG1eWay+i
N0nXzGIp9Rq0NQciH08oeClBTAHvvS89a5GjNY6mTL9epihjPWXt9APgeIoR5NUV
7q1J2O2tYSVDGtimWsk8BUgfA1UPoxesjDVETl/8lyPMUn5eBRQDDo5YJ+WWtFwN
X3DOgBsl37cobE1hhZ3MO/ieAeP+ZYl1JyYFk9M3LOXKh7SjH9eqfsMJXSQZ+cH3
ouOzgLLQ+cZMFLL7ARLmjmhzAVscpFnByNI5fAtIzhT2TVwFGYsO31hb8o1QKY9I
C3FIlUMjOAOKcQRfSADeQTttRiIJt1u2GIESfiiAbwRNcA8RqsS+GbmuZ3k7om0E
/DeGWKK8RFuvRCcVP++8QBHRzl5EjakQvz2S/f1Nv3yOnNzuti8UTVRUTCs74Z5P
b8kHuOy7ysk3eDEvVlNf7xVtTYqa4VgQDPt1JookzD+BSZH3BLSgLI6nTZ3UR+4a
cS4uUgJaFlQaUPVCrv/J+zZjbpiRAle3a7nvdBciW9YTYnph4041EMOrwkREs0+Z
PNdTy74sYZwztYUovXJGDPp99yVASMi7ASb6vs354tSlMrC1azzdVhGpaFJZ+W8+
Cbp4e8qgQibGwRCy2v5EdVRxeVAl+vhyf5WjWOHNyHdbkF4BXOy+A5ZF1Ztyahnv
0ZGA0YxHn2tg818xv6G6oa2mYDREUA0W3ZmEEtIYozGvNlUjqnftCjwtdgrp04uG
Y7Tmxr91eUimRDcrffm8puCp0NFykMZ0QAQ4mn76Uv7JS8tefYgKr57nAi5g24V9
6bKFqkmIz3NUX6ySBucpMpdPx8wULXjO+t5UmX5LENhLC/S2ofDRSpjtHi1ehe85
/FIHpevd01pWWrQXvEZHA1/E9PpOfCC3I+DjreNbVHK76s4obsDmJS5m4jYCMo3j
c4keUnV8qQiFQYK/8KIHyp3BpVkE7+N2WIwf6l3NzVWExvRyvzlsvp9jRezDekbd
1hwX6swpb1DOusvuYJCNXKGIa/MzOLDuo/G1dB9pcedT4F/EDiFk+Pswu5iJYUDK
FlxUQlBXpAvpszu4s6F6HOsRA1NoMZqMKuTqW3xHJPdRHkAez+p7aPemUuvZRrFD
HXc0z1P0Vq8S1GvMSSP2e3fRTJ8pDGRjcc9OrFZYVR0b/DwJtk3MC2sRQEy2oUCW
QWdeEuqcYSD27y7SvZJEhL6dOAu0mWjLRvS4SpaVtEbhQ5nSc/VH9LlAhAzQFSLB
PAGrC232jTtFGmE9+o+FgwWvHe5/vDU7TV9z4PEghfbveEOZyDdDjsnoNFazNQOa
P0aDzK+B9KQJwhTTRBH501cTq5PetzMOGU1qgQkhtRw06anGPN7cuBEefobm3pJe
TflIakhvsDTmOVdajQEIjx0BHnScNXuf45MP0DnylfGsy3Rh87wHrupYxThi6Gn1
8JDVzUlF3DMIMS94GLxCvSiM05htO7NqvYjSrLi9X85Vl2PytecR3qZWZ91VjW7o
9MTV6PsC1M1l4bM76MwTPZXT/rBzeBGtUApfbZLMjgchhsSQYmNZijcQfDqjiQ+c
elz5irihDkvkAyGvnsxZF2iro/SecsklzlZ83N2jdxRlbrijWc6INNfSVI4ILHMn
zTD7oeu5cDL8S0IJw7YLIQAxOdztmaTv1r5pjFLeW/lH9Y/F1TjTP7ogwEy8yyfI
4VwCQSt5bWAju/g5Doo4jLjxKIZQDd6TMm5qlIINMYJW7ghTHoEBMAN4jngLsfjj
rBHpUvyWpYGE6nhhiT4GvXgjB24tP8looO87bJgqlVjGyB+Ujuy2Vt9CedqsRqMv
WMPdjt/K3WBuSn2BS/H9yY7tXcQk5LGqts/mHBIdkDHnS5qMPoX5U4H+FMrIlZMB
iRR9t2qN83V+H+Krhx2+daqrwB6EnUjk22SRrmcGJnEkoQMVdfTpu19aS6g0Lisl
/kpSJNM/dePwUNI+m9c4QQq/vVy20DhfjjcUjMP6cLyjNHwivrPAXEoAb8cbT46S
V1xwlpUm6qJCAkpd111VfiW49YNngFNNfe0Ggt8yS/R4trqWAZgHdkJ+2rTUOJ+l
XBKwymp95BxUvelSkP4cPnBeXjkCzV5v9bl49q/gGdfIEIHyHLKK+APpiPj7I7gx
wZAthybZy0Rmhhy24sMEbaRa/okpTjFY9YtKbo3NlK49IzuuzX1CZiJix00S3uVu
PgMi+fTM8mKscAJiAImJPd0XG00nwPPS2S1SDlvNmaKRdOkcvN+cClNrfxhIniyV
nLZK2NrV3DM6xTDkGnoC2Ux23emFrilYs3TFacek2Vixtplgn7HR5tAaPlcjBEdu
iG2gMJzVCOEQtaVHCWsJCkbHoYNqsN/1X1l447IJMEA8T7re36FNKDiFxHvdP9bC
svjq2PTm3YEBfhlz/ZuHkIbp69JJOAtRggzf6WoHS/C7fg2IjfsrEx97mOstc5yb
KaxCvs42opVSTRO0iX65YePBJA5Qrk2JHO4AbtacJocopggKLh+gwXzrea497fY6
6hzUuEr92VVC3gtIv0XCPyFKbKZ2OQ6eM2ZKi1htUnsKshcdH2u5MUbUzNVhTDcP
RgJKRsCpLKlienHwrZF1VE4unF1ZXYyZa4UkvovnS/NLd2kq7kDiBn+GhFgFzYSQ
COkXtU/DKo1dVu0aYqJU+5e76wsukz7yZoQXi3PrervLOjHqAYejIIOlW7Phf3kw
Cn+YkqN/+j/0ib3ZKZFyb1qaLF7Q7JdjzwgiC4gMxVsNpkUly59qk4ObkkL+B5Ys
noPRNDUE/OfKzwiEKbLnFhIpSBT6QdB8VK9IuqubMrjypxHVEhxwOLia8+YUEBjs
zrPqbjj3sPhrxBOxvJUXGvDsfK885D2pd9fTAop6hqiU0IDFc9p8lItMjEshaWi7
/TnOYiKNfHJ0DH9Q9JMsXp+DStngtJwi0I0gk+d/CiBX1dkzjDtazCqCMA6PSRHc
l0AnnrsZcRvNs3hx/WpiNncH5syoqCRy+c7zYYXeGRvBxBj8BkYEJLfHmEWziFYK
T02AVMcgy4ZklzSfyh9Y9uhdTdNdEJeBSCLUvVVsjPba+KygMOry2IO5QJL+AnXA
fQMLpy+GZC/b99QIf11nErs37wwdQujkkj3xJV5901/ADqMYNBQoab/tvG9isgJo
ORrXLMF1NuIbR+uQalTJATWZJZbq3ZenWDRyXZZp+b3ZZNsjLsrTLT27NMHekm8y
ofuPf3Y1ApOnN54F5MrSOWPxswz/WFNaVklZUaVET+OLav7hJswWh+YYJrdFlgCA
j+ZiA/FtwFdjWPMcqXeLbgayNBGO+17ebNedsH9zYICImGO/4Mo/ebvR8FbkuoQ3
t1O83hr3Jt2xz+X/SyCukDXluHoV3YFeZ+ZOXsvvM+5PqLd1lT/qi8Akr4Sw/cQl
GlaLS9ISzOP6MSlKA2gDeSp+4CCZkE0uF7e4WkyLhDOK1zgQtBl/edy5pw6OPIJr
PlBKB+Po/PGirqZBF0z1bmzKEqJbwDIW+zFBU/cfav4VQ54wUZCiwNE7bVFwIfMF
+NbLjbFgk2zOD1KXGz6SuPEKkbTd+7qr0jodYG3v3rrSchNMg3QbzYkkjPCbx8n+
NKOakkOGy9o5crlo7KSnEkA8l89ZL9oNIW/Rn7+EKfg7N3B8txUogP2ekJG7ifE9
nckc3xYwYYAWLa0T2ndjuxmIyTF6SmvYSuR2utfMYOFszCaDme02HeSaCLHj7KCN
QVN+gWtWXiNCv9krE0JWuJ46y8wruoMgm5mpHA2I/9Zq03IxCLYNF7xcsDzUK01c
8eS2O+Mx+gdgRIEKy7ObJx8ne7m1m2LdfPtQW4+gOTBhOrggcihICiT8qG9zxJst
uTrrgRJgIY5pYvDRLNIdZi1O4lbS/wKye3eLE25Hx7jygIZY83wadTCK3welT0xA

//pragma protect end_data_block
//pragma protect digest_block
QQs3jY61LCHop0DrBcxpBUN6ERk=
//pragma protect end_digest_block
//pragma protect end_protected
