��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�a�ȝ똇���B�.�Ue��[�=n?�2g�bHf.ӛ���]��:���6b��$l@��k�Bs��C�TϜ������ʈ��������#)����S�� , ��G[�:����h�Wx��KSEAP��� A�5�5��w>v�Ї�Qg����+�&z��ay[���v���b5	.�Ȇ���%�C&�Q�!:��^��֋�w�1��.0Lâ(���l�މ�ɍ�F����b���F�.�C�ɾ�Rd{�oc$�'=e{EsN?%�}�j��H#� Vl�B�GҖ�8`��u��I��g��}��G��YBȋ�甁�l��oM
G���wi������]�%�l (��|��L>����d��5R�W�S3o^P����6�X�7���5��������_�nUc�eg��6)"k+�����t�V�!r����H�_@TC�8�eᄐIv�A{�b�-)-0��&��z2���8���T��N�`Z���>rL��z����yG�� �Wz�*@H�$��Y��z�'1�?�2��sgp���d�"�	[b��q7�V�2bQ+&�I{�������u+c%�[I؆������ы������|T.-�H�v�����ڡcNT�:��V�u�T�s��y+@�r+���jvi���8�iH�'L��il��ub��p2m�A�o��9���k��$�Hr]:rLf�r���ɦfGc����6��P��S���������&2��[��n�_G����|�	��E��W۳J��Ή��z�|�I�g���j�8b��P'��a�l����S�v�d	ݡj�Ɣ��P�U �	�?�?Ƕ�^	�;8��uRR{i�i����Oi�o?2��c�Ř��K����C��"����M������":67Mo�y���1��>�,1�������7D����q3��x��r�����Q�	 ^ۿX88,�gv�H?W-�˅[0��{2P���pz��ϴRͮ�K����?[}�Гx4��6�X����� ,�B�$X���yn"l�N��J>[�5�������[�
�k�N�z}�&�#�m�4�M,��X�b=1���,Z�Lbϧ �e�/^�^��9�T��2�OT�i�`ES����\@�(���z�9���v�l�]H	�U�%{�CX�Ρl��w�������������}�����(���Swk�E��ϣ��Q���f,����p���<�LÆ�V�>��B��l}���;��Z���+l�5Dgr�0�v�
�84.���¯xM<Ѭ��&[;�G���9f�1Lrnl�/!��.��M0Gv��j|�VFν0�8%�P�f��+9���׼��F�La3��\�Z��L�`��TG��`o�3��䦎?�A$g���r�yY���J�T*�cL�aC��1oݣ��4���%�3;9�i��qz6ǂ�߾��6�CC��GN�����V�����ʳ����i�����d��o!�A.�_��ַ-����%��7�hIq��Cq�����x����Ϥ�6��Ph�� �+L���<Cy&�*���b���0��lx���Q��f��;��;D��{9@!�v��Oa�F��-af������TxX[cn���1
�����E�f�����[�����l�P�к]��V_<�/�!��;/����\"n��$�d	��uc5��H�����6x��ru�h.)h�T	ͧ=v��
ύ��~o����Y˒�- /I�%��앷���F��a��X�AEY�ɳ���+��P�ٷZ����
O�fn�����ҽb�ojap�_�\���V�.�[W�􊪹�����`\H�h��kna�޺��ћ��Y2���I��bu������:�����5��������t��͐�y`YfH�]�\��5�[��Fx�ybԥ'.��XH�����(�5�7��Z1_�c:�_F�ohN�u�]a/�y�s%;���ڢ��p��7��g�?s�
��/=>T:�+��0����Ӿ���x{-;jf.Ї�e_X�8��ԯ�C�X�w~�zItj�3$�8B
��v���n`x7ʀ}9dm�T�@9Z6��t��� �#XD��6K�x�<[�k(�t�Z��y�_�N	�$�\*�VE�4Z_a���of�%T�J1r�	�f"Y����eQ.����w�F򄗋����Hd.b4й> Pb�y��1����7u���8��9]�u��\�>�'������He5�?v�c��|��m�H;NZ�+P�@�y��v<.��yÐOf{9����q���crѮY����^���+�?A;�- _Ws�c�z3*k'Ȳ��f&�?"����_�6;�N����GnX�����4��VR#iݱ�A�Q���g��/��*��A���m�a��T�_X勻�R쑐x�}N9�~Ԑ�o �p�:�;�I�F��#h��t����Piis��NO�v�nF�6��$��F+�#��J��Wq�5w���Z؞PN�=�Y��M=h��NV�����Sr��/�ɨt�f�$#]���x�`��u��_�5=kN<IwZтП�ؼߖm�9!Tv��b`?����~����l;�\:qIDm�R:�U�0������G�Y�XCs+�ߋ1b-�<��,���`�n�+���ӻ�#�Z�|�Z^����/b���rm���t���q��Bq���\v����	I����^�5�X��-�U��C���	��
��1�t�
L���5�0�f:�B4^P��{lD�%K��M�;��-��t�p-���0p���"�d��}v�#^�������	٢�^�Wa���l�5� ��&;���j�-qƶv֕)C���G�3fp`��@���^����DTa�m#�Nl�V�l���������PO��Cҏr�-�4��2�9����"�N}��f	�3�F�������TH�˞ <����(�n��M��8��a�)��@l��;ʻ�c����Zr!�����фʁp�|l�"�x�\=�N�ɰ5�j�a�nFğe��ۦ�/�b������F��"q���ɸ������	�N�ge�\u{��7�G}䑿��h��j��>k���5�	�GԹrv���V{�k��ɫl�|��|4_J�{wK���L���[�7�~��^��t_��alE	��z�R@��:_�V�q����a.Ek�f�<�PĖ?YHЯ�N�E|������:���&�W��E�<� ����:Y�(5r�g�2���a�"��l�-L_gy�v�P��Ց���t�7����J�*�-�/Ť;�/�i�	�R�E7�	G��clI�I>����3�z�RfEw�ޒ
P��l�#%A���P�)׽0eʰ�������P͖0��ݍb�%ZE>��8�Jt��I��r:����t������.)�|���߳�G���!Z�Ed%3iz�o3>�� 	��S�(�2�Vk��[B��0��?�N2�RV��<����B�:��kv�iٯ����rQ���⺘�͆��
낥�ݰ�7s".�����������7�[����9=�Z���cѬ�9>���6Eeb�槵�TwB:D9<6���n�߫�P�7�d����*�42�U�/<A�����\r&�;�V�����t?��|��uY8����U���bG�����\5^ �VN0b�]_2�i,�3�Y�Sg��®ͯ��B2�-r� �ah4Z�d�A
pDb���T�Y�'��jpI�'�ߑC���&ɴ䵄�|&�P�'��,%�d�nwX�栄�i��MB�,l/2����ݯܧ��'�s��/��so������L���T! 9�B^;N�����Dky�-�P�ѳ� �L7]�ӘӅ��Wب;C�m�R�Z6h��*!�ȵ��3�o��h	У�K��Їy�{,l�z�%͕{'�����+���6���q(i�*R��fA|�ߦ6҂lO��m�yR;}�6|���&*Vʧ�Pt6k�_
Sw:�<����v+yZ��HG�UM�-�R������'U}�b0x5Ɵ�-��;Z��8"�\4Gn���"����@	Z�>���K��8?mY8�鍔6n�J��VĂ��dx�q=L�X+���-�,f���=UPK5��}�3ҕM���&��2sZǼ�ıD��phv�� �/�>�������[�Ж�q>�7a�a�:%�k_hm�+���:A�)���A���u�ʶe�;O
���T?�Ǎk�;�I��J �l>��ePWu�j��g���D%>�H����C"��Ѷ��DK�9LYjn��?NBv܃�ي��҇P��ɢ����ϨKz�D|�y�%3���_i��U��<Q���7`5�T�^�l�r�l�����aaqD��<��ƣ�������a�������h.��3]S5�}�MO�C{Q�an�� �^q�F��T)��;��섿�}b��,���fS�<��0Vd8ގE6�����+�B�/�F����%�MAz�����U�?�𫯏ڪ�wG���7_	�U�!�H9*`Y��aP�^-0~��$5�#�P�ꎕŕ%M�%n�y��6U�ʠ�10^�BK�O�SDj�.y:E�E�>� !����Qu�������Ut��'0��ͨ���O��W�|1)�i�:!�9yߋa�ϑ8�q�{4�Cz�;�5���cK�������/^�aN��w�"�̒� �^.>^o�m�k,B?��� W)���n��%a����O������a`�]K�4����(w���o�_���ܠ���u�*!��O��)Џ|�4*Ou	E������%�����$�2��d�z�l8���� 1�!o[9mQ�ӆ�� fY��+�����bƟ|Yp���^Aj?�2xfh���Z����z����]s�l|آ��޿%�������V� ��h\�4�&��^F�=d�Ys8�3��z>Ҳ�5_���-�Wg��,ōi1du;�H��i3'���F�2<��kэγ�O�wv���i鿸%�GE]&��l̛U�=��e6�]Q�� ��E4�^���zEx
�e�5�����T�P���M&��xe�2=�!�G��S�T�s��a�yg,o��\ր�8�Vc�$>vk2�
��`�?d ���Ùu���L>��������9���_�=�6�bc%%�o���]��.@��b
��*6�x�D-?�B�&M+	�zY��O@�*ׁ9Բ*أ��UV�Qu�/���E7u��g�:{�]�%6~�!���!Ͷ��}x�ϽcFʵ���n*��G"w.Պ����@���R���#e�BY8S��^��}���,��w7�5��B<4���LE�d�Lt��4��s����΋<��
�L�4n�'/�'M��9�K���^�e�(w�gL����R��g��'��"�����G#&��Ck��٘�{	W��H��G�L��X�:����A��)Z����4F_�9yo@>E�������P�����vJlJ�Yq�fg��I��x'#�.C	��R�Њ��W/hZa����"�Z�m\k�¾j����r1�[��"�`�[�������B�$��ע��aZ_���捻�Q��-�D ��R���K�#gr�m4�F�d���_�W*����=�N�4K[��ʟnhR�5�ie��T�-\��Nfi�߆�1;��tr?g-�A1|#e�;�!�����o������`0 kg�GeJ�����$If3!-���t��<�O4D�`�̾���� v�l�]���%q(g�׻1�G��#��,C��!9��C�8�&��~�	�I�b��i���]��S�� �����|p!V���A.<�7��W�Km^m�@��4�ٶ�HE���?)c'@����'��A��}��I�UQ���rĆ_�ӎ�RI�7���O7����9��B2۴L� k�yHgLa,�@rN�h�P��' &ko ��S֙;�	��=,߆�ۙ��������J}��y�6^A0`lE���'��;^(lbq��,�b�]��R��U��A�J�~G�Ҫ�e�8)��G*��I�J�6�E��:����Y�EĎ�=ow���=0>���Z�1�B������+7HK�2?�ݵ=AT�8j�1s�Ez����I��<�-����:�l̕R�� ϞrjV�2ǿG�P~��<K�&F:������e[�,Q����p�u_{5��$�snk9�=eL�+L�c��s6c��`�y�Z
CK�^r�}�k?Z�
�?�)�[�re��0>� ~M�L��d%�l�6*б��;+SL;�13L�!gz!���N=��xe�x��g{ɷ%�e)	zrU?�K���Z�3����"�QeMa�<.:�iC�O"�=�ܥf�ۗ	�v�����տ�I��	� ~��k϶��$q���2��ս&�{)�P<M)|RLŌbR�e:z��>K�$��1I����N�\���#=	s���u��Dh���?����􎖣������d�����&w�?����zhӝ^ȇ�I��k�h��$e��}4�Yi!�@ �ӂ�A�e�'rq9��M=���_� �[��� ��Ȼ״�{�UFK̃���Fk�55H�Y���e�r��+����v7'�Q���-�'z����2�1�����^�f����&������� ���fQ���~�"Oi-��_Ԓj�W�l;[�и��lR�0/)M�o�p|���C�iJX5�e�ۈ��ۘ�2�	���<�áV�1MEM�k�Ġ�&D.�r?��C�� [R *����.``�{�g���-��vZr�p�h��^6V#���W�/��پ)��N�Y����
��'��˄~�ĳg\�N�5i\F��ey�4�:�5�$��M���22��)�.�m}8��ˏWd�k�f��ѝ(ܴyg(���ݒ�x�mh�J�5�i�`��> i\uYd �T�N.>G=��E��Lb�d��s������C+p~Kg�w�J��Z|Ρ>#ڋ4��'��[���vw3�OYH��Dd�#cr&�Z�L�6����ϗh�>�[+)���&D��-m	E��ʝ��^�C1��%�ݿ��[׉�;%ʶ��!��T�,�M$�3��<����b�ɬ���J��'V�#�\����Ҝ&Lq����c�]J�����38�z6ם�����\��]-�՟�e���T։Ȳ_h�/\w%������oK��f��Q���*���m��<�E�Q+p��w��ˤy=s{_#M��Q�c5֔i�9�F1�Baf��n�ItހO��;��g�w����	���&��@�	C��O�H���4��'�l�:�Q.YRE�>�;�g͝��o�=W������&�OT���P�sX|=��w�[��򃙘q7Oë��E�B�0�À�r.|B�2i�}�����d@?��d'����h�+֠��� ����L�e�*T#a���reVco�d�"A�̷J�
_`�B1�Px����Q��(=݉����fg	�2���K����\��1�ö����%)�6]�
�-����:q�q��B����HL%!���/�}
�0X5�uaZ���I��~ǭ�� [0������9����ec��)Ñy�W2��n���Z�ne�>'rn�y��zĦ��lDu `y���탳�F��ڒ_�l�]f9������.FD�]��Ha��~u��_��t����}u��e¬c�����ˋS����
&F�	����>� �8�4?lc�i�M�,c��al�i�R�`�,Y����C����j6�mW\�e�pWbz���Ψ6175��Ԛ�t��C��7/�y�{7~Ԟ��)`��RV���/�3�Az� �����Z��*�Xhr$��!���dNvS�֛�&A�����&��'��<��c��J�v��o%�����<2{y�'���Ys�v��������g͇��a�p�v���װq��.���r����Sf�C<�!��p	��=��XJ]r��59Y�m�ͣ�%R��<؀�n�:{���C�J�	�l>��L�yr�50aW6ʰ��}�\"~���ѷ�3$�d��ojip���յ\5!F���N4��Iw�"��~K���%Z�p���F2��xn'V-����L�n�\���6Z\2�QU�'�r�Dx�S��d�4���S��W�����}�j���Q�]�A���~I����c#�qD�Sꪱi���u� Xߡ���v���^���^����W�[�h�9��C��V�4Vd�{;�Q$}.�i"��g 5 ���4`7��f��Vm�,�����2�Dt�E�7�?�#��1�i���&�<vd�ҀO�ʨ�Bu�9b�t=��c�u��۳0*<�Ɋ�����F�Σ9\L�rK�X�O��4�6�L=<m7��Rcj�Gbkw�R�uoa�k�7�?��'���(P¹�ɔ�S��uz.�ʦ4YV�����rK�A��@��b��(-�ce�H�ތ$���LO�羂��`�|j��!z��&�a� Jj���[2B�r�kċ�dϨ