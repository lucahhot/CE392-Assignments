// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
0nGDJxPbTbStNKk5HPez1x+KGSlofPZwoDEvqYwm9rEQGXllnBkcDSnTGJnstqtI
uUrc/UtLuf3YY2+rb2dTbdHr5iWCk2VaRrPgGrbzUk7tyAmWag4NQbZreigBLDaL
I6w8zO4+KiS+kIKoI/sAYNiY87ugailWPxn70XJBSU8B8L0KXLhUEg==
//pragma protect end_key_block
//pragma protect digest_block
aWijdKiXRCL39nn4Q4etyFXVsb4=
//pragma protect end_digest_block
//pragma protect data_block
c+hOhPS20DIyRh0zzotjl9GxeLeOiGa3gzutopL4TdBHwYnO9Kzj7vmUaNCauBmG
m2afvtK10xcHaGKh3I7SRzqkGGXDqX+SvJ/gMWvHqXt3gmqmiuqSlJ7KPwfK0S1S
TGOxyYP+zybwPCRZmq5kWEXe0Wz3L5yMM1LZfYZ5yckrPqyCeG3dtIYwrsW/fyPA
D9afc97R/ekJwY+Xu2IFtqFlTGSvPLnMff+Fw80jc8/fOw2VaG/HUz7zLQs03udy
0N3aEiSk21QiSwdy1Wm5h95FNgjPa2qDaoOhSeGSILKifOzikcmACruOaNJdoRmO
JCibdUN+txHb/DN3ehqS7dYHvgDtI85kqbL8dhqg2Mi5rpVYD3co2iZhjY0CYCKa
GCphvgPNn9GM78P9kw8MxMDeZuCFCA/yEM56/38HeDsXkCqothW4d8q0P4Uv7bq3
A1GFU9V+COEkApRs7E8+sJRthN7g9PrUUokeF5D1fhqk1Vx/K0jCxUnOHjG9BNa9
mYS8CRSKivv7k4Zolyr+bD9LXthseP9kSouf1Nbqg07znPN/tvnJ/JEOjq4+4rUb
9Pf1tb+nP1oL52RDp5fZU00Tlfs9S0Rc6wcJy1/dlLOp0U7ujY/P4hRIU3m5OQ5p
OKDHDVhc+wHdWauRDubtsxP4e8NNDGmL5CDC+scAK7acEgyhublyvHxlmE0UeWcv
PnBHTGpZb1D+EvDI9JA49+pGKAzPCKvpC2TqF5q4QYWBRUFxNFDYILePb/4Y/LhW
GNE3o34s2y+4dDVpga7XZpzaz+fhA9x9ClXWMiyI/zfwaPpzZPpmf7vjl564BHr5
U7zy8OH0Ew5EuMZ9htMvVUNPWZJ7TzSXN32u+2kM1W8AL5bYszCJ3FwPKzhqXULm
mn4zTDus1zZ30JMl2gjuYVWLXVzl7UmDbD15GBeXyZcCfu/jPFQxl+erF2lCLYla
4Sb75BFwHLIRc79/+7jf5h+O8r7coBpY3O//xyrxsecvxNA3jp3C3ZJW8g4HHtuz
hzRIC4Mghlavqueh61ZAMu9qh2tALtPqtL+zp65ixUaSF+d+NoZ4afBBx6c0VA3f
U6ArzRKss00bh/b8XlWwtVNRz/Q/sCzXOT5Ub+vQ5RV99YFnJdj1mpyBFRArArSI
8WV00DZ7SS/UaXvLZS8Kbx2FBWK1LLu1IKDI8hJuK8VAQEFbx3aBiiK6IegqnleK
6Ch4RPg8YgJlIpa0sFCDxlBkVeihb7Sd4o8UuyIplp4PxU03BokWcL9N1qWTiNGa
V6HmL0B5ZxtQSINsuPbymHwpv9ugw0lQnjE5FcmpDIDkZ/f/cN2O9Gcac5sZ4GjW
IWSsf4vg7twxfKCFJEihKQ8QPlyyec7GsDBdoTrvV/7sx0kQBC0yLMB+zBrwCLpF
a2N8REBeOLehMUkpsL597mARofVWMiHvfxsjzWf4X63cVEwvogL//dyhOFR5z7t1
CYRYjMcG5XYDoIMOQGJIJoL8CjiIDD+vuThpJ2hDxsXsBM/mdNqh1M55qO9N8uhc
SDwyzEL6lPQEjgalDCpctBczfeEN+b5ThWJsFL31LwpgrzgVrdJvwI3YWipkxFl1
exCddboVdYQf/pg+j920/Bj2EuWzfb3xV0uO0Sj6QelYZ0ZPhEep+JMpErusIiVH
QfdGvg3ZfaNiuPgrVw436UEXJhL7jFssS2C7lXVYbGqc5x/msLIb8L5yFlzbyxBW
phJCrJGy/+J0z+L4bUOVONyZIe5ZFyPcw+kKv3z5CpXDK8R7f27xLWHy9izBggg8
e1FLzVlOBi6K86Q5zgvWGFBcJhaXhN/PvQW2grfa2AoJZTrnOjv9GJEm5RH6G0AY
cF/g9efVCLVggToloY6V9nK39KpVci0QdJ2tDh1zJIMpG7tc2AqQGAo8Bf4/P36Q
9sfpA17TEnhA0RoQcDPw42cnZjOJGG4vH/ZHSVOFqtVH/BTMcmV2ltUUwmacuds3
B4esmscsOaQZLLFa0M27euTEc+FJS1wJrujaTFVxZr32+seVRaehXxfVSZH7m2dE
v+Gh8I/WEOX71y1Z3/8W4317Rok6cdA7vYndqU5/S6VIaSxQQJLwjWAkXJKn+SzF
CwWeGRr4x6IbQcEBkZ1Gn6YghSRQSsBJQMICooCz5tfE+Vhs0a5BsCjvuJ3iU7f1
wvtrtaoyyOjkOa1bvth7gkbtyBNPTYuqkNwnm2L5YrG410RApGtNowhDjCHNJtyB
jVoIh5HdoV6eLUXRQyYmAVaiL7lZ73RepL2WuUBsGWLXMOfi3GVyIp0SJrdqK20Q
iXL6ZPQ/7ne1uZtWLKP3dG0LQdzljrrbfjaZAXruHea4U44UQFpQOnWjdKbtlKYQ
B3dnkTtkcCJ8R6fWYgP6h/KRqkCIU+kxyQh38VKaJ6ue9XN8YmT9NLQMLtKx7+e1
0I/eegt8PxnoEOOcp8HfZ9D7ZA8p1QUhQ/1FcboJ5uxy+XaDCy6fa+Vd4aslFknA
ayMTCfxv7s0MagtQQn8pd+k+3o+OOQ02SoaDvvcOAJApFb++1umCbDVY4IlfW5KD
LCmVhnKBFY40Eq/Nt5iZiDpPb1iOuhilP1FRwhJTslZBcAv2zokHhw/QzdizYa4M
o9L/dAXBOPU4Qf+xIKqDmN6gs/LZ6OMHNzH1i76xj46h/y02W+BazjDUcqSYtsxW
JYPSX0e+MJWlEoufGXnFvHx2buGyZmIznwTZg+M1jP/0GAz9ND9EQK0mpcUwKryQ
PRF6vjSRfKEwWWc//1czzYqr8B1NgRRl0h07hLA+UBOr4ZoD7olMy2IATs+wt8sE
UzVOrKsDyFC8E7j9LA3SJ2g0MxzPEzqZmAN7aQO5PAYkc8BFmhgwCW/MkG62tnC6
wPtRQYSuWGlgpiF2c4U4NOavoJUT9xQ2P1UVTBgsxsVI9dA4GZyEtn5xqC7ucmQj
t15K6W8w1NFEM56gJoopQY/ex36DPSWNVy8lg/ccPeTJ8lukB9wlQbavVFMPn2DA
cjLZOsvj1FIsqgWSh1ddHrl2GVQOqQldCnJS7vyy2MbO5TGE7vlg3oCT561Dcm2A
iivjFm/bslbSYypm5PA7uMjfNT4LLD50StR9yhWSp8oYqiN2fvWrCitodeolUpm4
akDvED5isucCu/WeEPyKJFhEwCvSeXpiFi2FO5khSK1xBTcmUD7aY6xXF7309QV2
WH4tRk93DfBa8NGnfQL5jl7TE2yy3X6EfvU2NHz0ywB7Rfj3HLQC7ETnVPr3ESMX
v0l9oZd1VoZQTVB3tOqLeLMAbrkUiQgVMCwodUFmoilwJzvOkzQ9ag4GwdFTIzdW
A+lVnSCZPrsJrVz6EgZ+5TxgGYi1AunUggzlyrCfK09Jgpqmybm+V4s6ApxhrZeS
9Dk5614n2AbM5QoJ2Cn32VlL+Feu9gM7UkxqkgoVZvtgk/EDyXzvo6fGzTjYtIjG
7ZtrKEfLHIE8NoyIz+f8/h9mi4jesn/FrpheZoYWoSxX4TW/qI0sIxzQHhDf6YHB
xzHMfBFNbJpsH+3i4zyacJZMgu3jwEWdJf7XbyVvUDozPsyZhfjd+PQWX5NiaS+t
WDEUIV8+T2llfVGS0O0kp0vTxbv5NgHPlE7Y/Y7ZIUukEyWv+MmxRRWBbKbSpkFA
rQpKVxcb7TvilSnebvAfXp876jXN9QyaA0IuHoe3RqLg920STW/aoAYe1qHSKOW0
aBbfbIfhTwER/GwtnUy/9steame55BuGIpCcRn2YjsLorBr87H8yRyAfNUh++FNS
yo95sYAx3ZByzsO9Q1hRp3oGmjfPZSMRmfeeHdK6QgWM9M++fUtpCKWKyR20Ub1t
LfphnJ6x6H3GFtuWR4tEP9yyivws6oKCv/ErlMGNV4bR1DVU96e5SUAJ7AsmLai1
8gfSp1vnxu9gc4E48hhDdUX5J9NE0LiAWnaWiJtk7DA7yrQ6rHMd8G9dmPcIPBve
zNvF8MfpakpYOa20e1o6DctLa2bjSttXx106PEeqbdXOACfBnDM5RccojOePvmEC
esnIQUBsuciVb4xE9JrNFv6pF8v1wTMaJXtTv/xoaxYbq8y6A+UFcksP88EnrU78
E5q50kJvyP4TvPLEjdDTXcv7xpwKIsKcq6Iu0TnTEF/hpUcS2dFRVv8DBHMYuRuj
UVr2S38As8Oj6jt3hwH34eLveBTtxPe3+w4rGtXuSMMZEZeg5uURApViyolCSsFx
jtXRNDIQNjkrYRBRbUV1eKS7WEU2KhQ11sfvlV5ZiCE8Jjz5AmWQSL1e0+ujdGKz
Bi4YsxxfGpVQ1jaFjruNlZoc/LGo0li7PkKv4gJ7Vf0964KCAO7/54IKO5UAgcOk
DNNR2LXAZEC6ZvdlSUkiQ736tIIj8yducF2te/sERPsk5sZiuGBOpnNnV53H3x0s
BMYyiD4PRNCDhkdAkz8SuKFNM/fWUqndMnpbgWdjieDbvK7I2AIxEckgmnEELEbv
XlL+n6gssXVTo9CN87va2KYEnD96pWd54DOcm+Qhuct+tU+SjbEDbgBTs/RTTElJ
ATywsS8DvdigM/gdAvEYcBGTqvwPvbxvFm1q5j339jJ57B2eIIbyyFTKMEFAtQlJ
7iufTKj6p2PH8tIJcQ91FfuLcIQHjwU9LYx5u8Xm6qxlt6vJJoHIyByxvSa6TrnK
Cmyvb/4Nm2nT3FrGuDTBO05YJwwMcKtpK+qb/KWZNBNfmocAEUcbWfhP7Ex3fwri
seJrWC7f/wCtlQafENLxUS2tffjfFBh4xWp63gWW+B46iX6yUXhRzZs9rNxX+6JL
cmnMebApdNgwphTYNDcHtn3oyh6Na8ZEZICV5QuyfMV90Eg2s9ZNRaBfes0AVBJH
4MJTKLB3RXPvjKZs4zF9gFu+XG/xM0E/fluuwvZOlbTwWTWyM2Y/EEvpzpKt+gUp
P8b2LkgfpbZjH21i8RsLngoebg/g6HNalcERrvryWiMZ0NVIvjR/GQD/9IgfyoAz
wFMMdjbWDQg3sqNKZkTNm+woyU4++FupwtU10U6H+wfdLakj8z7QkO9s80yd3dvB
+SIvmuD0jHb65GsWBoY12GUgDFx1DpuWi+52tZU86qmvvsmhSEZLUzhusRaV3nyl
W/6pfBKZHxhSKglkweiBpAwvzjlXPBKYsQjHTwnHXanQ/+15zOiUAkXpXut2lc4e
d1w2PGWOpk88l8EwVGeC0zMomlQxnaqMhIs/nOQ5fMqsvm7CKYdXJDiJdTYHFNFJ
mN7N1Q7c4qwES9uyAMtRSUFK63kJhX+2tnb51szixbGNE3Ri8L7RTqO4T00o/8QM
XbdZqFVWj/ydCirOBMzbh+pDBQ41eoB7SUJh/pdzz6QNFlYlla/0SefoW4dLSKjf
TETIURmhZewFj2WW41rxeW/n7UuMhzBhvBw8jhhLlumhJD+Xxe84mLpEpNsHD/If
HYSlZ3AIdlaTP4gSqM/F77Fb7PVaLIiwN1At3j8f+pb730SKLHqWuZwWgmY7h3+C
/OQG3DjYwq5Y1oDzEtnHMoi6xGT3n7S33IIS6SuY66ZqbOBIqXuthIqiVQzaHReS
NSx4yu5NQxh6RTF2JurXnKSYJOJ0AcfqglclFIXDxNf6HDAnKqpvameUpZdDAjKg
vTZmILKQMLEcXi4yMmUdnhw4LlfLwRJDtA9O2+LDVpWVu44HORySJ/AOvIRXFQ5e
mUmOPuwafBxz+Jrf8MPZW5FGs10Roe5PjGZUSmBioJr5zfrTI79ccKT6/PfeBE4Y
k0UTTPnEvbEuAPI4PnG/TekB8qhJKEU4elr5R8uN9QPHYDxBW5ZKEWH7csP1E5LA
horOe+IxRY6wfECCX74HkNOnxXlXtvB9IQW/NbsVhsi7RVtvozU4bT/LlS6vs2t5
RqlyiCCnMiQrof2IAC5zIsYqHeOzg8LMiPC5pgf7KbrBM4tfDde1pIoccyvr26wS
D74TZuEoEHjX9WXxfvVyiH/11mi6CL+28rIdmRGD8CRdN1LeH7m5eFESxDPdLcp5
7qj4VB0/MZewrYxChqO8Du0SRg2FBv7a5bFKAYIc3j1+f5zxm4DaktHYYn5uDXRe
+jWhMa6bBQXaIATd/vMwPv1/mlsB7BLDkV40kA5zGocQ3xrTm3JCCD4hepHwQJyG
e5HoN2cALOAbkwBQPlECZ4FCYgkcUsy6waKx8dsKLWMXe1wsJJrhmpLeMYJoG7AM
16DOCizlD/4hWt6ddPdpCF4cr8kiEof/3WzvD8n1AXTvMMBdX79fRO4724DON8Th
hvBhQCCVQttLmrJ2Kr/DkiNFI8u+ZAfiRbaHENBV/1v0iSI52X1Wzh7U6lhSWl82
TWZRv4scbVahL+5fJc+joBFR8LepIpZ+FQOan7V+6TgH7zCweTogzeD0ikCJ3trC
jb7Y40dzt+RIyEYKwMIqH03Epum9V1nyD2NVygOGGGHoLLOuHdApwGjuR8HyEW0+
chpecf/0aPnvROW/w+EVXh0kC3DtbM48/ujYXpw15a9abVvgZL4O6ro2tSu1b3GP
P+BvGjPDRRseNtiDcW0Xg5YvOu1wi30e3TSENH8PvCGNN3mlqfUYqzCXJDWyV77I
I/9CGQjza7DYgjPtmcKkSy6EuXRnfJqtf3yNLTaNucAo+eWBC8OoxbcuAE+Kjdcx
0MSN5OxLTxRzhtF9H9uTbDsa48gnhPWIpGlTCMFfbqNaC2C2JvyfKoLzORVV+U/B
EfgcS/S+LzOajQIbDqYa5tkTza3FkqMejtCLU3ikiKpPlen1yui9HBBVHGK+3qTh
f8Byf6Z3dEa8rXmMSrTrcj7R9xIo2ZuA5Kl1FPDOLQz5YVgAeJbfqcN4ClCGZasf
OP3n5LPpWbiJGtCSKS2dF5L2FfNlhAO3z4yFuIeC7usjdACNuWM0cLOCqNYRsFco
CQL1mt3/IPj/Ehugtt2B4hEqN2s3xdWwq3DmAdZxM60SWd0rSuvD5mxU1h7T5gL5
KJ4gBzwc4tLGlblti+WST7bjfH5PhYHFtTrD7kwVrEorChJqms3tunNuogpNvLvI
lnQJOfJrqDiZELSx9iwlapz4SDU3f6k1OGnaiYgAQjumVS5TKl3pyqi61Gp7FFAR
PukOzlvrYmylrL4kEh2mePUQv/yQZ4bV5auTVE8+sxfuTeLeXYGiSSiC+G5HqQx0
o8TetBpzQiy0OGkPpselzKi2MNz2D48dTsxIiQ3I7n0H9LDXnomdhN1VomUZYczs
wFf/zbJwBU4RL3T0WruFb9U1WFq9C2V62ZCn58/gXzFdwrBBb623Cv9KrRdrmGEY
77jcvmMrAVurmZWVT15qLkAzcQgOTtD/tBp737sVSKHCsn6fB6JPjFOz6US23sV4
Vy4/RsLaRI8v6StHG4nfWPpr3qhEE6cD2CQU1v3MWLM+gay1LZRRrxm4TZ9vbz8P
Gycrn9+4ELABb+aRBFnEkwB5qWhD5axnMvsyd2+f/1BUQoajkpJMP4yWn7s2o/GQ
UOpZKrQ9+cUg4hlERvQuCMFpbu7AO7C3RpLBTW4mXxW2wfFOdlMsuOBgOHCFuPa8
lXw11DWL5dbOzQ5B/szTOFSXndSC6x+k/PVal4lfIegHSCvloGol9L3kKvREonWy
gOAoMrBCcCl9v0zOCr7ZBnxw/HlDzQyKpPD3qlmTojARp96R8hIP7OUDZoWLKIHs
F5sWEPc7qD+HBTahG1GDngxJIjzOt8bVNMERYFMLJDjNheCPNVOXcSbpjKh+xGRg
GMw3tp7GOuT4CMeDntePt1kAgO4kqGiwUwJIReOIt/vLf4C8dOYWivvUd6J3MGu9
yAsjHVk4VedHSEYnESMpA9Wulzbtqshq4zEhER3TGPAU9l2YdgxBfuXfdxDUqCKq
+gfvCZfpYMzqPcq0n1O34E+h4hKvls2enB+KXWNK2Cfdj9e8nJ2QfOpFX1IYMjt6
+Z2vsCwhrypYX7cfNiQglEqOMoJ0LkQLWaYjcTlJBw4y+8YSed1gieARLxA1N23p
6lQPd/OlZORRByYh+o42IC9GS9FHPOupdzPwX18EQw/YX0RvbM5pe5H5jMy24DXj
ztEUsvy9Yy+4QE0xhQhAI4ezBN9tLa7pZMv7prXIttqghLIb8y9MPpYVCY/1Ih+U
4TAuI4OhVHVfjqghp9z6HPFdehs3VKWras+/1wxbPcGOY1wWki36EXEX9KX9ED7s
RXEhMGcPayaZGcv1UiEH+KW7UbTE/sGr8jp+Dum2XYANCmxHXjbtY7QwE2r5huWA
UeWtapNJ3vH+qq9+AG/rnoYuJGQF2FX0cBzrqk9loSJvyHXEJaDRathD6qhp4S5H
gRtKaTdcFvDnkfgfKvtVvQQUzWFc8EjwylvJgxl3Tttf3Np6gfKeQBjoUytMEFGU
GXTKCSpAzXY0QmeU48hP/McdluBuyJniJIY9h6ePFfEy8YqqkbP5pzSIXETRM3Rq
D7y1tK9jGMDEu1g92xy2h8NbO2irpSZyz9k4W46wjnjrbNCZwZX/hSiVr8nR07/q
CzrRLDy7WrVC1qPdrFvrzLiuZngJLaBqGDTJwpps8q3xkDAGyI3U+0kVyMqNB70a
6LFf/nNu/JN1bAeKSKk9ltfXuNk99u7qvgPa3eZv7sJFn66NlUUY1zI1nK8hosRg
PDrX4+zYTU6gDeKuiHyoq6G6c+YgN1whq2xnjw4itYyJtGqE1DK8C+hMqzmC/Jqb
HQvBKqtOFXFueu6/FoKx91sPD3l0TOicAkzU5tZU4++KSGeOedtzktGEIY4/oiLe
eUJi+oYt3+o/e7tZ3GGjaZa/WiEuQcTeghjyS9zU3YG2HU0hafz9eLPHYXRcFzkM
dxg+y0Rov3C1Y81UJiIQsBxKd23y4cLxdF0ESDn9t96/RmW/jt4U7iw8iqgUC+vb
d14fefry00HYE+U9A0TQEfArdfn4cCfR51o1idPBeu5Reiomh8ORKRR8u3zrNwem
eslGqvLQydsRPVFrPGWxgx38VNvxMWzWEwMpBJ8JmfclcjpadKSabQlp9A9x4TtG
0j6a2XyxmFq68WNapuBYAlfsBAlR592Lum76SOcqvLXraUnmmQjVuervSnMgN+cn
T2Uqqz4Q/HJ+2RjCyHNo+KwDNb/k+4YhrAJYjJ/NTrZ70JMTwjoH4J0GiAcyKo9Y
KUADSLTvwSWrF0m3dqxPD8skM3yBp2Dqt0UfMLtGdmLcQ+po9Lg693TfDYq1Q7Ev
9Jcv35sr6FTg4MB27MVbpWu/mBbY+ca/4tkjGcGx4FTDW0ZuqBNBuvluXUprt++9
M3e7fjx9MBZcQpoBFUm6fGauzxMKvJ4jO3g2olj1bPzKG2pKJ4zUkBVwg3tXcGKN
x4JiYqFasSeJ9ZMP1s2RM9J1qB3j8z6buuJ6K3qp5RIpzfBFWsmUxLJtL1OGhP0J
j4ZqX32DAFaQL/VVXS1OvJ5o5c9USMMUXiCG0dQPIJpSsP1cQqtDEhX6m20s/QcH
5Rz8uD7px84LRNhYRd6P5jASVtLntZn0XqOZy+h5JhnkmfR8q1o/le5tcxmn4DY6
1aCFqm6fSxQQFO3st3a27Zz6K38MbmKhNO5fnOgk/Itx5xVHEsu8IpbBWmJtu0Sd
n9DZpcmiCPARgRwogRajeWm/a4rSkcVI/dFFELi1FhfrjakQ3Mw6dQLIRzBPl4AA
M3Yp2gQvaw92SGsb00Hph8MEMjmDiGMDGs0yI7uWGTY456J+pGZDu5pNm7nwOsbT
KxSKAYm+J7gN011p6DHK1ovJSa/UyPqzJaldE2R1ABjvBaCqPg3M2WBcmWZ1nT+l
UmNahw8W4c3/XvD3ZPK4KLx2+2ULJ7Yt7JgHzj70j+Ke8kXdCAd9wBiAM2Zvy9Ck
klPYZe6bNbcVCPM+yfFNg1zIgzCcVjnNCqfDVIVSVLrY0WSt0QuEKoyG18wyG80t
HjvgZp3/baBtWaU6F/OGLeHP+VCM5YKXfMgNjHfWL9Nkab9U6Lp83lenAVaC00Ud
gB7R6aLD7tMiJ6UmOOUvUnZjfYVeI9SUveiS7haIMx3ZAVJlrJ2di96fL8yPJxGZ
MkMMJjjoUFKMQ+Nbrt7vuYQxMRKkTMY6xQxmv/3//quKSN8Xln7WDcjZr46CrXGQ
AJ0GUuy5Kvkp2h3ctkunnWIJh28MakITKg6K1u52vxMTpVWlHe4cUUY7fJ7dnRAX
2inFYNTxTKg5lEqb1QztM+62mTcsyfZmYLqD4xaNJuT43zOlNRQxMG3AQfp83yVF
//DqpML5r/CRW5LxHnCqSsmNqSJfUhZoBO3WU1oMxKrj4io4vrDpGs4kpcA3Nu+I
jIU4Adr0VOcu7hAZidFAjI21Ae3H3/ozPVDROvs0CK1PVfTLQl46zq2H4q+V7qyF
Tsl7TA84F0C+NVBAx7zxyeMv42OKTUPO7XMTHbuZ1uFC29yprPpsljhOX3i+b7+G
LuLrJm7hN/zyrgWlaf2u8TevNl1agQWm91JVNqbtxInjhaw4b8OSOk4CF9wy6LB0
Uw+CNUIAGnAGyoLZ/TradQ2LLYIf17D/8SCGzPRtF42/EElbbzg6V2MUgQGqX9PT
ZvFhLbTri7m8rqKAFVXx03uD07Qxg9ZhIXItza4BGjSarqYCEnD1BQ8nEjHFUl8E
Etm9Ba6KBpn8MLr1lQF2Qu75iHGuc7GHHS46LuxleesKhMJl8S3wyh1aZ4BMMMDx
WOOhskhZewMmPgfavsVcq3oUl6js1HjaFaUBad3KF9R8zmtPAZlrFLNR3xjoE/30
Ci6Dwki1UYAOxGh7RzdGlGatouEZAtRmPXpRltRYV1MOEhg5Xal+UT4c/S1nge+H
zajUjuzdlIvSSEyMuQ00aIVsbapJ71hrJnSbo1ymVV+clDltFAN+2gGx7gmIfqVo
ifveC3SkuFqdQAL4oMR0LkxoxQ3C7AlRHS91oCfjNVm2g85OtTlaRIvuaoaFRHzH
Cz9KF+QQqyH2Ty9xLm7d4XQHPk9NtLBoAMaCVV9XgTn8j5OgFiL8v4ibkUD7npbS
Tpmrtrr3PhZdpDYyJIfkodTdgWSJEKK356enMgCcLzvD7uqLPQBs/LM3pGwtXhdP
OlCpisVwcd3XC+A1cVGIliuS2N3VSBG7naz7RVoUFCpuTOY76uPw4btvSMTghk/n
E5LvUv14BxodMNKE1zdgLius+dkgcyxD0zsIp4YAkg0MUpZFq4cdiiInP8sAXLwg
iyoAc9a54nULe1NTL9ix0vyQcz8WanT20IGezDgNYd7WLyQwoqGeerUD8l66OjGk
xK4UeYZRxjLkjGnAyEyLbRyrgigjYzTS8quWY/1jgtTF+yTTXQl4At/rWKTsBeeC
VvjWOmZX4o60IQqT2NxA3lPG3FwfqKNGPQ7tes6V7yjbV5SYeLtnDTR8E7gWmJSb
3+qv+6p/G4/sNQfeqBE1RKVWEyQ94dIAO8h+PQRH8IAjFJ29sFwHiY2/p8m5NfuT
tfjIatslD8lCiRtsN1SzsH1ealmbdfgXGlZB+r5z4gi/QMOZgxxQwnEDSMW44SoT
1PaX2LSjDAXov8J7/h7RcTd4+iuVKdrI+Z20ITiCYFTtD3zubd+h+sKk/lDY/Grk
GCCUtTPgwQcuhbDQSse1/2goY/+UFpO3kmjSG/doE3AZ32o5JslB1ouARSiDwjMd
FPgkJ1fZiYr+TGwU3pU5ZFS1E61gNLwVOJo7b+KF4uX7QBU/FrDg2C8LpeBUlWx3
k5LVrgo2J+tfkDjPCrRWhCAckDXwTebvi50Ps96Sr/D14BFYSs/K0JwqJOTv4onD
QNrAC1CQsXvZKsChLiA+W8nuYCVP516J7CWXpKYM7rihGRiVjDOBDKBUOeHOpvqG
7EMiu+tMhUZpxswe1D+YCvuKCZeZ/9q7McOnM2HVnwVikHN41mXMm/UZQgYjQrTf
uo5d9L0jO2d+vvGZAKtjxhNIl/GJbMRKKDt62GWqjizNaTql9dwLvkuBH3HZean6
+oQwht8sAS3O3XI0/X8chEZPe84+cKtIoGPcymX1mMfs1y08vKckryA01nPv6Djs
E2ainM+ig6/SuuPDQvzx+7be6kDJ2YPuWLxPo/k76DlezC+0bSQtSi3NypiAYM8G
/ztFZpm4afXtx6DAyffESwExbHnevwfDI2W0tf6iBBS2JVzZ2XKrKxRFhqTmivZ4
0tIifAggOJQbnynAWw3n8sx6huvT0lBN9ZKnlpJgzKq4XLNHWwd3KxZJOUXnEVqn
lJscggPQ1VS0wqWCK/+BisJqWFfxwI7gk96pTUmQqh2+Pjd6/qINxflNgPHMqjrw
uewpNPgwHugxCGZHUXgQ0ouMlHuiOSJ+xPGxVDQOUsTnEEbFQbn7no/cVnLZyLz8
5E4ZI2elt7cPXRbEhWzXjQE5dYdnEvmQiWTSyzkiZ7gHkLFXL9m93TkHWLCYry/6
uufz0Y57ID2m5oOth9naxkI2MP5W2Ph2qY81KmobbLb1wU/59EOBH9dwn0U0Qyac
JbbtCqLKNqqK0v2DbJK+6EVbvZ0hk8RZi8d3liaQSRn6MbG71V0ywuOgRX1vwxQ3
X11qnE+84CLsINYWiDeccIb5kqJ1qQv1ZJJJHxFuIzOgcUMykWVKIRIkG/gFVTwJ
EEnAJV5KaeHw9Wy7C/ZkgZAvs37FI+aNsdn0mTfK5zZl6PGGlA9oPVbwseCVYRvI
BYOsVqipcs7u1AuDZpzNIp/gbMAQJbEn1xW/+DIHoH5bAd9uFv438l4adqz4UsOm
HFms4jmAYNVWQjmQ+uR82OqjEdONhJHrHtG/agA8XDEWiDFgZ7ZZ5VEakposcYu4
gwYBo2hfTXjG8FfCFXTnjOVAlJvG+JKOoMg7Uzm5fR1rhgiHhRW09+gI1ik9kaQC
AA0mN40wQBWkOO2XCSvKXGvnGCa5/ZEJJYQO8Kugw0ml86oDNxXMntIqkRAhsP1G
j5jdDr1vW8lP+k3y6QqVNcf8iq0w++dwm2kHC/g7QyBuj6PRsTDm/j/PK+K5u1M+
JuDgFP/fW66WGENsl19WDDTSg7AEPBCVjME3Rpk83ayK0rB8vc/rHNQnTRS3jYPd
fMxqKwz4v6rZYkAfzHMcwYKNA5HyvtZRIHJoemXHF4awlT6nPq7l2yR3omwzdKpC
ujYL0ACBd8/aSCxwAxr4lKpKlOGDkXoABIhwWw9vPCsEjHrtYTajbj8NhpCJ6ExN
Cam4vw1aW6MI2KYyaKseLCtN4bYzv7BWNJQccdeaJbLcs0s4G80qXTlb/xjQOCei
UxLNNxpJP9n8gQwqMCiaf/2GMK0MzW2OenKHocx2GIVZ8XPByTfR1VQ1I/S+uH/4
LinoSo6BIsSBTFAzRx83mw5Ifneq4j8ksqG7RveQkHD7W3zYyM7CKsDcYiDmcGjg
lgCpyzRTlHbHLDfrISgM9sofMZAL9O3NMNUhK7TM1+Un3TeZc3KQHLGNSH7M92R3
YNKnYr9d0URaUKv4yRB8lakxcNYhcJsSgRKm1db8yFJ2C9ibGFiIQ7od5gC2XfjO
Mi6Nehe5Qrn7MZr3Zl02UusA4mNumkn/6oue7mHR25ltanaPv11oOOlHni+n3iqn
ZgViArY7uvbPuAYyc+TJMJR8+wuWoJoDdIg4enq1pKroQurilgUyv/yT0cKRJFm+
XlmUeqAol2eKtASwOW8zzc9sVsPgu4PUCYZbRrFZBS0eqJXOOoncmNNHqmvWDYab
mnhkkGIUE+EU3bpr3hEKtK8hoQivEcl60q8m6g7FKpyqFR5qbtEvakRKP6dIuUpN
Wakwu94MyQ060JA9wdLmKUY3+Xfjqw3Ja6dqwW+AFlGFLZeDbmQysJE/PqVRrZz2
Ite+NgnRgUGv1kAokqcwaQqq9I4cw4ATnigF3V5TqmEWdB4QT/ssVxk0nLqFYqW/
vwZiKIjGKJJx38E7Eh9KxoLnL5qKfIUOQLn8pBf0jb260G09uzYaNgHzozo7AuyR
fcieDzqWvz3w/zQWTWa9+y7X+e4hBqs7MUyd9W+CxV56HQgfbzJvCtP9dWO8015a
uKQk2tOJKhsdQaB/aHdZTdHlczK+R+ePQiCeQ8VANcX40MyuTSu6N8YYarC++tr/
GCQ6+9M5eWvj5YmQ2EfBOoKC7u+uMlmnt2A0cgtnQ4qqgBXDInbjsY1uqpe2U/qr
5KHsLTlJUaUqxvas+NQ2XP0PLA2dutk5wxfS7b0x8rlVm/CCzLYKgT1tPyxtOBoz
JD8pFhqbNlL607Tnho7U8AFyWdBRpz+v/riAZ6SHrYXP1Qtghu28SPz8lHWK7ccH
3lxzeFNo8a2mMBCws2SSWotNM3Af09Dzp400fijiqJcJG13a92NVl0t1w1SSh+3j
8KKN/NoYLlBFIFYycCmo+81rOp8xYb1EU0IEmxGV+EEWvcZsBmc4zAA9uy3GnyxM
GhLP3a1FFZzPxM7c+66Gvm2rj9IHFLocB0u1dGHnuRVdP9VF8vfcCaoBCtj+SVvl
K47y3ksZmgsH3dfua/GEGIsBGu1kZXsxXJWfOh4fJd1IYg9efEfR+nCOAS4RnAF+
1J+29Vi32zOziOKHIGIczyhIWAvIyjOANBVGAsX+4/RrWU2NHyDe3JmhrVDhva9g
FgiRopwkHgnepVvi2zEXYRc9GoGcyJ3vHDz0Bhku6XBgSIdLg5BOshgAndXfivkE
8x58jCD784LWIOa+kn9+FhW6w6KXl7AHYdNg68KHUgrHizsJVq2KBXvgspF3Xy0R
U5GioX8Vwif5uS/OHQ3SSCRm/+yMayJvYUJintaavrylV//jtI3knLqvVJQ0p2M7
KZgrvW2sCSNDKceZP4tNG9Uz0hIoyz7o0qiq6DrfT8jA/Wq+2lrjBBQllYSsSJpj
uvDGxX5ibukFPHsxceGJstwztfOUGus8rp9LpiBmIrpHGwjORFU/jjViHhaNmPlq
OoYri/Hj9+FMO8cFwP2VhGiUROCTmg/rl7QqUQnBl/iam4PJepiyAw3kiV18faIl
x4YoYAuzGpxRbibbo2IbmSkNrMK8Qknbo3Xy5K9PojCjFrZFT4iJVu6kKsdQndDX
DJwxQfVaX6QRspLau3JwzM4ZcMbLsJEpxybDOwDhwbsT5kEHaSKIPzlEqyo99Nac
nFar7NVeY/rCAtOtcWTQACe0hk7dluKTEeDuEPVnijK1FwaTfbWhP4EtVc4aPFMk
+iWEvSDGml1dEFXSKHDFrk7NySJ3O5aiYJaJAzhV8I54fVp3cVGFuGeQC9YcgDCV
7Jyttio710fulhLSflw+D1TcmWvJpx82j5SqxUKsGCkF9oYYdhMoapnilj224Rnl
dMleRQ43ciBnDRAE7mAVfs84jOj+VIkxnDljf7wg9nohjNdb/zhDPiHlhxrSOSBo
gGNBLQHMcxgAdfkXXXktaIbWEpTaoVaiRbq4o7DbeniTQ3ukqnl/aPNPchMPyhqI
q+bERoHd3R36OJLQ9IvDX6qIsySJyiQRf22sSId2EM/rR1u0Jr+Bn9+WUA4FjRn2
HwPY1blYyn4BZ7sBNGrUPOo9cVcTmQhaYXXzx+YVCKjOVqpEDb/zT42e8ircCCxs
40Eth2uWUa+So2g+4oiEg8BA2xhKelO1MluvXotpqh9qLJFOvfMGycu442hvCIE7
xAq9wDJfiOj4VHqwgCGciqNVYx/Yv6tvGrMhkGHV+ug6YHtwsEnX76NfH8q7eXE6
YnMd0NZN8Cns7vm1R8wjw46O+AWbWREY2LgN2LQk4lB0z2MsbPR2AVmxYjW3MHyo
amKqOBENZWzuGjo0MIk58OfjBIM5d29O7MrVK1D2O5YMM0RX2/na0NX0w4tzZN4+
HRm1WuFB/RHvBJ6U9FhvhRpkSMc8PTI5HsnTUQ9k3+/JA/3UZuSkJ1rLC7MormI1
pMTHhoaxj9bCTxbFgnD9Mr47KOoJI8LXujcdMGiIKVQf1i7du4coogtcameAPq+E
15QIKVgAl9YCiS1koAYwMejGCW81FNCyH560GKThBO5+AgR8U/5amyJg1Fzuvbw7
8957KhrtBJALR/wOP/mpgmMayZHS9WREID6/ahuwpXzBM6ATnGvwKMdHx0qVYABa
c6sGtHIpVwbNlXz8FwU0rZFNLKjX6RFgKlf9/LGoxYD0EAOKUBnPihaqQ+43szAX
dl9bJlStZEfZuxRhWaMMh5NdTZAMrJ9yvH4UxXIFN/7f+Y+Byz3EO55xga5AOpnI
XvugrZXUsJtUPiSooONc8h3xIyZmd8X0Dux+KWROFsnosuX6+1sK/XRx860I4Hwc
fZkIH8qBY9mnY+QCCn9oYPX0OjRX2XOJIwpEoD67kMJYt4qJj4ZM1VW4GVR1+hqV
qIvkeNK15ZAnJiOq7htcSuIsD5jZ8mx4rG16V2r/BMfafyT87K5WdIyAm/AlSWGW
V6wm7CWu53pF7PmEk3OUAh3na0Pg/J0QsXwRDo+42fV5zKZberJekYRprd6v61LC
dotW2w0Tp8zJVzcc2yO9HXnDlDQGRD/iQVVS1cpelQ6oaHHfIl+GOggO/m8Rx8E2
f0FqGuN2jqh1ftpqhDkMeyIegVMBlRELc9eKgTFQxlNOG5s1MBi0r0hptCd24Xob
yaDsHnRJi3CSafbhDHpkeiI4hCycBV/clzj2svcFcQp6To8Vo92U3DD7Jw5oCb3x
axw2ZRi8Wplo4u8HszUR48KajbEpVgYDd4DchxTm74M28+3A3bc8bAXtZ6kPlLTD
Kap7+oJfc+Um/Tr7H7MortJBpyHpxMS9ywsDe2t1q64LnTWpHoBFhskI//0+jL3t
ZAr5xLNF2LXp5AKxHg/ByKAsQyAFZyLXxBCTkehnTv6UYFSrc8I9y2/5zqisiLg5
EXV0iPXzzzsp1lAdVR7BlNKizlhxeYlmbJtIwprCvPyEvUybjUDtTiwhEB0b6cVi
D/d1dhpj+ppbIOKfKl+n2VccbFP151mVh2yUEE5IspwD8E0YSsRXAbgO7oYLA2dG
sWV/RHsAxkgQ9Ro9FRJ2fgtGJIv6YYuslvTaZ/FIlmzahiDFGv9YRrHhtoCA7Dc1
bFxUe69Xu07KLvVisgK9Rj6yDNH4kW8ab62s+kudKJ8Rq/aGBC/r5qaM6N5eGXEf
PwIYXJreRKGoJeL9cg1DCGbn2izTt2tYJJQVi+R0YpKseFSEENWd4n7ugSuu2sH7
UC012wu11TZ5kY//7Tt/lTtXwbGsJ3e143ukj8on6nlL19eZgwxPHcOHoZqwY9ES
epxSNTbO8r/IJHgK1jny92MhRjpWuMZHPIg/um9YHhC966bZJXj4CxLGKyEZn0lH
ZuF6lnZYWVCPirlY3AIKc2O6suljAzyzooi1bbcS4/amN3CDhIUfD5ZY+6Yo4RhM
W2in+8+2xby1lYgkNCABrZIcLLQmo+hHKcmnhYP3qhA9wNIEm7/tj41dqBMVC9Q3
egmoNxbuAGpCOaRwYoqLu572oyJO84yznD7Yyid1G8nCljOnNQjkFhFJxVFvfAnh
IB3NgATRh73NVHnKwfmtPXVmA5tXsF6hUEstlBxFKatPMj/t6XDSmdesfToj9RyW
WeDhgWzXtVq6xXMOKTKyredTUsFP7DrVLz6B87G00361g43lXIUOOnrj0IvGFqS5
GeEqZvJqoS6ZFiUZptVYeOXdav2g2T5c6UVn826SRJ7htcZ5GMGmXSxvorTg6R2g
UOYhyHOlU+aYKn43vwmXOQqpgfwfC3R7deH8EhptHQiQkpu6wL8ROGwqHDERl1rf
piHcCh/9umDCNt+c+Hdcu80/CuUP4Zh6JqFAynBstPexdff3lOXbHA8ZBFRBnbBy
rvIbCKy5W96OGuJXfDCpZ7vAbnTdEvGvAiyDeiDktgH7AF2sX5XTAA/ZfQ0cz3yc
PqlSAMJBYz24VtofUVHoPMWJbgePcs6pkTN5xzKH0nx2dwASOipoUD50GoY/frgr
KEpbZJGxXdrQ2FGycZAhHHgvf8CFkfGsecS8OT0/W9f5uLF8Pk1cEgtjZ3JMut8A
gdlYFiqJuAG0WEkVvsIuzUttYM9RCIR8d/Bylv8JiDX6KezxCPdZY/jBpaGzc64k
nnrZEuVaDpDol3VUS3KtVeSKtdVgkQwhLNS4rTU86JTtFceG2FYA8C6IxfPnjxkx
MjpKMUSmqKWyg2i+lDfaxB/drN4UGRt/T9cAn/S24v+PGp3QbJSmHDlD5Gc5dZq9
632HKEg7jAFrsJGmIjX1sSvCSVzHtTOcd1SJo11jfNQvH/hkC4P5DviT3uec0AgU
drH4Xq8ZyjCehh3VHCTaZuoMfj0k1Dn25maStNYZ8eqV66anfEWqbZdr6nFiA6XN
ZgRZONVnbItnVJfXDHhVEfwqKi9Ed14N2heyvIdbdFhQtwF3al2Yq3zvxdr9h2SM
t2piL0g0oTFCf90mVRItcJwOGHgUz8BAWcnZrnO820z7YWJSGHuoq5LKWEyKOf1/
ZyUgq7FqyP2GZYwAAiHfvNKaMr2gcR/8PSkJTLUhqSb6cWfPB87v+pbHPDVCCe3q
7qP6UiQp3wi7sXYHkDJRGfq9MXSjJGLnBcbMePdGhfPnz1F+ff7oevQhCk3Mn6tj
tkQjJcvsD1VjOj8AnbZ5K9uxM0Ok5AAsKteeKItE+kP2Xt2kLTbFmIBCH7BN3G9r
YGqYaN/5qP4af6ljlAoa0Gm7PgEqjEGYX4qReW09LrkzTyDdOaGICtUra6JI6es+
j/F0GnadzjvxLvoadFjoUEFAk2wPmVnMFkVAlahlDMfUswJPV+qiwEmr012VFGds
v/k4NjU0jJ2h31jf7+uBcYWjpjzsG8honyHrPJeSqpE4UcLa+N0y7yupTLph6r7j
ogDmPxfsghtT3m7vhGiw4C1eVMNT+vPPX5fy+HCsNOc/NG5gjcxQrkLA25WnWzB3
5vyb962J4wpuPOSqZSTqxn1qoDlaCs0pdVrFMXkHCX0wymwiYt6rHUsBUGkjlV/4
/4uSIoXPSwoIJsYvDsvgOvF7ky6DFq5usknirhNcxbz8IsQcTrt2gZTW9Nwq91oe
VBVczewBZEHt09PTxMzAzYGC04EBBiCm9tvEFsiap3rfO7rVBSMQoHITjUYH2HfM
HAOC+J1eJXSpMsgkKzw0BHe/p/V6HaYi2ZanFcu1LU9LhxvuweQhTcPqzzR0Byqd
SAgJKFbUtqUOOAiQ4tLCCnMrlPYHtlsjsAZOtQtO1wgSiU4qto2J7z+WUGiEDSoW
1g8CTJuQOMPcRYoSQJTURVs4ZDW9t12GuIsoKRiPyJtHz0D5EmDgLdd1s+w/FWjR
KLaNPrjsZEBbd2Mom754ExwuM9e+Jc/n/96bEc2ZQllYyXufAQWKQuoDdbBXCQRH
MWapX50r7bEAW/ybJRoDKab6S2VfpN5wHyNCr00HespCfewNbpzYHOKOx9Dax7Eo
YY8CCymkHINwfgJiLtasA//gsH+lFsLfk9pPw1MLnm5f66rW8Za4BhkInwEZbvgI
LnlgskfIcbX7RMOCBWqDHfNulGZNf4F+KYiJ/L0O/5iAxRNbWojHjE5il8XjMePU
UkeZm5INzzBIB/xNogLC4RPfjSinJqUZNKrkGZ8zIHvImayZeKOIMtpYMqjE9TuP
A9D1W38Z9hko/mm5bWxcu8JtrmpMnDPK45Vsj7KJlbyJ9MNrKPDnFS4srFlJx245
5yUBob4S/yrO26lSZerr0RRK4ksETGzv4PM8rMqPh48SBzEJOZQ2wQ9SpWRt1zVH
cSg5hsx9AHtu++77t/h6Fk5pjlCw8tJXjta7+9fR0gbAt1BV5wIR8TT6pik5CNFF
/gimIzVzlISudI358sRCXhzHjRB/LxmHqbh0HiXUfPIEb3OEX2GEnK3MurSAXw9Q
xNvOTtHcfto4zMgRQXmh8LZJkxKzVjnRJfzPJVzYjVY2rqZTM0AxSZeNYLctPku8
PlTbFpJx9w87JuP29T47vFbCrurYak4vqkY1OMe217g6SOnhJWQcUGKGboUFByCe
oqchMBLkVsa4A0+8beSdCPvQr4nZ2r3y1fierpOtzVSv2MtkmryjKcqGnzSoNUOa
c8BZZULdX3Zqd+WRnyfHSAlgG94cpM4AVRadP79YQ89j8AVpKbwvzyPW2sCirpTU
4/ehC11JdYRF1sxzuVAtNtBbP1IuutX4lN/ft6UmLJhsAzGmKT6S9D5ItCOFCSab
ctFyDzhYwIInr51HKaAMmdc8mETblT3bCVaCZLPU626Qmg0Loxn789eOqJifJSmM
iASOj5R/iclZ/dR540kKAoY0Lz0maXwgovTtvSRa+TQ/WoWRaqsDv45nbOYWG1LT
tc3RRkETD993Ka9v1MBWox8Fvx8PzOEHWM28cz+1BmREkVLcUE2IUg1zY19+m08V
V+5ZBMScTrZ1FQdiIL4HDsglifFmVeVyH1wiqWeSS8RUTpQCagUllUuEKietndoV
qpW1wzbeZSc/8cYbNbiV5qj5WcYz11l7Otc21Ffkyh1MWgR4E6O4My621FPE2vb+
kt8Ns3ysJqVuapvP0vFxUKvl9ctvRaEbb8uYALMhcOLEGO3HHP/psWrjHPh8ecHG
HyfrZSzOW78tr3Ixtb5tuNRdHcI7vLDlL2xrumrhFMIshnu7mqvmyH9cOTNg6IKW
RN2wcmiVJjHjD2wd+LBI0SbatBvWMR1YZxyHSdnnu6KAKPp7vYnxFVY6SqsuG8T0
FwA0LJ9Z8VCS4Zkcq75NeKRZxtcqknYT9qKzLVyuTFoGqOX+0JZWsQFjv8ex9s06
6DaTRFru5iegKkGSYKkqxMqbfUSvgpPY9PKkZEYDqL+Wc/wDYv5LHo8QGjNZ/h8p
jl2Y+5hfulTMBo2io+gtO2iecXUjQ9b4zxQYoFHXBGIjQdT9tmxYjcxNQlw8oirh
NapX+d3K+xgJF48Wg5/w5cxdAPm7YBKe3seMdfw0y8/oR2OW7X2+KRLHrzwDsn+p
lkXWSFzDzFFmZEnTAknLk4AWoBymYNctDQhngkfFXTD0hovYMCPkmNys9vs+1LHP
vBzye0TTehoCi5lNgk08FUKvV886PRZrY9pmZpKxIFHhBKEkUk7QpK3AG9NfoISp
G7f8YjYlwCh8sTZ3Nf5pmkAy1NYjtSSNOs+H21sckenye0XeH9JWrmrMwZEhOoeR
RuR4HKbYaUzOphITksr/+21hkEODrGryKTkYnOhiqj3mv771a9Zw6QdJlekbemAq
sIOZ8YJPSdefwqsD4qRAniFnY0DASKZSb0XBRf1YcJ1L5V7M3PWZRcZUY4NmwMAI
cB224jcLNyvOQID+fjLQ/fGxN2QiSfLI/F6qqhJWpdL2rJdXNq98fsf02DrO1UsO
ZgYD71lW6Ti01/WG4O73YG8/s30ga7bA5beN8yq3dvpomP3zqa0bcOfMwGIR+QCU
FW3e35MD8DhDIBz1MuEEBSbfvH+a5mxP9EiNsPonWCt+WQPcF3Kmkb/stCY4UxoT
f5EPjPBxtc3X2DYsiPFachekhrMGGiHB0zFu4ejTgKuglftjAehy5Qvw24hUWowJ
g42UZ4wVMTD5CAia+5XwqldYNdiZtB92JMY4j0sFO6HAP4duMCIfObH3DPWQ70DL
JFlPb9nWpyCQe+HVKu7L3WG8sPJoBvI1AZYthCwL/KOGixmurcG+BLl+TU5RRiAn
QZMAIy6FW9VBKtq8tlIB3TLjBkD2GrWNhRC4Y663oFAgTBWJFY+vsWSUGXjdjzas
KnuWXvCG/BSSd9fLl0Yy/Uug42f/c/GqIxbCmaDvRke/24yVItax2IkZuw3UaYaq
q5NDi6XrrjKBXS2wViDRprGIf3PtMlKeNSyErISr/al16C472/+m3SMf8cTPqpoB
rcXb+x+TGjQF6VZ53uCtyKhBt4eASncukP8n+Z9TkGsTkMkX79aW8P/7UaHp2Mbn
qQS8qaanudPZiQDE8ae8hHrP5QZFkfE2p71xna5TY5HgWO+13nwLlgltlS8g+ayf
VTbLD0fkTWVoe7vdJOga6JQds7uEtzb8JDEFYWSgnEIlBxl6ml81ErlvDt90UtjE
+MxlIUd3WIzCORVTtqXRZlK2eBc48NePUCDdcZ5XRucIUzEajQYyJCbQPggtMd2i
2P1Ti7Kia1NhnRZPp7R3g9ruIhk1IbSiOfbJrfFV1OCck5W5E5OjjqOOvb785ubM
cR3Vbmh6LLRP4dWvQl8QCqG8vfGOuMk905H/LP2q3nwPlPtb7NmtTrHQ9y51Ktb4
ywYJm1xq2beWZu9JPmZWGaYfitwXoJXjO3nf4TxDmITUA2dyIC6XTDzvC/CvjqyG
pV7Rgxj9YR0tS//a2XXYET+ExrkHro09RPpOz+xUtQnVpziAcH9nJh2236e0TDXD
roF1PzMPSGcyJjtbcmnGPLZvJW9+VYKfOgKPc5GnOV1IguOqqsFOK0hNqnE4dVov
LVaghFg7R2hO1USNcZdiCUxk7ZqIHpIEkHmtzSrLEF+G34F24u5Q5HG3httHvPSF
/YQz9qeejlutzSlWEN+l8Ic7VOVW5AOYDMlCkV/a6ZEs2WTscYILMjiobRl2O7Bi
nq4mf3Oy7rFIPTN05/lWPpOw8o1AL6z+tIiFYuAxwpE9oGrlvnaeY6UWi077G+dk
j0fSmXtkxV8KslfHYOUCQwp8duRJJkfg9niPxRKrVRNjNFR9sP/t/PqnI5h1iko3
Al5c2mNHia6Q1F9zE/do381X1gggK3WYE9ntZblS7KLTb+bgZdzXjK3fGn90FDr1
aluou3Qdapz1tcAFpWlrC1W+aLPxFUQ7NNwoILsVlFGWMcez3UlpIi8jLDzG4FZ0
m78tUaK2dF6PEh0OvX23DwdvYgeaSl0OBhmX/YPyY/tzAZVIZQ7PJzKk1aM46lzr
xj920c1rp1DSJ4N4nHDbDom8J155HRmNOEboPbozam6jPOkL1178zarUbxYD6zDS
WcKBiH7CwuwMxY5/NpeUxkNRKCL8XsazEmeMD9zF06K5IeA3DQwPAyzR+VMatJ/X
GTLODmhT6208bqctmGegvZUW00pViSw55S4CdKjcvy5GIDRdcDsFfj81k5uNOWLP
iSWH3YEdzq+/tr3+KFR7uPDINy1ckPSpexcSBsReBhhBjArmMfOCV22e3Uc0Tg5P
HqKUKsUsWriwwLNZHEc+bigicl3/uJIw0JRBIVLQEmW1O8J79o+P17DeDjuqebkL
c/8Yuk+TPXh/xdSP0Yw5unmsny0kXODPv0BuRTiypLNoYOxkAsDlRSYRlIr4ggAH
7byahYE5Ep/2uQBOzd9YKfUvR01mKl+aMWdFkwdaYuXZPBTZGJXdV/ztAOMX/6zc
u6ujUB8ka6avrKdpdr23mW4VN+lRK70RNzaTUU6rdbZeIUrtRW8P/7ZmWhj7CitH
zwkHw7R6354uLEhSlTTHCE9QLmKYYjTvLvckUUzo7U6oK3cYfkS6ZTWC7DfxbMCi
s8EIWr1VmrAgTEVaOnYyGKwnqBV9sGuD2/ce3wvqxKwtCy4mDsKsuhdtQryGgiBB
/PBjEUSd3G6aoXmpnYEzZLCiijxkSp3WTfZA5v3n9VISO4FI8RzfLIRIBk/68MDI
hez5Q+98HuKA1OhLYkTXa9stMZa9jTiutNijN0b7ClUhs6OrGaFNSbK6W+JsiGw3
rDnhHCMjhtv20BP2gyiITCeV84UWjAcTZ1BIa2/MSDxY3zYXui8sA1cfWG7K1Bi8
+R8ErUWDMrOPqKW37cd5TH+EXF227iWWLN7imyKv1eAI/hmbKbrmQTA+K74Z3dEi
4jjGBTZH0smrAP8//ed1G8nJOPQ6T60lAauQN2lvOZ0HGqL30yaDynaJHVoMi99h
DKRrFNHakA0qIJoOVP429/NCIokNYY4Me3qAoMNSj+I7AY7YCTULEfsOoM15Q0bo
kMgI7gZF6rZc/QbAdoWkw347WnwslVjrHkPqgEeQ9/LdoMRVhCRQbmguFOZlHllQ
NQD1fRzyb2A4U2llS6FgWxkNkSg+aBEB52xcE10Mu4gOkcZWDMrsuuUcPcE2NPnG
8eKZJl8tcvyy+p1Mi4oqhOtd9dNDqQOVk2jBIs95vrF6YDL1ARUsGmqTv6a38VPA
4xBqrnwhWXvvnUiZASXVzkzwB1/92yordTzB6v7pc8Z65k0vcPV5fi3eYzE5awWI
6hoExcBTpQNrKULEg4NNgbVKHAdsC0Iay9X08zBDPCwLqS+qokkcgTIBBYluvL97
Qe9CUPV7l9oxr9ucLYCxg+J4h2GmHOZ487Xm47eM2xfRPB5nOoK2rlD7SdMMSieA
jHXbLmGe93s1J3wv81j3Zk3taHTZ13MJ0NBuSFI5czIXMl9C9A2Qc2u0j+ReDTuc
PSg20heCb+UhUHt/qGfq2G2O6e/y7MYlWWDZ1I+CpSiUdjqhXCUqcqDJURiBDqt6
kNBY3kZvbskj/QC8aX9L0zSYFIe67H5M4D+NZQFfoQdm3AqDJNa1ecxFJvoY7kmI
5AZVVwuAa5H6GAOsGCFYjHCxeoKHCfj4HPJp4XdkjpR+fyF6P9H4aIawTbdkP+5a
TH90UpiNYBM2ZN6tCSkYmuRryL3X+IcSHlkQJ/gBywRELLXq5nyKnWuTkFJ83Q3v
+PibvzfJbfak1pEx1LSWmt/M50IBN8eflgK+5nE1T1tAb4dTmar8G3rD5jz23s2y
G6K/wUP3uGzRiHvrscatrzyIHBePe5zvZl66Ew+wbE80zlg5jSkIMJDg3TEYZJPS
dkwAKHM3xNl1Wi0DwQ43arDmEbSbpVCQK+6Qdf6hYjfOEDkCWB8g9PSqU9qlQN+T
7OM9e7VBRa9EVGGONGfSRZuGLKasw9q3WljTb9e2KS92gsJOR8fu+fxVzgi6vyRY
nqsENpSsRx0c+4BcLwZcPcTJVTpDSgKsV8pxZHBtczzi76lmG02z3b+Ohc3eTRaY
9gFfZ/XGtiOwPHWC7A2540m1HOQ1j+cDadbvTmVtR/vBpMOXBUJ1i0JgcNXROAek
unLvK54OBW4HAUdmM1mhxhu34lPteDhgaxOFl9lxVQbQhE1911lKaILkODoFjefJ
GjaSndn4E3NH8sxGB3VPsXgVKWyTHBtz4sZttBqiDTjgipuHLCZlK2JmeLuUwpoQ
ptTRQo76zIsO7ojTWukJGrg+OBqCJfOeJYuURDBeg2pqWl3e8oGcwFyy0P2fslU4
J217GvEm3mFL45No4TqhZG5Owd9DEFj6kKhT5Km28QyCOXbFYwrXNj9PHWdy9vfZ
qOKjVE7f4RaHyvmQYQ+4HF3zajCa77VhW4RgA/1pgoZkl1vABRlet9R/+LKYS00H
cesWE/zQTTcFId6ScbF/tUEQX85K8/7J0X+myUIS0SR2ycMn3sPRajTXwHP6bNcr
4K+kdulHk5u4c5j0lozQJeYghsIvSthUMyJJeRmQjNEQroEb4m2vlUj8WrUQqysp
viicENswjGSWyzh6TL29vgxKQ4vE1ojcMfU5iNyRtBawZjjV5XWxo6olk+5ANtiS
eLyP6JrSOhwpzU8ZCSyf1DkoWqawusm3VMFlbHZEWkfZomg5PfbT8XDr6DIidkqP
PfkaxUSq779eCNb/R3nOB91miTIzth88JHkIfDPgS50KNgJUJUUrBtEjntVnw7Q2
hyzQQ0IOxGhlbfVJ1VE7tKbZ5xgKshAJGEOxzNrzNNjd34k+WTEhosZvuNMvSdN2
L4AeeJIuQXrLPjIwWHc+xYIj3YuvahKfPzgYJxXGG0auqhwMT7rfWWi8NHOcIERx
cW3kom1fbVHiHk2dAT895XoBn8mUqtpVZ9GnzB+zzBFxtCzlCmHSSWmBsXpGD2RG
qC3vim+OpIO3uLiX6arGqwNdn0zfsjQwBYhOV1z8lwvfapBCzMbkwD3RX2aZ9sV/
xoQN7KF+dInBkXvSbMrvOn1apMB9H9gAVs8eBgSAv2Q2q2647DtWS1RV90FTPkO0
QMDz36k8OwR/eZ3THQLpieA0CBcbxM1uAtDvEnYeHwpnE8c+XKS5Zr5m3U5HD3xZ
3CCHsEUFooDEK735nxIrjMqDlg1avMGPFsshu8jvECk/M6yRlpG7cEcmwNSNnA3F
gl2JrztTIawzqrNqtK5A4U3O4bWQoI7AxW4/NeJs6ZLRyCVdVSNqmLhZA3CPemaX
BVyfB2vy4x32Bj7ivb0tMMpC9Ht3M0hVP3buRQb+z1HEvgr6jEnjeJ8Fv+bupa29
fSNhSWeG6BBzo/W69b8sdud8HNLN6U3fgUkN2alNieVkNGD4B9nNGL9GJph/sV1V
K0Wv++Bbh4Hsu9R2k2GsBMLhEQHIfhDF8JfrXx/RSdnMQnTld6MqQtDr1q+Yl59G
/PhPYUAKqd6N7R/GYM+5x8AUBai/0Ni05SlE1rM+cchJQHAXoOB1bwnxweHNBewK
QW/+8YGz343MROULRvjGuGn1lhMJclrPPy6imGN0cgiwKJYxihYwIxSbHsd2eo0B
JRnxVJffN/OFoKzVdBUlqF8Q/67yorlcRjJ2EH5rK3flgWoReBRyxVI+FXHTfPNP
JyLB/woaeZX5+hbB+zTyvKQDYawPUI6NIkANlrXt+xdHbTGb7DU0TN7iWt5BPEy8
CkCWPvzwe93tPv8mLErflys5ZKaMpgz479BFv6g9j1FXc0x7hpxfENdJGnSuR9ZQ
E8hffZC2Pxeo4wB3pVN/gp9DADH0Fvhf/8exlQH6MErR88hk9R6TWZz77UtLb0Xq
MU5eWDXwSop5x9v810FJ08Xz7MRt6mws6/VqPC+X8WI6I7ploxJWFA0fRuwbC6Zk
7DDkLdpvIHVSjLh7pq95+RtypNiX2exhPS+kg3KttFufBBFfP3yjQPR8WvKoCebP
RVorX8hafiKbGjmBI3iz/v4Gt7lUm8pUvgcXUrz5iTo/U5tCzhf181RTfqcPrHHJ
lpFebnlp9bTlRUuucKbnVZ6lEwbitbiMYoJ1DzgvZCR/gBpyvX3ZFrdIk2G8PtEW
1XE4fr4Bm2oXOlvh8n0hgoa+a/8IZN2wkFm3DLy3xLoPEMDSejAo85q8DOrUOEGF
iCFRd6ncN5Hp54P9myD2wgRRUZXznMXD+yu2ZCXsX2sJXAZ4c6MGY8fTbh0ak+L9
gp4N2hzWvOBf7DP4Cs7h4r6Kh+4mnecbS7NKc/70anJyWEz+VO2+oz1Cc9GqKJxO
DR6ygZ+dlDNtqFTqLra9t9gY3G/TRMPvAl7EchbY8ExxJLfAs5nXyodTUBHeee3C
72CcCXXdn55Am9WOyCBu+fkZDY3Jv8qmUIcn9qwn6+Fabp3lerPESyCPYcwtb751
i2qAp7btwBnN7kim9OQkBivd4Q39rGUsXZvLa4vgxSbvismqxLrfNIKfcE5RnHR3
DRchorBJaELjM1FckmQHXuOY4a9Pqw0vSiwZaRkrfXCQnb3vBiSCYiIqsT0WhIzK
f7RqIRh0qrvlQBrIRJD+AYwydiu+8NIiuAaB5AN93+2IDzLcuEt714Rz1Xww7qL6
a/el3xYAC/Ku5OgwElJv/TwjZv2sJElp1P+dyrw3fUrx2bnNQoDrVEWvh4SvEewE
59hhve4HKp8w3MkptxRtcD1HuK281KoFUqcDEva7QFv9z4A7QHU0FU0wC5ANupJ3
X1UPp/mfcI6rtbuLk0TPx1qwxKHFIGakblFgB/1Oo0pjz9vm4+7S4iFQYwFojSz3
DY/NcWWROpgjT0zSOvGd0LvwKeoDUy0tfaPHiObh+0zmpzVE5UXRpNykECE0p5YG
MslluL/xL3RwimxhjRcryW2eUNUGv52VaXjGrRe113cbhKR4NWAAYpRrfe6WFLDt
cpyh59wmDlsRKSnEnQa2coxsnmD+COd8E1mAzIZqW5Yu0nPqL7ALVyfdW6TZaV60
Pi3Su+xxsvGeoD3njNeKpjzYpWglPIDI4AlhofVysAI6ycRyxX4xTE4XkcBbMhfh
5VJ6fHdwSFPKrhm6oNn5W2cdvaBzMiSihgdpmEfiUTOQw1qnX10IcVIYDcbGM2y/
zuOq4R3cplTa1UjNSKbE9owRE5YoRZ9ie9cFFMejv4gjnOZFWDsNnFsZO/WYrTTV
AOTxGZllY8zZYrnVaKlB8IEVfCnGQJXN1V4nidi4SXzl/7xyorGVAoRn1qKs7PbT
iJ6ml27rQoRQd/O32YY1J8HW4ZECy6mMLFkWWX+vVM1e3hvkrC2VRCPV/EGwxuCe
47nBx1N49SrfHHF9iILTIwrQlnhXWzG/OBsmQ8jWplRewLrZkZWhj50KYmQgTW8x
1MlDOFzcakhduofNsCODBetprSdPRbPYX1YX8pyfF9yTQ6auMD8ueWPfYk2fCeIz
LXlnZlcJ062N8y+E/iqvtRbacgKWCaASWhPpRLP4aGlU1MtCOYFt55uOCDCjGJhw
Cj8znIa0domAILl2Z3UihK9O8bnN9Wc4DqtAaTDh7lmvHsFR97zpAzA7HhXNfqp3
j+Agm9+51e9x3Yuwl33AYoNjFhFS7ROzH+qIJFVoxlCghcdfm50B0xDLTbqc53/o
IpQgUUrTaiT1b0NYM/HNWiP6K4BwbGAgKeBT+SP6uNZmLScgx/Fjl6fw6C3VkCyF
QgftMqqjH9VNJfmPx83oxOFmrvb5JU2vDx88DjGAjJnuqyAVVIM81fb2MdXha7sP
+g07fHUyP3fmbD3p8+YnO5Y1XrlkX5GcvfKfXyMSEHUhe4iaghQCEhnHOE81Fjmh
lWl9/EtsRkDCe+iV+vFcEYkhEnm1SX7Q7ZCI/jhPmT6Cdh3Srvx4ilNd2Fa5GENd
5lSO4lrr98fsPwVD6baJQuQzvy8quBx3DkDBIcsovOyKRcVJESM2gOttnSt7Vsb5
68FM+vD0nhdoe2jDR48E9t9XUfmJ27I6iuWNmp61uFEEt6CnhlpyqhjA6UPuMabn
WrsxxPcV2urfryUM2pla1XH39NiPPII41f6a26vQQaFLT5kfdteB9SNxOx+37YBU
yW58JxqVI6nNDo0EaKzz67JSt3KiR42xU+uQzxRPt+Q7qkxFJ+rkMKe6VEFdlNNh
0o3PaBVdr6y+zk4kSDmxgA7g+apfBsBOtJG4O8X7wv2GED9nOBYLyNCVnMOfopB5
tSKMx6BhQ3m4mFmJCU23toFuHz1UAYX9iu04e0A8u5Az/AcKXjiXOV6ZQSZptSWg
d55SZGYCDUmSJcwCVRrlWM8gV2NKv7RVuW/oHtrALjEn+oK+V2J1AbblVnnlSosa
PhoMU34vHVA8cevBtq4bqugogL1R0BDb3r0Q0wM34e3OWO7dYdn117iP6Xg0rDrC
cX1TC9vHJTm93mNzjYIl8AaT7kUiT6Nrp3NEfNxAhG4GfyISeRDaPbkQYnI+NNLI
8KxEJ+gkppt6lN5nGKiEW+LfZUezC3pHKfABMkkf37/PIAKfL4Tay9SYzcW1d0Fj
fiAkAW+6xZgVjy02hQY7aO6p3uA/tlkk8RPc0QNB2du96omxxTlXI4/KobRL5ZG+
w765fe6DFAAQEMWX9DehFZFa//OjBVaSSpmJcaiueM15tVMBnE2TKOYsWKP/NX4M
jHk1qK+sj4BMr1zJI/FOHp1w7DWRnoVXZ8TbLoNFFnvvy4vBtGldTPlqTpmbcuxN
TpmAjK+Y2Ubm45UuehCdARjCIUp69Qtm7bqmn2cmZHyXhyE0TWF3Gk0XTxxsznJx
0/hVInOSQH9WL3XZ7+Et7SXzfUfhkXd2hp8i5JiK8WmdicxuVGAWb0BtQ39pF7UJ
fCzupNVx0FbM+W/wEaOVhpjSFZnuSkPo9semdJxPwHUtCjjoUOFFX9oimUzxQEl2
LaJOyPQBJbbAc/UOVB/eeOu9GC3ak5NxQ8TWT07vi/jjBsmLopDo6LN3wRno5Y4c
5Ub8VkLlXte4u7T37dSyh1T1mdCMvBBpKlySISCkXpvCCnDQUueUvr4t0rCx05q+
6sdvYFSLBKNRjpnDl6IRggZ4H6wzBuPowdN9gmrV5UIQRf+YyomY0UUqi3US8Paq
r54hWfSd1C9iiYfC/NyB1GTJrDs/cmL1QNZYckAM1/ckvjja9zQX4DtFkxaEoXGt
VCaJ2GcrF2aonGeRaL19A1BVimfNd1iv+Qib1kWzx749zNNY5SJe3ziqv94pRy04
LylaeMExU5OoNokmmSFWfXLYDFyvF46p2Pd9aNeHd1Rs3DmsrYrSGTqO94Vy2+Bn
pSdKhz69YI/8K54f4Iu1NTNeGNPMP3LWTa9njLRPRopVD4Vwt0Tp6VgHA++R8q44
2BaOpnk9wSzVqj0SfSPTspluy+ts8X0adJRbiM4tP6nYvekS2GdrHdppVGpdErUq
6uwT2EsmCY97FcBnzytfIzkDvM9ZS3jL8CS7mZ3pJwKhAuzYjRhYhIDSBsS0LDyF
gH2Fddr2O1chgBCo45Sm62FEedouVKEltBrJFlNeFkzIF2ZLxrLNoIc3C1d8xNmG
QyPMll+OP8IhUHpjoQf7KFdqOMrc85+oZVaC5MaHelvah3Szjhq8zFY8ui17bs2z
wAUbPmt3zkDEVdVEQgBHBNXp51/mz729DWm3u7REayXGwQAtYuDJvHCIj/ZHzo/r
4N55q837muH9E8hUBllCI17k4EU4l+d4WsoWQHbXQzzU9QXSobQ5DQ4j6jPoJicB
z5rZccffCFV9gTWUCQBQKPgMUO3JNc2iIhLTa1u2L4cRFfQXFS0dwUgRRCyE4sYy
ZjW8tENGCvcW5OXsY57UmZuZ1xe3j2rwXbAQQ2W72aaF5cUouPD0XwQQLrFndAZb
gMLHA42Z5gEx0jorXsktQ2PAk8o3YfqI3n1DJIOGntIXhtr6A8n+GgJAZzvwrf1p
1N4s00NamCB1GnvBdC+5q4yLED4//DiqssQ5PPlOtWtv5ci+c4eoCgQI86TCYpaU
ZD1H1RljYLkpUeY24Pwr4Tm5LmAdJnNxZyWLL5R/SRDcF5ChLCEfkq+PxsqDBuB8
0JiKQcI5eJT33dGP9Qs/XAMlLb2Bb9nyvmHoYoJBoFUoCN1qdrmYJIllvTbLf0j/
w7FVTx9VESkXwG+gKoDre8BPoot305OQp1nQsmNrFGYLgslkVJ3Kyg1NmNTfe5Ig
iR3aipDBiu4O9V8rhbaGTupXwZrWAzEqmiVcO/YgR9Ap0RjXJL9E8Qfi32k9Ywyh
RNXE0caPgl7LAyj9PopAEwtd83rU2dQ8VOul79O4f6pVnIWX/3ptl/xyqofGMIP4
zEAlp3spw4tqpPNxuLFNHcN7KxcQSLsiECOGbmuaN+baAK8+F5kR5d1mqKLnWbA+
zoq+ZJSPzdLUhwDDcsoVXJ+yZnw6RYWUhUAWeuNTYeqZDjT1nIRX0EmGhjU4tXka
pcXP3oFmjpAHQMtCslNm6Pr9cNiu1aD4iM9+Wpas2ktK5FVch+xspmljlrJUwdiy
ywu7b7BMJD5519QMDMsBYrOUrixK5nUfOfibcByZ6oDUzT4Lv/5xOBE3Ev+dzYXV
f+3JtaWyb+yl8z0yu73wR14fB/axVwFGo6fZdTBvqj0NuujRJ6tkemoTwtpoPH2E
5oJY1bLHNPcg5XGRFub1VVG206OSJx2zW9mozl92LKytRiCEkFd4k409O5fW3zD+
iJcCjxGukbKMSfWbDm6h2GhqbiqaETYWOL4grhmrSSAv+qXHzT7eji8BknT4J76J
0CCGFgHdLtR5Ci1K14oerRWeZEHC7fzAdhaOCdZGKqhdrcfy/kUiz/wbaqgqlsVo
jR7+QCzRQ67pxP3BSApf0+HHavbYYlUJERR7aW55yhd/2podGWaHJ1uV11faTTMS
ZaLOFVKL2misNyZNfD5YD8cM8mo03WjjbjjTKNj68fdVPZ8V3h+KLKxhEog/HbXh
Wu+7Rm4V9f7e1u9kDRhB0VaCwkOxofXwTtMeVZslGALIwWAcBFs95zmyayVQq0to
qPbo2HZaMUtgvYbNxp1Ulw9hx+2HW+yc6hPPeaS6qLrpQQUrA1PAbCn9jMvNGT+F
ZgCkxz2p6B1mnHlUuiuD8AFh0LiNsSI809yK8mOpaVcJZlfeZm+pUS7Z01VmlWW3
Z9t9DKlwmOjrSneFrpb0UtOuk5slbZv9sjYy4zMXlOkMwwJ9Hyeeb16ExwmE760f
2KYCQcIQGjAUTj0Gc8qK5RG4iYzV1Nf5Q/C8F8oOr5A4ZSmk7VPrY2+7iGoBAfDm
735Y1NmWOWdKCemMOQl9ktem4aPdutzEdWaJZHUVnqubC3gqKNOWNpw0ap/sHvX2
fkp6Ot3CZKt0JJnmET+iHmVO3J/AOvXJCih0WvVGVz4zFxM/Eel+z5EcJSqrSQfG
L19d/AblwAWsJVXCVSbWpCFB65vUnc0fHf0TxDrLBZtenJiQVFzi4evAIorsOkLQ
Y1Uj9jRK3jRNV2VXhqFCkrhSmmJKRTAeEWBMv+Y8ovFqrP86JmIcN3x0n7ouXsLH
fmKkRs9MC2oH31+uQmymgvLmujVuDH0n4gzQylGEeeHD7ocChXJ+gk4S2R/meTAM
Qb/n7I3x9uU8tf6E7l5jGkyWQgE1HDNk3K0sgLRcFQpZCqvP/FnnQeM4BCtwwbjp
NbDYxSD62kZpz+3B+dBiIxkq1gKOP30S5GN3NaJxI34bJCg1dyUqbcgoAxDrrwKY
6KHGSDBno763aoON6y0o2Fj7PlLjy6DLsCrG7vqipuGsiBIHmRAkbdfP/fhyiVjq
R+wA9uG3IzDQCUUuF0KloFEx9e6jLLYbnABGytTefIBiMi6+G0LLBNw96kOLVvU2
Zy0mAvZ+Ui9ESztv4gI6y0WA5GZVRIQA/2Yzyd+ui9u48acWx7BL1rDefFIFLL92
/+if83bpQC+BuMvjAwnmv9DmKrGdPyBnZuTSWF1Mr0pFVZPzA0+eJeuKZYH20Rth
DB5RMni+r3yuDK3UzEc1DZM7sIj3ngYKKH1n00vB75hOj4EpRWiGRhK2riH4I8bM
eOcuz1S8a1OOUDP+ggfpxO4Odq78wS9X3Y6oNz5AGHZrvJpifWuyRdcLY0VAvQu+
dbW74W02sjB0Tmq6ZrjpE3DqbihnJma9j6ambp+dAZyK8DGhbG+rfxkGVDmNXIaL
jio1omVbmiB6nVqj6e83x7VQYbHpdt8uOBiW6nUnq2JJ3feC7g1Hmmntq9nkKiGH
6pY2uIpuF575H7SJs6XKN/QFU3bHwdpIfJ2AvZMhZlhUycttzlwLeVNcubL4xUfM
+ze59ahjcXltPWragg2X0aH4d+AsWHidbAPGQTbiWqR5zsGDR9K5TEPL5DzYu6T6
pezWfB8bsP8N16jYh6gQbg6FFqXstlOC6hVE9roW5lYzN4n8K8pyyiXt04oH0F5B
n6TVkqUGNRDCyaZvGA52yq6XYBQQnd2pj1jPdUXt3Ph+3OwzKH16551wQjihyTfc
0gda929gG95WCxe08jaeb5gPa8PNjbC6+3dRF6vYGSaTafxe84U/SpM0HDuVeF04
Y3xTaq8JusXHXosI2hFmXjkWD7nUalxF9q4g14p/ZpffbKmv+53DzXDZEWr8Z9kn
DePvI662FvNKrq2mHNv2f2lmgoeviVcojuNgGc+iJkMjeTnU33nQBMioUmSNPBkg
g+OjXTr4nfTjAjUfgYrCJUN1eK3QHqfssEbYA5Uv99fAAZaQh4KD9tcXrPpl7aZH
f/jHDSG3m0kYyyrxW5gdFitkOriqhHOty7JVhfwXVSVglrl1GOUACx1MzZD+8zm8
eMWedqSk6yxJyP/QBETcsNFriL5Mb/nxsudpwZ5RFv9V1QuBhhd9A5WK9AYTO7te
bRUdQnw93OfrM51i8SX7AsKMXJ03mua8B6U+tytmdQTNRX0dC54oQ0UUpRowoREy
+5Em2tt8b/cM6EvGe82XR3xF/XB/7E0RKyW3UmzgHvrPAvvKIHxATDDBY+qvzpF3
NJsDbXpABPed7ugIqLJH2khw6s4Mjknk5FI5yLVWvDF67f8DLCTJydGPkFLqaeKb
o6DryaqVEQiljJRtPB4adxBT9JDhvoFvPKajLlOacugcEX55J3kHNHdQOBaB59ng
613mXegsTbGzJIInBOKgUd231AZJFn8/psJybz4wiVUv+OJ9z3AgYXzDB8bx6BP1
8LSVBgjkpMQftCEP+OBDpzIhzAELnjDZolKq4EvhUlMJMHPxbv5yKyw17pfawCGa
+GJkHUB+TgBI5pNJNqi9vmoygmw2jfUeGPLBUN/TNFuBRYh/L2gcmD6lJFqpXcZN
shRgILlaNI0lr3+LMq4fOfg3YufG0wKYv5wnGl93sMGMznBZn4hp03e1QxjLCmrq
5bgzXI62utijvjpnvLVW8TK1aNDaGFKUtUygKSkA08sqjeDuSB6FkrgBEs0A0pLh
zkDJ41ep1K/oFHCAmTZw5T6Lus8aNjuR1VbmnZi1zIpNAESRT67zycBpIAyv+jgT
TspSZ6UdQIYhnkXfUEE6kAkyaiIEoHdGqtpUOxG1IADVAU4BHZ4NCC2pme7AIkFT
fkPn5Cztm1hZXh1Uk5tsCtqOIoMkCcQBwu4VH0bi1TlCKMHbpvWOB/Kp13YwHokK
Jozn8xisEiCILVBuoFoNEOWkDwmCx6QLTubO96MOmHKAnb8JzbFlJt+K8svDoZSQ
ne40SeRJpd/zcDECujny6iQnBtmfk1nEfTn8sL9ah4ZbYjDQHlzz0CccjTk1a9Qu
WqRfIy3QhWuYtP1X6dwB6LuIKcNEeRy1eTvAAXUbteDgVK9Ah6tx07Nxyc77YEEC
WWlNlUBqaVmxZICYNQSa235eFWjLHHhCyeY7GXZu65Wfepa+dPHQPEaUVGBAzNn7
pgVAM9b18LaZCYTIHfZFSyB+WF0h/PnOAX4lF7DO0ke9WlawUzET69+FdvJNm+Td
6lyna2ysMkNymQzp5yGE4WxIQnipsNAlsJI9ehkTDpiW49QvSkQOpwvlPKLwCtbX
1kdqmJqTkD12U5oj8mYafZm9ksqa1BUeKw83BTV0A6ejqkUj+C+bAMvJRPWzrV6Y
oM1aj69Ffy45qvLFJahTHna03HvUTugdwjhUQXJyfE2T/XCfHsjNnyvOZoVKQS2D
oYdg0UND8O9Lz/cInyrci+zbpOPESVmQtVsnsJDCFfHIaeqzEIfoIwWZyZqwL2Mv
I4thbzVG8J2rhL3pCaaHMIx+uqfKyWHWaZ5qk+J8y3HfBtfJOYv2MpfCQTGj310t
coZUkCLZB2CFH0G2Kin969OhXgavcbK8Y69YO4KbyftqG99wwWmSPN7bMEd8GqJR
WO9BMD59gjIumBUHXXhIkPhJKdKxsWaOxA5Zbq3WjRYGZ4w4t5fG0k7Send5JG0I
De3HwizvPeWUaEXr9A9T0v/BV50Lrknbgp1EOdycIU1LEBhkdgXxLUnMTc0fU8u0
w1g/uK7bCa16n/3tdXPuNLz3QpAIs7J89j/qEFd8j+PLWdfWMzUPB9Ad5IA0M84D
3BblEfGHX9OI0GWvtMWVh6edVrexfUIKPbXTPW2+4KmgWrvpduTYvGYGHT/IIbID
k8PaIQwe8HzT06vmWDsYd7L4VUp+KIvKSPyci/qowdX1yhZLRoiEH1I0lExdG86s
cO2WxJsAWe4BvMS3BEqX3rrF1BT5Dl8dTSm4eBXXj7Uwuu9VNSbELi1LyXcSlu7O
EY9qDGl3tzghffwt5Ojtlv8qUKyTRvQvRL0vSqaSgCQi59apmHTldO26D90K8gR2
1WIjIi5ye0et6+Nu67YKgVVTYrPO6hTqynwo/377M2vdyvzgSE7ogLysh3J5b6NC
2MKFWntOLT+Q7oACuyG9GpUZ7IBBF2AviWIvHpti/BQ3TLjyYR2Rx4ZDqtzZ+nn7
C8wZA3SEPGHkGggpyK/cRdzpcFrAZoff+xh01dKQvrD1JNEPwFJtTaA8wXY7QVIm
SIR5UK12Z86u0Vr5+RGAiMWeJOY6AYWn5ykTGbE9F6/g2uILjI9WT52I23EHD7V0
1gh0lVdwlXsBLahggBhdXpn1lo5w7/zUBk1fpT2o71hdwKzsw7skha5q5ujbx3H1
OG1iLdq5j/vEwi/af4VNMyD8PWPm0SBEVJ81iN4BlViMb3M9GXGiiejEX4DqYUJx
L+1mkt1dAjxkHg2uR4aqh5a6LB956TG6sami8/wdVbI5djga4kTrjS4zKJtQ215Q
YgjXGqTW/jQ0pmJ3X/+Wyz7tC7X56WMFxvCTsBTrTTDyJCo/vR6XFJISwGmohuNx
+5+LuW58OfTHfXpvU6K8mV3TJqBQ6gU7xlqMYimuomvA5sPJ2Hi+oKSojmnF0JXW
p5LnfV/VUvvX7Jl0sN2HF8sOmxNpqyU+hpV4fh9E3cV7QTSmUOfo+oWsthcJ3PGo
1svVRA+NJzuTa5OZwEbhG4saarI51Glgtgf3ymj/BLbHVEI71fRUQsOVh61ct/Ce
mMICm5NuXXg76uwVUUPordU2BD6dZcORvDpCqPSsWWf34m3RwJcHvptvTNnrHKiW
d9LCqBIEtRItv29psNc6Arv/0CvtbvwmPA9dHaR5A8snZBeRMMOz6uj9e7tjh8TY
pfGAXoxxftgl7zpi22Wna0/BaIW6qX0kwjT3jg0n3/6E0jA1xmr4PEysThGDp1Qn
rcfFrJM+DHylqd8rF0VsYQ1GWmz2JwPI4j4gkem5UhCavIj5zH6+vjMR8YLD5R+u
IiCvEojRRR+3Qec73rb3cH42DZE0AQbJjLG2jcbJP8hLogErMLwWceLlN8dv65H7
+lrM5CENRbs/DSpk5GHadQAZfTi/A4zmIMuZQnVVAcf3WhwU7EHshsRP1i4v3g7p
SPUT4v9rpEqdGuttjmc/6a8ipVzRrmeyG9Np70Uf88BrBdOJuIGJjrl2MpPfY0BL
HhRulrOLOLANVv4QHPq7o2jDoy8T3Nn+beoh/4Q71ur1anW8bxx0YriQhHRoRvnU
TdemZycgXmICHXP+QatDQZBlAbXPFi8XC6yywKPx0YAUTud8ho8pe1PMUJl6y37X
dOwY9fcJhln7KWIDSGX1KgzrfRqwAasPohELVr8SU5y0Tr5RgCM32pntaXsQRIGw
bi3quyxBiSJODss4C+B8rGerZvcaafe+ldIv1o4sQj1AQzte+Xm0WtieoI0WOEB0
T4CR8eNrrnTnv+jQuWe2VhMc9Vh1Ces72ew3g4oGSVmy4RkbtgEVWyqK1IWIKkm7
xFSLvKtKiYC1nRQFuw2tKDcByRVea9fEAKyCOYqJb0OMbr//Ei5B1n4VzfW6A1o9
pd8/MZNaYf9wXle6aQOGrS6SBhhmKn2k6413y8MLTO7taQjn8NdFlzTDwmeDfsXr
o3VsjKRlpMKbxtUcwh6pw2F28RnHkVFh6+F4S2DHuGxDs9mokmA9jnnTZjRORZLe
pxf67dhcOZoD8aeDIXOr6jlgoGJ+p18xQ/Jm54wdmgEaDXio4IvRJZ+0TvxWWaQN
eDxUNnERfAw77Q0bmzAJeSfPi8ZmhBKW52o69wDqZF5l2mD2KHQ61ZWaNCEwjaCl
+zHEucyuBcxlsuBRBBMrIeu5q8+Oai6cXD+tiKxgpWILDBQwt04Q4ia2lW5FUyoc
z39F7IM53ZMNCnR3WwrjQGLtt801NSCrwTkurOUj8Lqbtq2vEyQFy3zbrFW/wsht
yDgLfvzAzO6oeZ/Q9ftw9wq7KvwBOKKtHJlwHKg500iDXZwBOBtg4zd8sB8ggju1
kQV9btabmrvIVPPdJEE71V3HzaKXBw/qw7dzPqYNl0gfo0L9nf77/Bj3z7/wDMPw
ddXxo05X6ZEk1Rl6d2tttnYyifzobvEMKSiQp3yJw4Dml4s4IhYTgXuAz85s76Tz
nqCDNna8yhmr+/HoeC8YZb6HWuzfnDI9Lt+xNkrKGcINh7lzHnUt+3/1cNq4CiB/
JCt7GfRFlYftqhqThLkG9ejK1zF9ZHTz8+I+JqKwsUYHr/DZqVmjqJrNsJAKEH4J
2xltOn0m2wBtzkmRrN65nQ+vi7zMS/cAfJCxprS0nqnJHEduun3Y/LGycweMxYrD
Mhr7a95JZnwqmIw62PuOfmaAA9rKOBt9c4Dzj12e1gG0ytbcaTNgYQsvrDkRCaEn
hc0TntIWdxNfYN5SLBcDSUSpg4dzx4bS3yoR3TuU7Np9HN+SvESFz/f9oDI7uqeQ
5AOF5J5gRIe/mtziDz5O++s2885U4Z6oLn1qEoyyww/uqhWFuGonyz7OEwIY/OOV
wg4VhygebTvDQ9Ab5eEHe0JpTlGfCzytiyAriHEs3h3A1ykF/meRZJ7luFwbefGb
MrwZcKtRkRUYC8sNhg4nzNxt6whM+qEOZQxxVMxDsYEXkDh0Ecep5DwhDO/ETXcF
G0cLlKlVovfH+JlLT474MXxa9BA67Ccu0ZI9mmAaQ+VYofnZ+HoN3kBNSBV6mkO+
uW/AZxlbqEwwdJuj0YkTI0T4fkJ2q7tbS9KNoGDWebR87J8BCoY1m5BG8du28q6D
PQSjTWCSsb2Ozsh4/pwv48VwEO72gwnP66xW8RwWoOkMeVWUelVp5+OaSMIhIX6V
gar+2nhCBJrA3G3VkuJkH79/L5NEXBvA0iZDozttjTibgltgjanUxt1qE7KwMXWb
kGCRLeFrnd+9wJjNHSs3Bc0yrq5fCJYelfWMMXGUphfaINpxbXS/VJYOMQK65Tcg
1Mda3S7o/n6SCMnsri27eNDLpkrhjFTXNwO1rlGl4OKRE9HuQlBODmm2SSytPaG7
UxThb7hgSJMkzp7TziVXhCcGk/7MDjIwR3rYBwH3ARoEpuOgBP/VA5GGr9K/+gvn
xUXt8oCJ5kOiFLYhg68D/q87eJN+dmSvgM5ZOlOkMb55Oa9sVy/URB/Eq5MzlaaQ
JphBM9ymMdSVs4NSMihV5r3udnA45X5kE+RaZzyoCsASxCbsy7tK5M7q8dnhkikW
gla68GlcB1H6CNf9NJqQW5rvwBbBc5I/gXbGdlL9SQ80W6SAdV9L5FHigY+YxOsN
ICqzO/IFN17n7ceomMs5rvYv6A5QwZEAAjD4D/yvCQsO5sVMh2PngNA8tgl7/5/Q
7dPqppJOVzN4ecdZN4t7ViK2IGfWwmiuysfAKuoDFMf8gbwkrvkAFKfpqjCJILx5
I5I7/VcaGGmcdyvjLW2Kxcd1RnNKfY++OeQGAyzpd2tAFq/0IkyH+3hDq2BV7kuC
2EkYroTCKJAzs2fuPz0rQwXywm7hC0xC/NkZ76UlrS8ugiGOQT09kDJezJXsDVDF
+giFMxAKVrXokxxAoAFtpQtthaweObtVzXmm2rJMDmeevtYG7XdTTW4T70oAvYvu
Zh8Jr5ua8srR01nLYS5VavF99MaGXSsEhpOjy5gXI+H+xi/3x0fi2dIqarNUe9cL
caUcbJMhz4baM/0O4v1xUnQKGKtUVqskpdLatw5iAp0QM8hfhN8PgKFSmjNpVIYu
TRL+ZP9X6UWh0vecwu6LENJPNnACyAf4FyvZzOdxWfHWCUYweIyaeuHcmrbSH/wC
tqFFSJyD4MjU7YGfpFFKZyn8dH9WJgcOr4P0XiWXR3+RGewI3ioY0ufiPJs6ueot
5NXy4LpTzfI/ifkcQuBm004e4/ouheC85XfHgJt6sfLXPNip3YWn5rrPD0bhV778
0o0+e6sS61xTqMk3MsZX8BFK4C1SLKma6fMItEHubQScGMIxP3kk1etPUIhJ6JKe
hovJhkot7O9xh21n5ctNAQw/nn3ho+HL9h7ExKciungQiGvHdZuNZeiGI1bbOKwK
NQMiuiEU3wlKl+L7vL6Bd+PBl9mJlPUhANgTqC8/XNyDveM9Jwcs01un27PKd2TT
IU/hMXwd08y8+rRu06tLHAHKoTjJgo24c+YCE+1cgoDiTMZWN/K8GSY6yrh9aqkI
qoUiHu0GWShoPpVtIhcLpZe1UJik79Ly5wDXAjAsSMuhtIAus7/0O4reMzHeuDoP
QgYTH78rBWlboksUU3gzGD0h4bwm7a3RCnks4IEHkvS3ENQDXFpOafsjNn61ZrHs
0fL735dt2l61wizhQYcm3pq++/hVpfInw2qvb51QXi30UhB1pjdO9J2yyDeAokfe
x64nZ4G/HjFprInFS6pYZvpdPYpB6ZSgeBY4DvnnjU1w4HqdyNA3uisoXbl+1wyz
v78H+AqECY7FZNsxn1WADhABTWzovKlNKJbnh2VrCVveqpYn1ThtiBMrPtXVUkjU
I+JsgBXgq1BZdqi5QeTwBEDY/f0k/0JogrT+lnDL+SKwYIA5I2ElrbcFIWDekhlN
7uxhSvu1n9pe6u6REZaLrQD0mmE9s3QFH6Bi9cHnqsB7JcIUm5P1uXqlf9dGwEoe
2nycNwfaObXgWkpLvoCy6MufZ7JnB1w25a5nHRL7meW4uj9bKoEbgvvCTqy2Bk4j
HN//BnAp2xahR8W5+mZowJlJzFUllGCGoD5OxpFq5+1Yf8GVnrOr8Meue0XLXopq
cntUBmXZqqO5UwvUxjria84a79VEAj+MnEZSqrbnIAPUzpXrmNpgx2edd27FCGLi
mV658MsXgP5PvIPDjB7aa6IepMP/fHr5R/lc/3IPyvB8QvO5JnrG+JdJ40bUM0kL
bk3jS+JcfWqZPaJzYpwvcaXu5JB/YAMQarknPkBY3xhkWJDMp0NWjDc9KZ2OxAw9
TIWUkJKrEYnNSjBrdptO+Ru4smrTMi3mdQdF2N9Lyatl44fPpn3BNoBcUWDNGeQX
BJH8SxhYyy190eTCAulknFb2UNjECQHsu1eC69iN8dHauZMScOrSgVTSx2qJxjcY
EtRyhKKX7RF4xAdrsHumcle53BLoEjRqfoWpjgTEb1wsej0nU2vc0c6OUr4aIVTq
PEXYpBqVVMKGJiSVwuyfhlFyglLKW4PVgLYXh7KEjFJerPrBzkHn8bhhaQDQs06u
OCAk/mnqPKHAo1AnojjIHs874vIZZE/XTmrUNDrIZj9fcESrdPRaDOS3T7yg5pkb
FF2QoanXsEfZEwssdb/9xNkKfNRk5Zi+F3PjrcyN6tLv0Ia9GQUjMcmaa0l9jaD2
Vp5AN0XucmJGZhNCPmvb6f53RVsm5IYMnt0pHlInFiJKH3s7Npor7yaHgZwcgf7w
y7YTFxHOdzD1lVJSzDXDkf2i3JCpxjvLnQcHJqUbHC/TxtFCvn3lKP9D9Rjm7vcR
8nfGQ/DrE4wRhLYRCjsrt5yMyHhshkRdC/h9Ak5aNyXSEJZ4ZleB1Tv3/vgGJKXa
uPIroFyHba8ooSsq9tfsFai1+qCtGtNOQwVLTELsDCaIH4iCv3A2TrQrjkhM3pjQ
kml3Z6QBAWmiXYqYmDLddeq3kt8DcpyPtmWM2U+T3RkFDIxspBPd061MdOyrY31D
XMghZquiXKOcX4NMl7c4xc2+L7L1766K7C/l2awZYorkTY6KUonmPeqvAsku/BRM
YrsexM0Chk2hfKR3z5VLO9tBaY1ppwgdZMVAxovb9f3fKOoyxpM+LXdMY+kuQIzT
E3v8hJtxiecHWdcEDBdxatJdgxV7LjKkrYi5NPR9nPlKVrB0w4yNYqhoPwAW5nct
xxXPFr/8lHnnupfrlqFbpsnee+Ew8Y50j8PjwVM2xvut0vAv4af3fDlDTVvcXtKF
Oqs7g4kdIS4f4brF7X9fIu1DJ+FJRqFzRHUdm7aXLZAbbLAUV0VAq38fw/UHMUy5
SSXfntBj1q2ww/GvyH/uyinuO6+YeSY8pYcXqI+rNrzWFvKMLwmrb+Fo/tib6Tjz
R6/byVAamU3UMgNoIBlZ5sAHIW9NH+nv4QlF5tHtszVQpHKxRUjSDPdsiDbx2fCE
znjZy6oa9g4J81B1GzBz9pnlDechM+g1BfuQaNvZ6SuCfteOTxppZelCxGDRBMAn
NAVOJJPNaQWyZJ/vBNMO4mbkJGp3nTRQ0bbKHH32bttlH9s465bXDKbGWBNaleY4
ePHIBJ/x9ybXV5NOfLR61+TWHcoy/w3I16qIF/eSUetrno/S0urMbasKA5TXvumJ
UDeivV5TBoQiGu0+c7b6Ul0pNFHi7UcAzJ5i7qafqafiNWAvow7ooFlI5fO7RJP9
egNMakn8XCX4Ylsh3D8DnUMxwi9ElV5W7Tq28YAg4huJnZYKYI4tPOc2lKHlbpXV
xdd72PyRN/xXJpeX54Gl+XIVjUjsOTq8TGL0bMgKZfL7OlSAbHW2+2YC7aXG9NjY
9R3XgucRRvBA27d4mCfdVcySV3gA7N/hUPFcqFcF6MhkbKDAbDdz64noWMl7FuoR
GdF/OZdBQVcMn1FDau0V4Ve6nISQqVMiMgxB4ABaHvrMqXE31pd0cSnIXAwo9hGS
+xPli2pNgmM1Z79vcNkrz4O5EnEciL2vijw0+ApJyUdv4A0NZz90VjNNiPzkefK6
U0PQQfTtHzziOn7STqUuGyuINaN0nDUPm36VxKYO8ZRYinf7Htr9GrW2IZuIynk2
aadBSsJTP8/Apdpj7Lh4QzOlsn3qKJPnlJkta3JTcdxSx/0w4N6Tg5l3VSQMyLiS
+7Duh1OwpOIi5G+bNUUe/Cu7+8+wRTjQ4y1u3pHFra5+VBL1dFgBag9OuKMy2RIM
BJkjy5yItGJy+vnAh+SsWv/GjceemoVXINIUGj5dLZJoCOueJWVLew3v1VlWNtFv
9IBCvfnZ9YB4Sc/z0kGe+yDYQHfKq4dDEtc/rFb6uGerlBKQWhyBlCgsPyQDsGlu
8JGE7zkZD5RSWIm0xcj8vNJHtzE5jemKscTIvSVWkt1y2iJJxGuWTQm98XRojXjk
FEAvKHmC0ys7u9lsVgxJXIcZNnB447w5NBOSqwom9l5LPWSNirHWmNk9Jx8MkXuo
CSQptxVU139JcpOH6gVXVsRVegNlVXbN79Re4PQvTHX/B1gVDqMXYX3Vq31vaqJO
5WMyVhzF4Dv0J/5xqsDzFgqyPWaAcYyPKWNiXITe7eZNtm88pXTP0w2mMp35afM+
aZYzurLcNxesQsd1axtGXyPiBdtRXdoJkv2OaXQGC/9cH0FaQkbNRbz1mL/KC0R5
/d/kh2IjF0KrdCdNvZDweBBKdUcjyH1X+v0Lrlifboe/JsLz4M9gfcRvkFY73WZ/
1fL7B80CWq9m0E4iDO82E9EAoElzB77i8dDpd97OLTnS/Ds44ufKPf4CySum/cEm
3bTRranLhXSVMpNs5qaASW8BDwhXwjcsT0XhAFCGwsZ8IGPG0EdFHfkB1Q+VShQP
1ekC5esMBRpsPUk1P0SPlhvu3XNQy2aD102aDNS6NQ3Ff8lNuI7t4a0arvH5ZMdT
IcOW2Ri8Xi/QC0enZAwSKDBi4w0UIUFQ0i1U17VC6lRDV2CDKWueKEwrWKGEqsNy
zhBK2xC+ojvMqROx62EiDSD4EkY/PvgEkBlzDLvoozuY+orxUG2o843teiRDKos5
B1Q6X2zkAWm+0jAM93bsyMjXyocNzoKKC3dU1f42ugAiP8GFRagHJiE25reCH3Cq
P9XnttGIlQxCx5s9rTM98b8wqXgME6Q0JK3XLXMAYS6HNDWTVv3lOyzeNE7uIZwc
hXJzuKKKLeEXzpxiTMgmH3jMDwjvFvBFYQexQTkdGw7q8jEdHyp4fEuSWJ6qE6qJ
qYRn1lhWyP3tj8cutWE9m2U9is6iI4yG+ufEtykOX/YO2U6XQ295m+tAwt4L2vQF
S/LLVsqFaW1od3K5LJXPEaaT39UzRS4WVdjBE1btLGvo8WoJqgejcmW2IIjPQ7G2
sZt8IWFJpXwp5e7pq4BFoqGUvbitrUL5XVYVZvAbj6M04Mnn4YgbGh6vqDNWTWup
dNZ/d5vqE++ZgaA40xvSR2SFFx6Z7B4KnM4JAPplJvvKGhI/Ddaxes7EYWCeLnv5
dkry+GaLe+EPdGIPlg05Erl4g2tSTL3IZGdn1K4mSQFcslL813rfqt/K5HaFxmc9
PxF8o7R4M0soDBvxyRX92vDxeLNxO6RkNojKPKHToD5MjRDK1zxjiMb0cEHhtbWO
p+Qj1pxpC/Cu+/TL+O9iSytEAlKIM6ONX6CnT/udTqlhlKJQ3/mVlf4PXZhFHVTt
eryI6b+uIFsDK3nLnwsuii5e0g/UEvZiGJVw3UTlN2Gf7kxQQUOjZRF+s9gFp6jc
GMo40tUBhnxJTLh/L0HeLfPY9I2Na0CmB7qLQ8xqp58ElDN+HPehkWD8wnVoup/0
2HCVPXrpMAAsLrA1Z1/26rsEvEERDF2DJjUpyN2duXEMG+3EBuA8Y4Vk3/N9zZ5D
HCR7QwnO/7Ipml75TnNM+1DLIjLZ66wWgngQks1pWwnYcfiy1u7aEIzUq77Vpkib
EU5R4mPzcu9oDkZYH7fkdNcjyxdXbzWdCEk+pt0uJP5sAVmDu7a89TknaZYgieRr
jh0linBluJcsT+OVGQFlq4Ex6zWUfOJ6C7zLV/2TQMlRxrXVGJdr2k+hNly/IehW
kUFvIqOPcOjIh1rDBaRT2ElCt1CUJnIyZy9RfocdrqNN6o7qtXtmDkmVeG5eJ3H9
e+8Dv3xaAfEtUsFM7TA094c0R9Y/MXQTTh3VA3mrrNJn2SnHaCqAqvK4CsQugAh0
lApwgiT3h7YQ6gBhWbbe9O85nThLz0VdwQ1WKIZIDLQJvjJvUXCi+9VbHueFCxUk
SBsBrhJPVTaKL3U5FxmnAP6B1L4TCO+A40mprLjsVUux3Js+E03FIfqdE3f678mN
Tww6PppcoAusWBbWR/E9nLkAolbKLOXGL7FrfS9gvYrhePy6xQeSz2HYHCu8yUZ/
rEmlHiMCYGeDFgL4KBqkHNx8snxDG/nhb+2cPRpaTVaCjpaOBlkJdjsS4syH68sV
jPLzW6R1QjvkNJlgJAXQi6i8Gq8Aw7NF8MxkLi6ANuFhYOIs7v0pQZxQNWABb5dQ
eavskhFNE6KrwC2zK8lg6S3Rw6uqrftSSQS5WnWPRVgbhrMOqKQGW+D2GHoUlJZQ
6H/vCzXviYksTZv8hEGWrCqvYtMdNOua4OB1PJjHiL39ltnvoqNqHDd8N3e35BXP
QiOTGFLUFyKCVhl6eIhj/F4JC32fMQJfOO2cBRbtDwG7a0Ww2jI5i3P5rTco8ix3
825UWDzjpleMsy1cv3elT1Uw8cZDcdVdrsv8SdVo0HRht0o7uACUtII9f0QbFApR
1kPpFANopJxJlxCgCOPutR2lv9t/DM9EGwaa5PwiMJo8Xe5yQmUjSNEcx1irvwsh
lFCJoFC8qNicCob0sVBbrQj9CNITLvuB4Rruuiw+6xwnfpLsWypex94dmPaCsgjV
GHHkHtR+4kIqAgtA3ZeW4Nd07jHHrA/OFQsHbzWSx5DW2mrMAo1he4KnKOBE02gQ
guEzXwgmW2/x+6DyVV5/jFvOdHA91/zMzAVo9yY83uWSHCn01vtF8cWPrPXMtpOM
+/P77GwIw2utRXZKMCEgRXOT/Ar4SZfHt/fF3sJ5zI3agg2IavrnsJFlsl8c/luE
LS0NbcmumI/7atTQKBuIRCyXcoC2FFLmTkghDmjlBrgbtpxR8HkvGSh9e+tluUT0
zKsNFq6jkglNYIC+4N/X3tqa6dNnSYKIvrkHFoIzItDFs7hhfxL5tzaV7iz6vnnm
Sq6ZYweiidi1J2eWDXKGidgG32uaHtA94CW0eluQHhTNJKliB0gUwgjuMv3kIxqV
/vgvZu2M+w49MCEbbt1PYp4CdcQuWL7oglJwAwqXGfI8YvecPJC38LzTow7F9RQl
rMU8+0craRReM5hRs7oyM01KDp18EyUCfZrvsuCa1/pn9njjdB9BImiSxgRcjzu8
xHmKCj+XtFEwd8fZ3GHoeoiH/PCBoa5rHI9EsNX5LkR23nc60QS1+wWpJiAsfD/3
uvvTId5/DVw0V0TEsqn93qBfDF7hCt7YrTvyP1LP+jJRs56XXM00z5RvLYU7OcSk
Mh7v/+T9AAP7uDJGfUTzIXSOo/hLGKpF/ID1XUlMDKRNFUQKIyz0GXf+Sp+IhMNQ
nRHBz1F6ZmT6QFzZzwe3qdjHZgNc/lxMpTNwRM5UE1+hJ4hG6DjM3Wxz9TFa3hFz
3DA3XeCpRPBR7+1OZ7pp0ILCxh98dstrddw6m09XxoeHStip8AxjST13SUEK+bHk
ldO3YxOT5tT5g7nsiP5mgMi/irC5nuYGfzm/x8XpEcMLh0shdq17gAUxzNnxhE0g
eTN2Q6//R+N9QongMnJH/IbBc1I2eHM1VZMIFSgK676+LtZd08ekiVSjVeS4SY6b
Z2/8e7jZlOnHBo8J5w7g1kEYoSOeLCf0Je584Unyt7v1cBtVnlmERmv3sOHzwiAp
5RjA8UlR5X0IJK0gFwKFexl/jJIfNHZxi2W4pHQl59vMySGQhsXiDeRl4kA3TMAg
gUYPKOrJwmyXaSb9nwPnYn4zPnzFaHVByaKnKohHDiwSfXG6TGfKDycjeIU8hMq5
TLVWpY5kKg0SH6jY83wWyeQefzKXNv+SYinv7o+HNJWPqkbfMfp5SvJcjmFM7nuI
LMSc+8qEVtNNWUhQbExtZBSM/cu5y61ST/2vnfpbKwHjQOKy4xtLWvw4IK4a+KTr
08XEqsGmo7sjZJyCNGoO6qVzWcFN9L+0Lnf4hyeP8obe2WHHvPG8kB4BDbgUbMv+
hdE7rN6HxXwo7GzSubsnRRoXXxxifJc2VBFz67Iqrmb9LKyRbBJoHpzvcqmUS84t
SU/d4usrbUk5ghiKHL5W9Qg8nqtt41Q5gATksIAPPPQcJQU309izLder4OLCiIik
iQRImMP4LoMLRUM7Y+rWjUNGytvFHpvpN7ho0z5cV3TerJfvv47fxUQ88R0yK2lO
RFLEmHTdXSSP0XPk6rM/XZkLxqPcaRn3oXoyGI07dLHv4pMw5nZB/tSQPGfcsJJ/
jz1MR+aDZ37KmOt1knvE52zfvUl5O0/ZmrcuYjDNhxpDCidv31cz6zfhm5OdSpbi
/7ozQ1b4LW7k327SfkZkRdH2iR4WGO4PYVBRlVCY4NJA+zP/CmcIo0+J3nsRI1+Z
6gfhT7PNaeuNMYSZ7hdRicK1rW8Ih47nNr9OB5MMcTc4MyJyOH3EknFbLmsjqjMK
4WE+/xbtPAyugx3IU0/nfNflt73BuiYnvnnTtoK6aWDJodbKd9nme97EvXxo9uQG
AbZ6JNTOr11n6AqCMWQ604ulamotiogPUVsQNmp5TrxSObqQSzl7cN6vrG5ptbY+
dhIcqZiyT2Yj+zB9phgQazwSEBhpyZxQt61FrWhiRXFPqEG15CbOdvFRBCXp6+8o
e7dHAbmOxufepJPhH1a0fgn80QVAVilTQErzUqNeTS0xzMo6h+URyOi1mEloQxim
766+vc1s9zR7jekT8F7HZaTYTDsFYyah/GI/Wpzynyb4OxOw8TqLJPJi2Sr6WFes
zBFVS/oYkvjsLqpsoQ8lV1p+kwOpRtMBuYoxk8mTrSkApUWncd3qQ0V+lPN6NW3N
Y2hVGuJGu4JawTSC3R9BTAGnR7YtUUQVoPUFkQRbxo6I8+VWPd9ui8WqPLygC8EA
yZJ/cvHOXS6nlNf550QjRN95wrMoF18qtOjNG7DcKw26pMh1AauwLNvSJn2wV5U+
+R0g1TyRFX6+V+/+wZKeGAZURrEhdo5kNupoJAENNx78acv1VavLc1umRD6OiRSf
gRDGru2kZcEfyk6ykPiAt22t/fwD91BuKDVwB9mR8Qcpx/N+Jd5EDjMn85jbKXow
t8OGbpIDbRt0BgdFFaVkwQAxDbQ58ZpAj8Lic/savoJtBWTx05qewwUtb8PZebfa
pnEascD7blLeCM3UkNSClau+Xm94QSdC/+ng3QOru/GbnnJkdsVE2vVHV/DM6cGR
ojhKtSg62dLPHbEnA3tMYax53rIZvVEdfm5NEGa+ZoZ/k2PpQQM3uMHlty1qjXdy
RuL9e3SCXjoObLAQ1VqnKQfqnbdGCa8ps68IldMcX6bCfLKYOgNhPWcRIuZCQRMQ
elbHQcJ+irnO0bIQdC2zAn/9J7Vt3UfhSX7vD0OoF8pMMmENF8Bn6QPckYYYGnvq
7hn35JgiaMSY1nHFNxAh24hTgbXb47jmMm0bu9qIt6FI6mwpAw1spCYHXLocIhjF
kw54EjA4CAMQ3zJRUBi78isFgJOkx+qAXlt5TjHc3qVrNMg5UgRJ5fnb3GB2K+5i
abtaGXBOO6MANofqMNhXRs1VCKBgTtkPcfkVaN9+pv3xGWZNCDqj7pogvsQFgYL+
spBB1pOqyRx1WrK/vNB0Ix62sCnR61uGEmV//GrbsBrL2Stqg3h48NCDoSh6rgnc
3XXBLUlO5AupdGn4/Hm7G9fQnEGJrmtIQkrxsKCmINYMjGTur9YJr/lqCNcxriIC
riXpXsISojoonwM/x0uwMK7KUbV9CllbtshUodz9IlR4muXof9/vRHfyBMvpmAX9
gzuDMsGmfeOQNSX9v5wuR7X1+iNeotWXFdXROYfD7AQyU87Z29WPAMGWvn/Zf55M
F6ZIf90b8CFbTaUxVVzW1kXKw8hrB2ndh12ik4+JzDoLVASPcvYzEl0FfXDzhgi7
YwxWKhrU0IoUk1ZCx+eeNphMJ+qN4TQ6b7TCoW/qULV8gt7GYcdundjGDtrh8OIa
dtRGUTXlJXX/JX0YkMzlBpzG/j6eWqrUeAfCOnTyr2gsCDkmI7bfHkrZch1uP0VX
afr/hhhuxl+1rbsQLS+aLkrVu8euXho1bfbrwz85KjPQPbiKdALguYxjQ90Y0mVR
rVjuyGZNT0h7uZKwPNwhwei2pSgmQMtGWqdC/8+P701v2IWPhVzYY5z/6nIB9MVG
wEmXuYusf1jtbrCLy+uQv2eqsa2KVPiR2RWBioYZlMZd6YCr0sKeUEZiRjqABhTl
/NZFsPmnINOBPYVfhCSAA0Kp4B1trQ4PR2DrMiIGAJoz2km5KF/AXtHZ6UwoVDLK
rgW/kHbOW8kO9aJ6Y5skYd4hp5IQ9gr71a3JNw9i+4VTvbVOQSZBX8gow6XJQY5n
wEdu6z/SBdtOxdcRAPYneAeBMqOCDOGr0+fwc2dMEe6yWzOTP3kFX3p8/X0XC/s9
ky95sYxePi4Y8nP8VCOwh5qy8xCHFKV0ULJQZ+1m5d9RCuPNpLzvy/NDzAZXztiz
fIGbkhbpubfD7dibm7xrGWc7K/K5v2+suv6YCR2khgsNwvfPAw/eUxHUTVwRf35z
ckFG5GUYWkCd9Qm4WL/INPFbKb+OfiQMJVdMuI6rhWNqKMhQ7B+WaK4F3xrIXHX6
bJgUq9sT9OPE1VtVRKZJeu+fj1DJQyP+1PmZjhJ2VWAhmXVJ/t5mMU9HoVNc+el5
bFGQVOrj1Uamo+aEy96mKf92iiHopvRzv0bsIA8JfFyG5nKq73fG/7/3rSevnQ1b
/vOsILawOSfsM/E0XZsZcw1XbuYRZ1MUbHTqaOdYihL9btKpYJWL/dZuAtqkPfkW
WqZGm+ne+1yX5R3BaxLmL42iVX8K86dODc+47IdlZTLeDv5F5X+zanw0Z1KaRHMl
VTMAvI/2vK6bd5+OeS/YreNHGSDyrKf8hdb/hlELL2rgQ4TE0wqZ1zl/4QKv8D9E
EhSh8f9rvmcwmmY2qH45OXAA/xFT2q00MgZ6LQ5pdtlLWECS46tCa5d8BjIjkZeX
14QqGuWq8J4/FTxbMB0JafJKoEq3n0C2cT+BINIClUQ+yRbIM6wa+POG0eqY5Yrb
xqYmiKfOlryYmCmgdlzkM5uNhTKrqtax7gB+aowF/4FGhRnX/BbwoOcq1OF2LHwl
msDTkofs5KUjkewUidCFJVlaFPt0tvhq5gJ1j+qO7VoaTZsiAER0k+lnZDMMX0c7
oZ/YQomZc9AYk7f7QtcTlbIGjmv52HKfddzap7lHdHGbag9kEKLwZduUnrPP8kkO
1asmjlar432cCB0Xk6mCjJFnykmaO0pLu81Fp5xwcpfuBTc+jAJT0CWtS1X6xoed
l4ZIyxSEjY/3nFcYJ81hs2eOrNJ0sAp5bbFk2bsO6TYBzaJ3irMVXv1d/QDpuTqu
ToHsXhkvPtt8/GABjrUkpfaLinKtOvnkG/TjxGi1vonaHDfA8EEMDEQAaxjzIRg7
eDATBWJ4cvaISzh2kvb86CO3T60PsHGwWyprTCX3YypQOIcbxaNt6b36rxSLFt0/
z2GANYn7yd2scc6UsAJDH0xHs8HCEPk0m7c3pcADAFZE6Un3IsWY6Oq9so0vR7bL
1ZFWcY1iDJM52OeAFHcMjDRfPGHAyKJt40xYhSUNBFHgaypauoiGXXawxcDK5kEP
+qv7C2HcmugsynB0FMeoP/SOwUdaaj476DAqtzvF7NJQV2Qu7wyELCeMIu9r04WO
YuSQ3GryxZqOSmHVYJyStkT87xX7G6X+vNVHdx3tmjSn8BBeC6SD92wYZsseK+zs
KPy7AeXd5/NUA3A1ZSRHxik0KW3OrcPzuYztOcL6vIkMtVPUJSA0MYv3keJA0QBw
zrNy78SXhpMw0gMlF+uHkxUrsQO0SscQuqOBH8lstgOn24DHvnfonrQ8tmXJ9rmR
wfZXJ8DyucHgdpKFu2278e5Mx8jsBa9UaEcGJuHhxzxfLatBj9WhK2BWGk9/rHTz
EbsWGtkbROsf4GPYTePdsDS7X0azBoCb0+SqJJ7uCI4e3xJYMsW3kQ+D0zn9DymV
Z5Zogl/Obx5QOObPNNT1jX1pwzgN4mZwMgmO/VzzWNnYBHMlA/ob/oMOcEbdTwND
aEjSaOrcdamdknkEkJmiKAM0RznGw0QR7UGdEy4RO8SRDQHnhvSZsMlhu9hNkkQq
L6ueFbYxbhsGrPnsXQCdD0LNxaenPbfO2GMM4+rOLIyEGbNxQwLyf9+/6Fp0+Ct+
XNdw2jV8vQmiDR8B/7nQicYJvh8KnDwin4V5ayh4f1G6o9A3OFZf6kSYwvoh9JDt
LmcDhv6ZwXa5nVt2wlQOM2FQelmV5TTMXNDoEHQgrGgcDRABVzZn5120UM8RAmRb
NED5umu5KXkZzm+YLHJtDGF9frBJqGxDaLv4Gq/f70exhEdf1303gB5t0/gfLflt
LMjbkeE400rEkUH3EaMprLwg+rI0UGOzRnr4xxzkbMbhDjSsrxWpTKynX9pwR03l
zKOrrK3ExAiDuxggKbozgq+Ou812TzKxF3sxCrX2EtRp1X9q9h/dzkEx6bGqXx8q
3FUCrHN5jCcpGuS/cNO8deb0KvFe6FOEmPP3w1yz0Y4GQCcmq4rcwZdR1KRJJnsQ
+nCj9fEOnOM9u7mOhhsCuWnIoBNm5Z1srkD3J37v3MdAUvU9GWYxJeJFap6KpCEz
cREhYqUIDsk2M3kqQlbWaVnF7/4ljeCPbORy5RsyXvKvxxrHLGKkh+JxKcfsRdgL
OAPeU4kxqbxQtSOZgfs1qxftrokAYq5dPjhar5OvQ8tpp8Nxmc+QE/J2JvkQau7h
RgSaJdBtjTfAGpoGHl7ya7elzmmqkpPHcj8ShPQ7I4eFw77qpu1KwpNT1KOa2tgl
RrndPSVU7YS3e5MKJczVPL8ugj2dnA7QqMXwYEP2CJpDWCIbCkeWkVunue7HlnRz
uRav8Li7cHIrI9N7xemucNwFDKAtIJOTNRGFl8oHc6bApsfBTBB6Ec+Xyi7kVEca
RSSgsbBNj7g2AGYIUt5uWrr0woipK2/IGscNQuFtq3FNX9NSy6NWr9QZYgZJjhZZ
P4gNfrr0ZweeUwrJw3tlNt6ShrvF8iCytDrb3G51vGuf8khDw8hbCZ1ULKqENpte
a49E88+SEd99/d5//7dhMV7xFX2q1x6Yms9XoQ4vRjj1/cZGQxUBU15JqhNRuSo/
4uC/9eKmuIpgedGiXhDawoP7+X5jiSbb0lpvGVBchycJp/8miPFYdr3FTLcIlQSJ
cm5QV/YF+V7+eDntKoSjCPKdD2X8sA0Te3tY5uCExFZmlkXox/d5EtaNDBc9tBzx
3e13gbCltfmXFCYxxmOhtZe30q8JOum1/cKhU5hgTqHRSAKwJWSpKAZgJfQyKW6E
Z8CDy7UiDOVYT2y3f8rckWy8bPfYNgNvd8Ci0hQrJWzy3At5g3EnfFN2YShUNXR8
Cx6QnqiILAyFbEffimErcRWzILcro1k01D7i5wXGJMJj5wDD0RUwD2u87rhvoFWO
DbqOVhve1NYLTs+MRrnOatJISEEi33Tu9mm2H/of5Yl+nN+3oIbKK4oWLSTAD8uH
Dujgj7p2NZXpg40TOPcl87WpVa4unW4xlNuYoJde8CxYAynIIpQoZ4opphoLuAGY
l8PLManIcX7QV3cH51YqG7GuZjlKxm5ELsDCC67kUoM6kbOeUg7ZuzAku1kmHXu0
r/+e/gGp38HUafztMN4IDKklm/6UA1XzOAYdbCeFWcGI6p0oaYsrsXHlLJZYtpGs
1++AddaFIVpjaRzExIWGZWOh/7EvexU3nElo04Pbw3u2K2XGHhTV86yEL+1Iqgol
iQRpk2rxH1Vp7o1pWA+X6hWC97CZaEk566sywI9CEkuBhklhlRVEsQLsJW+Wtpbr
scqXmjd/zgBM70ryq0jDFC/91YPD4BC4WGOrAMIOzH9eNeaZ97FH41prBA1fcGQM
bw9k7pKg8Y0Jy/3STJWp6uG1mlPHGuN7mZWDiX5nzi/D9es5yo9/oLoBleTEt3Sl
NmnsxMJtnQce2HQMCu/WPWe2AfftT1sALK27t8Y1AYpFIdbMHSwmHSQ/2GZ1ux4t
HkcOGBXKSvvZEJpRo27pXQbUiswUJeTYbMd/s6+j/Kp1jb6ifeqcT18qAe1Tv64Q
CqOnBF6bhtpTfy39gHxO39xhwZhYNIqkh6GSwAsU2ULKdaskqA4AIKbB5SLaGMUm
OI7wGjKBlA5CfzmIzyofWUSHOCQMvysr8cckVuTUcffRcFdbAd62OLMczfW6Uj88
KAapR/k/5yG92AWi7PD+oj9odEhuGVEhkIaZffQAAV/Xr1ZSghc7tJGPrsvGpDc6
EuhAXaPh13aa28Sd9zBYgcUxdqpRzwCHqT3D5UYsnc9ynpygIFbXOKDcNvwifxQS
/JGDZtpW29Jx6QuowQDJ5VDBpYGxqgSpHOx5HJ72AZadcY0vKgaZfS7aovCMFH9U
fiW6fM/Us9lKv0FNDn+mtDEG1h7MWzSGVXmeptYF/UPd55lL7YyFJQUSVXg3+50P
F7setJk7+rGXYFjeFRSVvYK/oyIJUpXS7FWdp3vNqrjvVTlxghIhAawQbqO6S4k3
cQOTjL7Bbb1J41+C1Kppa+tbG7InZYpJBPu33/+itwZ87JgakkezJZatL6c9bpvi
Vb1t0IPCinbaluoBcK3buLXig2i15E2ipoIUITSsgMwVK3H8zKzKmBEHuIVFv/nf
Ychj1q2YEEQ3FWZBc1AODpBjNXmICTek/GCuedOmI5+MQKzFTl6EBZysWXWlIE9O
pioMF6SEUPEwkn+RYDP3VRVyWpuvT7QBJwKwu2YaOsAm4WR0xg+YGolfwnBnwFdb
uOn78poxJARiX22pMnkAb9xKDRPZNt8MoaYh55LvX9CvWIhdn8GgGwMCZnWvyi5s
LO9L9+mAFgk9MyatRsYncm1S6LZ6ntp1+Sk/yh7X2gkP8gUO57iI+TJTnv0qVHnn
VVw6X8ED28049xbb2KoeKeuWniuV2Fb6UXe5G9ILsdLzeXR94lA0dJHr8/k/L72W
slnJmgnB0YdcosbIgK8faQrACKv4wRCgQ8W1RAHj6CYHnuBGsj/ZbaPDtVXcx4hA
w7tHz32Ex3GyFWIphpqmivbPZOGEwtf0fEF0KxXm9iYrZrwiapcW7ciEy/x0SaJi
ynB6AjyNgMl82uV02JLJF60+Yn/H0OiY+sHLfpRUjyWfM3Z8HtX4l7blGHNarPhF
3S/9QBxgRq+3nIqO/TXhCy21DvK9/YPpPGPYrZC3RcNwGM/kJ74caIAd/0oglTZx
evmiYyvY6eeuEu6QusOpLwHsWDfI9+qjupYVXXFbLl44s/IiGN1PjLn8/9iAfH/0
30CJEM+U1/nJYeaXKDVqnHFaHhC8acaYoqR3xmnIb9HBaLD0usSlEXxEb7oXGzTw
jCr/cG9FY/Zg4DrEjd2w5G6U5DUHFO0H7bDC/M2sPkqPDG175eeTIhrUNbWxBeBj
HocRupyUyt4jt3AVP+C5Ceiv+nP5aNatRYJRXYvuMQfni6Y1VmKzYJGY709NuHLr
OjtLPvtAdhuX1wfZc7j0tqhsoOzHR/himbF0Z070jicJc+W6UfuXYZF/Cv1vfwaN
F77+i2cKJJHa6PVaNBIxlRJX3CSBek2kbWfi/WJDhpUNuz5wwj0fRbYiqKcX925f
VfFxXU5eoDl/VtI5IuCxHR26LoATSjJAfLXng+7H4SSSm0v+z+DEF9vKwPozzt2q
NyNt3sNfy4DO12HgdJgxVnOqMhpkoHgpy0oOFT2IjL8VzdhTAqopHzkLciLr5piV
cH3EWNruyEwx7RKx7fzUUH4KJjdhv9rmRDA34/FqWKf8X5FktyDIxi5xq5Esle6W
1wRGhwJH2jvf/zcsph05Qvg3lVYQJVY9TdidLqcK9k+CyW//7XPysGyw/w+2koQZ
wkYCaORC+vDmWUJx8l+RH2D0fwF/zCp8BI3B6sKWYPxo7niH76hzq+SpogkzcwTH
naMD9GWPl1O+BPtJC/FfyzqPH/esjvuwAIKLqvVEuyN9MqlgpSGQ0qQOVHO5BNWg
KZo5Vyk9Gf6/6kCiXSD1qFEp3S26a4vhrVbJmnZwafSzWXih8WnAbfbb82z9zava
+rQCwWrwPAUnK1Zaodk5GKBbFbQrz+s5n+11monS1gRly8waSqydXeGUGvwPcLeu
NyaPM8xi7VEvkUryKNfiW+fBokcRqcgdmqOW4Th1QnN0rN+YHZ680o3aW56zueJW
G54ocbjlAVqyAOdUKyJ9XK/vMT+JzFr6XMkkhQvvQCQkuWPA84Ii+KewZdDnd+EB
aDGu7Qh8C3K6O7By1dkMgo2N/KIygib8P7UKhcIteuch2UFb7OElmQ6reIqQ576r
B5egxbqmP5JHCnOoOasG8Fu9cnhLjr5CSgSmnZHTc8QGBOhG9lkl97L9S0SGa+XV
uBUgS1i6eV1m1VmFn5XYinUzjjp0urV8R5z4OWDwUJXCUOIO44fDNEXsmSa6J4zj
U17mN01Nv7mEXdJm/Fw7tZRtiJFPYdaw8YEqTnI07kEDAFbObtAo8EUh0f55CWqd
7SZhd58IEyORBhZninuuSbwsjxIRbfDwEsfhB5ytrytznqD6ZWLLt88S8JElL+Od
E+a/GW0u9n1ky+4azkMzmZ9A2cDKOp/Xbh8aWuyBropfgBC1cKyPcl6cl9S1ljmt
1VRclpSNPSfcnmMCpo9YIuSOu/ivO8CqQZ2HEHWBsqnVse7EOR/3HoOnkfBE15bV
Fp4RHBsZYsjrrEWUvXyfe6mQ6ZV9jUk/mrEo+6vXClyk0d6YPhSq82sGdR0Rh2JE
mo9CZckvPeeq9pLJNrTzO8Gt9kWp+WTH0whsk2fkcpNKvtsII8205Hess8kZfJa6
iqYYeikICUFbZnl3FMeE/X4jTNtSHg/HtiFcNa6+xtNz0ECbs7et+2cfgkMXDZCC
eDRCjxP9LZ0FHUM5//1CG48u/UHyqnJApa9bNM560cZ7U+UhJju0A176Jj2jwqKw
ciZyuq6LN3rPMbhKKeUKPJeKAMAn5LGfNHXheFCeGF+AKCLzmPkqhYtMrYOs23E9
dRhx+eQI/v8E4QplL4FxuEUl1HFzT6xY6JvMPETgKb38BbWwRwtFnf6cIcIBhx5M
N/a4yP1j+aJo/hkwBthQdjGBPRHdGLYtbfoP80vgM26YxwDnCLUoGsSWCwCZJ4vk
7IH9ugpSy+Q7KDMHN13tpE5Y3qd5SZJmjgu0BH8wU8Hpljsl7Wod7oLK9+CxOnwb
E+vOi+AU7wqf+CPPSe2MX1tQI1/o4FlJnnxnc9y2CsPd7+6rOEmRP6yHDeTDkc5U
inwBXwu1f9YwyWiU7SqhaVJNOZfnzPI+WuIbw1i5VIpeuDmVgbaASakjEetPtqFa
NwrSv+C+R2rsAL4Kt79pOaIg+SF5O7MrRhubO1cA3Hf9rZevF/3hdhdqV16tt9nd
X079WkYqKrqEowrux8XY6PgTqli/esqEULsKaesVSnfgkquf9uRy7LXV0qpb17Sv
r5rWy238cA8RtRMkEyFhaxIAfjeG7/b9DBglyv+sIGJ47/dCEuNCS7yhBq/c0ZTy
7B7DSvV3VmWZzfSr3GwnpKD2hmYHQAFEued0mk7cmaTcWk4N0MDpm9K7O8e7LoP1
M830xSoPLh2qdbCPoBBQaYW2kUqWtEJuJD1jSpH9MUqiKSiCJO7u8nMF80aIh/7+
ootFGkke/qvrcmXFgkSiEkOCcY5ebdLXyC+hoNTDNBj2Rix20D/nYT/7X6fb4GEt
37rnftq/WjdF+FzhN0GJE1Lt12+qV8ksG/MgUf8uNfGI/yA+y142EAlCSx2w2boJ
2o7kpF/dR5RcgauUb1HXOHKfsfxMnfemSqBrEY2sgBJRRKOLHvuY1SOdKWYpJwkl
0ap/wVjFpxLV/Ijg4b0D0nrLCIAgu5ZPeTwqx0AggIaVNXasC3AuGBjVPz20OMPc
R0Sq8PNqCJ/8Isw5RYs5NjjrFBkk2jnrsz5f21KRRK81W+buSg7kLyQL9S293vVZ
lHzEcdhmBjRJT875+i7hT6t7+hBWzMkf+RaAWjkBnEJbnkkQBAf5tbtLnjWDrqEC
q+p8nknNzQVb5tEubjhay4O71+cb8+0Lapf5d4aeGQ8MePiqoDwKHeezn3gWW9Jd
oiIc0HaTd9EJ9p8wnvCoEsTJvOALBbi1lw+EYzbz0tiO51CG7dQqXclfDt+epZAb
Qj84kxr9OuKXrKXAMCr7kx5oFs2JTqvjutnC4rcP4E2N1Wk6Eo721v2Y6sRQjvhG
7FhdPZqabFTai7/xrmxKE/F7zA4BeaYA/B0oUdUpkBOuJcR3fqoTthXGdxT4zp1I
98Dwc3xzAoiYj5GdVa3sMawvNpvvucjfhr/IMe5BTnlRfb1foF0t9m1UhrWyLj8r
6DZW+mOZuz9GLq/c4+hh8mmJZ1wAC5Cxth350FBe41vb0Vt2INBN/ocbkJPFrFPW
tmLxnkGXfqgd4/1NhoDbDkzoixNPCHuax+F+kurX75vFtbXv8owPQ/PP5Qwqukiw
2pJio28PzZb3e+J+8SDcBwzsZjOow1QSKXk2A+E5R8DRpPj2NcTQ3IGv4tiMF/4F
GtY7DLxXO2XJ3cYxNYk3hm9ylzIQUCVEZtRXmtSbUEgg9CJ0mRLRxfER1W5HeHa4
db8QXy+jwFluG3o6H7ssLzyiBgsoa6Rjnd4uPZ4b7dh5FJfR8/0WA5Q8m4aIYcVV
8quwmQg/saKOInih8EeLegPZNmQvlLCp6QK/nHZf7XfyPuE1rSB/wAVn1NsEx6VC
pzKB6r5DOk/UGp10vuy/5+5X8G6HeOfTtbmZzNxzYwEJpbQ58OkXioMuObjT4xGr
F3R7xoRL+Omz4koQXk7a4jSXPddf40X7LqQbT5OyFgVCsEfsqxDIlbQ13EmVfgEn
LLUe60tfSWUDqhGnIbQmPva1FCZvQ8HWtOJT214oJsO2CHaxDuhLAVDAC3xInQSf
cCGYIQ39EIMu1if9ChpDJEcn/J2fdjsXojLMuwH8qEZj5N9PegJJ4gAJIji+bIqA
jaLavDxZOEng1PSjZ1G0mM+I1CbbszcSGQnZlPuT1OkOexH/WIxL/k2UWYlE1gsf
pMLhqX4H1PoSFM8z5uqwiFhHforFOTn7ReofEYI4c3ZfSLfN+kCuk7Joa0ZgHJiq
I4YQy8SbiCmWtzBl84cdGLRdsqzDgt7yQ0IGHSbOkOaTMVW3ohfhgifttR2pK2vI
hDuMD+RnbQyYE7I+dAWC8MLEGCc4OD4BWALFu1GOdDvw8VpEg3Up5Dfo9H7AI8S+
HXovtzxqlLsFIxzhf8dKnUkA33cyRjN6+eDY+xVQZjh/TWyQHnhO8ie1owwBnD38
fD/oTUA3XIgzlgTV0Rh09OeaI4LEajBBoPeZ2vQtJ8B5Et/12fxIhx0kY93isWXR
eNiBxWiAqLasY09Ht54K+Lkx1d4CYK618rVtjHmtaPB7boxP8iZAhI7sZHmxz8aF
Sq4MpiKf52KdszuQUCk8fGjtXbNGvPvZTB3SbbgkXBVAsrvhYeFFFz+XY5yS6rSc
Gq36UhV/hFyoZdk1y2lTqjfBgdOwqktjgOo3E+YLU6ahCBo58LWINgP5tS7Wa5g0
NLIlTcU7jwR8W2o7UP//gPkFrY/VL6iSiPu00a5PnQbtn9dfFnsEBxYDBvqyiCBD
RVz/6Mwqb1U4+qOvAvE3vqKekVTeHs7ZFleJKtuEqoGeNrtboE1OBPnuOB7MyEfk
QrMPYSvOkbKcbwXXAY4CloAt8XTQqaH5pa3/Wylf0GBeU1GoCKhZEoDExyoK/Ykb
RfpTqlLPh0bfqA2G/fxA1Vmg+jHQoot41/FRifWlOJjyCJUvPVOD1h7QgoXYFgjJ
I+CRGv0sXmu2Jm1PJLxA/cjNW7Yszamp3F8IF7j35E1D1x4TCu9Ebw3K6SKgo8+w
i47mprGVvzH2x1u2Nz2n/ajk9DJsoV4vNJuzRAOP2GEL7eVkPnWG7fnBFMJUnsi4
BX2xI8KyU4St2KeUmUowrhvqgvqH8E7xVaeFajph+ZuP/IN/+v4s7YArbbU54Tvr
tjDe3L4lfKVABlAJx6B+sxnBz0dmK7Efa5zARNZWnv1r7Cd+34Q8nl2r2WvKZg6s
jvC6ru+2AV1kRfE7Llz+w84TdKXukxKO7pnymrEBgTPLpOKJYdrsLhFKu9Wxd0+i
ut6KardJhp8rxdk38cyIG7cNTLOrGU7Zntet+OVLjuaEkAruyC9AbVFUsPrUZ6Td
2gnw6p7/mYFLm+nYmKvyEgMD5QM3gXfxghmZ8pPA3ek0iY/KMf2iixS6VSzlp2o8
ppmbr/wUG4JVgaCT9qM/JHJzAr64VNGklY53J6CLthIjzOEkRAZdLnGsj8VoMlB+
DJ5WDjpeRILKYbsPTrhRolXcn3R14+WtwjFZQXm4jBkVmKhXHRp1jFt4Uz+OQpmo
iTOIlu+ubNJxbx6+oq9ZvuWrQ93L/D7ph73ggBLAW6QueZXc8/cnWm1t/tO21WTr
7pKKRG52Y5uoqziyvp+5kSdnkyHhQ+SuhXUuuQWg32OQmOTU6f+XCBjholZOf9Iq
y9IAWkofjmARbya6E3M8KGH1YeJyLQIc9vIXGJl84v+vhUslobxZ+eSpX8dN7RJH
23YRi7FiPq/6G+bkmcODJMCuIHDaypkr4XaO8BHAC54M/iqXUWKczesVZ4uSDobm
5l6I0a1gUlxgtA83In4GGX8WvHsxu1HgRyAKHuTXhlKl4ZIl4awB/biq2/4tP8YQ
q76Gpd30cFea6+2wsKm1xXKFgFJsRsXgGbPo8cwXQew5ehZu4eNd315iYEx0r4V4
Kph7+SBlrtyuRtXuJkBUjnTMjk2dU64XtRiOUncdyWWuRVo06G7nKBkBb1qkKjno
chSYqnVGz34oYTYUh/mXUUCOkNHgcgBRO8tvrS9I+E+mCSY0vebLjQoY/zJJkpAO
RYbmDfazIWjuRV6+EVRi/wgLjvBu/aKlDSBw2JMXvlo8pLr6rXSYv4WlAxtfQPUQ
QupofJq4nq3cMOw0xImfoOoraD60mmt9RdBEsZzltUZSEVHtT8sTjOVy9ofTS7GL
0lg1AxwWX2pGALLOagioK+uoM2kY6tcKGkjaZbgF17eIgASdTiQSTY+Jg/ShOdM7
fTOGznlN5EAp5Tt/JRSCa1Rs+BGh04y2chOfwUiwqafD8qGd1FqpYrH0nO8F/TJi
DZplz4c7IYOKG08EL37eXzWN0poW7x6tUo2FJpIQMxEZTTzzH8KbaMKkNa0JyPVe
wDfmFkI9bgwmd1gj+GIRmuAKED/7Pgn+AWWKH6hrAXtdG8Bv7XbhxPLv7WmzxFOO
TMWRAHTeueQLxgWXkVMNmKSm+Ihgon75CyC7YuuJhen36krF92/FFE68k6oZXuGK
/DzAbYJXwlqSm4fegj2uLgc/ILQaHJjQUb5aUag2k1AU2FJr1O93qBsuBj689sSO
4iAEhyzH/5uraoffaa9iKCEdXy8C3KgYNJuTC2QCGqklSyqa3V60L8kRYgLMsukY
DEblqMG0+SLRQk5K256DxqNC9NkqaTYm2AJZkfY+znbocf4yCTRYEEYvqABmCABu
TvC17E9q6xRWtbMuAWrPrd9gfmQrIpwnoATCqv4QV9bz2YVPK+PvXrKTv7dq4jfZ
27ZFPWSKbYbSwkBzs7nTsnkPYorTimfnQVH4JK6ggrIjTfucLRLSlAjcfdqkTC+Z
krf1Q+ua1NULtDdT2TvrVjJ3YsT3HzH/mlg7XffPkDP0W+4korZmSm6xV7vsC1Dv
FKubnh1kUK2WVskwjiN1IsugY9HrcLvHOtrPbOzVEsb7svtRmIZF+ZNIl0CkmIRv
97dVCUu6xj/CTCUgcENbSHk1EoF3oJi13wZdESPMLzYLGyFhp7KQZBjvCwMbXRGl
WhV1Xvu8ufP46vaHNwe92Heq6W5F1yuamnrzCcJblnFMsocNPFYUl3QVHWtPXxxa
HHb+k/S6z65RGjg1lwzJ5utSq0YO0zWYFP2y4xEkrMmqH9tFQRt6gbLGZy45Nhag
8DEJZUJYQTlNbzTu4bETEjF7RUVEnZpMLfx0VjaoKFeZ1HLb/0Ef/NAMAdS+YiAe
7nuWF1mfG7/IQLqQ7iQenH5XHMQhe3ylpOxe7cMiC4KRwy3UeTZHDUtz7kaYmJxI
1ORMxrlUAS7Y23p9OrXFWF0XYpfyFip0Wx0Y+6RKHT+0+NyNXzJisqC9j9yZRmbo
DyqFRMDjEfVl5xsL+vF2Qf6tc8qNzKPCWIAHr0WbUeMDfCzEjCkl486NVCUvkiTb
tY3EUvTRtLba7YBugWnL2mNF6MmxhNmhooWwboxGFTb4yF6ncuGg4j9MmLQmg+yQ
xgkpmxkkQgw4q/fyazFhKK07K5mJxN2PwEwJo3+dMAn7yfUZf9kWlmAhMGVjHxSG
RSMqKO6XdtA57ZhiPRUVpQOK9cwTjxAcPgcFRn4A/C9J88pw+fbDAHM5ULsytnff
TohOPFvRQHDpWTvGIqM5ouYPaZmeU7pYUOL3jNfFnmkWpsIdHPyLAVXY+fiTY676
U7uFwzw68b1rVnqb5EY4sJgOAdASbcdBA1QmkKw6FtS9eS4az9xv7gPZwQx6CIlc
hFpYo9OJuqiqZj3Nn0dwJJs5qG5ceWtGvirQElaQM0qfeMjC98ArGbASiYhgMxo1
XWY3H4FTOiJR9mGJKaROXiW+KWdNxoe6Trbe/7ovioq2bFop6MGYtCyu6Jm7Qkr7
XUrSAzWkZCiuL1PWVKaG8e/J6r2fnzy4BNiQ9iPPyPlNHBMbAZ7LasVcYn2dRjzJ
Lm+Wj5R70dspR0VOEWonWM29IFb9nOTWR+yRvME8r63r61QHguF/SG/K4flG/3kv
oJo6wSxkThBcaPCS48daHoMOVo3B85o6RxE1zGLMmkEReX57ihfBHQpxK1sRNUYE
6tOIRW6aI2RV1r5KtkhCAbLpgtRWrdGyQZYbc2pWvto7hpTGWtCqzeXohIz0HZ5k
ILYzBHbIpSNQm61US82N2qkRjXypeTdFF9jhu5LFFAoEvoZN7o7/huvpX8Xq6ZzL
t9CQgNw9qy+OHya0T+khUeOXqIPZ2eCmvmRTJzPFiZOZkN2ih9g4BI0QMyzhpBTP
Npav8XkygHqVExL74ggeTIkt3YaVkL6Mc7gn0Kjkp95m22h6zZkyLAZ1kMBmeqDF
t+NVS65sZKYcB2Jb2g0Du3l0CBkqPiYRXZgNzjxpEp68CiGRRZ71CLUgfxkC5N5s
m2LqOuNewbSWr9WSqaN9VRHxnJjs3KxhF/AdSWGwQsMsyzGtIwGXSKflWfNpygDS
fxRyaQ3B7PlvPAFsJxSke9SA68LLVaX9RrRM8b7AtVP/zo/fsP8oINGuzICms4yi
NTmUtRXvvASiH3bOaZq7MT6IQwaJpUps0jKv59PB3AGQDEnGBtbLOhRn5ZhLGQm9
CPrx0HRsFlL+kl7/lZomdBQ6RESJ39EroXPg7gCnL5qBN4O2+kZaXprSXGI3rZ5P
5f/Pb/nT7cQVBdMishcnZjcWp3CkfRbrXVDzYbZRB4yrL1+qjI1hCVSrvBDIYb+e
VJ+phIOIrGZSQZR8S1Vi0BuAuyw1AxMmcbG64sLZdAgLFLqKaaZrMiXGQGkW/hSe
Q1yChrLb449BGbKZswAIJeIApJ3iS4xv2XBi0sceUtCMpltjGNP6VbnauRosU252
xvaYH5DZwb1QHxdgjapYPNUapyCl5PJdSks+iKBN1JtkV/P4h4hegKVCngyLP2yt
2IT+xkGoq7tr9tp0l4nnQskTnptGOlWpysT5UNYVKwerV/vvKTqpmC/8Ik3zQrAW
e2gqFotJ0qSohfbJkJuxCf25N4D+ukl13byJP3YLyf/xaBLp3xEHm/dVRe13a2bt
TU4ND6gk03b2RGGDn7hD+yMz9b7ohAYC4u2Vd5ngttOREx/igcH2gq6s9ofOUglX
RPEpd3K/9Snq7FgYH010S/izxbi1LX25pp0JtG/DCcxiW/INuN6PsTfLpueglfoT
E6bidrqCdSw0wddRt955TkYwyiCMIsxmZ0qJTTmUueJi+px7Y5MZhYwD/2a2ThIX
g35v9fjMofGJmtqZ99wY5us2E5HI3Gek4qydJkh12NkjTCsc8pVJQs2RMpahTcsD
dIAVdY+C+IpbiRO/txXynEJtm7UPLoZdMN6O4w5AAwL++9OJxM+/tPgsDSm4njw9
5AsOGVbEtd5n9JjGcm5adPHFp0LRVlPSH69a2Wo4QkTrpKLQmP4g62FSWvto88Bm
j6gCICfxNGkMtQBShgfKbeWwDlNFR5NupdfvRvZcnLn9zuwl2XwZevKKX43FV9tw
7FnN7xvg3sueHM0ZsEVeszyLWLYeRcrvakB6LEanSRLzNxI+azHebgzD6Qpy25An
QqyYgO0iV7C5VcjoZnnK6Cbqpant6qPzGRKdoM0M2HRhTft21VR3FaVk0k/fo5jL
EYL4NPGLIpAtOHdio/ksPrwJnL3i0orxo0C2xoWN6uWytfkakLWJWRHv1LcogZxH
r0gzSeaPbp/zWEluvkmBOvFyCl9E776F3ZWn2e0XydMf4T5p4zzpXgx+IAk5o+kh
MKjCzmpHG7JtOpNy3VhFmId1Qz/i+0Fuv8UtXhdDtGVnTcASK7gXM30n8lD1eOnb
Kr/UZkgswVh+Z4JUgj44b4s8PP60sEV8ilAt10oYrx9UTYMWKhKbVCR6L9NAYPil
sCxyDLRt+X1xK2hpl97zT9BLBoYQwdEWXWENJrLZ9n4XL8EgU7B69+XJd/pbo8Ev
/w1Z3FbfWh1a6qutgc5649GFc4ziiESeKHip6SygQbyLNZMrvgTCNAjGPUcoZkVg
lL09lPGQ2SCfnCwHUrqbRbnJe8CJU5xEXOvHD6N/LCM74t7K0m8l7UWWiasYD+T1
QxbkpWsjuUxVYyu6q/nCcNuc60pvG/MegR3cSLDso47foqBeK81s3Cl46kIsXn9G
liRZWz1CCdAN5B0i+yoS4PDj6+srzAwaMq42AncYSu64mEnPEdZMN0m8FLR4BX5Q
zH69YFR1kioCYP9BYPnIu3zthwpAy6sihDQ6+lZAglBtek3HtbPVJq1r9AA/rO+4
3OY5FL5xBQJVql291LEpqKUKlP22cRFZuLuScW/W2IwmCZ7jfwTcHro/gRuhNELx
n+AXhTkmS3ky3SdjoHHl2pjnsLoJPqYLwgoo9bOFceP8iLJMzOOZiSPQT6Texg2f
t3t1vrWE4+aiaPzjv/VFCN9tLzpmoFxNFfObVH4HC7HNnp8usmWKLNH54bsJsPJ0
4oarjwhday8FuivjU+i+RHueh0eXWzPuwHVmYUWAAXN+gCuRN9rPtj30f2EIgZda
Yj2hzQ78igxx1vu2lCAZhdVaejS+dlT0L6ggtd6k3w6fzY05VM75J/TwGi8YB5UK
hdJ7SnEi62CCFrR1Wgdf6bVFKUxdV8/XQGd0vdw4uS6WnHEwzY8M8TkECUZ5/rvH
JtJWNvqEpzZ8xWQsSfaB4rBHdsV1RS3H7+0UkDNGqo+3vh2DfJMRiJdGI+13CPdc
lwxAwzNMajc7kbV7yw9ASkKwkRk367nH8bHMI5iVqBQZpJTbGGykXW96UL4YSqpq
TJ4uilYIckfRIyWJVmcyPo41mWFbBPssBeiaL3KX7cD7mIOiy8kOwX9J5OfbxTpm
hRN/OryGgHPGDDJbMRvywlf4bpwMyRVfmZVANe7nFB7cSMKtoalD5/gU5htD9RTN
hld4JKRu6zeG9JqzHhMC0erNBdOiSXZfmLNAQUOYp2drpuDJo33z79vJJU01oKLm
wWMEFWDEyPaxIDtN3T4+akmVuaJ2Oko0EdgmeaFy4IeeGRTj1VjAUHypA/jzVhPy
XQI16Z1aa6HzWWfVmvNthqPclFdcjDawRM1cZF5T4wqmBlQpp1haCWTq6R6RgDYo
OWxikuA22rW+YDpjZpAUD75hOrK/6ZA9BfOL3ccLatNNIARP9vaAdKk4/ZTyx0kK
3+xgkFvWwQSlySx4YI2+QNqkZNQa/D3WiMPYCLeQBw0rzebH/8oOtZyCq07QcOl1
2HAFwo984s0bb2jbVoDYdmjsMi9EmbhU2hN700ftlelqTyD5wSft6uunARTMO5El
MzQqiE1qXPGV385n6gz9VPmeP6GRBtLBJEztgFL+qtH3qSdxfbCdT48aMPRva62w
JREbM0nYYXcTkBQ2PNWW7WCtemNb4kIKW2Ficc5/i3jX1+jW2sS2UOf4Lsrxr3dm
sDTpACDnrU2ul8VGzDpAxoIw7TMzFYLXQENME3QT9WderOPDipX5EiiKB3xhyo5Z
1LuqYghAq4HcKQB6tfxyBi2RtzZW3lE9RheAEPDZELtRFucJgocWYWBmQmFaoDDp
D2CJ3fmOoAweICVhiri0KmrE3QvR2L0GzzbA2/J4CPtWijK0ujsYBUAhy/i+kmSE
EezQm4CoHErE6qX6hF7OCdTyHUwFWeDXlDgYHONt1rIiVVOTVahiSKELq8KL9uxu
bUzrKZ6pkYkXwb9TICpjAavPhIHEWGi5kt5G8ErPk2BDo2UC07zbXqDTU4oM/c4q
pQOR/uMKcgxFnue0OsUAKihVvDmte5aJzdCJFixsSl+OGXR3Nc+BWAuA8N56JPD7
4jbhe3FITYEVNDVF7Z2Rg7o6Ynbt9UdXWaM3Fww622sosjWDZopCdDggyQxjocAu
1NjEKhH2WvV4p/Gh+ffukhlg7ZaebjSjjLwfIUwcPhvMy0rkcMVv350sQ1ZK+UN2
wgBPsTG1quNT3V+N8PBfor49SMcVjeOLX9QLA2U4VuEKrmefQOYhjujQufOcGIpR
e56JsngtzvLpAgSnkXP/Xc3VaGLmhq8AadyUlZun1xJK7/FlXfjfUGPfJbRD3xqX
WAwIxr1Yq61gT8LLN6kUvPn3nDztpgBkKJ8QLgUvYX4Jg7GLg+x9uQvAA+GbN099
skL2MCH+lpPUiajQkUTm+LgVye3U+q4l0VgyYQdz68B93iHAKT30Q0k+0chWIXzk
yGEvcYBGcrXaAX+yvwhlVkTuORahv6QNuRW1k3oVioy20N1MZjYL7AVYH/D+jSQZ
oZJEUu2D9I66M/eXjJ+b8V6gFnmlR4J8eRzdNyG2Nw4dJWok7gQQUlEvgCpAjYsx
91o99OR9EU0GgaXm1kQxgTSbBVwZmFzs++jF34fUlXBGIo8QyFozi5fhw//e629J
duT77FgRcRgDor/wSc2pKFcZIy2gJAJeH/S0pT84xpgdVKVgDRJlX8ptJnW1dkLz
hbwmcJofGDO/fbt4hk1WnO0LLSup2u8qUyY4XSPwbodOGX1/jO27kuH94UcRMdlp
eLe6DcTTbB+illM2KlAho8JYW/vXXpmSG2Tw+0XCz7z4dTiuuq5YtPcQ1i8YbUr7
a9A857PPOu1W6fqybT3ov7adxqXdL0pMGrMnGGehyKyt5D+iwsXaqDnIMWPmoyD6
akdmB+2BJ6monr+HHvA+fga6S2+mgrVGkoN7pbt8SN5kuwwR5c8JLNH0V9MOFLnY
dKcajOgH+T5rfltbuZ0RxcMi5NOJnrNTGpBwjbQ6wu/hgDlwlwtcZ+PCAnvAS0Hh
jS7FaEnj9TPrVMjyhL6qiC5fw4ymNB/szKqYJ829QG1FVjyMzaX0qnrdjTWVRr0P
62bzRru/wIQiI+9sH+Fb3tFVkYxp102lw+mboi2nm7i8Pw4jQ5iydnA9P2H3zqAi
PW+PvmLFZfLJuSpnQB7JT4sqX+1AG5fSwvqOvhhHYd1xaZWfAp18jKwcMSlFtT6L
AbpcLmSb6SCOEzrX4xGwmpS2wzBHHc1WAHo1appWfN7d8deVuFmb+mdihO/0WjUG
DVC/ksxiv1RvkHsO+vCVrZN8jb1lBsXI4vHKfq+Ojd3WFz5U29N6bQF0Q8aNov3F
qHpJxFxRkcgd70BHlkGEX2tGaLjIV92U2ruiUuVC80j4AogXihNZ2p7j0I8/3wdA
pxMWLDYe7lhOEnhabOVcTUgyHQYC5d68jIYeNXbcw+Zty2jTZO0Ov87YDy/dy34Y
uUDuICmBU6lX82A7ZbRGQQObvYmlfLKflDo/odqzMW7q3y+3DRbt0ClzS9l25jvT
hU/mj5kdO+A8ZyEfFfR7EBa/MTdjGHMgWuXrHgs/8VTcqk3bPSCMrMIG9V7ZrbmE
NwrgF1YoA9tRSL08xOxge4IS8+GxC2wPIgRuIc9B8KjW5EH4iIR48xn7cB0oo1gR
dbvWVOy6VDvwRI7atzm/VXhJB5KHV0jhVquRcoWSK7B+myynedH0RSuC04wN5iiz
u2rcGEZZZxuvHouJDXjNpgY/V9g88jguBp+bPOvWpQCDCpltNPKGZzue13x+YKHs
+dahHmRHqXVFsuQkG/ctntt3RbvqilttHaUK9M7xWS0T0hAC9ZXHNk4Ggm4Le3Bn
H8KbKIq9JaDlDppalEbB1QqXdYhidwgZCAOS9NODzugrEfwHONm2Hx90w4uV832V
n7zs+gOmCDmrDIhy20O/egbGXx8skBvMx36J2wKNJjf0TSfRLb1AgS1u8/yZMt27
f8YyUYam3lVSfYt2OF6wK0S4kzw0IbmjaRVskuwxHFT1HiLT5olTHTKABG7W+6A8
h61kWMWfyWFeaqHXto1C7mfdUwumbyrIRilVNONa3n/nE4cJuivB6UXBCcZGLQpT
0Co9ZmEFc8G7bH7Q73CruOw7X0aqli3uTsRGajVEv0xQkIQ/pliodjikwGZ5fJIw
wwdG8SIW0msPDjDg4mqyU1qqGv69nPutNs42OQOuf8g7f0skjbnTW795cfL2Lwm7
QQW5N4wtBFYIVlt9pKQ/8OeaJqtWN7Yct6LkhL8QR5VglYTnaWExTGDCVSTlS/k3
uA58Nf15cepo5dv5YlknTIt40uuV9leq/5sgWTFeEHfX0J1WHLrdUfMvQsIhk5fT
QtEbiG80ClEHUvEGqSjDifHObiHeVGK75LTw6VdHfUQcTC8b+4fDwFNRmcnPvp9I
D9gfq1FobXWiFkXevX8vA3DXdFjp11E2TTUeO0jGmpsos4qe4j3a6rddbmJmOz0b
eMQiYdIuwj5YWsD/gQnKxmmo3ZH32QhQN/l9DVOcmu1hnAWMbo5tUSARt5S/Cif/
PajL8rCm/yjCi79OYg8tbwdVzZFGnwFNt5NNRmYHLhK568mcQgnFfHgBLIo3jcdj
7SGk53EVobF+QrhJes850P4oA9TSNZuoqycvZp+hTfZHyQXp14SyT6gcH/flF2Ii
BDg5dbEvFzhzz1SZFVTTkzHfS+81Nwl45ial1uKHRUAKFCLVVB4qpPcMwOgkC37X
GGo+pKxC3CrW50yZwmiuH0Y0fk9uvF4376G7P4j/NJOtH+GqU6QuFVzP/p0SkGp8
kGTbotGoRMCTGCEtdFFd1KfdN2QfXiutK9ARPCZMCgUNAgSabHeRg1cd9NizNsMj
2+SMfKz6PqI3AWS1eAGPaj9QrSx/UBBwtcSq3TQVyzU57JE5A1rIkzXOQIRkeJmM
IYz6iUo/t+W8DFWu/sNLG77tssrSZmMzbQqsHzZ+2hAd6YWtI6Ewtv/0P75e6Mql
3wANga6Sc2SiduQ2XeGBk21Dm2aEqHMYi73wN0+sn2ONySPB1DNT8CDWUpbvf3ot
BH6a8ZMbBak2zanXCjTsbJZzTIA4IFjdBgLG/XRpkI6g5tyNb5l7UKnqZ3bcssJ9
7/uHVGPrEAOPBvRGxGf3IRggRSW7SnuQMpjMK6KBvQ0ZlJ0QuPzRhF27tpjpv7od
OUUGvOiUVzlrRLMilURbN2oeLAScVbr0jCGuHUplIBOM3E+Tj+iKqkb0wkSzItTA
kIjIIv4eoO1fm4X96dg9etTQwHsogdU8nGUD4Lzc304egnKj6nfIlGaz3gzPE/fI
bSTKENEbKfrE2eHBaq2SuqT3giT835LjecPu7WuPITtI8WFTY44CdFxZe6Rxau3x
mdexH6Bm3jYuZz0C04X6+PST2qvB85xhAcAshXCfjrCYhhJbxGtFqQP7sF9PoFbe
xtE/PIKFa7z+/ERGIWtm4MpWS2TN8+SbVtPEePOJvchsJgN+xP8AJwU+3sy9VZv7
vO6811L9HPiRFhcgTr0nkyMZcYvZWZdLjIgsAvDMCxNo1pGkOe7r/1YfKuB87ETA
3+yGOUN5a4kSaNvxLQYxdtXV1PFapqeTX34T0oZAywQv45hh29uyKWMkan0BSDJ8
g10rXi7d72CzBI3I28BYyEoOnQHpWHE6m8RzozghACQzy1ZBwny2MihoNlGeqp9r
6oZFUNxPQbyCDWiMPilVFScJvVoQ3NYjkOKORXrJv0U3oO4865sigjs9UaNQBSA2
yBMY39HFjsECUpvthQoqkAMIJ8cAVml628RdsgaUpyXNcNXxxiBsBn+DIvC60trv
a6MZZAKKkZBhM9wqUQ12gEr3p4MPSUGZhI1YP4ZkEpN5ThFBk+RCIvWSbMfQqWPp
L7YRil2P9WKCUcCL5dqC0/mG+yQAsjgOMzLTfHBP4p8IcZbv+M7owTt4i2QDjjaO
wABXaHLL+bZwna2aw/O5legOtiRMohIs511VyB9Z7X5vxwvsvKaCJE751uEE8B8p
fAnqNuESa3AGPwKK+eEUxfQ0Fu912Qhjas8b+3hMeh+LIsG1yfCTwZ6PVo1twPjz
/6EYUS6R/KVYZgA+az7Ll+FYRbV3uWUNwXCIWHWPkAJgwj/V2LqK6Xkz/spUeTXY
qcKHq5h0kwSmo5VJHHys2xUIBtJYEs6Sw//gbS+6LZj4ZRMeWLI07eMOW2yDTpgx
1nv0Bg9diXX3cXBDhcV89qVTe7vPV0kWDfl+N3KkzTyK4AImTnDBvPnZfILORLg9
U+IQTCm9mx6e+NElEQOUbdDWnwbJ2OIOkF/pI9BU0SjLafKsMGwWKBfmEs9tjeKZ
gtX+XvhBnGOxhcNW2Y7unfg6XAKBBnYADbm/wxiRmanKmldcOTLyflh/vMn3GM42
o8ZfLsmINPUGn2cO36jfO7VCWEa+AImFpoZ7exQ2WfuI0fRHwccGoK1PW8eJSw8h
tUXX7izWhQhqlsPuyyk95Mk6iJzZ60zEzEcMhvewsrxnFy08h65LcNlhUKQVbZ9y
XAGtsZkLaBpeCzYvyErRfqbXoSEP0P8Y96KjEtslztgFBQum2kuTA+xJ60zEmJnx
slvvrz6IOW5SIR2bY/hb+TO99eRkGt7Q7hElJOEkplDBP1H05OhMXTJIZjPWVFHb
jZkADX9HsXeMWS4eP0gM38q+xhXNm+O1NYi6JOQvzIUPbkAeLwzFs265FXq7r3RN
X0oCqsC7JaPb7X004XDUDuia7wMTwP5GjokQ5g1eQ0NgpRA/v1SYVK9Tlv9XgGBK
CDpMIxnXsg14hmLsTn9dWunGNXafQCAr9lkrQ+xGOJvJ8zYxsfBgvVaukaTnFxXq
B9CzDDgnmuz/zrrilO3L9w7dFWgDCmf+WL5er7tLBClu3wsD+ogBr+j3oD//rrzk
TzhnlONMHMrTo+gxXpsPSMP5NV9VsIsqOXWrenWQ4dtqd3TqskY1e17tlRlW3e36
Vg/xL3uAjbujVeVLau+zRXQpYnqJDbtz0YVS/pA9ed/4BodFBjYkJJWUVy9KmhFG
JRosfInAGoXhf6OPViZpkh17N2SNzQ78M1wpKMoYDKgYeXBWdPGQdQfIQdtMLZMK
aFFaq3uohRPSYuCX/NaWI0iLmJmfsFdlmF5CYkeiqAHQvsL/olX9qAoSOP8Dwyfg
5qFpeEWOOWmZ2UntCTMRLouoM1IvRnGg6vWaGV8VFu/+R1cwpHkk7sJwSCHztJlS
mtI+udGngMRK7uxud7bn1yNLxJz2JKjxYK6U7p9w3/yXtnin65EIxwFVw6X9kLuL
dAe1k4WgO0hSBG2ycLXzB/v9abx4eBJep6CnzBr2xyNR3sV3CKiMHYS1XEANAw3G
Zd/syyCAyvlw26tFy8RdR3Y39DXLkih7Xx4/C+lo0Gr3ctHtFrCtVNZJeZ8ZoDl2
oCZs4NWFdxAKUm2miXoOvYrSDolAgmDHUxxrI1wKPcIaLa07fZparzaO5oSTNQU2
aA/sZulGp+j+X2oXBc3e9xqHkw0yvfeskZBAiM2eJdhMW9o7wKr/G6/uksK0gRKB
vLgA08FaljpdA/nkVG2p5sCXH7QiTAhQxAwvDJtxsg4x/89AShl4qbStPLYe+E0L
8I0A/o+1De7l3DF6OAg5Gd4XonMzWChqtwmie+YBROmVVghp2w91upZSFT+XWR2z
/eR9rN35U/YnDvjB5KjfnOKmIKafvaNA+On3Z39YPjaHKf3giL7q5yixvv76bXfJ
qVa8VcOTeNnUWoRJ8ZvzDiBLuBgcsAXXKh9cJ1cGQu3tjvy9mqCFg5TV77NRGabD
Dser80gFTDKd3UoFQefCog1BxBh3PgQ22CEg4hl5yETTfGHVKj6urPlNuILUpzjx
LkN03HWP5gl/uqHSzJNIUEZjzY0lgefcOQsH/pmERopaEsS+IsvzUF8p//Iq8OKy
RzLc2FdNoW+idwSTzi5Xd9krPKIQq+ZIWB67340W2v6Y6z+lO6T2WH10PSEMV+Tm
Srb7LadQG4q8nk4YZk8+lqS2xAuR9WS3qG/v0s4bbfAaUTx4wGcccGbrYP7MYr0Q
aW1SKX8Yd1S61X5mIj5spgnVqEoKIkKS07WEWyHUfkPmsctZ6r9GqlLZ3JiE+MUF
rqJF04mZFfA2TgdEDGve3FSbuFN0YoXeaktCdwHf9IZoXt2vXU/0tLuaesOxtQaU
VyEFmyR+1VNtk+Cvt/BAaNZGtOxjrvcDvP9zGI/in47rdWtwFcbH+KQgpX9tKxil
Tc3vb+VkiiCuLv1pLJB/2IStYnQCo7dxKU5ZgwIBc06UYp73KgFAoLlVRmQp9zy+
5WHRE8N1CTkBCygFq4m3vr5nydUnNXvM2FU6D4huB2G8KasKbVwiglvrzmLthw2q
V9m/XkR3TpJ8cTVX+KQzpb4fn8PeLDLU2sGiz/6bxRR2i300gWGuVOW5RaUgtvFm
6kaNJ+tzYQMUrKhA2KpgWbaqcFAnDmIxVhqWzNVc/HEsVk/g4q8WKoCs+MRTB+eT
cwsy+oU4JxHNP3Q6MWwaLS7dGk3GPSojuasoTXQAxyx6pvyvOfwV50loNQ4V+1T5
pot9rgyy/MQmddZXObJlDKBJaou904vKlLAR4/EK3o6VbGSlAduqoe6Y+Y0ce3cs
M54Y+MJn7bOS19GqOwAFeDgeAVWH7eAGcZ4XqlgqRFtye081VTXJQF9Xkdx/eC5C
E/QfJiZFWXtewO7NfTp3fW6u/bvraPbDWESrsD/f0Lcl80UXHaQ5Z7kqZCzoJn1H
haSyzKA0h/vnH9I6x0IJNifQPyOZemWdwC0R+v70bT4FlCihqT377aH9h+zV9yy5
9Kaga5UqFjYx0cMbAXfDrr4La3Qcbfskp7s1Vfy3VwRCaVqRQFXhgdt9zIxO7G61
R82FxqTWpdeohjk5iYcKdH5fLC8LXwCDDn457EN9FItWzImxDaX4oEg8vz8f8srd
vcS3oL8UzZNHtmm5Vl8mNBsK0VDeFSIQcOUl6UZm/w8Kb4KDQ2cSItdTRGRLO7co
qUUQsaCsH0LH2xvh0p6KZnusfw7i96FeuMF2gudQTqvy5DMJWtkzZHejVph68MPp
YWqpJmGvQ4QsckHo74XwyKV06L1Qeso+vGNtMtG/QibVc3l/KvTYy8AII6k8937y
yjeSzl8p0MTI+4s2hFmKL9JxUOXu9AE0ekAGelkRGNClntI1vgWnuaTOy2AC5iDO
bvDHmFRNnBxqaIcV0f8Taib6bwkuurll+P9i1xtvVfsQXdmi2nvLsDuYVbx1r3MW
GSyBXL5e0qEQVkylR3Fiou7qtU6L25dxyfs2Gq1plT4rxJBzEq+Q8oNE2x7smTYZ
sBXW3qc+6NTfW0WsDM/vQtYmmWvaVs5D3LPSGJ4R0hHIzh2oFH46RisEbmW12E7B
ltszK/W+nvQ3TDX8ZSn0bcZhDybG/ZOmliu4ohE+o6DfGVGNZ1fvN3yEekP8QThr
LULO2LFXj28GI+mXhneiiU8uly8uRP9AuhdFbP2jhKRGssCESIzRIV4K3Gc6Kclq
Aza1hScnE1kF4uFzoP76/OAhqz6yZpPZyQT+4jSUaDQBd9u3xF+orBGVUdfNQR/0
YwEv7Cko7edqCEI2eHbaXRn1Juhq7DuicdgT9mtdwshSL5wYSQrMlDCVoepYzWQ5
JFNidV9x4TY3oCn9RhYqE7Qro/6YEGmappvYAQjnO0jyItC2f/rYQtsam9qyt76p
iGRRnZFEXxLw///VMbyctSIFjN2Z53nFW7MelJ/U0jLt4KkdJH3tIEK0xyRTQ7KI
JcVIL4RtkeJ04kbeANLiqy6U6v+OwAJOIkUkguXbkDLrJCBMQflHmkNe+zYmNF1F
YtEf5Fqw0PRcqmCXePRxdw/NDzXI8vRjF65Ewv8iuZVB1hU2cZpYhTIdzIfHTJHp
LkaXNUpg/pIwCnkrDbY8aF70BX3jj+JIGEP08kwF5Y3T006rQRNL+3X7G+HUIxYt
L6ATASflWseulPyjrc7LJvNiLS15V//SYpWKh6WgVXiCExUVlLHoPYuBL6IYiK+a
YT2leEkrlBQ3I4HqpSuG+NVp/GzJhDRHIg16SsHTn/oY5SRtyiAh3/bHtez6swTz
vP5StkSvNjzsYUyeJ9aOdwq2KySoBhk5pTGhwyBWWIdw+4ektnMmtMJMTp+3SEOo
0lV1PUy2tNxMILatb7g1DDu3Jpu1ep5g0mjTUELtyiz9a1pbRlH7d4iNvmBwpw26
jgTplfh6wN5JLYJjF0zyd8xQBoS6sDxizeifDl8iVaDySh2/0lK7kHxkGSCgq9cO
VqehvW3RiFyu1jrv6JAjyRid7qzAsfpvX/Nk+JeqHmlWCq6RbBMam9UHP2q/0bEL
fZaOFrV8NTC0fd3oDgMldVM+FLetd06byYcnaq1uQvt2QH7GyE4xKly0mbvF90q3
5fjNWHU3qdwx16XVuB6PbJ/MtcwBkN51SUleNIpta4YPYSf459DRPABep3+05Y/S
+giI+LxKIOM4HhjS8s+lBy7SE6pY+HIXVF3uTvRGz7t18vlufGyJBRRTxdzPRS0R
JAdiDuaeE1P/KjBhH1GPODIFxRGarOSFL/YExJ/puQYjAUaKBZNNXa6rRdjmzkmB
OVxrq4oZ5FbUR9XHYkn5bKxYQzvkZsBNydVO2t0+ZB01p12SUgcWSanwzPAPNfyj
/sMkzXYkExD0H4QyreHdg3raXNPmSkzAY72julxQoCgL3ush4L3g1oXaaDX7L7zL
DBFRrdGJgRNnLpAxyQIDvvx2nuhqNqvkborVPIe7m893VL0P+UZFA0SaHlq/doif
v3i5sBXteOxaGVvu+JlyQFtMZB1QqlO5Z7vPiywikyBx53++kH80mhW8bdIGk86l
Yyrw66S1/+VYoTw/+gMo1k6+QQdNags+Cw4vPMDGVsCYRCPzPpbkIbBDqaYft3cQ
NnK9Jgdaclb8k7ZoeZm+sZ6RAdjlsqQOM3cixIHpowaxAyyOQH0LHTgvgOmMdUKa
CJjDIXnFKohK0GSs79CDsF/sHYIHzHWCLiri7bK0sI2fr3JgE0hKi+ZG7/h3K7Tx
ZIek20+8NxUHJUggrYV5GgBliFsAqKSkXH7Se54bZ1V1KcnWgxyfTc8lyniw91sh
y/JE0eaL/kqtjrr1tbCqFEicU4LnDh9KbEsVhfV1v3uFwNUwK00y9/TOsKMmOehT
l6/zZ0veNTUUn0hA9xicASxXMK1z/6RdHTWD7xzjPbB0LSmh+2qs44l982kdNe2B
afxpX6EtSFm/VTSR9DcyeDjjPVB/JKYgZtHHbqD5lzuFcwNWHLmyt1cXh3Ejknr0
igHyCeFPI32g0PRf+iZU7Z7qVGFqBOiYRcv9iSg594vJYbhKqFF+dl8Rhy3pSGK+
ksn+SDGq7MREEufG8cGxfIv93Df0JWMUbAp/GtxM+oXfOYrzRHgre+W4fJLb6ewg
lY44q34qWfvrawa0ha3TNio9D3KjN8DE9ZgrLU/8swHikO5oqx7RsFwXwenreCho
VODeFMU831A7tS6VCaG6ah+Pg6EqerihZjST4OVprz95rbQpyoU6GTRwE/6uXtrM
mbWITPYRpkgnj2qFvelPHt+2tC01J9bxXBoPnQyLptO4PIRJwZfsu57ffARHAHJQ
tDhfcjMvUFSEn5097RlhTzXx38SAay13h3SBe4gvs6WXF1HGUqioL0vL8qqfFtBf
B8CbuqC94YSR/A7nUe4aSdfIxCgDxl3bDZ37akRqc4Zd3p/iisx1l5AUSljDv+xj
GD9eyi3yl4GqsuvDQ8nz7Idk9yL1hJbZ5fdciTAsE4Y3e4jRuwc6C5/HnXh8hQ0R
7vOgKqy/4I1Rrt6O7LorZxBAgAtP4Sx44FpH+6h0vxGzWieWXuu4JBRel4ipY5hG
/yxi0GuROmvmdULr0WTVFk2AtPEoDNn9ZhE36Yj9Z6Q2XjeUx3rywkz19sia1n4R
tjQW13sXhA4+4UfVbvtv/TbdFIdtDhX0PjHl1Ws7vPIJOk/+fx8xdLC0cliN9kiE
xh1gNUi5fDYkzv2XaeyirFvbWI/ecNCv3I1dHucsAutrUleA9s7Rf5uU7UAqmNgF
L9C2cqVbThc7uo9TVZfqsET+M9gSOJ4pOdAjfNKQSkZ5P69clanUqM59Nws9bZ1Q
BRwrtJBX//s/Dfz0xoK/JtUlchiu4HZw+HCM8jHgR9pjcWSGVF+TbTJpPEFNeEuQ
VXhyDu7lTvA5fjiKTszsHFk/9YCD2WXyqMpwn7qazshBUyvvjLsfk2Y7U4Ck/1CH
OQJt5w4TQdG02pCum7zlTKsTcpVjh+Wr+wDrRGjopDWcTTZMo5v2wmkrXQUQIH75
ZIcfcjlM+Gg4/AAeuKQQHXeJ5ZHRQ1oZQexxEudZ6d7m2KVgOMdcKFq457bFnBKh
r/zupBDP/gKjYqxKwN3oz+IiA/RCVOBQYlc50Kd88SMDhbfhzIPuOCkth3LkkrgH
T3D+1pxAVvJpEpl0VDrbh/+JEdHottgJgOHmUdsx1Y8w0KOb97H0Dsvinm2vOKTm
sxVYO4Ie700ldLc6xR8wcwN03UJesBxsPU1XAhfBsRvy/oYWK3gp8j4KD3uGbS0P
ApQnBKi6jusWw6jEmvoTJPipNjFeWgSzIqmud7eY2al4pKmFJ+P+9yuxbKJRFRKZ
UZbJtJ5qCfhejCEALVZ3D5It0jYRBWe1Wit7iJ4QAWY4Y+0Uhrx///ZUbukSjdJ8
ceP9YytRq7aEIfi6N3vCcc4LjWl1P1ZEnYhI7KMQ8zZE1LpQf+FPZ9jP/TWHhIjG
wpzQPcKLfJv+mYxCSafzLRA2G/d2t3w1mpR0VP0r+eoDCXQqovpLratXZ7iv51CU
lrWeu/SVHxUgzxQgnCfe5NshjLDLUvmO23ivRDrVJI9JVWYQYa4XnHTG6nb3HS6/
dOdsJ47Nt8Cf5+D1R3vvjpsPwUtRHakbqJrZoYFpZvMhUEdwCFLAzCBr5VW2z9iK
shSJdRbc3YXSfvpmTOoxoeeiNLJIzrJBChsEK7urFXbKO6W5CFtDwn5y3p150phw
pVCvMUqTFM0s6W12UJeKidlS79W9zL0N/M5EVN0fFZQO8JSgHysjxvNhs2FFvbe8
okit+26iw6XYspJ1I3O2BHQfWm3dqjm9ON96/FFAhshzIdR3QGoXpce3j+G3IQFO
rxx0Iyd5sHg1j7YB0zluHZp+gUYIHD2P64vuoobbhLe8C08mTg8VWeFLopwRilqD
/ObXxlNj1xXwEz0SX/2Cn6iMz+iu59ebpCUAbdfBPW2GdjH+b49d7UtbZGo2OOzK
cwTD3bOgZujDJt8ZqN9H5DYuBHnH+ygZg2KAkxRIW9OXwoA37Lqyw++DvOUC8bZC
DBKeDeZr6WBPqmoHjNYeDV21ELLfHePqwBWB3jTO9I5VSKQTl5zjAafpcpm7Wn3V
k4F4E/3IkP7eoODBR8mMQP2WHQdkkN7OmKtA+J0iPlHu2J9JfXe/wAET+XDItpae
x729n1a5WGipWrCDhjUL49LqQvGAaZJCdmmj1hJxMBgkxA52d6N7haa76pyKkNim
MsUzlD+TV5WVnFXg87PbNxatX19AN8eGica/YhTm2FddlQ2YrS4cptpWCIcT/qo8
lWJBL7wmfaxJLTDcFzVq7JKgFm3yhuTXA5V6OCgtt7SMw6XL2vYdGzHT8bn3OEU7
3dQdkgYoTbemZHyVkxrQp/en/tQ2TnK+FGpfKosIaX6NWcKk57TOhvipDDbCBC1j
NmQxQRgOPxM5ZKg0N62DsWbpEWcYRnM6tqGm83QsEqsep+dw8qXXp+uZZ6tymCpj
+D7XJHO+MeFw+6Sb74DuUOqzZ95XFG9lBeRmGSOLaYMJIz0tK9Xvaouw1KncNqOa
A8JY3Jx0InutfccEUZm4qV3RVkX/Bqp7cFpTBoJXBBmN2iRRh4OzdrImTYlIRvdb
EI5/x5jC6jTWEBUIU5MTbt5UC5qM3gTcoqCVL3d8tkGOnaNcrZXmd4HCno6ek7Bt
hXL5VH9BZVKUTncKjGgJRmbGW7rOpVVAvl0HCzac0OCGYX4W0oGH9auSe9v09Dga
IzOC4FdSRJkzkN81pBzjkkF0RHJlDsPWETlpwHyuUriH/7vNeAMZmy92+oqiPZSt
QIqQbc2QD8KrAFij6gBHjyZkeMoNKV7ShVNEpBRMqiPSh4nt8RL7xYNluY4h3OlN
i4ncj7E3C7dmPRqfOafADJXYSa4/UAkgF1kRyB/I/0Zq6Edo67twe179hqOwEC41
5TAANG4O47ctmO1DqpdMgchbOk/MhZ8jhartyKBZTXvLfi7nL0Tiv98l23HrQKvn
o+ZMsx1IBAckfUEf2MeJdfNre+xewt0qI2zN/n6Jn62L8t/hSdoZ2afbspTVdbKe
E1tCP1aU7fw/6HzS2q7yqM8iUS3Xbe8B2a1NyqPx7sXQAMVQhQ98cARAPED2Cu+S
oWrLB9+SU4/rZeGKlAoIrfaeQBF7wfgWvEqvqlMqqlwEW/3GSyXqivHiqYYTn6PU
JP8pBylq0qBeijQ6LY2ZySoj9GgJ3qn/31h7CbqMyxZzm7Id8wYbw9R02eXcrAZF
/SMneYzKayzWItqGmz+gcJ/00jLaS1tmBsFLx7JrengNgC0/6C0o5rkHODTrieyF
P3yzIhSwC08D3GsxMYMIw1tbDCtHYTYKT0GcAMqHr48ZkWxlK8eMhKTqsLJQ7EGc
sySJJExnrvRS43NuMxYCa6ywMpYb7I3ZsxHwibJB09Yr7MFIn/80wZXGy/ziWZM4
9NSKen6STNVXO3Lg2H51JbjxoXTHuDjgyAcDFyHpJmYSmS4REG0Ktk0VTYOciZ6K
HrtcnnPPmvONiatHCnYtt6V4R/y9RcrrKtr+ZK6fUKulCCriNLMnHuisMrrb74Iq
wyVX4iCRqYk6C3Hihfh0lEbUb0ZJmniQSgVjjvhYpjfZGoZE5O98nXMgKiKs9QVJ
BdQydwQxWLNg4e/pzVALQr93eawOgezBqNSZ7/GCVKeJXgbN9RybIWW5R4vQlp6U
PemSqldaEeC9ZDoaj0TnKlT7seb0dsScdGaje/gz/L8ASGqfm6o1NA8lpOwVsNyl
RHQ4ccjPM6aOCkYJnMH9leqyC6fmdQvBCbRvUosqgU4u1v5++23XEOCrLdGAOPO8
SweSAW+0whHhZOasZcX5V/zws56vLR1D8F60+DOMBzp+NkMgPcszJ9FqnYNIc1Vl
I90Hhv7gWjBK+S3walVhcFUBCK/Q8INkDapLOX0bFyiwm0QfdLP3eDF5K3ua4X2M
WUcxGHl7wrCdSY6PQm5mZCkhdpcN+M3jiZdv8i8C4dedAgnoG0vpcJXxN4pVC6jU
KGnHdvLwqSM7Q3PxhYylbMV0gC26BXziD65zGgbVKln/Zn+45ulwR0cZFrwx2YAB
VnEFsxYvzzHJp+Uge6eFkJysE4jA2EnmRomqOsC853kmzhE/B3qirpjlmty8CLsS
4wIObZz717jiwm66tljY6OTY3XrGlNtFOOHauB9G/XLAfxwqDaM4L6ggBwdsGWV1
rmblxeUAn1bfbDawCvmvkNA3Hgnsn4bzL2jE427028n512deKG1pJXwbn41M11FQ
zcISeD4a30aocPyp/hI/2759Knss+WAHl4c7e8p7U4WKNtjNQHgHVQbPkqwLxopR
4NTubCZUg2JiupF6fekjxytJ4iOvfGkSso2x9+2GF4WWL6g6iHxH1dmfq92spiS4
G/BjKLtnjTL0FLVM7iZVQb5mxui20nh07uC+9IR2w/XIP7CMS9LSbd0hnWX9YQXD
1d2Ff6R9T2lV4rERMWVhzGR20GQtIsWufFolnXwfqnGv7sqKlhCFhkShg8MA2YnI
w5GvUsYTSv3ZIH6aA0zZVSaRE4G6oIusCbjn6PcWd//S4GohwWcxoyeIGeRbubAy
6ehFUhFV2D6CYP4lotgoqgO8fqKbonxMpgSr+92KYqAAp9Ci0k1ZKpY6kDbWRlSO
UjUbBY7gMrChaw6kMjGs8XERAun/9/+o/VnXfzWpjozeXr44jBKx/IRkqMF38igS
uEUbqa43zlzDDZdp0OIfcTQp2nWTdgA3nazSYhuZXTGiKEYMQ0D87ZnXQDT0WvDY
d1jmdFi7WceqUtmJK+BHKFzCShlVWuZELfB6uZbUPPiZYQAMX0k1DdUum3tuCElx
DBLv0NvcoJknEpNpKGonv0Zp/VHGUVeKwuNomx5uvDKk91z7QRjzcpxOznkOXLxu
koEiSGtPP5feCvv8mBIAV7MKLytlYscnnSXENjzaDxbb27aZdiL0FjPzGcba2mv0
s+7wyOEblPjmpGs3wpsflw7WCWLUIy7Rr1jZUGYy4m+DiMYkaDNTzlKrgM9/exHx
orMjzHISdo8BrEM5YSnTEc0CcEla5Yg1qR8Z89RAVFTdC4qKttIhPPtAu2U1IwD4
Fb+yTFlT841Wm0F1ZEU5Y9UO5lKS7MPEZ5RhF8Uir+c38EG0Q+BTqgvE4ZM/Wxh4
+LyjWuZxi5XxzeV09J81rorJo+CkGaL0bWnhpMpxcNDqC31LdqU09lUe9GxQ78ww
+gbx4tu/mcgqUBbdN0LIW8fEBBDQu/5etWUAfuS69hJYybP8k8c/OiNwo45ZL4fM
WCnkI0Pv3nNHpHfKCrq6NlNl0hlE7t4xlQ6aZ5x5CovAAkRVSh9S1hlsqiCzrx1/
XMMDOICL2oFL3idrS/xBkPl9fbTE6LUwsfRm9OT9CIawvxDfO+p0pvTXDSDQsCOD
L/2goe2wdlPl8Wj0cosOBki3rfEV7pNdv4Z1GTxKRlWkdfWuZFRbHD0T5SwIedrc
ieeuzaNg7ATC4Ru09ZLLWp45pbUK7bFJqa35LMf9SYvb0fpRxLApwWWNU0xnjCn0
pE1g5ZL43CL+sH36CPD/MuQjf0fgEGSaBzEyZ96FlTxJM2DKRpOgLIgK3Jg2oF3V
Apf0qNI1jcG75zidrCabiqa4xqimy2u5DID8nPOg3t+/fGetb6++BiHW5Y+pvhJ5
eQAkdn8ItuBlnVjJ23D0HpKPMhgCeCSYG/Cn67MMZTdi/isjC72M731BWEjbP6ie
3b2wQalaN+pVZTtZgvKIneh4w4vuP362G5IrAZT+lx5V4cHKSwPXJQOw5p00YcRf
r+oF6yePdQ/yIXyV0FbasH89ssw2rmo5RCbS9cKgidIkKJuP0MykM/5oWZcumkDk
FH+MOuuAVs54tcMTrdQ32hbJJMRBBEbjuS+XR3rkxl4o8CfGg6lrIsHu/mz9FkO1
XlG9M6cO4ERg40dqzyJlrkCc3B8i4b24xNMhWnvJwxKtsmI333kqY/iiqOX1Z7Dg
o2f81Ry01VSHXjTsk36eD1Pl8YwzJxMae2FXM5C6SiU05ukFsLnl5Sc7jGfkIsMA
RxRUCLhkQeHfMPijScEO35+z+kVOlwoP5anCfLp9keJZRYCUyOfONTqLuoA7n1Bf
rWgR1yhPQxpuI4rnEfYE57dFa70Qf0FOz0FEd37sNwptMR5DqRrtDqFDapXskyga
mCBFvoBKww4lFvFraZn/lfsgVcCJSqG0By5CfADFn195DTY0Ms6rI3N5CuakYzFr
aMz6ZimFJ9b6EemMucgJmd7XO3oLAAWQpMJd3SIYmmvA8aMZZH2TKnhOTNeW0/4R
CgiPPcyoSbm6nutHV7l3xdBfDoUTM/ZvYwBZUc+U5o5MbC1EZiraK+VNXSanodIG
Mp3kGznRqNk/nkdXvW3kgo1tYu+m+2UNA8mNFZNZCf+z+R+cFdzrvPEyq6SMXSQg
hlFgC1V311ZbCPCG5OfTRW8iB+IMEbPjJohSQGo2nEtfA71udmybIM4Op2k7w6z1
MLevykxh6p3liRlHdEDF02GFcsh+ocoD6FbDxUK67CZRZ+noErUA/RxqAnDZaf2s
o9e4+PMS0jbIIikfo2TW3ZoJlqElN/n29FN7pA+eAAWctM8WIV6Ciy1GFIGpU2Nw
wviuuPxYP/KzV1X/EzL1Qi2xgcjwr5/WmlR5sLUFXaWpTrNJnlqpcGC5K0QEqWBx
QnsP72imlhGE2XroR1nEzRIy+8rPkqS+FQGEOylh6GZebfJbUhM4vGk3+A6fWCJ9
6QTj5tewqtqhcuDKrN9D7XKegrF10zb8FKhK4OKd1dZoqNxY1T29pkPOiuFt8lZQ
sZjMknryXvHkCFduFywAKqNRGf/FHNaS471WkzjMFAM2+/7gJd0CVfjN6hQlIuqU
lM0QidWPYb5jlZuDKbrUs41nCEAMdUkW2qHBrh06IbH5BS90AgDRGeWpCBpKU8k/
uX0aoWNm5QWwz8wpQNSgObcS2gz4l4CCtt5hbL0Tp6EnFMmTgaLqdxsLpkb3D/Mr
8HZxQKct5JPqsInzmCECu+OOtvFPwOWP1dV+GbS6K2cUq7wF4iLm/sV/tgEXeqk3
PGgOekfayaNfjmwbV1ZP4hItLKSQzykJWegZc2Mr1yKlEWP3MREr0xKv5ytyNI16
p10gFvQ8WJivFYt58i+Onm/noT4IQ7Y9lZXSiacOrcLM/HSNSaag7RF1V3BZiTRk
mbzN0Mz4xUDhpZ+NmNvOLKWCMQx5WLOud6eK5XV1xGyylwJxZKQlCVQVxWUf9dwq
0tE7TGpxE8utnYZbddHktCKs45zbbSAFHHJL3MvcxSzez6nCzWPHsyTVgItf25hu
qUZxuv6KHMubFDXPxUB7Jts6NWK4QiBhkbtqjzfN+u1w8LcaoNV1ll1KA1o+2jFq
Pao0ZUYT8ns1F3bc50KSI3PgOtTiONkbSJVW6RLJ4+2fmgsbmtTsASb+7J1WJwFO
bkA7BvqqAdraYBKdyo3vQV4kt2P5lQaBq/J8Ie7y8IjAD7MiGzKBo4WLor5ANiNe
+b7hcXQfP5ocTHTvrGCTkhJjLYLjBqr1GD5dNm3LEsFvSmr2XwcCCoJMKitDX4fJ
jOSgclIFjP4dZ9vzUTph849Vnk8CvrPM+z1D4n8QpC8t4OgkcmppBXynui1bWjtP
8X3Ah1QKvW7BRhd7OxmlNuMvmv8/kI6BRpYE8O3ahvBjRFEpYWF2+rgZb/5dN972
UMJnGzT0D8GyAscKs/ouHFI5M1JjiYe9PCiG0Uz1j3nR1eA4TRTogt6wjG/DlWwr
I2KmTxw+mCKmxHynrwuM/VOXiDSa5i3PkZFuTeATFAUhuvqh5zHIDXGlL6QfW/ye
/Miwxmmt0E4ohHU+Ihe/2KUCz7q+h5R0cmYYm7wHU3sGbo0CYD3WOH6G0P/3eldi
mSJYNhqe4Groni4BEBWAkuyu7sorNYW2RCj7pQQIUmmE0s+Y+gTNXePDcmjC61OG
BKFIGzC8wvypqA1pPSWwtOghJIRvcgcXWNnkeHzFWow0M783dEFQbBdL/UztVXoA
FfSlgyVS2s1aAdo+F0lG1pxYJic6KClR2AlcQjNww4iiNAK6Debdh3dZllkim+Gj
tX2IVZWtH3e07Sxt46bzeYbnuukKgjVa3ZJnJPOr5xFr/ddChoNBH8jBKgwH9DFc
5Zf2zyzz3Fh1Ln6SAtgDEsjzKvcLOCUv/ZOBcnQ57bAb7j1SLMHPzyWOU8j/jvVf
zw6YQIwRzqxPZBn0swpWCQMQ/cPIsx4HHFZQALHtQD3RbKKcF65GGzYlNH/LmlLw
ol9Ywqw9ZrO14EFYCI9DTio0EGSUF0zv9NWB9al/rNCFJoL9dkFtou4O7ebzM4JM
v4kkzmSayJPrNTrRyMDjQhMoJn+5gX+G2kkoA+pq82Z/e8l53UUQw8UQ96gAtsDh
Lp4EZ8RYpaCO1qC+AKMhs+fde/VZAhRd06pn0aiaMdVXzG6hDBZorU6v2QteWwdN
JGKRn5k72UJM6Zqt9fT1f/O1i93nXAIWDAUxklGKehRufuwyIbPD3ZYITT1i3620
jf4eMALI9XWtTdLK+o/i4lpkjsVars0Z7XLv+oGPMWvsrTmyHjD4xXNJLaV8odKw
itQI7mXEgvN3qSMvSBqVJiCNwvQlqPXNkPy7GFP4oj4Cx9UKVH803u/Lf4whHkse
bBKnUC02QDNkXNLe8LM1Zl1uVEW8A+Du6g98/wOVxwpOXakd73Zmlf/9w7y9kFEm
bGa63Yp7QR8KnR8zRaV2x9BxKw98iynEGlFT9jvqqF8QATtbi4ojTWmLWenKrXmD
goMIXvUbwOveq5S9Ejs0Ybqz2tKaY1/ZwNn+2ezQfPyAdGKXiEjuzF0PYHuoCopp
QtZUq8eJyZ2pfkVVDKAhMjSLj/Twz9rh2HR4XbzvBl2i7jUd8OmXMyTqaL8Rgilx
MKyh4qo72LCt1Bg4MGE1TdzKG+q3McomvEkzkj89XEZLtRcC0Mi/qynbYCVVPHuS
/gr57o1QK5kQx5W5SADyupvPvXSgEIB2aWh8KYLJiauG6j82MnhbnDI2f7aZ1Y6s
N5aLSWZJZkJ9PG4wQ/Q7BWkGTDKY/dbKnKeORBCK4/T5hUKsRRlmtnHc0HOLpIlH
Fa1RhqiqGiupD/FQvL1beov7kz/Dpm9l+Pt/Xkk8048L6WfgMzsoCNaaURQ1xrW8
GUd/0GyJ87i45OVZsgexHobE+7Xtrvgqsd+Nr1KFf/+Xk0j/p7plRZIAfWWpsDK4
f1mqKonPxocwkaf3rX78ab5A2crKbQ9OnyTXrSuphbNgoeQ8XR23InOtd8ctlDj6
bDPhO/w3iMHFi8JF3DANcHrG9h7C9FbJ0Hpb8Kr9k7Ng29s+bZGcnzCMC42cOKAN
JkJJCPBQDvZ5gfOmfoUl//m20fCLpY8wMJKegPh25QfuVpc/N/OXjEAMRjIE8+As
7zs2EfyXFonWBc4bxn4ISqxl1qOsO+CeBS6S/D6/o7cQ1mTIElYxFgjsEKoT66Y+
dii2ECDEKJAq8jHiBzNbgQDQWqk4N7flFOUwtvWQPv3z68Ndmtp7Jdn6Jx2P8Adr
qbKnvD1jNAqaueZK1NFrY1W/LKriiq5tJjbK1jlfVxQGbu9n6C2u7IG8hIyWqjpi
QU2Om4ojhcJ26FEPG2UwygxCwQaLhbxPT57AWFVn8b5zL9LmnGrrEml87wIvUTBh
uOxxNOnac/lfFn6/x/9+HzoxE1f5fTLLE5ZGdjQhn4U8CeeIeMyXhXKt0lR01DnZ
K+G3pNFMf7rnh9D1DHdtsUysuUIVWH2s/uW1Ebraj1Rh1XdOzdvyg8aZ+lR3ouxH
tnTTevJNKMPZibpMpUNETqVw9btfMFPBWqcJXfI8ADp1ydvMcCfY5C08COCM+1jM
aYMJee68ZXBj99tFqwJSeqbBvsPB2ThUFYaAdrw2LJaGs2HeCWPl8WF3NnXpSURW
3C1ovtGQeDwUdAoOONu7KdNcez1Rs63wr7c6yFAI2SnFXE11mFQThkufGYLsDHvw
jnjalvM/hmlLpiCrktc/zNe/k+aGZkkcUGPmALqmy2kU+cgAJ5/XUvPFpzdcxXfa
x5B6mcqoxH2tQIc1yqM9g8PL1XL6de+0l8Qdtd+XBIuM3U9x53uo8Pzfy7vasdMT
ixLMF/oNkn43NQTT7YGVUukkd2P5ZwpTYQ5igRaQbazkm6W5MfePGVxpEBdKpWTr
qmdY6BpRC7VeHcAzTeGUp0lwVlOXvoJ5vjehLd3cCU5mTTYONEwcpOw+Y/2c122s
cYEuMZl11GykhAhCwiovoNdUD2XwqmufhwvTa4tJIDsjkc+mUOqul4YFRnG7019k
8ZPYR5FIEHBkxUsQ+gN9QHiQFVAfGnZX4tjOyuKVICmb0If6XxgasLDzNvQ17hHv
aMIbuuSZQTrTg1hfOKwTrH/Es9nW9I2ea8LHAovwaBM5RWq510dXzqqDW3of25Qi
VgJDUs5u7d++aGSzmB4otKafgl71zCmjnn6hoSDyT3KDFoE30wtjJ2YH74Gp5Kwk
PtUwkZwHnsjbNGXUqme8yvzC9h5Q8YwB2DLqMUC4dQIsXP8a/mMVZve+Fw+cSvkp
57ovQOWAdj3V9FvklG4i+TOrzsmHsUst21m3GCZgVzfrG8CrA+4EKs/9wOAJ0RCC
YrqgmD1akOTXkPvKz0Yv2iHTj6H61LmOMb7M9DkVvcQGtPpdqsVkhF2rOlbbMaMr
rpZ/Al/XnXpp//88F70c1RY7mCF4yNbvH8fzPwTLsVoMBUI6i5Cb4xkp07M7yy9P
12Dl5N3vg4lUTeWWb/nhQ8fFE6SVS5CNdDC2t+ewbgmT/aDxwNuQqNli/XgUpJg+
5XXG00a4S2nyCj8sE8yUhvL89IoEq1MlVgWJKYXkJbtvqXsD+L0KSdd/Ag1OrXqZ
Cx79RmX695y5IGZy+SmKYsvAcYXhnWRTxLYY1Rzu0Wwe1C8JM6LPAfvr1jDr3xvp
h++h0FpUnNBywaQDwUizSRLylAFUK16W43JB8svY4CKzuadfD+DLPFuinu8gPKb7
ym5r8YLd9i07swVFqF1W++LSHHmHSgTsj46fMhy+l4UmdfSyCeXSpXKJJ+Rqh62j
GrjIsH29AWgeHeNjNFHUrqngNRVCsOTps3K8FVHSKuTiB2CfL7hD+gZjRXn3HXfV
gT+ao/2qC7hxeJYPmkHnv4Iowd2y7wMJvyOfpXK41R7PPi2urMDQ+GMAuR32JYXZ
iAz5XMot6kxeDpx4IO8YI1o4NSOjNsSytZ83e6dTJ9AUSNUAkkwBZsEDmPz/dY6T
RJKJ5HwAH95bcAiWCtahArcjliaBbhCnkKhywWdRZsUuNy2taUeA3141A/0+niTr
7gxYbOZdKMRZnU1n3nU4joM3cI8eXg/Jz8rZS8DYF7qh8yhuGYRELwzCauVeXHI0
X4mTjd6nfYuHi/eAmLqHfs1lZWSMqMVKO4aWXRAt0/rgxM1K+GG8LRfjARWhXs6C
H1wpUOM4ln61KKhlkxib9QXut1HD+KSFXozE1TtsBb6rorj8Hqbqjh0ZWkbv38Hk
1KopQKc1Bwn+KatnlQF+UKpa1dmup+NUlIQzliwTSepMca0iwyH52+mLySBHBA0w
NPvBVRulfgXRyhL+TKIYIUUe+v2wYXu+/8VZSDK6i3RP0OpHkj2MrPRIUyOFU1NV
MpcwEOIUiANa0VDC3gTu5TJcUM1j1GfYML0e1hE90734AE5SklAS5E8Fc9hcEHf9
2NmdLKy4kJ779c5U4KUPmi5rCGTTOmHGlth2cJ+WTRoB/O5aNnSPKNJ+rX+xXsGN
DweoRiZfu+b+RrHl9oDx3I/rLeBMTvl3y6a8FoXoHgbzUvg701Usgr8EmB3lr5qj
zh2Ql5cuaCtKrXn59dBKkpGFNbdcFGDKMpsDzXqXn2Qrv+ox+jk0hckSgD71lxuy
ghMhrZiTP+VlBwoFClc1BxFVVV+jbc988AlSdTtsAR0oZ1ULLh9Axl43nh4+nwaL
lMd7kDN6ygt3hfBXQF2fWfAGYC3TyjqnCTRgtEGBrlygPr9Jv6DXcfaxxD+gqDLS
cppAlu6rSmEeySJPeT3nRwx3D+ZNT41abh/rjVcgT6B7/m7FKZiXxsDy6AIXNhvk
L0a4TMXRBswQRLHZr4Lk/L0i7WWiUxbCKugJodzlfiR6yz5P7OC2p2+qfE+8Uh2h
6rZRf08CZovZMQQeYfZPUTGKL9SF1f/5wEhDsoRk+Livu8bd9xIjqnoKTy3LiVmb
1cM0zhNGHqmHQnftu+hJjdGVmUSUrnX7b2+AbpOHPuxdbLFF2MksbkPzlLssmAbc
+ERFUoA6y+0n785WA3x4cNxi0HZu/+yNTP0YkaaZYpL7VysPe5H4BdY9jKPL0p2E
eq1Ooqvo4ntiHRJ8QZfzeG61yk8lhoWyP0dkCbjquOSeLGGilEim2OSiQqX8tmWN
zZ2FE38fiNclqfgP4X3ljERRg6dqRpC6mxY+eJxzZJBY408pLv/9Y9redl3M1qG9
aObeDCxQMpGOY3WOrNaWafLAT0R2aZwJhBoGRDV8Pv9irENxoYroZE5lUbohm3MS
zzttoSfNsdSCPEDol/X2glsGol0gIA9PcWrYWqd5vxZJWBCTmKfyghfyMwl6YatD
jkJAG1Q0+WMPv0i5codrdzeeK7/f9oM2Obttov9Y83EETgBoahXXt80P4ocYSaeN
MnMM8olV8C3Jh7GckEOJPuYzvKadd/AHzweDprifDydxs53foztVUWF5f15R49ka
rOqxTr+BpAQssAnBZgWexiDlUsWlomcGxYpkNJNJ0ikMLZwj3qYAMX4yoQf6AvpM
lmPs8i+plO7ejq6Czv7p2N00Edma2JV5oz/ssqmGYEUbiWV/OY6GVDH2BQrzPt8z
nNtxCR48fic/kvTXykRwo/bwxqYXqFx+NPK6TPYbV1munJjvQXDbvno5jNULuEMc
GYQKXQALZQgLn/8JgvIVDljpRPOw0LAYl/M5LanVa9uc8BH/BDR+I5k+dVmza0Co
IOdQ8Goe05vLIQ+6VoZtwdCLIljEUoEkE5DwdJglBuPD7sxOO4UAHhIYX4ABJ2r5
FkALLFSJevTfYqfW4DJEifv3DwE3D1ZhDHZFXarY6BJPWauRSSs8cSj60DzB4YLZ
kMyzGQ6YFl3b1wfIxnrgNxtLeTd1Ck/DrASa0R8game4ZgXCKsSnHC9mAN1P8t65
X97aLsQJsBA551IYCPCPuwD24iliIBxRzOxw5AOgzz9CeAXhAKvWhND6JuG5fl8R
u0mGjfHLaq/nuAS9/Zgesawy9xjN6ZK7rxGd3EA7qaGIpGqjKi4CvzjWZ/u0aK5v
9aIP5N1wtRLLbjnBhspeqApwak0BdwbCk3+7h7k6eJeL75Ubgyp6Zx/nczJnby5L
knvnzoVBOX1Obd6hztItpsax0IX081C9XcHxOU0FyPOnIJjvfj//cG/K3PL0/KuI
3fEWXTQN4UEkRYf7lIM6bcMPiKSwrbXRewkRw0jPRUvBvSJmVlOxrwdwDh0+LNu0
QBwe/X9dg35Dlm2WmIUXmRjb6bziQmUuUqbM7hFaOSYwIqNc2RGpkGaTIrn/6Ttn
AW5cdd/7gdVYxcb9xdF6j6013cn/kRzoIHRka4f+i/UrNnlw7HEf3XzfkIJQES/X
YLWDm0rj0PrQ4Jpq/kxpS79Ws0ZWODI3yWLi43q21FF86o/6XfA9DW9slvNhunzr
XopotvKkobNd/8eyAZpoWwp7qcpLPh04IzKTsSLosuDWvFgG8kjTtSoZ4wGSNsw9
YmwkHvtIFYeFmllDIYunQ9SGXDbIj3aa/2MUQRzsyJznDMonOQObjegVptyAy/m5
wTf03khhuMH66IJWDmfsSpkOZY4tRmhZU4zXxWXOx4j+86SZ4VxOqa2MbZThQCsx
vZppY74aSeEHmO/4vPWHVcDlwwHdFLr0jh8Y5H2V20UAupXk5q8Q2oh/7SuCXkcV
qMaZaAi9v2lq+tQOiiBevafVWcpm+OT7GDHvY7tA4UUJ9nSpXvBlt24IzzEhV6lg
CGxUb+hdbJu4Cd2kHD1Xr8cSNT9p4ZMFVO5DIpbtKeuAcXNYbosl3AGqsNjrIWqd
cNbXElCx/qGeCU63/GqYfLmXHu8eHB2T7FMI8JlVZ0Ma6gcAvkQmy/nT9L2LU97t
V3kVj8d9KpkQ5CcoVcahKla+VzKpuw70Ftp5j6oKYX3mOIgKtPKgvCklBUXDpHxr
OTNb7q6I1MwaLch8bTkEInIsEGuIWy4lxe/mNPov0l2b8W4nLU8xa2IHevDyEuHJ
vLQPqno/c5tgsECBxybJjimsolhtOAoPO6+vglzpgnhTjTszwGxXavQVMljXSNuw
AFkZKYhKN2WCPsFw8lUnoQCazz+vJmeY+vQOSjEt+TpD4qQZhoGBoAncMuP4mO/3
FsYL6BnX8NbqhEVrAsbEBpvNnQufsFxmMr8jgDAZTVnk8ffw9neg8qO2hQPGmhrO
JS+4qVzGcbOW6cCYP5WGTWxSu5R99pc/Kxm7BJayOCI1wHDxjT8N8HZ+mum3E7N2
rCvIL/0LLVPm8y4PdYHT2Vq3gSrrOhp+WJcM5A0u2SOUvEwXIa3UFOV9aaLCz6gT
5L7Qns2a7pDFt4mNLWRsOpw1P8x2u9Kemx2BE2K7JWim8qMez92BW3//jneMkYCY
KIx4ZtAP10atqiszy5tpRN36puA8J9tS6e5XEkzQN8vP/I+k7LKL6d7kP0UTto7l
BE5Ys+18an+e81Iasaac3/ftl4GA8wHLR6h7RHR/Y0nIFltKgVlQLS2MYTrMYGbM
WxtH9aY5Y3d1gvyLHHlPEr3qRvcW2i6oJbPqkfB1ABV09igwkx4o4Tur41OoUEw2
XaY6aJu/YQq1cvSHTx8hy3p8NjX7iXNRjxPXo2Qq8BFcnjgR4yCRZyR+OEYb8qQ5
pVw9KVs8HjQiWQtbl5a6qIG98hWSG2gkA/ztI+eiNhWEBY6jcXUQnf+EQvKxyN5p
Qjl+uK4kl/naM85g3vNUn26WU94Dr1Z39AX36AXw2gLh3N3YbF/Sx1490cN/71d2
uiWC3XWAvzagrIxZM47+KJnqmVEUEH2MPFs/RavspWCs3e/2AB+r6eKFWcjFoknj
25KKqsyLhlNU0nXUDDvP9yrkPaakLDWyE7o/IYByjx9+rp4YIGTbTRxQSVetAkkG
tW82qweYmo11Sy627xF9M/l51c5SSS95C6DOkOXKrX5SAUyu0Fcu5/gi9+hWKAkr
SOoK2OMx9wHo8wOVA+yDrsSybnyJLaGnM26pEobz8YHXdBTt5kI7D/NDp8KNH3+l
XHe7pEw876EKCiNk8sqGxavOIHhtNxpyNpZfioKyCdiHYaRLvE/XtMdOJTD/ehYp
LEqSyrwIfJdhqZcITfZ83Txs6hz3AYqNmyTK8C2APkjq3pL1m9wfTHVKhFdYfNtz
sxZJeaTtj0NW02CNuhba3x+3PUVttBIAlFqcUEknWIzmBbhdc48XhU1adksq/TxU
Ww1r81mjqpwwuM7UxKT1+D0HHNkW6KzmUNrCJpaAkdXMvPBGv0F23kf4Cfg2iJso
VLi8EP1ucYfAk0fwqBl9XvD9d0xQqX8NE+DC4QPDIGi7etBA+qsMPfyDY0s23sei
dl0LybujoRC46Dw6kRKh6Btv9sOGsQztHuehneu8pbcx7yZ4DnqMbUMI3EygTJSE
jZMKfAC+xS3KIIQYIC1bUcJxnXI+Q9kKgb82Q61KmKFFWB+vbpRwQpUKWIX3Y7vb
gMsHXqdUEEAZjk05UP4HBwYMG/7MUR7cIx4bKQdKGkmmP5PvVztFqli4XX63oywc
GWJXrewTBUTiNQLToC6oy04f27x2ztTB+q0R0M3vJalTXbJ3eRF0OxLtO0XDMZtV
OMU69KESPboPbllK5ZnEx6mzGpvhU/z3GZc+P3nCpTuUZslTJzG0azHv5qXPkkW+
UNxLmzOgpz8ss06yGDVjJdavTpWbKxE7AaX7dqtFOPqjqUhPEdF9LisKkHhsAMHV
/CSn2AMr9NOIAJUu0d3BGJHQ63Q157QV3SqBlvCIJDmk9RtwY8/te/CAYMaot8dq
6pIxYvaUqSSPtqthIwQP9QjU2W363Ij65eacER6uxpqy0Hoqdk2VShf6gNFVW2sL
HSOXZfdDLkfAkNBCEdQJXcuLEgo3GLr55JYR3kIlmSR4qUkfH+zCYFCR/wt2fT58
kOSPhLNZ5E09CX5t8+gdqIK8eLPwBzAdqPcx4ZpbCsmdXLjuMzX4mXcyRR5XxmMG
MoQ+dhe24kfm5IL1p5r26/hH1auqwEGTqJALpXeMukUYtbtkYpwcGgMsnOUHGeHf
BQHTRMeDDGFZhb5x4Bc/Zdz25+V53vDca4JDfgX/PtAamsfV2CdUzQWb4HS4DTgd
+XTjjjSOOolNl6mfTTPLxu6WZIoZjF5NeQZjVNEYDEkSuaYdZtPGtccq0Th/yf58
WGMxsh3dW1rtIJFfWmp1at0C3PiPT1PYi51nUxrABDJkUEWEiBgmiCa8FlGR1e/1
3VCqwSRjtFOGc0w1VKHgZPOQbiuaWxKsbWSXaf0zFc410asy5T6GRWGscyNA/UWV
68LFv03jAKzzNooIlX/gMraCJjTwezf/DhU/W7NecwdkDI9CTvidkvO2smK9qd89
Q6GIeODcb4OIS/rzy7ibOJLtWzpvRyfq4outFjF4EQYmDh4UTmM8ROgyX7Vbuooi
3yzongOIGIHeV7LlksgYnA0tjCwIZmalmq+AIuj7hTZt89SmhxYH0OWuE/HauyZC
S0TVsHRaXOEq1L+7L8SvOOG93vrYM6fiDbuy3afY19HhmatXmpdzS4BPRWn0Njzs
1spU/BPch2RAqTmcs2vS6PJW1QMOC/KA4FWE4PzS1kPTDsc9EO8YPcJujXvo+JoK
4d2RohHrCG3HCJytxYObALbKzcPwYoHisnvSRkB/lbrgnEXdLCTAFr5IpNwD3cly
FnMimB/Lb08Ny0jerQG95DkMsBVr82+Lpd0lKGRsdZ5fojla0w0cLxVPOBwK0Rdm
ue0+raoCi72d6fIsKkgWN8udp1hviQdWQ2QjKZLnasIJxcm6DaE8cW8IydQdOR3D
sYLJ6Ch2bZ20hO55xqXFNQdAXVt7u/dTkBtCt3HyIRzCHW9vSNSHwF0p+OJKY0qf
AM7RimR1YkoEHDKE0vjmyMuwpUTpRBq7v0j+/eoup7wU9jGpHFtRI7DbdNgk7xB7
w70FFC+8stz0xOdud5s5lVpf+qUg65IfOkuFwArQVIwGOQ9MWoGx8tQX+I3s3fbq
ZCyeYvjdumPD58iAI4siwU1otQKGMDWxBsH+Rutkbb99hmQDz4iEf9y6LZ/IsUHL
JPj90cuR7Xb5sfui/8dClzuMoqnAlL9fO8puaPap7i+rtaZLvQfk1UkHyoLPGCPm
mM4lbrfLOzdehTRCyF2btBIfsNOzBdaMy0ZD8zi72mkfH/uuKzejsJ5UPeIg4CSy
2QYnkitOH8KjaeYeREGcD7NlHOY3/Otje7RqfN+r9vmtwn3oP8lGQZ+TD0qbmmYu
tWqrWu18ZMt5o795VOcoXKwG3jsidth/y2mQ/dZi31Hc55t+Qte0eTYTmjwXoKRP
7qebmW24HMRW5SYfvNQm9z/oe0LipUAIca+kaXNGvg+NJTO4Z6Q/6z6QkY1ahbIA
UdCfi6QNUjTL+nrMwGy7aGOWHPnzdQqzIC8JRip1skrxPVgZBWClZfKzYpSUAeWp
/O0zydUXzAnRYub9uTMLGLldRC/Av8W1N+N3nrkLCWtLAGNQmUGq5dNKU6QwwHK/
FWLw7KbdJOVwXZ0+Uv1rd+M02Bc2AyAf3MEUG/6rQmmbjQf/c0l6r3l85EFCTkbV
7yC/S/ibpgAxWVX1DLtn1pAPVackBXb3lTTQZ+fJ0IkDWl2w6GDR5c50ISIQFHH7
lX5TRFpOrClReVMxPZghxUopqG8Wadjg2yjumDeTkWp+YummmuEWdekz1BDq2+XX
KrfF9f6xe23/8fqwDn46Q4FTz5U0MVGMq/XQJXvBF25zEEQfbg1yq02OghzwsDMT
21eZjFvqeTyIga7NtsYwkl4xVpH+FDPIc+H8oBnuD8samUezGZVpYvQhDX8sVo4l
DEt7zZ3I7MjfXr7TjrHCbp4Ul7FvQruAa4u5HwqkNjJuAFLZHl07WCvXSJ+FyaXL
hD5stR+mRYtkTpbSTtLI6pJ4bixUAxw1iWOtCMG5v0LuHoHlpOfGieGB3FecJtbw
XpnjaWMW0QfnFxRSdoqt9rcs2QgQi8Sz+hkx8TzGPW+We4J+In/lW3npDN4zP8Ku
Vbuf+gYRxDd96Rafx33t7pUVmjpZRAk+EtmhBi6yKbRQc7E2G8ECwb9t1U3xl+8G
VLWg/0RbIuMF9/JFdtBDpcCRZkQXAgwSDoeCK8oG1YAoMtf0iLuJ8uwOI1C/BEy1
5Ieexs9kVzzxOU97fpWSerEkl2TAYEOj8rYmg4+pyuzxgX/Cbwg8vjiDKcMbz3wj
KVRPznORXE0uFKemd4k3C7f3IM45dOqZY740LtINbNgEOi6OHMhnEkp9MNN4DKaF
R3vXAsAmf578zMy21QJmrh2NCHo2HWVVXaBkHUUI48KVAXhlWdRo/wf8q0fBSOL6
OJOd4hOk50nx0kYhVy2KC77gjUm9EGV/46hWpW1OburoZ0pXse5qgVFV9zgyg4sd
lcuEV6dw1nPKjZfc7ERESU7zLJ/fRuNGnAwG7DpOroZ0XHSua5INidji9g0vaI5U
gm+QLSkBlKcvP30zZPUNJ2jHq60S8AxJVmb4rF7Wh8/+KIzhgd1fN8tcIntoYHbs
rItt1b0xpLoS+LNDzDoJsU89+0SGEXdtWMJkMJw4IeAF+1J7v9AFVav7Fra7ZO6y
OvkgbRv8CPdWSIdbaPnaZxilHI8YSRGNKeQzFrQaqqmOb9e/EAUk8OU8X11p5L4K
A4UJLti4P+LwdRPtOngnqpQCo/huesRuP7y5MpoAcL9xgOeQgtGa0cGgeqSJXEo1
8eT8FyHR8RvsoG7oj8okAkFAJWiYIwz9mcqqXjxCi4cEbh9oAe89CgYNY9vHsMqj
f+a2uyV+E/HRYdSCOPG0/I6C4Xxwbyy8zWlAOwXYmJbkdUVMG+rwVibyMaUi119W
sE0xPT/BznhoK40Ax9cv5YtAgw3++FLVEv1xvFJXsflSa/6q151fAJ+JOQVCpKdZ
kd24RV+CADj7tl+8qjYQIwPSZMJ6yyJ38FPhfmpOs25EXg60n9x1PZjgzvJ42plR
51SaP7RLUWFVtUqkSl2dsaHiFfFUYkedttdaiPJQNymvGoNhCQNyRjZj2CHfXDJJ
T2O/ZOIZqx7igTUZbubpiZY4ud9r1zEnpY8fLJy5iwjFX8EINxU42MmiJQNXzcsL
7Z+YL2TqX4GS8elG2Vif2Sx4swH9sVdy7bgKQ1JNece2zbQIsapVOpZO6zPpK6KZ
FOOoglgeKAKyB6uRyLXQg2i2BpYJNg0oTZ1sOCsidW/l+uH/4nkfl8H8SL/UyyQT
qwvLms94M1i6u9fwOr/zAj65XPWCfRoeJUPapCstbW3pPuvcR3viRCIwHA30N/wg
d0Oy4j0eamgrrzOVbtRDODPsG7iO931/k16LEihmAkWc7CTQ3iS+FOSnfF9iT7zo
7MKcqV+ey6CWy6L5cjxU9NF3h6ngJ+xJS/jGrVTloJQ/j58is8/YDofAUefssnUp
F0uWSEmRVpQCfaiz5xUqdNf+pe72kU6uNbV/FEMseSn7kKoKIixm8i/UI3LL8HKE
fv7fG89xl5g3oCrT14Euj6TXYANMiibFPsrKdFLwNhxhXU5pppwRP5/3rE5qtILa
FS6lJ9hl+CYYRNIVjAQzQ7HIh0iz/YnZaDflDnlH1IO/gfuMWVvgpyZXkrSehIGY
Vu144U/SXIqiXuzy4cjr4vLQ447Iqt7nhaz7+09BGGnigMGBmYlCnzBKuYKWZ6mK
orZau9wX50q+xmucmkP8QyQWVH2u7g2rbv2rGShg6ivVaQZbQrxdGrv428seVmZR
uNtHkYqiz31TKRBboSb4UtWsJUcdkuOSWoq4pyNNeFQ8qApl4lBJoJGjrS2xzhQk
oJ8njqwNhkC3K35L3qShHDPalK/0wtpGmiwVokerELcaLfl7TISWZmqcBqmoAm1Q
SL7wx5+poAm2ACllLxBvmA+hiNk36ZwWlptonody4MF8YFTKa2Ja8/dodsIyOElA
eYZZlpPkqSaZs4LZ+pqxCHfke8UBFXHPPnTLgckaH7mHYVjfw8D0VUrLHd0OKVvB
/u3vfysxRKQi7N3Bnufdw5xrlfufUclxkpsHM9AW7KBtv+1EoIqLvNqvo9uw3g3Z
q8BN4MGMuQ8LhxXvUF9kaqxsh1z0fvkufTxkw+50M45+84TjVwLEbjP0DayNarDy
pVF4+03H3uHLXTwxbP3BI7M4jSTdjzLXJBLeHWl7uQtixFp5LwRqt1yiNQDZoObl
SgQfqnbcnChNN2/lW3An48gfca+EqmjqLr8DMbOvQo5+8IyAEs59fCINYODtS+rF
Rb0cU2iFLJRuronSyXjDI+58kdI90FZ5b85lM9OGhviHB4c646NRm8RdT7ernhlx
XXZtTk936tFkz0OypkCPSARt0HDDx+IhO3LEir5LLgy5w4tZpDnA+XhZEA0S5u0i
ONKvgnKcTOa6nm7M1tFt+qKNQt27DjegS6swuEbLKXDeq1uSFwOYvxxZqYP+ZKKR
gKoY3eb38QFpgRpTaEc/jEHVct2M6frT5as78RxNvwGiaJ+beTAyX5U88VMLsQeF
NSbky3qh2zGoOk7OGgtf6tzB/NHRsOFHDQy8HNz3Bor0FQso6ujf3wjMgAlOfRl3
B7FpJNZLEIxkQpsvP0Wb6uzFwPbVDj3dOurYa25B1DhTZzl8Vdb7JgLrQxbtw5vB
mDC2mw1aMvo6PvZj+vfEPHxy05kL1ejXEVR7Xaa1BrqTg86GbJHN8vWiC42360my
X7JcgHRTtr9W1JIPdl8W8D9yVdWcVIqzwU/m0sw/F5+GR2+4gWshW41NQ9XwALFs
mmIQMI8rjH8xJucNgIbY4LLRtzNGKDQ8jXUXKUY40PqK5nxQPRtpZ+Y+QH1tPnQN
dTQdbSFN+UehAdIlyI2p6kdmKmfU/ztzqWow52DiFFz9ooX/vpDnZ7HVy7NZ0WOS
trh286WMfGzBOjP/VJJKSnU/YovQkAloM57AfvO6QFwlYGJa/BZkt8te0vD8F/n+
TFon9MPVfk7ahMg7dpOoDRcD5lVXf8dhwN8cIHu35A2a1s5TtWfTkLJfr9JpHZYu
mvpUr5t1iBTtJ5U7R3l1U8p6tBt+hmsjPrMm8+6Hi+f/E3dflSGGeCZl0aDPgSUo
qXOEA6gN5SDxAXWMDfyRmEwww6WPMiNYdIv9Pr7qgGnHv908kMJmV+o5nI3LjJ1v
HMQmjL4IZ1cpEZMl1zg6AGU41kIYhcZpbxyGFbTnRBm1goFk2gK8wCDx0oXLMGHc
2oPijEfwpKcebWBqK+baXAYwN/lgWT5SLt9LYly5/UfTD2zV+Gg2c1ky9fxKYw2K
/6/y7uqMs/O62ooeORFoWLPvUPx7HQIOACoFrTY32QuOg7z1j3ZwnJkyX6yRIxIK
nfogQThZrXBKx0l+/Dv0+cLr9+JqA1KMZxmkRU8Rqyo/bRPkrjeg4yNsGV8Fp5w4
JjaUPC6kKNxjlO5DjCBbJtnE3khvNYkhiQjwgAUP/BsFXBMJrEC9eDsNgPLLha7b
VRLkQ4w7xwyh5g3hf4V6itRX0ebVp/eguAjG+UakbKDV8gD8mc+e7XgnWjOyYuCz
+3F/7dyZTV2X/J8UyeMTthvULriM32K21/J5zAu4QWju5tV8T++SMN1DD8JB3dj9
ZRSMQh4nDNhuy8/8nkslkNIyjoryzjtTjWiQ5q4hyPjAta84dOPDhpZ6lZT25UlU
f9Tv4zAsCb85UC+s2l2OoYpfHAIaFDsBj5+Izc+YyXwVesA83/HUNTiPlhGr94oI
GvFEikbJ6hOKVtcgl6/vovMzCNYLdi9+vEC6D9ipR2+MQFyX4fBmI1rxujscSHcw
ElJO+YEKohDpLkPhDDKU/aIHOG6uSAxXsKSCPeRObvmKg69MnqQo6BgVUoKYvpzH
A1RiqoQ0L+FZh2E6XnWNmFvu7LnbQSW7zX2jYmai27QDLQiuC/N1cO8HrOQkSYj9
V9VjoFzwKa6Nf+s1x4NQhAZwXYqbipJ6/7EG3dj/jIwE04sVP/K1Tnp/2CJ0hKCF
AgPMnZz/s5i/eJWhLFD3BlQmSpF8kUS524b6CkWk+bJ+RuPNF1jzLfpY/mb6GoTU
9ngsi+5kbhdBuxSNi43oj+O0BMjXuVwneXK3Od1MVGM4gcJyKopoBsZobxfH6SQO
yk6KFV0OOtFUeBT/9DkT8/npH3Me8um8CWP9IjSpA+rZ1HcrSoag7MdYUDOnrPbD
XYIk3UD4MK8lMjFAMThizaCyZxtM5ZEpfFOrNXBhWyDSxYJWWA7HOQQbI8xQQPyX
ChoZhJMTxQP9InCnvHw+llbBuVuk+CPKF5Va5h2iYHkKsOWXfJgZaPX8wh9NL00u
XaAwq24j0vOiOz7QFGtc4a3LadVa4kXRK+BmjAoYM32TeqGuMUsypXLHJLZtW/wD
F8/g0P0drOVMmuYnAxhIKgl08TqpHrgGlTh7FxNom+Hadz0QbYQVwdLJEh89tBby
4GZlb+9jEYsAfSFWmoQ+QQyUHxaV0pQwadYIWKJ08vUYTdxq3jNqclZdOVO/l5QK
cr18Gx3prlKHQ+3ibPRmrc5bu1XWd+4IjeWX7/1hQHugd/K8yWN3XC7WAfZBJvZg
tFP4rPloKfMY+yiLPOp/TvrgGnKlKKOGSWDfAERuYZV/ONoYCDXGATrGNKZYsN9A
ciY5kGn6JLjohFVPcqWjW2fTOHRCIqBqE8nAfpqyCui3lEZtgYK5LrHLbMdrgQqq
JgSKo+JKeCcBZSl1xe7y41nQB+oaqfG8LGnRTt9N/1cs/B0jkGTQd07TVma9njK9
7G6InoQwDXZi3ixM2kzABNEqTv+e2r4QpJ1bnOhM/Fv0sLDBSyRp9zyXcq+9Tfky
8MUbVXDKh3hZ/trd6loQvQtB2/YmR4WgVWjgcz8BwOastJI7MherEb3VHM5k/yLk
O+MwHZLEd0Xl4I2m7aQTOu1POvoMu8NnixNWlv6AUtJs+Q5DCXJK0CNYTHYTufT5
0SUrwgOIbWa8kyJ0EHJMOfl06jEU/F3lS73CVwXhUabNBoSVmmxjRyScremgNq7Z
CtqwlUVhx/wSudyroqr/cyZHaHIObnD8VKHWya8RHQsPv+ruehwUuMPhic/+9K2B
Tpc7ILMmqlhBjolKL9JXt9fvEiX2kIXqx5ucXQa+7xxY49TukvAWCLX6AdUGB0HA
deOK0QT6pg88oBhcopmxwmgszclQVspvvkhUcbptTGLqEosa/n03U/eteTsS58u6
ku2ToahmHQwxCdYFUHAkz72JFxOreG2f/scSi7I/g2Rk8ThiKFT0ndFNHyet+l+C
xDcRpvEu1Pp/aQD+zVGIvkHiqWongQCVhsbkUYAdfe3U7nSqLACKLw20c/TvwEdm
zHolhc8s2ZJW5OubedaI4ADTJYXP7HIhe9/KqWxeBZhbb6l8EvYZOVcg5HMrR8zD
nT0nzhtwFXk4iLDZIrRmMcYDBgOkYa49rwbaFN/EgkMKvTGioOwtXihf5jzjaXnV
0tDtQg6XBmSf57BEnVHXOKb0/6dkHe3jTdDhgpNt0Ehr23ocvem2C+hj+G7Nrtbj
pc732ujQLoOpUHOXYf1BU/98TrnKOvPPXiQWPiW7vH4l9L3TTtoTRQQ9VVXZwzkw
skPyMpcmVPHJRxZTt7271ArTaXpphyeFaZXhnFSUQeZJVvJgz6xZZSLvu6vgdH4b
kwWXLSDyn/NaKgHYGIfOPal2nkwpeu+qg+sln1cX+IynujP044tlMgDUCVT/rWlr
RR/EU1yIm8S7vtzcQT0t6B+nf4+ykOU5K0YQO2WuP8Oo66NvW6kUlUB9ucyeg6TY
qKuOOqiAXY121sLY08G9qy9Aj+UF7lHWcDP2kEwv2p8Y/be6YTVjQbHVvK6WTuIv
c4hVnqeFiAgnZbm26pQ4wV3MBhMbhQiz7wHuxABTvm6t2riEpePoPTSBbvG8LVKL
ZadPkGO64oWj1+8N2gYXXEbGG8WPa3HdvDQppmgBpSQjyA/Pjzfvxn5S794ZosDM
mZ8W0Zm2J/vQpBvxjUAMXcsC3uiSJ0t+HyiPusVJRnkXYA9JpAuzQM8ZN/E/6Xfi
4bD1tk+ImFFqYRTFcmKgSZZvv1WdVt0p8Q/JHyMEcF7Y2IY8xXfSC8GmoXn1f0nR
Ti7UePPPCBzCxuasBuCJPHN1L/6NySor2Pmc0BVzZn3SY2ll6qEZM0VM3NTAVIC/
PvcV67yxU8S+25IJS0yoGqQ6SyCQ0otqaanccVh3ZB9sQ2ZJWwU8w+GrGN2wWGUu
ab2hRGxTt3xz/h1ve2vSdcBgXaOlK/dj1IoYO65ngRnWofr6CMvJNWuADKjQ6Alg
HinBNkQ9CKJE4TSN7iMTh+NPhFnT0GoTXl+QzyUl9BFZkNiFT23dsUtJWqnMuGOa
56BXd/LIlajW1mqWt5ZDRTs54smpQ7rk3fPTcKo3jyG90XGIki5eNw0o82etIBqt
Vw9+By+hefFhMCt9mv1wX78+m+USTqhpBpwUxO+Cd9YYFzHxJcuIUkhFtcEUADLB
1Wr4B7m9wVd2oOo7dMcwwDvQYfDnSPrxQgaE5z+xibyFmJX5yJYP8U02QM1t0+KK
KByDObFNr/DXKmBK/J2/HazRJ8xRmjlK/zwNVXT7gNO8dFP3HGRQKnIyQXI3C4Qc
Wt4G6YDYm7O0sFg/rGsDLXgvAC8H5wGeVdI7rzXSvb7qPEFeuVPDeEBaZu+zAacc
frx+MaJQ/QkmiHlRh7UKqVIcs1x3CJaDcDcr89QwztP5e8ZHEwkRzzXN+q0cy74k
e+9WmCRtEj6oz/nkUSnkxID8ZBN/A0L0TYIbiRKJ2LCMSIDYmRW0jnHNLPvTtndy
kTipgOtI1xZA0IggBxS7KN8gogwCDw9t9+L+1A/tQUK8yV8jDdjzdhbNKcrZz02V
mi7q6eZoHQczQgL5kFN0rOLzEkYKEGkjUs6xlrmFCa3WSu/l8328A5H4OXMwHzYv
cO3iW4jdoxs7CNqwcbHH4bLNEOH1Vp9wqNFfdyn+cOh/nUSCCL2o8rc/7gEbsB87
ybzqEJ4KDQ/9OePrGauhmDcaPSnP0nRDa/9kaPd3wjXqRKDYBojqxxlPElo9oMnI
qV0Y9pTAdIoDtGpzp9dzom4xSo3GuhQedGuEXiW5l8mdt097HaFA1URSG3AHaDx0
FLUoHI3EYSD4nmxg2wbS5ObVzELleBxbOkQjcC9TT/lI2+yzUBIKk3VHoxtfH4k+
PTfS9s7Wbfwy2nGRLqie4IyuvX0HxOl1/UUzk3Ej3/fyhHLCOMZ7/dixcwb1JlOK
P8+T6sQ6RgZ5jqSEZJuckE4IP1T9QBdB6P1Znu8AVKBhcpZlQdlleaNwaKljU/fk
pC/a+dVg+gstfVay+imo3mc1to+LEMFmSr4EiQnTkLzwuNugGDcdTyJ2BWxsn7r1
6sbkum1tTnKBIlL+uuZz29hATvitEBHAwTpiPWwOdjXQPHtZgWZ/kd3SR57HMD7U
obbAwW64x31tSCc4qUt+VFsUcx1As4s/jnJKvuysTPypX+LyTxxTya7IY7Z/oRwh
/mXtxvyMe4KYkmjDvkYLbf5flKe3WYQX/wC2TX5Howj+RYam0XaIO//FEfAZfNln
ZCadQH+g4Il8kRLR3JoWulV3ARoiGex5n5BuJP1j0MK3PTc/A3rPjokHZ/Y2/Skn
i1odOlKRw15HFPU9x0VTUqYqpJRy8akMeC+rIJqrLaVX8B3bHXlhmYJRv6FSZr+d
n1vxiS+mkr5nfYuIAj8ECjS6NWWD5PezB1KLPC8TSxFxy+IC+BZfheMVArKTfTZt
Zbp0FTv2NCVs+g4cwM1dx5EEi31DR5vPJHoXt1eXF4O689m5jjgfZmrf2Zu7FfBU
SjBHopprQaIptVu9d37Mo5ZTybbEGml6OdcSv+c0CB/sk0ea1YojDEQurKwe8+M1
4PliJV5U1grgg7FEm8kRKfYHRDj7I5CtiRB8mOIdi4JQ5r3kuHJmzhtRlyas7UNP
ReyO6NDvR3l9SoIEyFQQeUfRHWpwaKv5p9t8J5fzmw8DXmaM0/ZfOPg0hJByJcp8
sHeXBo7COUsEcsAe/fR0k1dKUvLegA0AC4tfmkhEzAGPC9RPnonGM0trlD84EsND
thPGIfbxmOx27wESAru7MAF7lwmCg34x3mJFZPvDGOkcapOKuKu6oARTPd8LoWOP
SAoKRIJYnA+IQh4PziIBfqoSaPAau4yc/t+bKFFo4xNwj61iavUylD0p17TKUWaz
tb26ppxY3wnbbOh51kkeVm6jQm5G1BhwwyHQvLG733DwKD/U2tYsRkNyU7IAFBcS
25hRcgxSq6VvrqvG30VFTdKNKks8RYCtCsHyqKu+2Yc+oAEs1vLeUfBfVfkAgiGV
1OfpAdL944EVjQFmBwXJvV0uLm9iO3kyxHwvFGOb3akYGcts2duqrNtlAB+5N2dQ
xBi+FTC/3yNYXtPXbLoo5eJMMOuX52s1wKjkVY8ys0qzYw8g41vK+W1FdMLzimdh
oHNiMLei44v+gg0OWrkHUO05Du11Tz811/lhpBt5JmrZJU5no46zqUElvPYZkUcS
jdUh1GQhP/7rfXt6NxK46WjRQoUA5B7HKtMqGuql4bzJ/InoQtxcFIwjlplUXk7R
nR51yVwy3zJbB6VNSn69F2jn0BLh31zomX8wXt/f628j+WN/V0lDxh60lohxLalF
Jd2bLYX7L/4MdWbs5TjNrKXkE90ELW3L87xbCxrU9S79mSlZbZv57CJAEqELOfxL
EksSc5dBqYPKE/kXZPQYrupnSGjrpm683zh8vbR/s/IWcOM5dNdliRcEyQK5pT+U
EtOtXaDtGtCi3V3BPp5IQEI/KeG23WrulGc8QLncJkuvIIpVsDkHC1bQasBlGlSv
KtMZbpcH0TI9WZh7K4VcIwpLAKiEft/I4XHFzbsM1iU7A8cO+OUB8K9e+lIPGgeg
J7uMWddkIkH/EIhxYMQGfAHPeHFdD6bmEcLApHxx+l1ufDJF5+CdQr5kYX2iFrhW
PWkAH1o4yVo+X+CpOz//xYQ0tkfu/ByQktNK0jWICZX/UUutm51IXUzsGgctvzXq
sAUTzukVfY7ei0wP0Qx052tniUAhXhhMkb864tMlsqYGl63Dyh7EVV+IgTfofPZU
ZeqTbl/1hBQd6k5+0aLKR+9LvnTj0RA2ZFLqHEFNWX9S4D6xbjLWevsOlQgjg1WQ
QuMqgKPffwnrgl/73fygCPSsCTCND3qARs2/2WXGSdY5M8IIbrOXkQRnku6ZYpA0
HTjzJubPWeOF2FRlFZZSqxhIbmPdiHQN53MOLyKqH7IckH8Y/LcUoNFJrRDsU65l
/KT6NIFNgWoo+ww5tpS6ekRa3d7fgNbuR6cpKY0fLHQG/OrBm9FBlO7rQWOf3yEg
XRsZobDt4LA3wOAmAZSBLx5aOB0dNq0kWCGFNuyHsDZliSHO6Mh03oW7TwAb1mbE
1WWNRSGOIxlH0nzsuCZuHYx/t3tzkxVMXh9uL2/IzB2+rd/o3TYBV0xRxrnkBU7M
eVfvtd2D2a+twfgLlLXkYD/oamOlKojofNU3OImB7VKfunDpqJnjkokQLICTe4rg
KWk5Fm2DRg0isMJQ+biN53MLdd8EuSCRXQtw3bVT/CU9v6O5i1o8ag1Gp33jUsBy
tgGbq/yZgMDS3RWrzNYCXLA2gYGZfDeRd+IKOHHU6RIr6+K1KkBps/G+18M5vgCl
XNgrHNIUB0Cn1DQadg6sW5RgBF6YE0PTNG5D6oYvbyzO0hw/QyDWxXI8dntW3qMp
f1R9F2pN4XdKOZa0EZlwf86r8j+gOs7EG3K9f8RkgUPsIqDOht0HSb8iu6umElKp
uN1Fc3Wi/HWPRPPJVaouDGtt3f5LyhFjfSX91LMK9mKhgkGF9k7kQRAz7ED0ObC2
fUz0lx0qTunOmSWrO05qQVAZegleQVUra2DWsOreqV2Ft2r0R4nO8Qimfm22pvDS
WJO7iTZIR7z1JrwGXuaWF3g/7CcH9Ti/jbjht661XLPTIaeAob2kb7xT97uAerfJ
3SKEtCjh1u6S9WLL2CaSN+Jkh40ijj6+gpBtHufaGd5ZHOOX14WroOrOOmIdYiWS
S8tPAYp1R8NDO75F4LphVReB4CQTP6yMiz8GhixDX3bEqDQAUMQPF375l+iJMi6G
Pb3YYcMfPBiADsBH/AYANmTPxrV8Fm8kcEXE6Wv61flIdV7+HKkn6qKL7a71pjcO
SoCR1iotOQHhb1xuudNtP72/GW1WhmX0POxq7A4FWJGnQW4UCMoM+G+YOolwwt1r
H7BAu6N8+6akNgwcwKWuUOU+PSbpGANYLoBWEtJjA20GYkxHVBs/3ien0Q8TwijL
YDnz9CyJExC1+UOsWugY/fm/DDs7PdwF56h7NlCLiJxDEvW/qvrVsGjJiBSDm5Hq
79ssjyJTkm76gx5Na2UzBbcVrAuApkNh/cD0HOToxbvelU6Q5ufhUm9van7Mf7bZ
pZHIkwgrmz111kAfn4WQ0LEIG/1rSDta3Zgqq9QKOGWrROIO1TA6ip2MEyvduUF2
b6YHZ2kJMYAGZawR/G4Heqd8/lraDDIDsNlyKLhwg++SwbgGRt5Za0v/VpKQrV3r
hu32rtR0BXRt/VMUf885V0I8lvWjUivh6bf6W8YhzSItGPV/orCA/p22xVUyqzUq
PJ5hx/MTPmnVoh2BbB2qiCMlZEluMX0fvV/TyJh7g4k/x6gziz/8oHegJixqouUi
ktDe2LvDjfRryU2gcXnLJ8AqR2LZ2FZUJwPqtvVMypMkVFYrIhq7PHssU7X/t250
CVLFPZAB1v4T4FILjZcqAqv/qYUOUD3eVkVS5To1JUSFEvB7xFbXdFIKoF57IhCS
2A1ijNp2TvLwbyq7vz+catBe9atbeSjX73aTcALy+tkJ1r9tsOBCgPTTVGkUPrOv
guqd3xcYom09qvbn1wLXDLEjhGDMxweH7L7rTFD5r/2agPHbnGGzEDWFSEeWz2gq
4V8pu8effgbgRjxnh9nE0pCSfMBPCmF26nvfSDqKaYt4QmG5i3YllfK/BAzX18tg
CkJAaMg2obQcxHMz6rFQU6W15PBw/iyuJ/RNrF+95UteAZsMBClNpYhLXeFw4cOT
SOXsvyHRDoRsHKPilrHXgoRsh/oNPOiYsR/8iHysUoL5pr3DOvrOVE6TFA5+xLNm
b1fK/aZX/VIh7JpQcp7yuYXwDIpxhkIUz7lsuwDnZe9rM3rlJftzno4Gefg25T64
DnnpATnJKtWaoW/KZUPb0Y8Cv/7oLDbYfrD4naDqdnO4sVwE0+Uoke8j+qgkVPK5
d3I6D+7I7nm/mbyZyJD0fMAuF5etqVrbqCyEFlfBi+MnIWoi1dcXOVOzRJKrQn2y
NVgOCLmNuC+Ow1C17R0nGLlbCibmTzR9i+V4XfB5U3pdfmw1bt3kjYsR3bbM/8JO
lqDdl6HYVTLpfLDGdD54v1m94Mmob6qw0j8HQHmAA7QPGGyGjK1NcuBjqKJDaDMG
gda47b7ReTjlN08Yd8TcrEdo79c84tggWFcSMM8eNZyHLbaYc53B3Jtw+78HcIOg
3w4qgLQ79PooxAqjeMVUrTudLVv87CzRpttAVQz4kSA54vJAjnl98LNWSdkieufz
YBGbVau6/nTrvl+ZNduwwGyGmJdymxR97vmlh8Y2XiQEuhMf3HuUC8iwz50gHdEM
wVZ62yRnlily77epfhW5/ycPNTPu37LXO9vq2t1+ODhz+AygbPtbgdTB5OYtwib5
yZg1CYcw8ljcAS2Zv1S+k6RQxXcB1MtGMgrn7UQO5VHCjSlfDQQLzlOXSAow2mDu
euOXPtVU5TVAEWGP7QaB/OQ80P1MQ0WGQ2+rYVURX/pGxOKCg76yfh+nl3+ujhYZ
A0V2Y+W3VNOhF1S7ohFch8MaaJD94xF3nQsF3/Sgpyk6VFSg4+K37Pizf2uLEJC8
+AmH8vmW/BLRTJL7moA/+3AP+0ILrSGC/i7jcl+8vpA+ER9ksFz1Y+4CcwDU88qo
mWJs9HHo9or+PuTprB9FwrhAZ11u7i3OtMZiDAHWBv++pDMns7ybLETadhTrM+1g
5qg/PXdgi6AmfD2whIwq4NHycXl8y9+NoThZ4TkNujR3IK7fUun3Jh2TjZ/qhsq8
V0tWaxHoqj7c4a2/VH0wqcEabFkB6AiAZrMi1/jrYdOBgDAQCt8C6vXQx8dfoY6F
BuMwWfyZ7cEgV7wbSLgqDmIqpYoAYEnpxVGYPP36urphcroq+Fq3f0x/vfMxdfY6
LGr0I8+ptdpyEl3d/vq5A+dSdvLzT3dSZRpcjBCo5KRPVpXZWvPWJpr/ymZC/5Q4
xX/uyEcR8dHtE56wNSbVp9w6oVhEtP14NrC5QNjHj3RYaThihBuRkAsxXKgPHNJ9
A2nBZunS/cIoTSfVitClOxvAPiRZwsseWrkv2zzPBTXlsscreC2jcyk9kepJct4J
0gWWw5zz8iFlvVfWgr8f5C87OyaeO8K6J+4Kw24WkMSb7QawOZXDE1txYtkGNCEz
e2tSmtOGddCZY+c39cD15myUX8aI1N4ipwUw/gsQafm7saryNg2OxvJ29QIjEiqV
246ZnTGbccz6LmpO4wqk5IG66Fmz5+3GIA3BLuq0uKu/orMkMdmDCxtsDaEzwzyN
okKfod0DgVQA13MxuZJc7urAI9kKt0x5f3fQKCydAbZ0eEtNSxWtIdpiQ/wR9B9H
uWfkCJF5PLHg3e14ZVWlkfG1E52iU32mGTLzVABzI/AfJThV6JmfKl1cGKjEyp6x
qF9e7yHveH8XmkD6f0iiWk0Of8m6r2Hkr/r7s2oeO09zJwZFB2LhwQXBNJU5cbL1
UJ/CbU8hSXO+Vujbyn5kO4eAQa1KRllC82UMruAFH3zU3IghiodTE9TJa+QNPQoa
duGqNyd34CWQCgYWzOzcJZ7W2Qmfn1F9jGb/nIOCORoD3Zg/MDbHQFtIwmNeFPI/
JNxnnR3vVwmjh950iQpQb101MedLbELObyc3h9NCuVnXJ+eeDhfFiJPXgvz8uuw4
WHXxxPc5MUxXBpOSGcLt57Y/rEqIdydLjt6s9hBPctrhZpTuKV8fgBOZonC9swFa
O4rb+qi5GgzpB8xHZwZt0gqNu56wVoNfdjiQkCeHBfGZMrWWTrXYRu0GTB7Ix2yW
08NfcFYENGd7/N58JDJ/vHze0X14YwoMN+WVyNScV8kSzWUX9oYxqLziON8kX8QV
n06w76VKbfcQM84gAX+I4oAaGyhb7tthAabEn01sygcopNWwGh6F/KA3mWQovwYR
4Aut4RhpvA6YMeDg0Tyy9nNXTAMp+8/yXQpN7xdrBoZ4ZOqhd0S0blhBG9fYrdxN
dqBIxyt4yvq+NnHmbnGcOf6c+HH/KnpXRWVlovNrWFsuKX5N9+ObQQ8zKekjvYF1
QE2htFvSZmaPnNoEJYlOmnQ3KfYKb2GpF4V0luEFtnJMIuwfeMK02eyM83b0wA/g
yuTWrwtxDqDpmLCSGk0Wjt2XZiwDI2CvHGV9VlWmINX4jdCWeoVDJ013hsNJuTt5
kqtD1rOMCdl04utrWW0dV5jtwxiNTY5dFQPDyyfYs0PKgEObF/VqlUGG5xku3y7O
yuA/cqu9KfDmSLB3sOSCKKdoL/45VfEm601a1LQ/iuE7ghteUpqV34iaO03nEOHe
PeJRZfzod/QICiyJ0tcsGg+3fdqZpqKVsx631N1BW0ekbXYzaqNObix5StWD6P5P
U7AnZAR+RsDFfnYEYPEdhFEJeBwZ241bstUj3sKSTxzN1XTfPJpjSKB3FpOu0/1l
u+OMgkwBG6jA45UDgK64JG0AZBqKt43L1wAuT0uUc1n6+3J4mGfhZVFwVqvv10d6
SG6nY6ASs/+s1heYDsuWBY3hCfox6Zl9JRpPSuh2Qhegz0LUGQQ7Yry5yJioyoGB
WpC1KZR0wUzSgQ9af5fV7gvc7Ok7jkyH0lvQgKfI8qgJU1EmSoGcoH7kehzAnvKT
Ox8DNfZE4ibbW+ErQQdc4SBpDJR8z8rtNoai2ZO+vu031932z4nzWjHKkSFSnuHW
QdZi5rI6atKtTmNPtwRV8jfTrbo05RUpfQRsA955kDMfE12GbtBWprinjJEraotg
8cexjRfpsa6sV9me2ChbLrkNksb741PXwHcNeAw+Qx+te/V4/IS0xVkGZrOwOi+6
fhybF9QNLsUacPmPXXnYYREBQ8vN14E59r21erCYCsmMLuDNojFOhEQ29LIcMdzF
K0iWSFUo6kqVbk0Wzooccp18Kj5Xqq8saFF8rmDHsd/2yBWWZ6mP+Y5MACGUPn3X
2Qq8+25MGfsGJc9vxravMKw4NC4WxIpIXFhs3ZVi3t+Fm5gTQPSu6bVeCbklX6ds
vpxL2+tcRmSntuwhmks2cLBfKAWegwsXO/ZR1LnfbKijlVCFTN17J6w8kwKEFuuS
fhE8cjJzobxvfN+L7GCbs70sVR33oWNys1XsqU53DKNXdO5vMknqw22nCDDzSDDT
YMCmaqHhRLjJX9029YHDmGJOU6lXLbt1J1evgY9E0TIYVEHZFyDpMSX3wO0u9UF8
OdbMo19f2dSHZcsSH82fDgwGiBfnLF9eJoiFDoNlxI+aOv50m6mHQGtQeefDjNrH
hm23WHdrPte+mvVpl65zGYdoHT26zboEV1TAfxs1yRVc2iGzgosWTbjtVdicqwQs
0nYAIErqdtbLpm0x7s9ZQHLl6Mk/9SxI4UnMljgTWIZ9BGGia6mjjgQ5C50Ly5+A
QwzhLi69tcHUVv4Jvo/XuRKFpAoB2BKRyR/8v000kIaqNaT1ljxFhW2OH3RVRMh1
fMV5FUtmX6fu6GyQLbTNXPgcSxgFisx6XdzuujigNh6/CSiNIw/rUMm8zEGf3o4T
wjBpcgSuDc+ZqE0TGFqMKg6xBgEktl9JVwzAFYDpUKTe3/MQxUsifeTPVCyRN76u
uSc9QK2gt0Qt9CuxhF7QGDa6X1BqD/Kds7eHT/a005qUHMm1838yzhtsB3bk1+03
sstWcCZxqGv/SYRKMv6AHfX8EDnZRK/NEVFfxXD8orlSk6fYNFCRpG1BHtkAgbKc
YmbIR3JiEeVNrTwCVnjPcnk3PY5SWtOdqSx0991LnZZAYev2RwFobdSfEorV0O6S
3Wox5Y3D8UhfXUK39n2o2ato9FBCIDDFUUdv7rPWVzXmZ2MrYQ6/mP4JGnGLjQg8
/AE5qLt61dE1DQ7eb75wBsjcKrXCASXJ6cjrS02AQ69/yAojSL+Q9RCXMznBfF75
DZIRi3XhjdjWePIgwdtsuCqp3fRaKKKmZK61GYuiLqGUvQ2YURb8GbcwzPsN6B/i
UrUVuRP5rsq14HA+lgQvsqCBoMkD3EYIcVyEPZ0UH3DSGcvhKFxflQxTpVSrbsnp
36uujXy/QMsUuiOMhbaAt91HTmO5bQQpZkLPnPGuhk0BtQiqsKTdVYaKBZudyKv9
Ue+cFlAKHoO5VNWV9bBrL/XZNYFHf13dys37l/xJWDtxvCQ8hysm6G42Z7EUYYFe
4w6xcrr1Iv7OsTwXuH7ak0uiwDSQ6L4jF3kQANVzuqL5VcsMFWquPAPpWdhv3BMO
HAbDq+8PtM0RrAFdh7Gl6+XaVGmVRpTAPQH1tFyBwieAwtgSiSEuq7xwiY6+KMx/
119cZn+SfwLPQhJ7lJywFJveK11M+0Crmnr6t0yRk7Rwm0UZ3WcDbHBlvCuCy2q7
ZXvlr5uc9mi5f7zD+Irbfb3RCzsmybWJOn00U/W+bTj5RKSnorlqnbRxr1tKtw1j
Mnr3sV+26i2wLjUO4kls4NKGxcWTbJID5qerk8D+sg4b4+wj4D/Cumd4fG6BUhpZ
FOEnwuO43UupueqBXzgL38o3zq0UKQf4NcNhNoGMbBZS3PH8PVIrvRkYcr23IPgA
gUSusmuMSSCAmCBPxTB6vermHiQjDn+BOsj198hA5oygAa1tNY9T6bp8vZJhHZBY
gZBnWtaLQO9p8c9tZnVWkpPpN5FqXznMDeMNQfvyZXlNzEquFyoQX/I9wXuuZYLI
kZHnBoBQ+T1TF/QjXJHs21as4PQhdVczOG8r0OXhgiBM6dhe9RZWdpusH0bWb9Ia
DfM06k047TdEajMEviw7h3MCwL49eWKymNMrhHd6kKiXqwRQOhntI32NGd8gJf/K
55+J1w6+UxONffn0eU88CxfNXKLH93ke36XRGtYERdgtnlkqZVKeUu9/VrzPspje
27qU/i/G8+QsWLxR4XbAcD0E8omFTqgWim7mfy4O4vpHx5d076xp7pXRKumYgD6n
Nds4UfQ0ah//5Kt5/BjZytgcMcjF2/b/mqX9eznUc7CJGH1arxB61ldOuGVOe9bL
ivI32Q2hbB2P790RjxeZothFf5WydM7zJmqYLJX4li3p9bt8SFgT3jcUdX/vofcm
suMy/2AvGpfxNjnwa68hQtx7V19g55y/iv05InvE+Qr8gWSskg1FxMY+4cy8ueb+
dGm7bA6vC2/0/v+UhNHYjGLyXVHUo0/SBXkwMmCGtrSCwtrBFPL8bvOwM4cDg+xM
ztP+vIoEgkLK4x7WP93Le13HwzPFD3GV9gVbHPKFWCJ3LKiMa0mIv2f+RDFQ3Xrz
AxkZBQq5AL5M6ib/j9t4t2FVlphTjibUhcW6wQ+JztQcjf4IN0q6rUfOgPZqWhXK
7NYWb5wnkTJ5EX/ln2pf4vl9f9s6MD8Dl8GpL+Cd/lQX17lLsiol0WQrcPcpv8Ly
weZ2teqvVi3p0xOM5LAIVt8XLGbss14viDj8mUP/ZzVk3hK6NFbmoGAQuZbcCy9C
OxmrLOoyu5O2G6wocbJTET8mPEFOblW3rBjVc+I0jFPEsCez3YhIDjWbtH87o6A8
G70vmA6/T+gRhPpVgIVi0WyIZCvREuccVRxY5bjHIFJwv6hST0boRLwlG1lREvdI
EDbZOd2yAOhq+ktFpklTr9FZ8nM0121a83yfZDPdlgu1jLQWaNHcT1QhL4zQ0DA8
fAtyN8UEfVqUf0P+X9/WFX+dUdOP018H9GTfPyBaAnZfDBEDDKhbeNVo3IHn8y+K
u1bNvIs72B5bJqU2TaT8s8GBAfsh0LHHo9FV3lRdSmEqcPclF14A9GSmo2iKVTMf
ITNtyAyGIk9wL80jzGk0rKL0yKtNtulsxhcsF24VntyFd1scNruJJlk7JTNt7l+2
UZFMyNvC+FWJ2jQJ9MDLgUH9C8hllWwaxuGZk2w6ygGoW00OSnpbL7ow5eOYTdp0
hWa6nxmDTrEYcXerebgol0Fdy6aFmbKajTpdn9ieILkwRgsfGVMHf/RkMI1l7bAL
deMTQqd46uoxMYBO7dGOfBuf1c1mfRJaPdtszai4fjLgdJA/GkNfV4lPEefYsQEh
bv7xLoK0jzpHMYx7jATbSyPFqTmbDyFvUnvX6i/Jcjj90gfWG5zkygEayQBxAbwB
FV8D8xy8u6c8mR84T2/zLbJP6LSMasul3QJ5H5SeFO8wxM4j8fn2oWitN0ouUkdv
uLTL90iUD5v/5p8h6i4G0msa6gJ0A5NpHi5zESdARXXN/qQHeBxXR9a+F4nnIyKP
5HerPj2t1pZU3iRpJZt/dsrKkRulTZXvbDgSdv9uIuK8vAdmJlNbwoGtAhbcvJph
mVABUONA4Sm76idxjkTUWpAj7oXcvQim43O24IB9xzi3wghwX1BZCR1wEJoV8Wli
SEri1Oqh9RvODysZ4gm2KyGBRU7In5DoLhWm1Jrc3ZWMmVrrArj+fM3vx98kicDs
IrSxEtDlwH15+y9bGmNQkOrPjOuVVAHxyTsqmegTtAv6x5R9svYMV6msqOFjz/tK
oF6EMU4w4I3URvx6EQqYcBig5DLxUssWx4Tkv0MGL1EyQ7ohst4emoN97kwEsT90
5C0t8vyjSWFjUFjT5y9uTUZrntFL99Q2JfbvOlENgDTpN+1ZYdnMt9WDJO6XdSqN
LzjhNN7vCsHc8+KNz3Pkyc6YUmE8Lm5JT03+y9u6Z8P/2eRuZzYlRTVXqSbvOkjw
yiMp+IXYsRZ3wCpHszIIzJVaukcQyfT9xfs+jLH5H75rzu0k2AisGNGl9nprkbPL
3inx5pnorNdEGkkeU1laWvTzr8nIXCMI63swpJB9trYMqTHKoqktzipwRFUVOwdT
Nx2NsjanqWk6MRhNSZuOhOW+dhdCqGM11LZBY8thzgFeHHliQUZPT2dNr4tIamo4
vqAkbOZgUWonCT7lGFyKwtFos0S97ji4CqTHxHrQzLqERM3AJpAWf5XcCtkFPozb
SGYtJOxFhJBV9NCNrZeUfEmOKHerIRJN+r7PkergRKG/nVTL9hQfCAI8JSppm0z8
aHXz3FP/0eJtOqkw4MRg+iHkqOb6rqLjWB60w3LdDVsw4El67Lv8HpiUQf9uW7Il
ftcNTkDt2elkcIEPJGohDLb19m8xPekmlamuRi73itu+VUvxsEakK9w0RDL0ASdX
NIsXhCug3z2F/X3r2qIiv/Xn6IZj127N/ImP4nyvklQa/bbdqnTPdB1vsmqJzcon
0izvpQkzvHBJJN6cE28HVo938JP4eWWlX4fHJVT32mTgiFridKl7rD9vJDR2hsK2
HRgUYuYaur53SUOjWSXgxLkCN5pypSXfp1p4o2D7e9M+rCw2sK3QsnihuCKrFZUP
yaLbtdDmJVUWXO10A3CpgxkvZACWHCTCNxaZPj/V8tA16oKFOpbQvtX3kCbJNDq/
0gPgvpYlnKnnxCQ9vWtZClI/yxmHjSwREzAWcsYUa3ETV9ijLf5YRmXeHBjfh3CK
+U8f08BGkoD6mu6og2ZJkwM1vd52QpO+avRASJe7gT2YaF7jB0AN+6taUWugy7Fh
UnrnhXCJtsDLimSJcqR9gywYZcJ+eUE2starE0Zl3h7UC1o0TPcRPBlqXK+17oLN
DRzOegcrMTlVh71YFMesTkq7kXOu/3VJaTpzMXFM2DVEgUDdv+REpO6Rxy/wg33X
6GUWkOWG0pnQAnbD9tooICWDpywcTo2UFqfPhWxc5juKHE3dmPG68I8/SuOqoly/
9KkYxlSzmdU3L97BAnFOLfaYXvF0sMkJNV+8On3HIXKI1uOG6uXd1PGL2McO0eZG
l694k/npW8FqexPcqpQYW89xWZ1y79GoPtzRpw+PhXMM1U82uy1wubqB9QmyJjom
sJkrGdtB/mFK1/nGvZzwUx364GwBD5AyKT6KNnCYtpqSAoMhx7WTeGLZgx+b87rg
oRaPG/lwTmeYT2XWVHiP9SPAtMjc9hKGvaAKwqRul+or8UfEdH5Wt0g0lnpYhPj8
S5OHArGJWqthncKapRovzKWo65kZ/aI8e+IpGQ25r1/QzOvc5JNZg8KUcMQDK7sd
QFXKZycSF9IwghA+Lq/NwRvFgGJ5GkQESFLsYbC2+Mwv7I4zV2RsEmBnQFeeiM6P
30k+/K6DTZb1n4P7hy2hL0hjYKmSrBPU3gEgQANctzJadAnd53/tb/ibE4p7WYkM
wc2I1aTDVhiBRKu3mQKb3djm7t/m0ku5Y4eXkj1GJ6CMuYLyOrI1ZrWGDVxWv+Vf
K/S7Lm8JtycNas/JCYqIqXlYM3kIT+ziYAbhE6dF7qLwoCnZNbzsOxYSkha5FtH2
Cs60NrFrUtCLT6XNSkvKujAGD4k1H9dJWfTFYrJGBnUj3b0MEiycak1xt43DngqJ
mErYMpZGse/weWH5S2f3ZPXQyBMN9SmSx9uwRJoByb5vO7U5r8+phWsDcuBbvdgB
1/NUljQeSl6rI9sdLmzUOmAoIdRZG/W5tNAHnTL50QAd+kHEmEEzxRoAIBVl/41c
BPDmsD4R3gPSlhoU+7Y0JDL12zgaxIOqJF690aIPeueyJ7SnMOCr6Z8Jin/LMN7Q
eGhkPFweB6hKMSh0GfFZYkR0QyKEOY0uudlqM0bOTe/N6LoNWCSXXxyNNkZp8qw9
a4INC8iCi5DYlwJIErHDWdRO5C9NzzhDyrVAC6/aqucfL7rOF/82l6+j2x4mBIVF
FErskblaQAMhssHaXhSYtjKIL3u2knnckeyyd6Xg9TVVrfYb3vjQcoAPAVSOaKUs
MF3M8JnpwSlhdp0TUQPLZK1Hwbf67Ozzl4hkvqspCWFLB/8oi5j/PNiv8ML/kXcR
onMHP+HvyHxv6FzZY2mn1ZBmI9JizlQRong/8AxUjPxaPjtdVvuKS4+nkZuJazm5
+xldX878saWf9dqLH3cWlz2+kdeqD0i49Klqvxh32PxTy7YVga7WWtpWM+pfYyqw
qYS1K1jwRUkSjjLIOlvEAG0YMGbcOTtRfGjoekLg77LB/Nkd/UFvBu/2DLel77zC
x87oeU+tzA/AMVJqaQ158573GnsbbA607Cynl7naYKjfrtgmO3dPht5gS5MwPVZ3
cAJRk5jqauVndeuBeSxm7x5cL3ELExAuRzvwS04/FXus5mECMsEtHgKNtetWZAF2
YdX2oNm6nEowLv/PC2WGRfDc206BNYCrdG/Fs1e8HnnHVahSVyYyw+ueK6ul9JqR
amtuK+YAgavZN3OGGvh+JJafUQ0j/jWzrQdyal9/iiMOVbj85B+RJb9w2FO28R4i
m0TRur4t3rvcS5E1oICMj1l28yHaMb94A8xekQFxV+bz7F+6PLgThP/Nn+wPkewd
jiNpPiyBoyX9YYTJtaj/FHgk/LbTaO4umZStO7YzkWxakYv4lTcHOo1HXU6w0Bqy
JFvgUFBaobbiun7nbCVK5q10WQqowUSr8Dasq8VBLYqWPXkbP9roEE+IQclz8vV3
Do0OCy5IJ4as3xWZDkCFFV/+/QdoLHtuf7cnv3LTuKrXV17bZnY5cLmVQruXAaeQ
cAVrvsiswHZ1QbuUMG+e8ciuWaVd4brWX0VEo7AFsGh/GLIcqVkU9iSIAnlFZa8O
hk5um0q26dRneJ0RFDYWCb8uRuoEL6G3uUE3Q1UD8N8CnXTxseukJBbx47H1gJnp
XfiAvRb1YwwQcgYKnU24laAYO+m9hLpTbVpEXBZEbd7lv3SnVznR2NmW9ghKN1B+
3OnVy6S2DXhdhQB6Z7JhnQ+66WnvE9tBBZ/U2rfTnoFe73227rlWSFA1SrVdqvtt
zsivl/FsAJv6T60b8zydwt4nCVw5YkRXqT9LDW601xH7M+5pLG0F5Pp1hoG+BPuZ
VdndFZtE6FTRh7tP+S2FM8ZaNt0kQ4mnIXna8qKKep5VHA8E9hcH6c+vg9AcZ35I
MZEax9pHygUtcwGTAQbNG0B5z887zS3SE0TYg8P9RoR2R4agIc3nF2h/CoAAHOAj
8eHsQ/iQvp8f4gDVbanWQTNThoatiHEOQ+jVKqoOKsKacFISkHxfiU+cJoqY60O6
0V8CQXxbMiERGMJSJ8vftnzpbHmjRmmLw70CUnjLn3PvwRjCe/ceeH60skDuJa5h
shg7D6leZ8JR47/GG30eijrCh/ehsdL89mAdZX9/qFAtD68LVesjUB9NqbhSPZ2R
O0U0VJ5OlswEZufYIvDx9ldfMndtbsksnFME6SQ4adqoohOPGZOkDCZH2CxWW781
w8bOSAePu+pVpe4C/g3RjXjUIzPbI4qrKYQP5QPCF3XLNHbEC2krNfgHZOx88ZsC
6vXNq0too6zIGxFvDlF7fwUpmaonVlctVQWxLkuzrXKYCcZMHqqBWGJxND0bhGiG
mU8ZquWwWpZ7zhVOI7U0fH0+Exxlhu3HZRiNAZqahSYhP+uv0ci2igQV2H1DITL4
hDoOfS+CazUQOVxjb2sR7vqkuMRNaq/cZAjrQ0FB4lRPBCK2WaPhlGK329wed3pq
E3d4JUnllPvFm+Nik69hKN1z5PN0uvZOgHuS7uQvph4k5nWQa50xSgvHt7zbfR9U
PDc3p8fHG5MnyWLb9GtZUeALkmgm5hnsMqrdn9uwo32ihnnvqlWZCgHZVUzqji/R
hkV4oTexZ/VH3T+roJHQtZq9mjopMRWPEmdjxCmbrTg3+RvERi46IBYRuEm5RHNr
VvM8dbjuTWivgCuW29GSf8dDJzrNMc6Fmcz++Ougza/vmc8ibFkYTCHHqVuTh1LU
fvGT8G+NO/nfrIwrbrZpR7s4UdtBhpRqB6dNRVgMObZx1WFrucOlJ3ow2JugZ9n6
HHZIpg/nQvKK42VBZ8V4fYEzcaE6ygL+vmdHSRieEELKv1hbCZR1sFfQuL6VG+S+
UVk7CV6t8w+tF7H28/05nVp33mtEZ0tMwrxy3Criw6+sji+ELfc6hfApuL07NS0l
6Y6QobK9daL27RRT5/b3y2qqy5SSHjEHkSj4XUd4lC9vXcoeiA1/JjQCh6Bv6Z9o
Ie9Ym6F1dRiZcadVKHf42r7gQ+M/kRTdg9SJag9AOXi179kyrn03JUoglKqHDpI1
SHjl4hhdIzsh+BIKvene2RsUGv4kFXG2mIK+ozWJkiTvk98j7fYCVtMRAB2I+rKz
Va/peK/8EnDujNwA6/5ZZ+Ua+KdFi8/ycr2PalNtAEgXZ656JCNX98xtmxqmgrt5
2pxWltZlmw6Hm0MmOtFJRovzb9ZQRwfjUIcROOTIXoutucbY6G0MzBTL2MujQOBi
14qnDpMf99IcKQkf23v0PptHmrSI5wiY5CqMEAqCJsdOQALRNZJiwiyr3ATDnhe5
Vs6o1t+l8axiUDljQZ1gHD+6yGHMucbbQ54D9KYjbtLSSjoSy3RXw6nAoHSMYULd
wZD68WXxVCkkIWS6h8Gl2TOva/z+F+UEDoS7oxsgxBJC8IZeBKrS30TTBIa4D5Fx
5jdq32FSpbBKihWQpTsZjzItRkHg6P3SV1BIO1iIE9BO7nqd/H3tmXSFruzIGrg5
gTmJ7q2asbK8MzU/vP2B4b2somN5huHihCbVhH+9SFtOXrGWHzJBDxXZFfRDBYTx
fvkvOCW9BVMQweJumMzU1jgaZuBq7MeK486w7uBp+78gN5o8pqvszXybrL9ORi8Q
kCEhqGv6QkkthFAyeirAz9d1T4t8VSqZ32oX4KRuMCTghWiPo5iVD9UPScEg9wv6
9m26Ig9CO7G/U3v79iy5M7YeMBmr93+mqry9ZGhKonvgTwcSwZliPQZP2+VZ9tvN
5gSZPB6T0BSW5UbXk9dt3Fqqrbct/nl2YreS/bERBc9PsE35ScpsoDDZ43NFlTzQ
LnoeVUytMIfmo1OmdNsZNCx/onzI13jjFN6ysuKYwBsYml97VNEppWIP4I1ANZyI
/beFcQv83R32jZT8PoCDunTy9dt1d0ek67W+GyrWmntrjY/n3nVo+BOKZQmZsawC
OXcDSg00Q9/8rzxuIOeJ1c9/Gl5MnaL2mIOm265nCwHB/lhYgJuOqf3JT2040I2y
a9OzV4NWdBtWst+XNnxEaBTiwLSpdsWmxhkUR7W4cywNFoZDJZ0CFBq2+JIjRBX7
qoGdInOQL3kIptaEiKRdcux2jddWyqalle/6l3xhsPN23o5z3+K6ymm0cI4zopH/
jsoSnGfhiFNTcdnhejGbOG2bVCrm3dCU0AyCxDWR5f0ZQAJ4PTc6pOYlUeyzD4ob
Bj9UFDVyhnA7sbI1XhTYVy8ARiZAhbVlODm3wx1BlThopGlh887Yn1SS99gk9iv9
vu2jCMT/xRt+HC9gcRWk/owo+Gg42s9fMvz0eKlRnma9jjt9tvlBCcBEbXKZ1y86
pHpuu7bbJ7U/sIbROylvS3FpUHlznGvGxb0M9/jFXODVw+Vun513eL5S96uljiK7
ydrT6ev8iE/AGKHml4oo8732pSV2alntRvs3+pGTALZEQACtlFVJWMs2BFk298Ra
EY4T7rRl2rW95I379giFXDhEEushc/0PgA7BRNvfhL18kDJwU1RW6d0VECqpK1nE
YQle7kBXJYVcM9fNCRFTGY6UAuarD2uEiffj5hh9Dn9YXkE123t5Qvz5q8y1Rd6K
cGguhucdgymdsZjg+roAVx++LxMQCqf1F/gTqkCzVSQC8+0PolSTkfzoJQ1KKMa5
dHgHk51UngV3OY1xkVjMIuUJIaR0/YCwTNx5tjt50fgshZEVliPUhKs3VvSSf6Aj
kTvLhweg6NXZfEpame7jyerMSG9XhDUFe5oC96CBZAT+5zJ81LUPv7vCFLD+UlW+
0Yjj7GSp0HgemuX7m2FcuCjfE+m2WZkB2je26y5XWPXvSdLCnO/wAhzf1gI6iO+5
ZaTyv1vuptc6Eeep6bOzxXZTZh/QYITIlIFQc+c/zR3GcxNL1y6501vaCcn/evid
IoS0VRECeu60gcght0tr+Fe8GSihnWJjwVC80gGD+5SgdehD7n4USfFBE1rupScE
jH609KzTPeb+PwL99z+qf2SG1wOdvA587XFmSlkT4sZaU4duLiGXYiwt8cra6rmJ
rNjh/422LX2uS8EKUIj8VEAugTjlHs64ndHHX3D/zK7RSGPvpEeMURwnQ4KVXDQ7
FD4g1jzHymYShBiUlR/eg9eoW8EYBuERJi+SfqoDDuERkZMn1n3FjzI2q/CFf97T
U8So4pjWEwHgS/lOcejh1+jxNDMisJtWf0Lg38p29P+z2aZIVcCzKZhgA2aLbMJK
9w/9sr6od0taICMWHIwRDCf8F4sDK6Uc12ajIZKamU1O3XeEAq5rl1o6piNguGvA
1KZlmoFjIUg3T8OgVFw9UnHSyiKczw3pPdJQHPr3uMAipW0X9EKjW2H89By5bzGC
mWpMSQ7E1HnSCmluYKcCJCJps6XbAdGMVdyS51X7kSil92RKObCg4UF/v2SrYaTJ
vC7ls4iWxef3YdlQpv+QKZS70Imz838AP09KZFJR1t6WI4DjNx/nzFJvFDOOFzaK
QfC/2XnioBVOX8Mx+KP2syhozpw1iS0J/yzc8fCEURt/Z1zEqeZ3mwCYiGQIxzsB
oIty7LVdPZ6SnsUlrC7yK5ESu/uczTvOKQ2awKvrTsVX+qSn49jU7EeqaIIRbtdK
xJsnvofvHYtd85CUnInjNx5+G2JDCl6RgNgPFD+Ppsnu0zvzFw3V0XEgZygLzc3t
0kGyNdAwGzFm3EnQuN17XLP82Jpgm7zeUnoxOGybSA9hj3OZZwaPACuKCDGka5pu
Z7MdgruoUEdL+OvrwieW1/KVVMsSuoINtLgvCNuxyX+1DH7oXS+ya46mWiK8FPJ2
NBt+tpkxHhmMF2miLCMODvktjJU64Hor1XtrbU7efraM09tn7bUolCrTGj6TGtp5
yf9yKfmCZYkyBf0UsiD0OGMhe0if3PMeDDBAgmETQL1l12LwzV3ev/1bYJUN1wdv
26JX4c3kxGuufPgxHmgk+ft+uGb/ckHH2EWqnyjMnJA2Kn1N1us+qTxTELTIB0bw
z1SG/wp2TZXh0HS4Mm3W6PzD9iZ3usLKPnos+9/Sltql8NHzserFVvYwe6vOv9nL
6F6asYnSb+90lDBfuR2Rgq2CmGv8etXM6Plbc2LStS+K2D1ljyhDbKiuYO0lWjSG
WPAYTMbaebGRE3w28PtMjYzbqx81YLbcxGAnjW3ZYyK9THHcPjGLaXxgofoNrEcG
WpZs9/C00YGPDXuHtrf24KcEqd0RcqefBjCBtW0HIHaOrxLfeUqrBNKEBhaIKJo6
PpN+ijfrjKO4diZ1FX9iRBQdvRUEvVdvIdlAw5s766aTK+hhf86r8vCSocJN2x9P
+/7av/rEpx0JZEEJSyZQ9WuaVCKrQCjIhXeU6bkz34m6PNBf9m3xJN4QSsn9nxoq
0oKUlx+gg9fItS7P7vkCbRTXk6wBPkbNSgTllskqhmdoMDYMDNYmWY2ak09W4DeT
cncbwTspEu3YH/rFPeAnmfbCA+HBaY0jVzkGv21608thabrXXMMDhYQScAG2kIYE
QiA9BM42J3JUKOhjMqwhhPKuvgFBaXVHF0G9c0NdftGE4Ywt3KliN2/4hcG7abSi
iMRt5XVqUQ8LRvePbTJWaeSXcCJro8Rjo4vejJFDJH2iy5HeU0CpSI+o/Mr6yEIc
E6MMnjfli4Kcl5BcDFfAL/McBFdGiDk4YNFxfEutHT/239gMOaXDLK/u7p0oKXc/
8fgER8QwBvSSFonWfJJ55FtZpmQjL+mHjeUWbTE7YKDuTdhF+n601XnCp64ectKY
3sVt6cOKl1KHwU4hHW/n89yvgaEMahhezDaOFCYnJi/2kQAzEVHu+AyQl07czqGc
We79HXY7yUZEgiFzh16hAdqX/i19K6e1eiJhtmRVy8gTM0K7FdJvPvp/XJBFIlb/
vaculJS/L4WNkSNMK2G1/E4dVmELqUhszCisYzL4TgQAoq39D0/ttBcJcUeTg5Ba
AYf33nRT11Zoo9SXNAWRUVScEPCTum/zZzPHQfE5OKeaG+bgLa6SK81hm4ZGsA2P
y4TYbReVXBZ4LputLZW2Zw4PbTE9869NxasHqo2H52jnIhoOTgLz373Ynml3qdwg
eUBsiRRNckhXsTY/b2V4DYY/8n+htAbhv3vpO0L68P5+1jGEcnCmI/Bd7GaS/YDW
GcpJMfhfgr/JV2KsidNcgZWFRM6u+Jqq/FVBO61kFqdowaFLcvwcwM+8FqCawRG8
8G3TRkDt5exl01VlpF3pPjx8kcOKGeB9YQHXEtNg6xpQrXwAhcRbbHY8B8dTjups
IGQVc79DI7MX7aM1dQjroF3nfMGOU0JQZGwd0xIO77JURZ4YbCdDq0sw3T0BIH3+
Ef+5TMnPuFg5RBatpqR3w95iLC0N8Tln3NacmdSzkZUjefpFd7FLhxQ1fi7HNTiL
XHUUX1n7cpTpIClQmossAfK8voCJEnXvFXnVvmMJnKcf1J0QFrTGhSmpN43LQIRc
F+zrqdpcORsgkqxfrCoHWZQJtFDSpM2XyoNxOA0vkmeKbFsgjBlBMJUH4/kFz4S2
SJK/JkHaASnYJqUJMBCEUBnIepYG1twBRns6FdFMts5yxlQKqEisqZ6Uy2tbUf2b
iyyPiW+Qoz9DvkEGIbN7Yj3JL6paRRmC7UvusT34w/RjXQNaumCUtVpej9vJgMdS
yBYB16jk3x2VjE8SaaH3ZLf16WYI80zB1zkZJoCHyYTzDbSQJ9z4T4SBe7BXA0QC
ar61iPkNFxfYpuuSGxkHhqdPFyGj27EpaJpGYMjevg3yD+UFOKUxl1aooE03a+4A
7ljBApQnVskowFTIWEBuBhTgygDgXTe9WjrBGFgFAzjQqzO9k6I8TnfSRG7d8m/Q
LQ75lG/OFtf1g4FtuhfY7tnwxQtF4A3lT4zgblxN1sroDAXtsYnIyyCmPxvOz/IN
qhC1JB04S3hVnbg3iUfJeGykgtULlXtyJApenwba1XYGpPVC9lEfSdV9lmLvNRWa
DxqqXRE1dZD669zTDY65m19miWxKmQ5grs7p1Arvk6m5yJtRraruaxm+jihkKSG9
AKi7yhz2c7WF80k751W9+uf20FkdVOl9DTPE/fIdvdV81MrpGMnOvsJx9TOyEBkt
klY5WqEdNs0Lao/CtV13GGWXbKWDvk9s7aImEvA0PwmterPOMz6R3QLAEZ9XE7Re
kh9OSo9woflAr04sEJ4BbCfWLyfe5x7QpIVU0mIkSWnYPvp8Rchz27D90ANLNC47
rIQPqFVj/tKP5B2tuVLKWgvKxdqmSk279Qb4Mj8OQfPfOSO0YRCK95nO6E68XCcH
8OYHhsqhcTcPUZtD6YV9H9BErifGotpRHeLxUbcTUPWmfmBt9dP34bWBlay1db88
bkB1b50p3MvoshZzpR90hd5QB7B3I0aWvLl5kF7IDs4+HFqAXDnFb+Ccn8Ul0w40
bYUtAF4VZEGMdPtOCC+TKkkVz/QTghg40GQE49s5kjgn16moYaeyYDlzZC25ys37
6eeyz8N9Jp81BMLFhWvBzHHnWnEeIHiF0YSNQ3eI1cS7f0saMVs6l2uwTcLg2bdv
rE1uqRd7BCAt+n+cV4EYAdtg9iqyl0t1V8pVIXA4q1K6F98OCcBcjh/EYOvZIJWw
4NjFMHOeRkTEti4FtrfEaoH6bqAV/qB75X9ya6rlMJyf9ezhEV3uKt/b/ufR6rKz
GFTZjccANLrnf2DAZax6gRAfJgfhFweZz1jv0hPr2Pck62OiBfxeTXydv1FcR3Cz
sR7YS07KzmgpNHc69tly9zM/D/UfuxYUddsvQAIs29bFt4tAk15zkCVLWHWUPbrz
Is2C2aYyXwygBnRu7ST92lVHtWDHYBOK08/coSX59PYWiBN3mf+Q9+HOaW6syCLI
W/zB8rpl09G0Rru6J7lwoJAYQFyZyM/DygBisHkK6qDEe68/3twj72hijOuX30fZ
y3NUkgEBwMv09LRTIU17b1TDeXvpuBhoEjj5QggPE2/QCWdGeSdQsenc0kzkWVQx
z8J5tjzGCOPQvSuL5h6o3L7B0iEPwQLXGUnxnUKdsTAi7yJNWqbaKdEUME6lCC0G
STIPZ2K7lEjWC5JauXR+X4HGvz79EVtvh3QadFPxLjjzEM8PqMCCCyQpP71OydA8
ep4lHXBwN/Z0AmPviGSkKyeaSrWk2/57GStzMsmFE8YWSvHBGivzETT10sFSQ7c2
MEh/J/O8W5QQpLfEZMOEbKGabNtipzrWFCcOtfzxtxyDFnTpNVtUud/gXvO0hp6n
bbbXtVdu8dZM9mZ2RbBhORfjHc9iR+1npAjOE6v7mU6GQTQbBfmPHxUlnsP3yd35
XU+vnrxWOk1fu/bFrKiUYWAc7tUnT1SEI/qaSHCs3Hf+FpHLXhvWYYIgGLCo8ZqS
iHu9DuoUaBZEYLBukB7tlafq5aEiPHkggntPcPMuDnmHqpziJ8A29txQYTe6WxTf
Fgx/fLCQbu562UrdQT/XWcBQI8lRqx4703EuD+q6o/3O3SHNSgW10Aa45hX9ZYhV
Sqftg26SWuxeyvA4p+vRdvyry4DHgYNdRimlxFSvoYk373yoea/pMsU5OXOV7DCd
1G8q/VPaF7I4Uc13Qcdkc4CZFb9VFXqXPCxFHSEhUa2fBb1nG//hSLMICadrIF81
n6tqHu4C/azgAzpdt8iP47+V/IHcXlGKkzJ1U4Ez93McQ0ZmWgt+DjNFtkutwBkl
3xk7js3exIviTfrCs0GBwQlEXfcNI3of1l+s/ZosaN7roTDu5fp1+wLIS2Rx4S5r
/pUlqRyGXXIhx3wDw/90gcn/3gXyaP8FzMo+aCmSry10bv9l879ZYtYu12nKl2qj
KYqyQNNMzPhYTxnv1PA1zxTvoy5g/2lVTYXAqi4ubYPpSAzdeN42Nzbnn5s5BjfO
Dtc5MIC5hXQChrx+7DaI8RLXnHzThtKg9SalTjDrurNtImzYS1DQcRBgQlg7BzcZ
H+TJ4B06rpG/IXr45T7tspLC4AIbOMqxlPWVSXMhMBIvOg863A/xYfJfpdRV8VCa
vcz3YxtwBSTjSiz/4DzJYBjzw1yrhCSL9TNH9tr1Qx6ufxPeymatO6ULk+PSFWYj
6n+OjLQwPtt8vl2st/f39agN8oL9YzKii+HR09n50tCN7yhKtMkcA4ynrff3xGuF
yzGvDwE5P+a2dqG3EWiPUwt4VLm9DeeMTh/uvBhanc98xEAbZiPNgCnlg8lq8u23
BSK5bTWBVh9r7lyjbIaGF3KJn+v0z4q9nDsQez6G8PdYTLA6+iWxk1XiHRk1lE5J
X3R4186J8qNN1jNOFGXvmgNhc1pHRNH4J/NxVCa8unCOS4eRBCZmPb7E2zbtQmj5
2R9Ui6d6dCb7L6039fA1sw/0io9k33xjsfHy4SONesbA7nu/W8CZ5HT4z7WpLPhH
YOn1czsV4MbQKJy7ZFQ9+xRJZSdQVZaSidpNcwWfIr0pT0WltUMO9zRxVrL/DPOl
sItCDORVc9amb3mcgM1brgErnc7c0zczA6aYcLYk4xhmb7CIThZvbTJlA0XlnogX
TSIE6dz/f2Ji6hRgXUk82ne4CWz5DX6r8R9ZWEZb/UHNavHv33dlj8L171xpkwtA
zhic9njw4IJa8ZvcJWqnxOKLdGJRYb/f+acVYZHpNX3GNq01PmmilpVFYOzGpTfs
c2mymD0oGIEEoVUShVcV+xQkujuBekVQooCc1lTDxnvr7NcQVZEIP8ji2oSQsDUc
I9qclpIntK/4bCERvlT35mCS3K7YMmYO2aonHNnAIUU9fR0qVJJNfOPBKuxLIetu
wKcuyHXmJSAniH7lstcp0wf9wVMrv+7WPwIbij2onHuNy0jv7+RvtUe7V7Z+mDgE
yBEHSnf4GRlFH/QxlpLj+wn9muCp5jEJ+DJUqSwWYnBySWjnJvy/7V7n/0bhHSIB
GsN590iDMaJlUDqAtizGN93QssSHf/iNFgb47EOUnxaYJCTxEToBrheKHMmbKzHS
AptqF8sEUqVZgC+OPfLD/G7bv7ukIdQu/uQC4oSFVYSjqeELa4C9kdZzz1xvuomh
xtOmrS9Xao530lIxUX1WoFqtEVkkwyte3o/dAyDEQZyB7oydQ8ksSfSKZNGvFjXd
0AF3DGhnMCl3bX7+5uHMPc6Pd27caAhB19W2M8BtWEDlBO9cqaWMINEwQXIYyLzz
BaEl+dH+xtzoHpaO8DKt3TZraU2itW9/4dsRGn7ytXEQsqWi+vl+NdczEwzEBF1k
VnjTfJqpvXkEaxfiIKoz1ROoPldbYDQ3coM6VFah0MQuKfjgynS4F1x45fpFYBxW
tLZrcKC3E6WGQaKHg57zIueTVgN/cR7FKTgGa59tvv8Z39aWevVhrKKZlVtxowY0
9JoElpDVHKHR4lvEA37Izp3OslnHChUAmFUQ+9q1puenK5w8TbW3G0vrqiU70zwR
OiE5i2Ji5/s4l9P9xLWJF494wuKiw5EQwBxS72/3gbP10fDhcADKlzjLlrFP2rht
Ai0lPGNiajMDTFh41wtEz8glch/Wx6cyfyT4xlhAZxIJZupuoRBlygoS+7TPvGnm
Fcsy1AwZsZ6vIvck8hUvpIryyBeILN58N4XQzEA9bCAQabRRhhmcV/C6T8Xj1642
dwMUEu1k525UHRfZi8gb4W/cRScKCnR8kmvfT3GMJI7ONjnI1ap3JR78eAwHje/I
kG5qM4Q827PgT0GmTWHSSWYtQeQPzSWHaSs5WWJPJFav81iQ5aWEwhQld1neJZgV
5wQ0KtADKtxW/iDsSDyH8YbJmAAPu2fqN6ZCD98apeE1FcTaYccl6gIURzOKCxJY
2ks2XteBVlUaITZGAkFBH0uRF9lfOoNh3xG5zJQeiYwBQ5lSmyn5f5ObiSgbTtXt
Nwpsa/jZyRj9bhpcsSx45RApZUgJjClpk22BaWoqDqOUoVhtuVuT20H9n8knrSLd
cSC42/mrmqsyw59VVQqIXN+lAenbPp2PC/xhM+F47QoQkp/QNOtreRMHFwln0ViV
HNbC3ljoqtD7TPZNELlkNN5dEKvRfgkR6MpXvuZyH2g3Ezxc0CBI5O4Bzv1IdFLq
3znEgvT7xkY/ZTWVDKowxpZr7SivzTiqkt0fEa7oZJmfHhDERdO3F2PKsPlmnb6b
w17zet4YbSN+0SU6tXJ9ZQmR6/vnGS9J2Fta1g6nfkSesj9hRxYNUF4H5DsbjPWF
zSon+15UpzjroKVLdUVW4yqAvl6eLuwA88j4SZQ1H4T4xaYcILe90kYXQgCiz502
b1MIopC9cXAsF/fHl90m6NMkIbykDKvq2aOQ84e9otAbWZdb+Jy4ozuGK3L+/PFh
kfJQ/MeePXlEmZ1dTywVn07QHfIOW/IPpK93crDG1hSfFPXA9S1AnIc/pJkWTDjb
ounR+evjLi/ZZZcu7tNCbqJ6W88Le+PQrF2wJZcvsFHVeCtTPB+DMaRMiaUvJMB1
QZcaqTJdGjsiBp6N2VkmOW0phj9+jTUGIa6cQd9KtL0GQZwG40bRkgaScqjvaQzp
ZLCk4FN8DmneJF+qYaDzeFqjkbS5Cw7vI7bq18m9goOmyXLxMsM4We+rMHtz8MvU
g7JmInz8Jixhv0lZ2CjAt+MgpSefJAAiJbLR48umMozWWaSCF1WWNpzYj9K0rHy5
9EvxKUTFzMgAWfextLxiLwd47thClfzgah/mLNgzto9XAPthp15vz3aWcWEtPpoj
uIBWLRk6QXzYS/hrxh2TnhEl8PprJrI70CA6OxS5L4+q/PIwBrTn6RwlQdtyqOEv
h3j45Q5WnNg9oKmwB1jxf3KL9x8hD5ax6+/DBjq9dtbJ3Llo6nlnGlyX3NvRRm1g
YFtHRaWP0DyQBtm/72FFzIXvtMlrzLVFXAXCBhBapgyXJWhKI6F54zWoTE3ou8ky
HM9ohOSXVVDQT+9KclhcqEf/MtTndYQrrXGIkHEcVSCVwNmAH7QyIAIhtX4wXvjN
658awJL6IWuXPBwzP5KMyBz20YYPUJVvODFAYxku3NZpTPdOE4Fw4YIeBUDHWupI
FrL8NBtXlUVqYTNlU0VrePSS2iXmD7q3bgxvv3aKoHjEUtgFDuhbvyluQ1n2uarE
iW2zi1KiA71Nvh+d/lZXsfLmkpfKZ3XP2UPRYOjHnNJTso8UGkwQV2lpWChSSZBL
AXyZJzDGOqcOR672xV6H6Eanc0ebUmnWV9s5t4qi7tHolOZP1GhCZPIrOcfFkJED
je68fIssTZka+wemQGmrQjlz9JL9OJA4SUeYS7Mnjo5ljxHRtroFTOaCfwlJkHZT
EpW5w+dbWn8tJ17y3mBM9mwoi7wdaYL0/WBYbgF4qhWHrwSwl9ukNoRChFe+7RXi
iKeZIMXEnjsyptmhTPBbBuut2NQQDXMjHVvWVSZ9nou/T1KS4TtmfbEsICBcqyIf
PhRhhddd5wVkrBwiHIKUpT17Ie7jcRdQYL33/sZxWCsgFbWVAB0jJTZmnMfTYDZ3
vZXdQKvEojJy9uLRiI66oYersvD5mAfPyLAnQp4qpqTV7518K5nQrynr4YTwV5xI
g+5Ngh/2V+9m0oUY3rR8h8Bt3C6UGs4lzci0MkpnjfU0/+hFFiNDwiBIvg0zejAv
4BYexbNbiFmfrjHh1sTTm5DRlwMTw5KoHWC7SnAupCy6W5SLEXm54DwjkHprMYKw
YTHpfhbtDYENgyAigGMCxeg9l1mBYG0aEdYWFOpQ98r+HCM03o0K/DNV5vo89ugD
Cn0ErVRLP4kWBK6J7iEtS39vJjP1K4wqEA1DEWZL8QZ+UQHLS6uwg9pbkYGbzNan
Umggld1jdKxCEFoJGcOrW2B5chKNwYapPLrmDB3ii3a7oucd4cCMYWgmDnlapCmJ
EOFQJ5KEAf9sRq3ckwYw832ScG+LLQP3ENAQq0P6/dJinGxkvXcIlQX+uSBxHFv/
VP107w1eH8acNxJvAQebvZlhlqqSMk3Aukqoi5rJzyqCv7bI2mbWSvsDDUPyb/X0
vGGK+NcVoCxFlgkiwmq5DI4yPeoMMqNaafe+SO/JU7GARPNUC5crzZxA8VYsSJSm
FkRnwAWEZsofgnD6+s3DuSDG9Snr+uoWlFtJat33bIaQN2gMSFoy8UyTRxRuLwp5
bsrqcLRl2EV6berruiPFQW08U0794sIfA2789p3/FHLyvqfmI1oXlw4t3B98m5v3
fnIdgoornUWgU5A9hiDgUziiFKecpD9TByech+5OmiDcZv4WflsfN5XNaT7LMxG9
A0jF7F2gpjejstwOEwXhjr0Abdk2/6ckhNAEcGjVIAUACkfHVsPfSQKrzMLXoZps
EH2xD5ko0ATUj8Wid/YiEHjefTSKPBw8cyMl2a/P5KyPBvRVwiaiDy+YJExvsyIk
hoWP/TMbNX3xb3puZ7mXwze+hgmLdh4S13gXWqmfmt6Xrnd1bkJU2IMOLpKbCc3V
8/c0cwlchjP5wh1TwDgyVkyjm0nWU7NWKwR62yftmwP0U2ngU0vjzW2xhjMFnzUx
/d+Y0n/2VbE+KOkG7htVX47q9VMoxcVp50SPo40oZkW4gzh0m0duRbxmYCaW5ca4
qzaxs7350ROC7JoFu2MAXN1RWAXjbI37fgFZdfBs9gvrN8PoSoqZX5slJXfRxGrk
4nbftjm0T5P77vetn4wrq8O+t54rlSKeJ805soUgOGXkhNbqIHBoGuCE/Z9pbQJ8
CaF2h9i16IHukj4AFrh7gIRY1SenV0n+DFCrVmNkuLJXoNRUIPJQ8B6e5jf2VU5s
jYHRwlA9qlrcdxL8y5QiSyNzEHwdDtJJzOhsZE/81AwNZhWsrRUXi8XFfCU9t8tT
H+wvID5ZhfGaxd9pFGeOztuVR9k9JOZsknzzmJCtOtSI0jAeWjTm4tkm6Wq8DI/v
1oW4Ms+E1VJ4SFvyqkxYZwUwjVSKLrf/4HH183IQzsMEYWrWnWdQigGnytSdJri5
KN3JoDuKgj1IqoM8q5mG9tDBSikVaG239LlGSxsqXF1eu41TXOy6V/Z7IRq+Bw6w
cxlA1pSweP5TDC9BvbjGFRb/kdIezWRYf0WQZkyZardUyQFuPnNTR+8LmrIIL9Zs
olvQdmNSMpWIArLGjcdFlGsAqho6XNW4tmPsGly1Cvw2Gh80t7v7y2h0FppwTw7O
f+kvMoGThf9bPGg4z4EhfibBN1jwXkUFdcgXJCdFaHl8csY71FZT1TGPxRGeV74Z
c0PKzS9e/nKexLzpsgkPbU2jrvY9uCmObsERAPEEd6gN3t+9b074W93aj7RXpzWO
W0XxGNmz83jHcMqNFMvKvffPWJc+sSNomQT7oDfQlep+cSSVrH+L+LqvlqtfE4Fh
9ZBpFCqKCftg/jqD2a/3u4O6eKYDgr1HBsMdzjERYN0tpxaYSnOVLUUaxwv0KN8z
HtHAm0YDReYvXDY+AJdsRjfd09AmtuC/LWDFA407BtbyfEl4yVUe5dzYhBIcCGJz
8udQdD2OV7474kYY7CMGfApqn0GWuMwFBaxViYIcSbMc266Wg2eFDT2hhBJD/jPh
HUMj0ZjqMGGvfHIIrTPKmcqS2OjZX8JSIVjukPPx0b+SZ/R1Jcu38LXySLUcmpo8
g5CqnGqUNwwXgCvKVDjpG28BZ2nPJB1aqlxKIc6XY8yLzi4Xbbf2DQqHtMgZxu9y
oldz73xxw/Rv1h8Ky/ThSFfufNA9N6VgejEZ7noEkdEyRYrpYtVTtJ/p1VMPcKIi
ZcyQ+Ci1KYhm4+d6l5In5IJL32suPqVHpmnd9oGZfBLyDGbn/3ktEsEvdOM10axn
iAFd0gYWreZDgTbsaOEbMjC5NuwHaKb4x8IQqAuplqsai4dlw3ZWbmPAHzqBpXZP
qGRRlb7aqIWlPbsLKB3eG20PpfxclGxFqZz4H1R2bjGcrhn9oG+Ycwmg7Gubjh43
r16lGvIqehaubs2fr6zgn0Mm/9HUPVcPcFwAEv60SGWxPnBmE8+WnGVBrjJ8gXKw
SnkbLWZFxErPec1KgLsBeIL487zxNF4VYtJDo8k5MORjzQ3Ic2Wga73srApsULHq
5B+MUApwID7wsWFVc53Jg9DqXZP5zf/y3fjaXWFBZXqeQQOdO/qdcFM+rUaU+v/A
fDdHOhGJ/SP8WyhhmcZQNHRR4tObbH+fSIWnzHJmuaQiavYQ6rqq3HjCPlGucEpY
JRj9OhX+u0hTcv8d//0xHF/URo+wqk2/2tiMazNNhA9n1kLVgiihpYKNwL6Uy7TK
F7Qn33J0hw2k4oTeojG6qntEsfbgPcg8qUSUiNeRIZn06Z5pcwcrkO/NPA1hjeNB
mKpmWk99kY4LrtBEY9b3/mAGFuAlJ8s9/MM2sqQpwqZAbtSB72NIxqFojJgGePve
ZdZKowdacm6HuA7WmzAHf3ujo1QVQAPI85bEZQbb3rY6gQEgo4h+AnaA4bMq5hKk
Tl/MyHsPWtA4MqDkAR/mpsKivYNGVE3uEBKoibk1r26tYMnlpEbzVRetauXDA+so
yfuxgkB7tQL1WiIwIF+rQZRufGC1crkhvtF4k5qIO1iDCfTuv8x/BPytvsnvpa7k
T7mdNQGu37qwvVrLQd5XUbnYH37e1baBzJ66ttmt625cfMLstIU8wzAVMyg/9Iwx
tGrRohjS9iLXAIusvFQUmKGU2h5Mv61l+DT+Qg2EmhArwKUWgplvSSqCKfkf2AMl
mcsh8QvvLIZXapxIXaQhnbpAK9x0e2WIU6RnVkGufm1hdgMVXGeYJd0NSiSU0wbU
bXty5GqO+6yVRznFLZVoIr0Hnrci2p6/who/5DvqodgGWEmQnmqv3p14sblNMDG4
NbMrFu4/KAkPEpFsJkic+bcbbMnd6ZicdPakw/Lx+MAq+Wak7iaxjTJmvjC9/1Sq
3tJ92kJXQEr1ev/J603G/2lOPmqaMM0Zdm5SfHx8yFY0dazLChSoa5wNl1RFhOJH
2uyKCJesAy/x8quLU7uHKZdoC55qyvu4R8l6RzgI7V1wa5K1Z7pHvbVr7yey+ag/
iABEDdPcpPj+frtQvAk059eG7gEw+OVyzsDkm3kIkhLr0zmf+ipmxBeAcJxuQ4/O
EU51IpVOlgHvDzLwu4IF87t702/rAPVfuCz1dHaqsY35YAGiwFvOqXTxsqpa+t5J
A6kGqBCXUgh28W/rk9GYBlHuBd7DxmCAUBm5p6rG5D/OJimnBMTc5l95mP2QjCxm
r5RkDscUftvDLzWQ/+4HO2mGtD54Ffl/Jg8vpP28khip2Gcgs1MzNVhHOcS8ELei
02Tzw9JIvTO69YyBroQwIINSM7q4lSPzczemOFrLMBbfS/35czzb+SxkHla71soE
qEAydkJ0UXIYQqg0hovcZP+EhbDYWV4Y2mYKZfYGJkoVOscXnWDdtGacPgmrJ4bq
sc9iDwk8s7emUadhWC0gdjL3uHeGB/HIpLbCmJZr007BklwDYicZP08C+gNhrdFM
5Ep8TtPV0BMF1no2uXRQxDvYE7PI7D+WU4WyrUVo+6Z2oU0BgmE9bEgjT/N6PuOW
YAAbltz07uQauOqGajM2pYCb/GBPpCQ29S1zlMfRuqn8OPe9DNqPxYOq87nlPfdp
I+qnt3gSmGj2BCeBqWoMI5i0Cefn3VZP52UU2ucsnbnfYLf7yjOSqGBzOvz/ftu4
bwrLSyeJcCZuWd3bY6uvKNYD8bTcRXIoBzFTHehzdeqxFToR/7klR0b4K4QlsFKc
2Q+Zs7RD93y24bj1n5mdmM1562ztGLmm0O1yhFifvo4oEF5RQdKtH6QEkBhk+MKe
fXRa6NnHRApY9xUtmmV5b+us0ECjwcIgTaECGKP0yp00W8sd+VA+GzjU1+DQ8Lta
UcF4hDa/fRjZmVqWEJBfHtjxAUQOCtZCRv5SSl3qrohXhR5GSMHvpOQMUo1XmrHD
DKaYI6R8OIYs6KFSlnBbZkUjfiAMDWUIJSSrJTK/r6cQxErAqtDGqeNWpJ11VpV1
6FUWOamJb1JpjnUTSEsqLWOzY1oJK2TK9HxrPhEE5jYcs/WGeTTajuGoh8noG8vr
pcfIzZBUo3KmJOm85rtgzp0A1e/G2Jgrv00RNWuNnPgXpYJxhiYLfzzzMOLSRF+M
/3nCxGpQ3iIMtaz+YUD1dCe5VLYWGcZ7I1Rw/kzKOtEEWD2Hd8DNsrtCsvIHmyyi
pWAOeHjEDFW2HjAuAdeppL1G3Kqu6ddGDo5gqfUU5dAHrloRDbV81tSOhqAviKWh
FHhXRGsTHIUnGywmG1POunuUXmEq1otKlDDY+Epvb+Ak6TLgdSWRrhj4Y0mJLzJJ
K9xjhG3w/TpP9xJs7bnPd50n4Nfu2uV+MbmGaG5qu9It4FZ8VmbDn3PAgW/Adwlk
wzJAW37PXEvgOf69vONBmCnxwHhmMyYmazSHfeds+o3My30mKQJT0tK5MHQwcHQ2
w1U6MaYe94HizhfDhmVGWywkFelCfsAF+D5W+MkUNzhG8yJ8Ax3urAgO0ia5kz0+
qnRM4ihjHfyu1bxMRbtZFbMkw/mAu8c1h2lYddiRos4oIGO3eojpyeSOT/0t9ROB
0osm9oE/jPqv8kmIhkL1l+JSFB3/pSXdqFRTn2s5uKULjMRnQpco/V+suT3YYwRW
piG5zFDDvHHAI6y5APSNZ7MfWZCiBJuakuB4Mg/JhJmHUFEhFL9phuHT7foKsEJX
fPQnZ7OyVNdH0W9/X7tup+mbLS+1AfEpEwEvzdqvAGfeXbAtHsjStcxU1BZfibpF
3ktQaw2WTF7tKI9cfx1ftarHlxML/D/hzPEBBd9L45jmif27ed1OnVH1FU6NfJ15
d8PjNGFNz2f5ttaqK/MK4cMQMaDWWar56cOyrg7Sg0XWP0HLX4OY8k0IZ5LaUIOz
PhuKH4hh+R27lpQacaHNVgOwa8M+SLo4HLQ1axBvlIkpslZJDNH0i7Aut+glVoNr
EZxOB0CwBpOrG5036IhhNu1Yw74irCsuvnmtQCy5Zxx432pxkSzduevwgqdiGsMr
gz8AjS3K/W8Xd5orGYfFs6yXKaqHcAe/KL4ROpwaBQtpzTqb7kPNn6M5yCFAQr3y
9Kpso+gdDcfLre+PVv3iSluziuw7/MyynwRUWRUpqBEDMYQS/8HfPprbFT8yjCfV
5Umi29TuVdl92OBz6Pd9j8rqnCbYLqpBmKURjzvLHsBPKqzytTBI43R1YlLZDHVE
qaFMXP7GKc7twNqNd8KsEfDuZ1b8rkCTczVmPogevUQ9WHxldujpVJkaKCSG6q5i
2nF87XyhCm9S9+M1D05VvgeQzptGqlkFEPgF7vSiuChwetrEzq1yi+3Jj4sbTwSe
DHPY60uF7GfLrpj0seeTQx8d8nvioBuhWjGp31uskXtT/n0Q0mI0xTtiwYbYzmDf
BToqnE6TH4Y8TrOj2vP5itcQJHGNKD0kglKg77byswgzSvu+I7JYaoDt6a/isD0u
4lgIcky55NOkfoXEpfCrIC7ah4BSy0RHD6GfvqqlXLxcsicK51FmpHxNQVAM0q/A
C783Ly1ZWJ9VXHuo3bGjf/vSQl77MjQ1GWtSowuZcJSY0T2EqQx0q9jc/mSv1zBt
aROqNcXc9UbYNG10mDaFM0VbRPpuhl9W8TJ4z+vezX4ZY8GHlQkA02xuTrTeE9Pi
GFlanJTEiaU5C3u4MeqRA/1y5qPY7PblzBXLaSgfjam+Xa4g1xKDsH+sQ6MXLOzP
iiUkfkn9g/o6amiksfEAMjFxs/wg8QTNV2rHtOIe1XVBlqIyLDVeJEjGypYeTUAl
opVTzDJC/znE9cu7lNqdn1W1I44MM9lB6DfMG6X75fdnprBKxvKEELdm73s37m8n
niUqpXjQGMuEdWVE0hRbhvJkq4xaOoPtKxzMjX3yJrD+y6C59PAS6SvYu4Azzzer
/U22JUwkM70mdO/8HTLjYsaDPcpYBzyt35a5wkTljFFcZyuaBixLZ/dESdzkAnAR
HLJzJISYIn93gzrjt69wSFXEkwS4DRPk52Fivgne2rJ4wzrcUu+7hOfnc8vtyzS8
LhktaNgeBI2k0FSfJcFuUwn6UzsZDj3Lg7NQe1iotZaIJjnnW+8z6bR4wzyZGHI+
r6PLnePCkNjYDK2U90TKN71UBAYU/mKCw6ovRhXy6TnmGVsp9zqIiqYAytg8/Bd7
4c/c6YDoYzCvFKZR0wJgxgYMNczswE68qfc3ysolktGQUEQZ5410I6WLZegF8lvn
So50xU+tAWbrb2KnIBvWgfJnEULSLFxFisrQGsJE5+w0MhRpRDDpIO2anmCQTNlE
ADCFpkR7Uv+osUzLuG70XR+kUVIOwd0vmPYasqjt0wBSG/V9XL16rBFqsOdyomyA
Sr+98ALe5SmXCDvaHjgdqii2MVuYct28QLbMZZ6rBWXLnwdNbAgLwj/wKLwNk8uC
PLNJxSbpcLwCQ2FRJWPezUam1Z+pGfPk+8FC4gMMDYtWq3GwP3AiAn98q7CwpcTv
KCUATAkBSKl8QgVoFkKdD/9U++jIrmZtQd9wRuMQmyg5yt2YQvP7rPa+n9xIWP2Q
I3BEJHji0lgIS8D8ZQqa5kyk92vpV1bZ1LZYvSEdtpf0dUlEyBMuOSJErwqYFQWh
LM5JyMqwpci1TnDcGygZ/d3gmb20yDNBMMroJSj++R+D50E7NfkcxPiHuzO8U26n
v5b9Ss2UFenHEy8Mg/N2nItZiCy351qegSeW0HzOPk++KXm1DZm/zhxrkCPvv++t
ZFTUQpdih+rny+mNIVm+qM+4kxWuRm7jUbCiqmgZU/U9NMtDQ0ONmz8AuB0XgPmv
XQApaojEtWC5oeZhciYGsiFVMY8E25CQvVXEk6srStbAZiesUGYFUtuZP9khQmnb
I5b9JUEX9AGJL7+X5YtijALGegHANvq9YqdU9D/QHXcohegQRTpeshW3Yhhkq8JR
KaZUlD/nUTI5McVfjPsVoxA2EsMujREVsPs0g/9V0kwsZx7CQC/6e5YdlLNEmSTU
Hp9V/udTJF+8vq6O/cLbnW7tplmkBKdH0t3NIfyJ3dK9m1sapc9rCV1PksdtGnUM
UDTKycLqmbpX8dgfPGoZnNCFYtqvHzDW5w0DNV1WyH986zoAV5lSkeOx3VQMKoKQ
nweD1/XH2+ZI7htOIIwDmd4e8PRukV9VBo9fzgLQv2EdSIQNYqjNS4yrNm6VZ7lX
INFcfWZXp4axVM5xJcv1Ic0OGYfiD3yM+p5TkZ/NGKmTd778ge2ITO/EDbup23jq
0hzkZTlTb0DUOJ8k3VdZ5DApc961k1x3L6N+G0nFX6HAaisx0ITONYBpj0hXYAbQ
PUvPFzpT9JePgq1ApHa8kB14JaTI/B22YdIVidW5sqeTbF47dXV6Fhj1SMNad9tw
pwmcUHopwahRJYnCs0IIQlyNS7EQ1c+DUJhidKjTRFcTAvcUg1NaetSvSBrk1gsA
mdFMUx8vl7IVnB73rcuRfoLGiz60Wg/NbNK2Iw7Ag9Q8WNIrl9hAvRY7hN1OGC8B
X4GoU5I6b5YbQ7rYiMS1BZNm1MtL64++lyRpjJMhs/cwbolT0UhSrZ2dLrmkZDz6
Yhk2pTWYXJCQTA1/j8FZ2XicDmdIsmHrIqS++PXitxjiiqe6+rGgxfb61bzxFCtA
jSW6+9OPTzuGBdAkd1Zej+WsS6heIbbeRsYuuXlcQfLcHysMlhJuQ5/iNRTsaeEn
sRXOsplIOJP++bq47HaVo2JeUU9E71KEkca7sm//7p/xvS2uG+kNvF+NVSq33tnl
hpN1UDik9vsrvzFJ3YgVe2tq8gkUhXd3rPdtRi68o3lLrrtEfUtmuuzcW8P7xqz3
J7kPyjwnL+5QjxMjpSNqun3Gf25WIq4zR/7AxBYv5EMBDV1R5Yu/+jSIT5f7RpGj
O6MGNRLM5wNzy1Ea85MStnmcSwXQQkhGucWYKkP/24Hr40dfnX+kMocYAcr/MT91
XuD/ASdFOBHQz9WoAesue3ua9BVQOCc3yH0Ksm3DaYU/vLnK1IqFQq3Sy+zfIzHy
34Ah1KMiw8GkuFr0VMEHTSgnTb4cNWPH2yjV7LcDw9TNRaNo4osRcsUcJJ93/9g1
jMf/Dv/SHL/pbOU93bGqf29RUOSx9BAlsFRun2zM83zVcVHyPxrpJiMg/FA0iF+M
WhYOIH/XpnEaQkUCcE7Izd5/dLvB1zWbhclT17MIGrNYcQ9Nd8VxVarRMImJEejq
G5oyThpWuBP7c9GUYNo+AE4LcrxRKnvSr0ozhdfeRtKwLFHQQKyhzKnLph/W7FK5
W01EO155Mm28ox7RjPO2/im5+tq5/daQh0Yd/rp3v6EEsqFUmE2k1Bc09nCZqNP7
lwbta4DIG8lC/bxt6FimTSfWVD6wM3edcZCKNOw4sG3C1i2qno+b3zkRp910D1NW
14BwMsZqohrW35hrKr8JSSPpAk30QJXSa4n1Hzn24Jb5P/tMovYqdtq4zHViYYc+
A66u/nTDDUrOt0n3u1xWBGX/C5Ho4be0RzqzTKu41GbD3XFd2AZXEKOvO0Hqp8+1
S8TubGvC9aMS84bB3bVI6ctkaE1SIAwpq7nkS7NLW7W4tHciQEdP0zaCxkMf23Lr
1jWuvjo8usWE/DaFUrRq99CPBEWadg6BVf9oM3rSoN/U26kjHNNv+0H1sWOpQfHN
9XxbUt/vu68JDMME9msoMGvaWdhJ2GxsELl+m5F9kSKS9M3pIftWlKCyVRBnK+fs
zianOf50K0omNqaBcbGynuYmEGympwc2kU/aUkc0Xal2xwVm8mG75HYTg3FbNQUX
SdcBGcDpDUGA+IRmBtYg6aXFAHyqNgln7T8dD8BrJfELMxpyz3rMXn1ePe3+vJpp
SgtrntK0aWoEd29D1l37AC7wM0+1tPJi56aenY0QT9pMLUsG839IrIx0j4TLGrE7
cRJ2ETsOzUn7ciqBVbGwWQt+9K/os2a/jsYqZytkt9eBAPnBT98h+sYmBjhFBfsH
mpfQDC+bpMoza+M0DsuVKE77Bxyp6RLRfgGKNtHjQJ0PJobxtIF3PMiGT8R1Y1IX
6vZLjrbIc8jwhDY9yn4wblE9FHU+WYVu3J2scZYBz44+QVpHFS5z6mQ1IxJf/Hr0
DwDkVQft+Q1x89tCgLKz8oTPFYsC8KfcMLSdU7YG+ZYzaYbTYNG1Gvj0mUMm3gFG
byJd7fGvDlDeO01Kq991uw1ugCy2UUK29VWftUAWPUteQI67JH0X8mTTjlVra7w8
D7xoSktw4h0Vkph/9kLJxDy/qxPMf3GQIVQi/eSn7GCz99bODKJy++pkrLf8XJtr
gJBgv18jQiSFUy/jyfRQ8wfcYxrP+UqAIpi38kRlz7NGcbzv0o9Zm+a8zS0fiUWO
jTit0LBCObEYwN0pvC/h9uuT8Rejy7QFH03EeHCNFoix4K1y5D0CoxlXAS8YGCDd
N4xAgzbGXg0Qk8taArhru6oKthExwqeoXxh9dt/uN0WnTNt7EWgyLRPPNhQhoKPZ
1FMy9OMiJ6Ipl1SxqrJvQcz5auIy9EIzkg+Vw2V6AtVhkc3vRKE0VxNY4qT9poK/
m+45YFQPxADCyOcH1XnEyONye9QeCIiRTGREcaMMTuJlCjeZUVLxhhEb0bf1Bt5x
of92ryJfNIFDkKBPwSGsQJc/wvS6LQkTdIb4f59OdO/fmrrxWmwaqhLwhD243MEW
1XcY8WYz2E5QxXyMQi+jSBfQE/B3XamCp8CN1wk7wTGZqShUGaVAvrDDsqVzCjel
UKQYrmwSujJb7KiE03h0qeohc6jXZoa4FPo9uASNDujpKzl6STxEMf3kdl+zz/ZE
YhkunYyMqMonJMwpPdnw6xPCp0kCQ7BLZ9pOuBNpD2CdEo07o8cyxIfDiq9/K6is
9m8n4zjrUEoaZ0cMRje/lnsoidXxn5jU2bLh94g01HmEzUvH8aK/THAH0ivc5wTq
be4MIUUva3g81GjnXe3nvfE7HI6bRNRiQtAp2ykSCFaOoW/IS14z31d00951NKK8
nPw40VdBO8nFQ9603yOxFjinKzzs6ovIl5t3EDkWHI29q0idRnvolFe3EWOkPMyS
y05sEHxP+YoPO6kmE98ZlgqoGFwqovoVeCwAoJGuwPry10Y3XJQ8n8Ae2kpH7pWL
5e9kbuZsI2XATg9EF461JRZgxwOhEfA943y/wv2uYL9CESVsyQxHU0l/LL7hblPC
vKuhjb1ybVjANJGOclkbgZZGjgMFsIqIdvnfDvWxUacaqNdBvJKUmtliGX5795aV
S//Brc7aJ6RBt9YnGgil8bbWsgCNs5XF6+pE6qxDSA76bXnT/W2FLa6gok3RDTRa
WgnjBBMltaXYYFbh9213G/uvwmg/fBKBEhomlwdxXIvN76G99a3sjVm2b2ll2318
M+hedKQt82U574M91eZpOEryO4dSuISy017XaYFH+psmkMP4QC7JgpqYX1BVKv40
FbWdXo9ieKDyU8EbKhCKUZYqxkiHsYnlnuEtqfgQpl8qvYA49A94zwOnjgWcoRgC
RRZVy1pi50JRH9s726TKH10Tu0DIQ6PM839JygrrNYsMETCnZ3ARu1R/5CqPO63O
Wv3jQUxRi3C0K61j2bMsKnixIumWS5CB2dwMsu8vuN7ePBRw893bTXnXQxA/pDbO
U/U7SSEastQUFtUf9Cj5LhoLFczKkMOJewHxSbAgU+AqHcLcJ8ONeTn5ted+ltse
qjLPDlnZ1lOAO4HXZTzgAem4U0KpYo5IGl/rEufJ/pCsQXyl1SRhaItzi1z0J+rM
c1ED1JhZH2dGJ/j+nsUPPhwH2/Uq+bC0bop8OIfuDDNulpbpduPwlNWI1zKiASgk
NSar8JtXy6pFpdS8aNQxwjStYq3W2gnp6JDcdqsjGG3sJXjdZ8s5AanQWXLMENpQ
woIdQ6yBzolFIQz4Zy5h47HN0/XHLoCqsJYUouJ+751KEKamO7xDroqrdkeVXAGf
QFnmhT93HrMHHZr8U8XcNGTMFtGWlDEpvkVW6n6HcS1pEC8HsgHciKcYJ1jMQ/Qs
3NwqawLmrZdATNevdf3FXziU5SMIV58CEP+H6+ubO9lPPQub/Oxv/jVkiGmt5O1K
5PlSDLD7eUCdfdMcf5LaQQTHuSj+dMJnjpo2LxBjiTpp6mikAKZHfiCRjsAYxxWI
DdcKpD5RYQvNNzOAfMPDPENpIX14KB1LWxNOLARn8nIBoZBHw05DXQE9PwfMC6AY
ekkLwcChML9EzAlR9/nIySz12/y1KQVYkVaHXF7CsvDU2hxR76IFuA0JPTDJ3jUO
rJsWOLc8C9nybCz7UKTvtupi/R1oaXud/oCEBmXiQtX0HpygJe7GHy4lwyPII8He
hSN/PCMgzJ/LzO0KibVk+wgYfESZnnKMCXf2VF+2h3eYBZIonUPa8LgNuWKCNHd0
9tf3ZNbryiqJDLEna81oYqYS5iutVAu0WdF/n1CVe878BZ8I70ah2YDFZX8o2Vvg
UsW4PWA4fp/2uylxrZdoou4xSNDu0l+U43QVEdxkdUXsPGE0uFp9N2S95Youzhuj
la6Ti8WF5ToPIhNbpXxqznqN6Q5ZdFYAI+ujYbPlZgsHiCulwWImjk9nTejt6Fx7
5NUrsrUJ9suAbG+qA0zH/6eNe5HaKKuuF4ulqMxtU4zgDktLpBuSeJwGsqoy4cMJ
EpYBUUy6DQF0YP8iRntBanJ+m5i6zY5KmS+/CUJvp2KLyBuxG2y0FfcbsCTm6xeC
svhpZ/xZfSDwonqK37jxtw/abULYxoTEFAiSG+zfXfUDmvz1THVSV13XHmQuWmOz
TGCVcVa3Eb+324VwKhgBHnstUxsIZrUKuvwO+prqwB+F/PqIVvXBwfV+RfCkg3Hw
0uXF0Kx2W+ORKmL6FDgHtAZBMpY1wqKeSvkjolyHC3NfhOdEOdOiOv540AOzMLo7
D1XMkVvPgAJArSEE385TSySaoCURH8BeAiLLGRUkybPM1qWUWU54jq4JsrA11S/i
pGrWerlNygDrA4VuFYH9QyAy4W+16Vs/MX1qbFRTx2NfFnuqSJFJZ5zQKv975bEk
HhtHpb+3S/TI2zp3tX47BAgxRFGZz5ys48vR2D96+41CS/w3j81dMitO6ydcICS0
TZZx4m1G5BsP3SuO/WlQM8WITB13F3ml544qfqwfdVCRALGbxnSkoIXnu49kNuFZ
f6/bwA3+1y9MwaVOJj6LpEUYxaww+Uu6dEyH0mmsFDe4Rrn9gNLljpm8ho3563r9
NzY5GxiPcRR2QNJAeFDBmqHrNZ3s6lENJU4xb/L1TxckIsOnL+6dKvv4LSLoGA5n
eUNxbL4NbrbA9/HRI/pOqawjp6OiYmzQC999yBxxcAaUO54zc3aSz8jd/5wQ8d5B
eSVb2iVKEJ1TWMjdIfoc6rLNPHta+UPQIVPQZ6KPqSp5bSyz7kpYCs71GmC78/34
cDrFYr9jNX8X5wUQVQlYAxjJuqHoPZKaguiA/vGSD3izaY/QPIB3niVafvHlLOqi
UNZyrj56BxACmugbMgpaeFqUFlrLJT33rn+RCPaD4bNhU2HOkqV2WrIRVPmdNLgU
A+eEgCS5o1tLNzKuLhcgxYTvM4GbiVjFpp9arG64BXA6F8nIg+mv8hRe3oGlVTz8
qonifnRuM2SXNLk6zZEAizVTdKTTJSvLfZOYCudKRItdYteaLVM1lAq0EjI3H4aI
PCN87R8nG2oYKkJipPP1iFGnF01+wBPPOqF3oK7/KrCSFTnNfRpEmjNxtYoiew3e
1grlKH4ZZrs8mRaP3AUyDIfxWHkb3TQO/FjBSD2i0rOxg+WRNv/vjsK4Rdtlu08z
oTtp3644SA6YOH3dm2FAkQNBTyU1SFi2Mr16Qk9ElW8W0KxhMjifOgAEG4Jg1mR5
jdDNb51J+6tdOzJKpMJl/d+QPHk5ynVPyvfUwDwgUp511cP/+jTu1PXAMGnZv6Uq
jEVxSXdovh+hnvV5Du0XOsBvq9nmBp9I5kT4qO2HvQUpjBarTzP7pzMNSc+IfIoO
jOSZhmw2i1rYicTueS54AnOd0dRlY+cAGdcgliUPplLLAiA8eJkoJJjrjjd3qwkk
SOFf8T+2yVklYpEqrenm4dQpDnPEogMrPM8ao3/ImXnMpL1RvesIfu0eWlXU6Epq
NvNAL6XVWbtJv4zhke65d65hG1NOLa6CAntzOxVjovYpKsN1e96z9MZhGuFOvkz4
cH315wJuoYlx522gee3LSpR9vcew18C/0RPm4TO2n+VtDY6JH/aumVqfXrI30yAM
JySpihiFseHaoOnZgRgSkU2CGISsE9exsjiADqDvKiAdUGiYN9trhbw/viFhjuXA
WDSua4xrg56X1J/R/htqesQKLGhMXoPaBINA6I9PmNoaIGIvD3aOuqUen3ayN5kZ
P8XK7RpEdyF7TfJ5+gAnvt2CynCjWoWc7B7wyyWA/Fcrawc1rhFp8vxhEjAgP4qI
Tc8Kt/jilX01SeDS6RcJ9T4DWdEfMrQiyjlaGUz9Z0roIo7qEJhonmyx5ZIXH6qw
6HELN58ZcCfTI6GWMclf8rqpPpSAcUwKvwWzTogKD3Bvc+DjZ3o+dbilmimGPdOm
2QvCkG21dw8FtjR/X7Km56TknHqakbiLizZT8s8OONRfqhIPf1uJZZdyRGweVsA7
88dXERpM+6VRFjeOoVsAtYkZyw5Fsx9NM5fPlpYPeTj7GQeU15P/Xq91puFkti3F
tSlKYVktCpA6c/lmsnXDYa7azFK7oQ2YRKB40WM15m3x+NXFhqieO5tDgUQHiRGl
4gZV/dWxWXVS1JfxjkP5fKP3o7MtnSJUaVuy/OcSa1TF21y3P6z72AcDOTMg+Yik
t+kmzGBTAxzGReZoCeHR2uk33sT9+jssN4UUIAK/wEngYVmlKvUUH57YhR08MpDW
Ti+gFWxZ4K4Mc/56FrvJdfuk7VCYTHTAvgNcFOk/7FtBU2LcMTU41LocoVcND7FA
4jObX8ZdVFg/0niTf68Op78jbCs8ER92A50RrAGzmpo8irS8kDORyiIdW215+M/t
LEAm8oBmfwzDumNAidKy3kzPAH6FoyDChK1kRUchZQ1W9o/ChkPp/rntaI3Znr96
Gdo9wREqY7ag6lTmgRY9CBmZQsK6+Op5Pp6HjJz7XR/jDPIKcDh4RARSXYpQ6KBa
CHLxNnpp0MkN+lqWpzWf+L/LRewkyfatFddU58kKBqkmHMEi7E7+MOMrpSuA046s
1uGVjFbaLed6XZE5iKrXYw0bCIArISktHWXUfi21OCgfEx0mhgVV3Ts6mu27ur4j
NC9Aa9qbD+PrzBSTysDOgybKoceRQ/kdlMQIe/xsM3Ek8TCfOmNUpRcKx/1V19pD
Q6TkU5Oz0G4GIjGGlybkyUZf8+TR5/G1uOLIUi3Tfdi6EY35ilSM/XdPHFMF8nrp
5Ub7TPUmeKVfDCFGcALQacEAGWVjqVfQY01ykRIp8y/bysfMHEvEiaU5Pa8GJv1m
15b58k5bWlBgsiR0YkoHtfQap3fFHBXZyD+/CYDS5Gdi+dKHz079PASMhvmY9Rn0
k6s/G+L1YXw3w5Ya09hAxw0tXBq7Lf3L+jNGyvIjrv2YVnROu1yAWnw7m3+/JGw9
U+lXmkKCgRMjgDbCG+CZA1ueIilfPAnNy1Ttpf90YjidS/ziFHey8xiA+Bklz2bb
kX9BeORPGt4jvh+PjS1t6ZjvGDG7EecrcqrWLeFOZlcYFbZAAy8u+oqTlDpZgB0k
GBT7RhGterJHcn1tPZxMFSNlZN2B+JhtROnNDtU//ZG7fZwLFK2a0cH6EWDs3qKN
uO8PmRzNRSuNPrmKgZ4NmilA2hLv4RItV52NOWA4kjoIk4agMzi+wme0KwGsY0DJ
YR0NMAY3lXhEiMd7kYRXhbL/sZi3KCCGELQ5XOjuhPOxr5RfoN2iWI7HU3HcmTtH
I9uS+oDzDvtUhOJZvu1dm35NyrZ0OvjhYJnNgPxVUCCnfIhrna1Zpf4Lo3jvdp+U
9SxDcj6I//57N0hXwO5Z5zTxVdmbnBtLuBHiEXt4Lqx0ZNIhCjMOe/jbjiRHFSMG
YHB2Loq4FR60LZJy0qOCv/CM/YQW5UZn3+L8PHrUDC7q9w8uGVl283VeJ8vgjH8+
EIsqtrHGsfjfaW+EIQIPjs0JTENYwJKu+sqfyCU4aSZ5x5EyKDdnb1NDrQbtBq7X
wPbCC5YLTgIXmenUzYOFzd3PVkGP8FE79BTobMKetDVgSS8jELrLVdv9fIRtzfWe
3s4Kfn9DENGwfx83iI4+NEf+Aup0GaGdruhHxtWuVgoMe0YVNxFyxkAiY8sikMU4
7Gv5VToXJyDCjLtwVAmd5C37IrWFzQQy8nIt8YKizYQpRc3OCrR+7C09PFx4KlmU
ZZerKoHc5uq/ctQKcXpGpFrnk8OvntmUnxFF7L9TTtBNHbqgypYsPZroWjVSjSuA
UmcSCN1WHye3XjRlKWTtfOfM9Vc7cgzHqv2wCfLCe8U6Oujm1htola6wcpGvS3Mn
aGwKG5wndix0nW4HRWxODb/Y/YOUypWY0BnytVHfW897S3krcUkGpUpRqKeCqy0e
4jgHuCV51vBzOZW3DSjL5XJmJyLicPXncdJyLRArvayqATm0LCSiNdHJ7hAbJgcx
/EKdsbvgO6JLZ/JCJgGPKbSbeqJf4vHOZWrI/2y2zJkL6mLTCzcPHh0nsY0oj063
5QBzIHM1eNsgbe5FujZfcGiiMx4dtAG62uzG7rLMnxEuPbVrS6/6OqqvCAhsmiLw
7wH3tPxR5wGzJK8jr9Ua7Fv9ALESzFUh+aa+t7C6zRN80U+Ks8ATd9ZN/JwB/wII
HJPkOfjKZVJRp2OVq+8iYM7MoJhBT2aFlTTY4q4P9esy8DYc+w5viftRzbz07Hyu
2kzhn1qGa3eG+IJFMK/d1HqGM+/oC0EB5GLIzkhGtpY/2SNwkz5C9bK023+G7xag
PEK0F2xd6StEJOWFG93pdQstH/WTlBMOHM7JEUCKOEgmOf6A63efmyQ5/HuOI4xm
2H1B+k+xY3bVVd5F+p4B49Hh8z+1fD7+3nOylaEDwGRGBMHhd6U7fXjjdXIUxbAF
SKuyQtaoCibtepzoom14rDv/jLqrQOYpz1pn+ZIq0P3zfkneXsayVBUyhAzNnVnA
jDaabQ6iy/Vwntot214EIwtGp90m+tNfXcfuyuzOvNi9lt0g8pO8VsM+F8Y/Efic
HTuhGYM/RtCi8uoIC48fJKd/VptSghdRIR64MsEJ8q+k0DRkaPaonabpQ1yuFKYL
vCOnS7oHp8ff9Un52hYOOcTUl4ndE/9Qxsc6hROKpBQK1/yjBUhvi8J38Ms6h2U0
UigYWHUiDDaHj1sJa+nmEBnONrV0r0ngfRnfdwOVyE2LKHNF3eFbXglSfAekr885
gtRS2rAl0lRLWJwd7Lcsvtfr14jfRLA2xn0PfPLsuwEVztY4lt7/KvjTtX7K5Lww
h22OeqCWtfvNC3NehzCL0I0bZGmV2s3JQplJLWKtbguYq3OS3DnsK/n8KSgIaf1n
aKDT5K4LyblfZtnn81MQ8O0//AN5lgA5vKBsqV9TRD+7YuXDn+R75PaBas43gJ9D
0j9rjTDDnkPOeQ1R1c3M2egBoP1opGJzTkm2VtbYt8iRcaqAZ3Z2HTeOvIDXUxRo
NWOZgUhWtLw0BfTOEounHfQDx+esrEQqQl2S+rPbTG6CY0EMfDuvIFDofPS3bvBA
imBf0rw2hifOODAcV+KT36NR7sbPioAvtsZYtUonk5Yf0LvwaTwQ55kvBv7cK+9x
+XMMrcVPiUOBBeG8gF1Xe1gtyAFrKTeYes7V3x+4Z6ISOpRmBopMVklQ+diWTnYM
JilZ5AJcLY5EoiAyAosKmS+el2r5I8Lt/vkl+6qjYyBSMT3m9BibjpvOiR7Qz+4E
Hdjgn70VWuXWuT0ZPSvDgBRqO6jhxv+zN3NJxdJhnlpXfXWw1xuaGRkD/4BU2nDV
W7HEbTGwvjSxvzjjqA3lIQXNO6tep0AH20SeoP2QEhvcQYUl75TIFjEuJ3Ii6MRG
pu5P67Ns8UKKwnX9IotpKcrH2C2suUAL6g1azO9GgmWyfkijz8jdbiPK3XW0Uz3n
NLWSnKh2etdvAkCvqEAv+kcFNa6i7tzH7alDiXEGQ1la//J6HgX343IU1xVaKTdi
DUSkHS29WUU/ByKq7F3aGxJ7WKmjeZO9GjfBT4HB6hVReHf10nmt+qBXqfDe1mFz
rJHEN3UL2EMbshntzEAqbFDid0G2YF1hQ+L+4lT0WA+oJ8nB6gXwrX9DuSVU13wj
PWF8Jsa8mo3XVO1XNwfnGQWDKBzwknSOsUcH+CzX57/lyNytKXF+Vv+H8r+YFWGv
83AOvDx5IDyAwjyGqppUBK+WfW03bv0W6Ex+Z/NJzxp5FTOZCgUPe+TwWjs5xlnQ
xcTTPHv4nJZceXadRwbNVsV8c9rZlZaWEy1XYp3xJ8mu+BZ7v3NqengYNbq1M1oT
4Xtt5okakCdq5ZDrKLEUuIMEuLwrJoniqUUStEV5OzYHdyni1qSv3GIi+c1oQKy7
P0LenOu2jo+zjDF1jBDT5gDVTnj/Khpk4FmUbP/RI1iGubD9IxPISK9m8aihHTl6
eVGIr7ek70MJFBmMFVHDK4Evh2nFlKgUETpWSJg1HJfTjJbdVu/jsU2u7xhRWYIN
0BMx0RcrRPwKv+GXRzsWVB8Z4oVxALu16RhTZulbnI/y/jJl5WON8Mb6Fb1E56wX
ngnquwCNiKmb7eRNN2Ibk2vShOH8p2uBMGvjSuYXgJjy90GpwRtZbRv6t0JXHgop
QSsaipQIXheYsY5ykBxVdJxNN+lin9Kh2CVWeelrOrt1eg27JFGPm01qnowG6V4q
azHOYZAAM1bSEGQlZFjpCf1PGARkSuBt/BQEcmnXkNLR0M/y0Dv2/CyN9ZSTbKTC
eGU1HfrmhwZkVUBysCcJX6a4tr3imioGEIQxoJReXuo+wqTFhdWa7Il7pGNnQN72
sHZ3j/L0vcWIa+NQ7urnNVcNylUF6xYQp04HYuJ/3eCRi/W11uwXGcd3wynSZ01X
t7vgwE+S0RM8vcTrEpmShhZi4QfN7P4MXsJT9rYd08xRIya5QkvyJZ6xifFSwTEf
NLGp843/kut/qAwg77Hsmb6Wb4qvIH9IKNwvdy4+9dk8BBeWNbUNOtTTwdGHC6IA
jZ9rm3PoCHOZG/yt6IzQi0ui6SUDKfhftme6gIX6V+0b8okJcnbCXlXpQWaoiGAo
JdFCAn0AkMhjVS8vrEWK/o29tY5aH8wlvC+je9m8qHKg89L/i4gGVhHMqKhG5UWy
I5yseS6aIIpJrUC5Ptd2o+s1pah2xt+wdS/sAPmoT2s=
//pragma protect end_data_block
//pragma protect digest_block
XLZLx8c8odTgUCtpdDAzW7ShvFQ=
//pragma protect end_digest_block
//pragma protect end_protected
