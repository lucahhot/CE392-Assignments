// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
wbHsaXHQAofmu6HTxJlKO7jyJkw7A5DQ4FxI7ds18j5qeFezvJVqNIbDavCWTNHq
63kxNuvfp7xDRewGMqkp2wjjLxiy7GHtdPImeZu9MGswl/CLUj1QvnPIdv/nHp01
ZjYa0P/tQIJT2NizK4dymHZiKuzF2iaR5ag7jydKS7+1oMhLplHPjg==
//pragma protect end_key_block
//pragma protect digest_block
QQh7QV0OQViCiUVq405a/1aWszM=
//pragma protect end_digest_block
//pragma protect data_block
yFon4mubt3zz5XdNZAz+vmM+PBKZbZDdwdDSTe1VMjpt/nk3aknt5M4gTvI84CBk
3GsR+qzNrilxbw1Eh+IAIjZNqexT/1rgYJgS2TyY8vTAHttQiu7u5uPjLZio+2Tz
doQz0JvXzmH0QFrHHlrib4ycOUIcSOSqdJdSfw7+pHxDxVZToUVCnLZvQN9EDker
1qgXtzMsnSp97wRLeWKdFdM2oUJmdS59DAcDsHB9jPrlQfSMSw2jwbSpJwr1+XMF
tvUeBwWX39WWoy6hiSRRTXUyBhgmTnnrDgb3ISMRLTsK1cgE1A/niL5M+42Z6NeC
Zw3n1PtNKbhvIlAgnwXty5Fa+Mky7uzNX62JU0EJXJGi8MH1omD1Ug6bJBEfHeNr
ZArHCuuJEDPV8UCTwMFgdk+kP5JXkivqa027JJXF5pKZkGImwzsAVh87K5dSZAeg
R9+EqjrHuewocs/20/EjHahp+FbZG4V427M9wHi2BsEZIb+MPF6yrh+y1ms7kIkk
sqU6dm5QZXcmA67ZhIjLCK3UPs8mapITHeNJgom1IQzbLHe4f0b/pNs/M4RbkvLz
/JXKxEcpjNNPBuOPOV+emImNWVmvX7Zf/ZlFJz69JLWFv20m1lS0nUCoiQ5xUokL
mTjaluhXQjh0jzd4BuVIBtOWZJJv3MjZB+L5Vdu0Ky/9DWJTInLPaQ6o9bDzZsVF
qNJ2CSRrBzkTQdl/oWGxQioIWxiIFGM1eSVQuNoC6lvcBzNB1lQbsLnXYcIj4d1d
OWTDNPOtkfykTu2Z3iuFKLCUH/qc04zlNRYQLzjxvCqmJdxz2z0Pd4XQQUZKzaPZ
Bb9qbQgnzgZO/vjYnUpVOJdqe1qDndqyec2PGP89eaR+ufS/+uOwOncXmPaarJ4a
ygo3h4mqqVxLHUALCSY7CWjcxBWwaElcBg2KPbHV7IM0k9NZJAd9cDLZNbW6FDki
OJC6noNgmdNUIw21Jx6iATCyH1oSJ9VW+Vl83Bs+6y7VOhzv/0Z9PMLvQre84jXh
prDUtDMBtunZv3lP7xZPFvdAD4XLIKPpWCdQ49Cpn4dmJfZidNaczH9xIj3F4fAi
w4pDece3amKSwCViCpyzFRtLpbqpaYNcfXu4sc3SA++LiosqpXzf2+jd7DNadp7y
d9tFfvbw2ni3uA3zPl8M0MMfF4XVZXEaAf8HoTMN4GwmBc094XndweDGHQia2s0s
7C1wQ/2HL/bbuVQAKjONWPE2GD+jdogeFZ55ddRjTnnjL0R1QT+XDjIKTV1Kal9t
U9ehSIldtRnMPR0Ynb0o6P4Rt+5vttc6KIZS+U7vys3rZLvZLw/soO4PDlHa+gSO
WnzjY1OWdNwIsKSWJfPltpdHYMEP+b+0r/IGs41vpWGISxWHy8AhP/FVCLdTxnO2
jnmjyK/xhgPgIY3aM55GDc6YomO6t8Llx+P2nTnzY3FNKCXCppZ4LvxYEK+V3L8l
XvAmX0H/7GEUr/aa3x8ctqrHxj0R5nbcJ6shX6JLYq7rIUFpKWpgiGMR+lG65pTT
Q6clWBCsu8hC7G1OWfys9kIVNHy+WxnliKVEz4JAeKY4t4OwU1TLpPXH8xwaz1FV
1/TBm+eCpHHk9GOPUHa8MbWJZOLGG+P//RA5FKopAwutbWaPsQa9YPMRaEiTnUWH
WG9XLpwOk71vb8yxY5vkddrJXSWTzXfp26KtlxFsGeDYo4xNTlj92Dnl4J7RXR0e
Mlescm/hbkaISVPRCvsRIfkJFmLuKBVG/UaQGyoNsVvar+5MjuIkQ+vXgp4FR0wr
VAJThxG6xuhjtYcaBq5E18aqELvmaTKFgp0TL1m/O+4bCZyO055p4whD1yvUjYRu
xOzw04NHs0H2fovMlSH2OZzHKPqLwxOqBWJfJiXJJMmymHUFTFfaLMLNg1J8NoVR
2TBOREBSBVRfh+vT8s5vhmXDWGUTpHprVAUEwJtwMlP7fa9QLPea6WjVZuONcos8
X1dzDuPbDRVssh1/ByUwbGJvQ3DVu/elvQoBxqZFIMHDoTC2YfJMdu/jnWhAs43x
1Crp0Y5CkheYQDECXEiezr1FYQxEGD1CgUp/K1a2AeXOZu8wxXvZY60kiw0D8/qr
57GaGcqAye4yKzt2mLJFJRVOKhHGx67mupKgEYpLx6GQuMcUNW/2KudypesqG8vZ
xZONbPweiNNNh6Q1/ntpvKlO77wZQXDNjClRCBa8pmrnU5TmCaqi9xZJPgMTDo9R
l/4N66OkTdMeuM0IY8HL411zlvwPivFuesEWMDOy2mDDJPEgwHbi54iAbeVma2G/
bydEJKuxLEZ21+G590T0GrzIZgmmb1dgq8qn8d8iEFMAkQRrLreNUMAR2jBFPOx8
60tUK1d6cdHL0rEz7T5bexWnsF0f7Hsz+9a3xyeJvyQxIZIpdg2pcKulC1Ru4Oik
M8e474HURMku5hB/k/HqX6LoD/zzasveZ9dyC+L4hJIdH8JpIEDpTmTYPsmmxYKL
DxoE1akPgfC3n5Q0fArGGD6AL/djBb0fIIIhVHzyWMAllfoBIhpoex0WLdrLhDLS
15oBECOR9/7QK0jn4O4FzmXBENfziEgK+rWv8aYZ+WrrQSLSvkuGXl5vP5bR8QgG
Qs7iEWQ5ZYidotUMdv8f0R9KDtdRVv6/QGxWq9s6pgyZBzrZeDsyT5nZQhd2BaYb
yjDbV+k0WhiWOEELjQW9b+DL5tNFVq6oWr42YZex6TXcZ3+aALf4fIfzcTdOJmiI
BQ0WpBEbGy2aA1lQLWoJpu5OfvnhxUtqXi9Y680hi5RGxhwQd8pO6IrYOuCoQKsT
3dLiRVJdyJiSMfuF2HMWsJfx7QKA4s50KD8zkynQpnqSRvJKP/YK038ATZUvEecG
MItaKguVwXY9pIsSPpAbtVHxRt9ZGeI/YfhOs8boCq9FHnQLgayvvIfW4scl02YB
z8qbt0XIPYaVpLMq7McpV/xC5AbYg3nnFuhmG+KZJiMcODciOzbCC4ryeiOYG8NL
1J0A2JxKqJ9SDnK2wMPUnSXoveB9NQ+gxqxH+b8i+tnDnTPi+nQ4+qaqXgWjlkg3
bLDel3oT30uI2zI3H2hjFwF8Z3DwOw+tJAuykVkckTxxJYMBRvmbxToEF5BIV0fg
ekmjdwO8TRCKPFIK7t8A/IL/Vo0+6F7Xr3RSj2w0KyakgGTd+bWPs2G/5lDltkq2
Hy692wnCG5GZju3WVO+WQWD/b69+LIZWtX03pWAxWRCavI2MZPZw9wtKxC2IGWKo
hqXTpetAxVsLZKgEdVw5dm+gF6M7+orcRzhjG3J7WRx33rjSqLNMgb8Qt+gV64co
QC3vXcqmyBvyeNwXU7DyOVdrxEZpxv7dL4vVZvnjODdO3kWDq3bn1pOC/47Vpbai
3Oi4eg7n53kg/o608lAVS6JaErkru1vintGceXzpdr9D9+sHs00WsFRygC+O7Trt
CPn2K9tcv2/rkvQAEbvO76PV17GStTy2qi8V3mu6epw8rRzVwCY62Ka92TQpalP0
3MrWjq+aa0FzI6J4t04A8aMA47aUTcDjsu7xYrr3dEu83cqLfCo3kT8HDs3mFSl/
Wd7wTZ/F2ILcS2/mnBkkK8GKqkdtnZsEdD7kPdcyxYPMPwPBEJJdN0k2krn7v30D
hhnB8RgRlxWPv5CwlEkAa8igJsm16U38ouYT6tEZXP0JhTbmXCkwWHEzY2h5Zi+j
G5II5RnbB5lZAyiAMlqBWsMyxSY+19UQhoTdtY0YxnaC6+FqGJIF8SbAVARFeWH2
npPsZH/TesK3oCTqUGWKA0FRMlBy3+ROCR4i37pjatT1U59KwKiDZw0lj0Bc1J+N
ycxyBy3aY1TGQ3adPaEyAzJxIEgfpT9ZkVGarzp7o9/2TfgpM2Jo9TCaJ0MIwqk5
PQHp8OJMqyW788AQAmIr4P5luFHvRTkx3yImnfaRFKYDIHrQGJwQ5d/+gay8YWyY
QsqZ/6XEUXBlYJV51jOF5OWzI/g1Q3nNLFg91w8F7MTCWLbXhYjYuBHnsFYHn9Gq
+oLXhpAUVV80SfFpd74C3o60IKCHZHsDX0bbKtoEOw1MCuJDz4lLRrmuO6Di8slo
WRmWsbaIr5423tuvCZrjq2oUCoWdyi4seOsibtj5+SDTQNtNqotmGNFJUw0qOhfU
bGa8QZbyb36zZZK1Z1LU33XO+PHUDZ8tKJ7qxFtNBYNp4K2jrwjBVV1rtJN8oAzd
2INBbhizZHybjjCH2MelanJNKNrL9f+xXDRrI2fRPviutPo6BK3Zv5tf9HL3Tw/S
GYZuGT3KrfSw/3NKyu9KylLDbYpIuuFWAEUZh7f3ryBZ2SPhfkw7O0p1KM4wc0wx
KWngjEpdtB51Pghm68+4OAzZftZix/Vbuvz+BRfIBO4J91DEVVcgKIf8U2Avri/a
r5xl9zAKh1m19oBXOL0rpSzRED9InVixr+dN21JbSWFWTv3HZHie43IsW/tzx1cR
lLkxl/i1s37PPXyNlzPte1Fj2Q0XjXJXlIllCVCb8rwXsx9+9EHSlNJPqi78UxNk
a+kxDXFLdVWdNm8HQV6C5kDOnXVjdVnjBJT/Lsm8naLAnKleABeMbOnlyZjTudLe
tjO8movsIlFHliUAdRrudkzsVlrxZ3MsK/FfVM0uj6CxEKM2JS3F8qp5Grg8ck7Y
/4za2P8A7pSj70kyOqG/OfwBKfd0NjsgQgoHlrMksTagJgKEWvEWJXdehw+7bdRY
Ev1AkMhTyjrPKsNbDmL9TV/mWK7iblDiR1qHmh97Sj7jiJydUTq1NTonFxvN1n9D
orsaYHPqdLpWiKsqivPny6NlCSjDdSZYw9YUD+fEplcy+cTo59rV5MjE+5HP33Xj
PDVaOhszftZhQ8RkIUGlLWybdPmYOc1P+eYXphlKM9lvd8xoPzPdPkt5dEfw/OrI
8DJpzVSmOOfNHta2Ncr7HDyexPYczszgzdJA6ChFejpmUsgKiQSceW/tIQSx5vtB
bRXJxI/0pNYTsqXyDnZvh/Gs+Ze1dLmBYv+9ZgKpkeQ2bNmZa86xVfRafrr2SCyv
kcdBw6i74IRx055Ax4nwgP6HXgPT+3Adh4d/IA5HWEGL4ly+hFauVvbJ7QldGXtl
U39JVoigBhxS58fpiLnbDEYGoxK+xwDVkWDRS2leNUUNyWhXxxcdmw2jRC6MfAhK
PCScE8whfqusjdArQ/YQWdM5ILdBgVlAboC0fRjYdquWAj21WaTwwrGAFSgTplRq
WS5snVU3PiR49/8z3zPjqw9kTvrmel47N8Iprgn6Rs6N0HUwIqj3diUOWt2Q5eT1
nTBf1rjFo/2wDBL6w5gWmsWry4l5y906nqn+bd80baYWbm9pIBcBV0IvJk3mDcai
e7pX9DmxxknHWz3P4p0X+7pTLVC1hEZWLPhhlAOIu6AIut7AqGbcImkeATh3Z2u3
IAMWRO4V+haIZPpns+cu1dlSyAr4f5e1PGYnipxzpv03B/OeY3FFBnCqKa9kN7Ic
TbBLOcnEmtZ1jKCEgBTXXhUf2sEZjZGscCg1Koz0Wo20Z/mT2FQ17oyFEfRcSGQr
/I/VGkVg8kLA6B/GizhbJk7BLEf9t2c98a8DZObF2Tw/cSU8zwj4pCs65VOdjgaD
Cy+ZGcM+2otcZkASTuEUyz/DGAVwlW9QYRqUsmy5VOPpBMuVD046XJt3zFIKMuLY
ic6Irmc+756KKRjY50gj8jMo1joeZGJOX7cV6hEy9rIfceMRO71VW4ut5RRu+tyx
93X7acV3szMQo+y/dKNQOn1GicrerfEHjZ0VXp6KRnEeWFMFPAjWXaeDvg/9m5oS
Z7UeCWI2tZsTI7iF40QebAyIARunwgEOEx0KejfGnlxhJEHNKCemkOSIBVxORBh7
2l4/8jTHS2/rdsAtW0/KEH5B7o3NmPluY283jpj/wPh/9s15K3l41gCK/5vkpjM4
XAwna9lsi135VUwrLiiZEukuej5hjMNTYrM+BsAwag/cYsEEx3wbA9v5CRSz8+A1
toutka4dLKE0PJfkkKUVACWpbFMJxCFUMTlwYaGBCXLM5gmNIgpuwTKXojTJtogj
XHY2XvPUSKeB9ouToYcPVblj5Ka0k+80AJ+N3yPqr/5Rx1rn1MpTXtNK9jleg3U7
5MdO/lF7Jtt6rkZ/W4qpmrQoQOtcvldGuQX4rF9IsG6KzJt912IZOqWWzThmmmF1
iiFn4wmtsCyPe/Ij5u8XsFXhnxPa3eGXiHymriZP1Ac3xdc9wSEtNXUkE5DUx8t0
gXyNGtQFaZljXp8u01eNiWVT94/a8mzOGmACqA6Su4Ho64Utt8nhqxWsm1jwz1qr
Jw0/8SnOmAm/AcuZVTYbJun+BxWNVQgFjIEnC7czKI3cI3WxKGQdZdO2+zrBTbgs
bDMo+9hIpw5b4L/4OIXs435M3Zf6nqClEVVw9ucbvsuFw+oVrtQpFACXKZVgo8vH
CwBSF4WniWknZVifLysI1qxnLWzJZGOK2OoWRTx1aVb0eMT2SNkNoqpXTpqxh7Ei
RdDFPA5kJFn4AWw6CllzI6Fb92T2A+56PQmp6fIvsuqACPy8NbNPlX8AcXAKsAwX
NgVM3M4+XUiMRyLxN1chSklfZsR/uWA2Y9rFCrIY1ngPxhEWuWzVWiSZ5w2Gbk4A
WTVqe6V2opl1el1H/pHT3xfYoQ0YvUPRiKLxd9nOTXtXHCupCi/0sJdSmNWqvUEm
WSYBChOVCrZqJ8W/Kru0EGriQiM8YWLCGFQhbxxVMukZS3TL3C1wbp1Z7n/Ku5v4
zf60ZfCEO95c5azi58s+c0j/6esrwhjdZhSBgS6OC5zvtm4P2A0ZI91en/NHKg4j
SMzRVD8Yd8r592POh4dJgFkVKtS5uLIMXqthULfUBVZjNzLLRHBsNI0ZzT4B5cQh
DQAm/i510UyY0eA6e6FquO0IG7n7VJPByb9lD3AYmY0EpFgF5iyQNWGE16OL1XKe
eB4IjK0QTYQperERhQdambNNkNFhjesmC7nCm2hbn0Jqg+j2UY/WxKDPy0QCbRwC
0VRBHbb+6zPoI+btgmIBJi86ujw+VM8ZbLAmObDQlOGwuelFfW+wasPR6ul4kvsJ
2NLdp8uGtX90XUVzIHZ/6r9ulsc1GPRm6OrBl69aur70wkWuV3yvoxOjKqEteFZx
4wpzwGXUclkxvC5DhtYv16j9iJrFeNDoowJhZFQCXbLwH1VgdrFUQQwB1PYiPgCa
9MF2k51dZwh6j9MKS0KYX3GzVAHSt/kdl184LXIC9n5RooVt5IHfgWFeo/+FDvp8
d8q3MCEklvBpcbIuWINosJcEmQHB1ElkXKYXUBBI8h4wfr4PEJtwbs8q57djrIua
FUXXbWz3cWV6kT8zwjT0PQEX/11kdckHngc4VtdZT7+DJNgyGbHjG0q7puGjj5r/
QMxztVCDc1hPSkXZo9Tt3j7atXijxZv1TNYOO1KS91S5SXnYS0S54AtVGz01zluy
l9D7lkqZ+tLd/rTKkSJA6eiR1HBfa9JUw8zKrEjiGf2qQlPshs9L3a/Al7g6IXLj
AWMNQuculLZylrcNiz97IPi72At6gX7IqV9UWH6ZkG/IT2aO93a+sL4dqcS6Uxoa
PpZbR3PzN2vYFfzqDgz6dp6G4Ntx7gZU4Fszu2Qgs6nFgnk1VNPIT+CgZQwsanUX
eArpsorPFCQNokD0M/f3y2EFDMXkYxyBgjDe31xZnXFgF1u5Un9LygOeyhlsR1HK
JxYo3d/cfUc3yUHEj4XcvSlDlELqaShsp585GEhD03+zPWBxZwVxfB+1GGR+gueC
DAmoCkcunCHE32Vm4Z8k+kWjg2guP9ffjP/dYx/ZoAS6yYLtBh+gjsSZVvDaVTjA
+PE7p9QobQfptEfTxWWDJMOCz5tjozLG5ONP5Usdz5SEDIaTlKqqFqMFi1V1jcFU
roEcNg61UUBKlvU0Kjqa2fVV5ReLPCi/sumNhjxRfQp9SM2QU7VaNa2UXrpzE/q6
/3xifWgszyr/bglUmV2eOQ05Up5ylV55aXo9hR845IQcScchNXUBRsbs/OlUVgoo
rAuaSmDPbk8PMjj4aB4qb1M+AEbljn0YgJoKN1oDZQlI7q5BwOI7JUzBEiLfLjJl
tpAsL9kCZxdO2aW2oJzinjM4aBiiq/V95kk15V0y5DPHNkZ0/YyRj8+DK8ar3Lra
VT/gDOYU2ieWNWypdVBPlW6nFzZaQCStXy0yur8JvRj8cxwM/JwKvMsYqLjaRWkZ
XYIJFHouYRva4XcYy8cu62qNKgjDUEd6PBFEMOAprIbqYYjSekh7bEYuwQnydbeK
2/urAiddG+TzdkVel3ZaP7NLj8F66Jqkm6iWzt8vCpK33zdQnQDwb7nH9y4dCC2C
BpFDJ52rrRznmAKTTY6WxtboI2ilEB6OKqxNXjY2hZgBF5CNNvTHC8UQPMtVMRGS
jlcHqdkBHIzDwfNu+Q/7DXsyL+SXYkRWex/f2UYfdUGVtcknk43H/LeokStOIB8f
ilC5akeV13aA/A33587nkOZW9P+IykplEHVV3aIdfp3fANlmDsrqPkX4kFB4PG0A
9C/YMdKOp/GhvaqABeZAGlHeZaP6oWhQOtWct68aRUpOYcDQzxR7TrBpg28vCNWI
pJY1uO8TL63PpO5V2hWknNEkEBt3B41uErpJq9zb7lUS4yVoMPVTQJoqar3YVjZ6
ygFMGvWyxpNRx+a3P0210DGmKPDA2OxTMJO7pm2zpMBAQ0tUGZvDooxQafIUko5E
wY00elg5IpahBp4JkQT+yzrOCiB8RGHDqpC2MYKZi/ukIgAQaOVOZY4rNjR1zrad
WK2faNvmIs80j8q/6Uk9C+Y/EYsu5Uqam5myNqT8tCEiibA2ZSWGcJ1rInUKgF+9
sDVkUBzsIRfpyNan7L3dUqFviHfk61uZPftBpley9SOHFpy3QqSjgRGUEpNkoHTz
3ICoCRhqObsWxySgFLVWRUhsLaf3oK4MPjsKvv52fuf1ZX0Ncci4ISn1qG4SQhOO
ULNWF4omoNE+AZYRvA9Fl3MeUVM/W8eUxDZ9wtpwVb8Xm/HDAWLlhldvsFWd8lcr
ARNE4vPTJraJMIpn+GHnJxvQ6NFkKe86HqexYQt2Bjhlh2C/LMSP9jA2WqVIJ1Ka
l0JdzEGinoT/H2j4jDezWNVixj1V+VPwI2jgze6MB39eu6Z8wuA5pTbpONL4HoCH
oqIHJQehmrrNyy/0MP/8TRnyo9h3vrPJu2/+yB+1KogxyeMOA91LvUQJnp3MGSX6
/PVRfBFQhbulQuMG0l3ZzCQNs2qH6CUnZzQKrgSijCfBAIx8Tww/xf6Y/IRZu34c
sfBGgq4w7XSLHaEQCWaN3YTzYFsWsyicUI3vDhSEQ9S3z+rJwM8VsV0JQlOHG9bY
G0N1iIfnY9ae0CScAqLa+fguhLixVQQ4V0lav7VTFdfV/x4p/p5oz9lGTQabNGg/
XOzr2pdthW3MZo84VJ/jLwfawzKqUeQPeO11dTsfmUtiiaMHh+Kg9DUS7gh02OAS
r6fUoGx5ZTIk+torbmt7oHBwpOSV0ZsVG50Wsk3L4+VWhmhHbrmDOODf+mrEU2rP
WFrijWXG9sT0USBVhf0NF8POkSCEjDISdQAV3cDEt8ACEDYkE2jSl26qE4fFD/ig
Vo6dmOSaNUiiYLkXleF9m6M2pjyQ2wX5wNReVx6mIwDRtcwr6aLGp8qwmhsoK3W1
byI75hiKA2QgrIFCQsTLXgrcA8uDC608Zdit81imNfWayFn4A4FQ4VrYt5/VybnY
5nSkV4jaGwJPRe+C6khkzIqKkT8ij1x/KLTehW2u++zIGROcrG899Kj5MPJ7JwvA
kRiXXGfY8hhaPS8N+pkRt8NJsLDPUXyaoP9a0Hldrco7VI6I+acl7BXeP5s7Xdzp
cQcELKuBggzXgSSUtEZR+bscGOqdLPNo32z7RvJTVth3nM/uZNulvM+9ZUwGOTTR
D1DaSTuu3Rjku2Da57z33cEBIkZ5Gs/OPvclXipnhDIHJb4byS82Kqxl9iHzqYfI
LGsDfJUzJ4LzicgAYYXvI8cMyt/H1QkufCbHmBr6vTOEJxekCwFwQWZw4mqOAu+E
YXk0yTeiLmyq/S6rlLaunl/LVN64Yu5z4eXCbPmfPxUbTGCzq1W373SLCD066k1C
sk5ocYhnIa7fJqDOOcOLmgrNeurcf4XLsn8e7p01+axJKgPMCWUrvGYGWiCowFDz
ss/tzXe8Y6FTRNiSqBRARlhuhkZb47xi5z0/dt0WeUcn8pbk17xcJjJwM2ESXvQN
WCJf5F+xpbXzR9KotqXX4qVBE4rWbqP4HX/BICfLyEUOScxCAMoD6J/x91VhbqDr
8UNYfsabMk9QcroZGF7gC5E9lIhtob8IEGUB7rw9LBkMUj0jXOfTYLZ4jidfcdBk
W1EbOuszon1y3hEjkFqLRJPi/0Ix77Rue9yLpyjdePo0MPAtHPZ/bNSp1uye9VNu
CNMzCVzo+g/ayWo3uo0rc6D+kbJpv5KoGLl2zK8J/6MKMXES4I5n4u9Z/wgyLwPb
YPzUrw+x73cBWIAaoIs0c6ywJNXTL2STN+xFgqKwtDpnDM+ftULFtEHLHoK9Zc25
+jsrXdDnh9qEhwoUcf7tFc5o1M0T/JkZZ9xh+UQPb05axLvMbJYStBr0QY9oPo7Z
7T2IXrxidNTtp73iwGSPRDSYnm3D/GYQBUZGAEWCj2NuTFsCtpy5Epggl15Feyd+
+xDQqj/YPmhM5ci7nRm1nUOhi9DiqswY/kRA3VsXKMNF7nNPaRb/bmmlhJl0iCP/
A6BLQXIcNKjj9mGTfaP7EZwfsg2Lt53z+9jKCTcz2/wxa/q0wQc33EloGpcQTbtf
0GbcpfGNzJ8LM8HfomI6Bo6YV+qorXLO/7iXrBumt04IYthavYcKUSsYyg1gQGB9
km/WGC6zwhhE3EndsYVOFTJ8i35DWA9F1mowg7f8w3RiywcrFsCdiFou/ixh2nWB
wXF1pb6IaKDwGn45FgAA3QrUgOUl+gg/7+fpNM2a5yNBbjMHxWBEJQw1RQx1hhrj
BYkdCGwvPwQOOenChxfhKoiTUbGchBVXMfEVmSMYQCcD66uKQ5JCw0+yPRhSjmRq
6EWgKsVUeZdO0nit4CuPj2t3SKsWfRCU9jmFxFW8iEcKOsZjowuMY5NyMy1aHoaf
+XJE8XoMX/tOkxaf+YfesAN6o2xbyP7Zot9LGgLeBgZh0h4ADjbCcdF3x2SfktUt
UGAvUBM1NWO4ugHrYKELPv0EoqNArmX57pyMMkINOBX7TzuDtjrbikGEalKNLtJc
TpJ5Feo57lzQ2nkMES0UXcjBS+1T72KasqoXLAMqikSQjHQ3mKvFBDmnyO6h2NKc
vBV/US5cMu37fIu4yXGSGMBmtMUsEEgyFaAIec4YUBlukMht57lhEd770Opm/qrC
EwVNykobimiuyArTfScFsVOWlPOtALfc5gX/twQWDTyxkD70Yt685hv5XcEShNOq
srx07TX8Kk49q6MSWziejvnaRGNCfCMrGuGI2HFlOpPn5lvThnCOxDf2Ul2xE9SB
tev+AaCNYA375Ir9QZtaWeP7Zh4epXUbg7ueu5ljvlyw5UbxjIpq4q7Y24tyyIUZ
WJq+78Ac6Y1ilTiVGPFMhp5AlRIx17xvrVreDu17iyJWD2yLleUkwXvE7a9edtTE
jQC30bSkydrEDSR3UUtLtceVSx9oe1K5ZwLKRrsBVrR+tYQmw8krUHRNlhS9rq7e
A44/Y57vTG7wMT19C2+2gLkNdK3Ais5w7jLTIodSTMHqOrz05VF5G2Rob23chGp8
lr5BitLHCIuIDgy3DvWaRx/SnfZ8HyntcA21f2u5VXa1EU3S1SaUqVz7S02XU7Vk
tIc4hF75YivrwrrkJZxY5IAYGjyK+Ce5v1yI1wMZmxYn9T3RgqzbI0nh6F5KawE1
ttvbb0jOzMQZKxCQuEBjX1p64jLzHWb4gh9pgabvL+vzJxC2mPDtOqrC4Cm+gFgg
S6nBRLLrRIr0mVFxZDl19geDv4A2ajYC2SFlaF5XM2SmMsOAino7xZs8vlSLgjnc
V5s7qkRQG7hXxfUi6emX9EQkytxyOmqeR5F5YIe2pqaSCnBqsj4rD2GKjiZpG7T9
5cqWJ2DKfhEojMVhKV2KIxseD3vt0qS4p1Q93gToJG87ssoDuJWJ2smyZsjQDIAs
OVKSvLrkEnB+VWXSPCedneWdezvfwIAA9JHjo5Dzc0SjnISLChDF1hRZaVq9vupf
YsCDYo6TORr6XqR5MlWt5ZByg5bQPuRoZ0GkEyOoyOFDR1wEnR+/qVDLth67V0/+
hEFwFLyfO4XeEyrj+wvfSk9qP2Y8AfCCVMvRMNwN6hmyT5ygivtEve0LvhwnjZkX
osI8yFXzoDerBe83iP1obgu6BBvCxC8C6LNf37kCkxBXM83oSVhPWW8xy56p8GWH
RDccZAfAc2ivnOKIWuOkpr5c2vPjfz/WRkLTeio3bu28YpUZyVCxBRrQWJJO5gPH
nJMvd3ZC0fPDhyHZQcaH3qlD0xUI6dnRb5btOXQGfU2ftdFZ2BzUJxnMIEmyd2Dg
bzkrJne5B8eYDTgarD4cr6GfZd+qDb+D+Qv9wLx0b4OkxEsfgD2X4gI+6DvX+llk
JPkdMlhb9XMlTFcB1qLmqC08rtgH/1vvuGm0oUsIhrb9CDVR3xx4FwT/toDAPoRm
GZ/AdiwP6PBywgtK8n6PiZsqKE3EVXLwKhRAn3rDUYaHru6qbLXRqqkZOsylXr6M
txkNZ0aWJNqgNoGkS/qFarSY7qTJEtVu4KNB8RLuuiYkY7QayIGvwltpER/1h3JX
bXJAAMp9TlfQE/ZvEorQY4kX8MvxsKIke4w/VHrllLnNUzd+zoMbcL4e2oqiLTGH

//pragma protect end_data_block
//pragma protect digest_block
5f3+gX/5qxP58baREmV3KVzH/28=
//pragma protect end_digest_block
//pragma protect end_protected
