// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+sA04Vmpl+LhQdEcd8u/Hna0mKJL6LNjAz3QiEeWO4ehiUeU1TW5kMKopscINwVT
mnh5TD2uRVn4F+5NdizIABnIOlS7GoTKTXILn/6L869kns4RixDSvuItOqGlKBCi
J5NneQH7Y+pJf0W+BRUftysvb94uaN9n2Ox8mkZ3OHZzY1cuz2D2JQ==
//pragma protect end_key_block
//pragma protect digest_block
e0dGvlZflE5trdqO8bPa4tjdsYk=
//pragma protect end_digest_block
//pragma protect data_block
5ZuIUyivAUVggJ6rdw7XZbvh6nB6VTwvCwRJeBwIy6eMuk+R1kTeN9ASuHaYEre5
Lu5B43/VTzSlZU+XUKKXyufThmOopCvcsqhFntefnzzTSo+bZ3HhzyWj/C0PJfOg
H217XtMwJrh6Ol564SqpoGGaCZ+TJVt3rYPK8tVXPnE0IVyt9iLXcEQGrev6cCVQ
sxLl7hUaoR4moy8pHq0GsdPuSW6iLsIAXDpuGuuCodSOPFTmDh/6daksYxdxbvf7
LoaOHfdJl8MuttyjBUk6QrPPoCEdyAbgPNDEVuccYIsBK8svvBzDbUv4Q8yahcNn
ZOvWyIyD12avPWdoE8mpO1hTw3enPaD7aaEdnJdOzZtXQVEWVfLrST1yYZ17u29b
+6TeJ71sNKxCCCpSaH4pHbNbYJVaaa0IgHSxhP5TfIEBzX8GQd2Hs0cZ62QPNjKO
5ZFzMkcSFoShRTJfadmT6va0gf6Mb6nEAR+P3hu6dBF4q6beh3jWQxBETwtnT6JU
mH+jTYn4zwbwNq78p2PH0hs+ropyb4LgfNmYZTZloHUztc1Pex4hHH4HvyKrGLMp
WAqBr8jQlhodAV1Ker0eLOGgLkXUxMfHidS5l4yLTrUbDL9Y/VB+n2ltpM1FLaKI
abxpCusD6L2iYxmOqdkqccFbV1TaAZZ6yQPPgkPeTAKITlLIY2ZVy2wLnwJ2WsTh
wzAxmhhFnNeuFxYZwwx5JJs8OIJ779Aqjs6eBl/aSZedzRHWOQIiMvSBuaeaXIh+
tjlKA+yko9K+df5ZbvxvsoqEOBCMgwh+BzWqvWJFyZqO13mACSGT3DFNZDqtEwt8
2bUbarWmsXtfmaQ2qwC7EAoa/6fiaziHYLfj39UEEmyAwvz5N5XkHWqVPGKqgL+I
TMStNo6Mada1cN5BKSQgDvw2E6D2v0nE3Oa91IKo9z9LEgzjuL35FA5LwnuR9wOQ
SPO308PDBJliJoiA92+xRaGwiWGeuuXrBsFOID4OUTrcb9MlKUiIgy4IeEMR9mgj
O+XLVTpQW2ywEX4OJ9lifBrVo42sOofNtE0cQovF5MXU1ghM2FTG3aalxZCFkhzx
frRzm2D2Yd1yn11aJvu0VcV0eCEHXOSgBxZ1RsWbwSRIF4NZz1Aa21NN6ZUvXRGv
swPNvp0cHJwXxHuwiUXRnzu5k1Jtg5UHxvQASgLNmuJXUQP9FiP07GET4o4SiEa/
E8y8Y4IYhRAmDMqVjObUA5NdIxHBtQOPm5dbyzx//WOYloAsZzJ4wphBxydec6Mv
iGcUtnAyUZd1z/jQIQj3zJWl2boB9bmnc05MqnYDAcQTZfkORVYn+6ogxb33z2jh
KzfGDyp1tnbgeOGnxDa0fLu/KyYRDBDVLa5sy/AuZYRygmYUKYLWsYuImDLLyork
nrSNy5ljt5ykAO+luIrXDV08C14k8XwgZZVx2oxSIsZFfwHGyiPYaFDxooHgEPhv
4DGe8qoBcNg/a93d7+F8SPICuHLE9z28UGgxbhli003y7V9I4U4HzlVOIrremNoA
8n8DQ2GJIBPOV4Vr2T/2N7+PvktiJek8eyIdNmx3Osw1GLhZzQvjl2gvniszQnbU
JZaDBRjCZ1WRisZFq9+8lkQGO04ty4if+znlh6rJgEozezGxEJbV7cPpJa43ht+k
3/UlYVTFKl1by4o82w6IqUU/xdaBRqQortRGX+IIqbGmZb7K1pvkq9iW0cIgWCgY
+2sIrn0Tjtt1CjdkzDOd5NxeiPVDzWeZ1aWMUptHzo973irYNSJfSDh+9TPyxvBF
sOejiav1FUbRSS6oztpYR03nWXt/IQH85EKW9t8UN7UjUNLXn84+9/Cz9JFEfLyD
oK8VNCfPd6jwAZ1jeFeHPn2pn1Cd6/QiNDMVSteh2XAdstQwrJ6rJaMhWn/k70lL
sUjxQBz9DpucIZrjmBD7QW9vgIX5e7/dsYc7TW4n5DRHQbnQl2p7AXlX9fB2FWne
RoGFe+P4A+bl3C3LeSaplQcVkais5P6wgKxT1sgce6XwNReg/VVX92H02tCKtkkE
JfV5PIQgWhYf1u9xwKO4ZLGbXh7zivIRYndzevJIxLHXqpdn4OmgcZzDcsTcVyWJ
6WC2mImCR+TWMv/vu7hZ1fdlzJY3bHFc9ORmDcnfP9ungRMg/Hmri4efaJgGS+Y7
oP7LMd6MmB6J7lxa7pAo4fFqK3WnEYNLnwP8dbpysGGQakmRHa+xFYHCcz7cIDVS
qDIEWGpl81WaaphjGDgXfHx4OZts2CQ8WnW6Rsi9HeP/C9uMHm06bULkzc4sp7eQ
J7Zb8DuXQHwUVqThpQ05pZ4kLZ2DvbxXQDDZwHJeruPOBfVNWwHak/0JoXUo+Qd0
QcwDRvwaOdG+4wp3itkbg8/VqEFZT65qKoOXsOjd6HmcOqyoaJyU70LAea0sMlVT
T3E0EzhgGhNGzVsunCp+LhH1JvC8gye073uR7dEA4C7ZssfRHyJW7lJ+6d+Z831g
wSAPtBmFPT/7ac8y2E3n8OtYdLC0INC27GeEocs7h7QdBhpEhflJFCMP0iQjwMMJ
sVHhN9uYgdWt/KAed5SFndmhIYScWCBp+fVb792+8JCw0AAbFOgJZPFKGntLMexX
lcBZP3G+N5qFTpKaO/c0cMVeI5Dj5ObaMFdAPJkOqlpLtj9qztLxykvuomh14NQB
uXPCRWTfsUA+RILjohPrinxd7wl4IBSpv/G96EEiqOJv1bdJLPmrP5weWq2HMRh9
j3s4toB9vK3tO6ljS0/W/xxYfCl4i87OOoxMCuj2D5oqGf0SwbyeQl8xAcgh5hdq
I2/w9VVdBikI0UDydtGRojPAzep+yXPPUkczQ8t2tbOl390uOylTG6C1Z3nbkgIp
+uhxrOAQQwlByLbyVP/8OSd+mDIbQQk7T/9n9IfZzl45P6JfGS4VvyWeirL/VEmt
URn095I4F5jwU+atPKpcdlEvYEemfbycMXw3LvwIomyB+1JvIk7FkOFA6/D4a9yR
VhbdE5oAxxi/9oiKQtyHvLFix8Sroj/VNaxghMKgaugOKDrAnS/P36ujY3HMHyIN
N4bNf5c0bEPNU1hPa5gbrEE2FBUXAuNO9m4k6GM0wbLugui+fIrIuKe56g/AS6UR
byzRy6NhKijdI4tdUiWZXjkZUYgebhXZ6L5OzlAXyJdP39KtH78rajGvdIj/HLjc
00QFTyRyvwhfezb6CKqmkTEbAVe4TMikJijhPUF04ADTvvc/SBCzRWLbjEXGhwIE
sE7/NWxqyh3W4dQNecGfNS71eAbkBtvttoKJ9hP4G2F9FfTmbf4i+SdXTzL/y2jT
b9vdN0RGpEltra6UPnU71aOGmTMrhLNoG9h5WJF6hEjrVpnWfYtjOkX9CKaPD2rv
Qij8L3hKXr3xV5iTRv9VVssruUc1q102WQMl7LN1+OLCZYdNvwLcLVK2j5TdlKpO
qWKy6as4jzCBm8inm9hcFyzgOdobbtQVhJjxxBf5LdqCJr1C9RrTEShJ0yj33suw
cypImdcKujhfzdFidLVdqKiCWvJBDXzyrlBoiTKDFMesS/uv+yFYxRRy5ah+5WsH
HgYHyq6nruF5h88yBf4nAHZb6c57abliHrXtX7UT7OiL4RVE4BzWQbCSMQXD3WVd
sSlPphfVpOBcYSb55s+P5DwbdO4YOkSw3uuC83CQer20eoBeQb+WOf5XAZULEPd3
qMX2uSa6UGHW14GLAy4wIw4Q5kdjXPhOH4K9D/V0BBahDuSz7jOe7Q0Gh5aejGct
ALzXvJyWft90Bbg1WpIBhhtlJV7f4BvMwFGzFQ/H32VJntkG3iYEasFaftnX7AMF
5FyNjzbTp9pCECV6m2P1WCq+z8BmPw143bpA15ik3zVnrk40V+D+o20I3Qkdgdbx
pWow8f0H45gOW8WFGuh4bq0tQ9ta8Q/soUCNI17TrwNzPCWKyGHv7DF4zRnbEDSQ
hTX35M8iExTNePtWg1XsAwfOthhx50zfSGKrdDEz1scieAY5wRqY/Vkh8qfQ9umo
m+YXRB8cSgnHRJgAbasLrRKzi11gAZzLSpTcAfg2ijW0xz2NsPEHcapX4NdOA5UH
C1xblKU4x8QWKfa4tWEeKfikIzAJEtouLGLIxb4yhTf/RRBd5E/XvsOcY/oekAt0
sKWRE/uroJhlfCTre8Hxg88FJvFn0mhM9SoDy8dhJiaOnRSHa9vapZj/gzsAuwrx
eRq5s0NBCcpmLWBHunuzGLyQIBWCwCXedUjK/VU+rHQ4A9RGrnkmZ2loIOe/w64O
znZN+7k8B1xiEjQD225QMBGDZlZoMrULyjRSMdyceyqMAzjP3wbulv+cb78XiB58
Ctmu1oKO0Gxt5ZiUXx7TM6psdI93J1J0SY9myeiy0/ly4GcyFu0ZFeGVBtXVFoLa
0unzNmumtTly0/+Nvgx0mW3SIor/jTma+dY0xFLUcz/dQuANtBkXJsvrldaIBN8j
s7pjossIbteGG6wZfWKCtZEi5nwiuvG8DYsMeRM83tXt46CPl7eZ0R6qA7DsYODB
5P+PQApPYK/lB+qL9n+2Ny7McJvOekLOJkHhQ0B/rQDJN+OQJsDbplrE796eV+xB
RSPluEWe9BTDMi1C8vJvSbjU5XhMSs7+DochnpXE6OhYEdqFADhlFTANY8D9Fvcv
Btu8MuqVaR88ZEZDzL65gWyOz+SxFZjw52nf+0uk/QZ1Hjhs6Y3y/MSHQ6zoYVsb
W2i4Qd+90mdgXgQX0K8GLsuj8RYP9nNmMQxuAlAKOTaCRCh5K+o3Qu4OmeegSX/P
Ww9KtIdZnyYaCgYyB0uYiHMkDQiaq0QZwCjCnt+vp8UcV0LrotOLAv+kkjITG4xH
aQiaMTw+BA5O84rk98OSLUlT+E8M3iU4yLpia0oqg58UmcrQWCx3r1MNdfHesr0y
hp2hQF0sZNBbCXG/AQCupzTi1+9qOivqvRTrm7MQVGRD/CJ8CSM6SGbG1pmAFO7T
MOPaQF06zKIYQ/HCg7RStea8zv8R2Q2YGTNVQyzcA1Kn/VDr18NGBiI8D3OK8xaf
E541zPGaNopR52qM23zuWeirw1THBwVrqnrVpUH3ksOt2+uYO7zMXnmI5wuJqQ1P
9oYv7LyuVI1VFKnva+x/HwMxchSdeaRd+N0m4rZPyp2veLStKGCDcNmhrrLRFGu+
BbwXCqv9CkO07FkiU+/BJZDeovhPrfQSxtC0nAhI9+JBD/z45byZQ1+3swPYRD2V
AwJG3LkjsE7WyYMO1kqa5MHXO+kkGpgXdk5LSTm7Ipc8Rwg+vSviPKYv2mO/ulgw
iZsfOBnkMEJAwgL7yCUiFldYXBm6oSJ1YCgXwsXJlM90AiYD+vdudBLKLIKNCY74
TfhziKQFTW+uz3DBmw1bHJYSHdOaC3vwYnnVKLCowR0JDchq6ZkUnRTzbl+iMpww
7EBV7jVekowDTgHklCxu5+wt0+9hZIbHAGo5m0V0nvhr6Cb5lOiNwTsDPKaGXFfu
X/V/CTQE2wMO89yaiW+d9UogGdYUVZOk8Fa5C9qhBHem7Qe6TlWx43iaphoO66Y2
hPNMPAN0IXyZ7GAWzgT7ZpWN5+jDAq1wU8T07aBv6idwL9KNBBT2U81ee6mX/U1g
Vp4M+VXr+nWAsbWebIhV4BplP+6merJlS4PlpkbdLoEk+VEYIjCCChNNpl6GjM1F
5Duy6AVgvm20+1tN1bBIaPTiBZOGtmCPD6uBtwqKURPZBMmOTGYMBKJkL7O/PSGR
hVoAjDwusdTwpe4k1BTtlct8xM4HeC6oGvoc7wDKPHpehL7tbl2AO2bLfhXAnZ1c
etV+JQy4knHTDipMC4mkRiQjrjjpUB+8Tv4b41j5Uh358mB3fU+y8yqnZujCZROv
7Sqw9z08mJ/BNxoM8ASEzDJzFOpY2lECBNmbYjqe3Oww1Z2N2cdRDCArmdbZyBHr
mzomRfQCVnNGui7bB0C/xMN1MCGXgQwQrA7fIlWvHDvv47HP3Oa3gEU5PBizQ7HX
aMegIbJNOTZvesBujW5JLStek3KmH1A3ijB8xb2l40c4X8Ft97538J4vKAcyjtvY
VLXH7YvcruUPMnh0NdIKJP8bNWwr9zQrX2WxB2CqkWFoVJVeV+Js9ATNRmmEWZvH
yJ7Ry/T82OKyUxOivLwu7o7YqnbbQP2pLG3S/C9B8YhhRUxS1Z/1nJX83L7fY+qe
/jmr+CWqiYxx943SodEjxxhpAOpIfDPcKqCiqlnvRHf0+FY2zHoRZcl+G6jt0hpU
gCaL0M79UMOTY3+/xq0gtXB2jTHL0mcDZrBx+gXz8z6Li0fZ8zLm9b174kEFn2lT
t5WMfuIbBLlTDZxAfZfBBkyFprLRul1PH6rhLD8DfChxW6nAIdQzZ5sxjLwZuX7f
/XsJoO4Amvs5rkLes1whRBZGTgc/w0KnEs4VZYT90lwQi7q1/1hhy7Q9IoVRHuDa
sOZN/u7qLi+V1BZ1bkZfAbDrOCFqW1KPaIdKj50PLOUUyWoqTByjgc4rcv6XTCSA
VSfTVooMnQT/tKYhTHSGihOjpMM14UbBOioD2eL6vYIYHlW9n78Vrq6fxIbkF+K4
il8iEt76CuYqjL1L8SbFDDdKtOvEqrznOSanppG7MPs6D+dLodyE6afBhkvLwS/i
W26hucqED1iJvH9HKiiLRx571iR7Majv6CCPk8ebWC8dr5SxtHA34g9vhpdTY0R0
DiT4jxrKkrJIN8RImzfc4BNAHtn+CYsxfip3dnT5hsA1V+qXgLM/2zBHN6cSG27p
w1sCf+q+fYtwow0PJBpXPLvkjyQ0QJ6RJXThCqbUJp58creoLA9IJhIoXUwxlFqD
mMk2lxI34RzLPfqwyqSxpno0W6yqHTPwGY+mZ/llnztqcQaKXuUMebYs2Ye/uvlB
tDA7LQ5M+3v1k8fMPTNLYkjtT1x60p8eU12jWhKKmuqBNK+gRxhJ0pppIxcY/7il
9qzAunPTVmKRaZuVNIy7PwydWafzE/52oYk8VrTFrwHSRXyU2nRjVNgTcEjN0S6w
Ua2jWtA4ZfQambC/orMODhy+hY/O0VMoeLdFrzBJ4oWUJHHe2ak5oH6PpIBTPS/G
IWmWZRLghtKUv52+DTgi6O37nkBTicA3G98TpOkYOFYYyj4SSTc0MmVhCDnt/sbk
qmQsCp4y6nOF/WzVqM9K7/zb893T/TcIoXQ5xVw9OuBzcPeA3cwbG8oNaGAaxzhc
RhcC94LkChRjjxcvV67dpawTsW2Z7MJIkRT1+uFfJjFP2OW7NAwl/0gTm7OLF/00
L+rY2YFDYZYb6Zqd1mqqkLRoQIl3TZROnkHBZvTyE/j2cgeBHAdu24Wn7LE85rx2
Jy8pKO0n4Kn0T20ieSB2ARkLpJ5sp+28uFhh3KnZvomd2hYpMhtbcJltVB6OBHL0
rDau9LaXOsNUTvcYFvANUYFLwYO6fAfsJWWFwE4/KK4DU3L8pFrjLmR24UTgTNfa
orUyLr6UJt/arb6lvY4fLFQqZyZhqSYMs/gcAakfOnXAVDOL9VQ0xqOEIxQfobLU
Gog0tXmbRI5GCAstMYf1aWxQf04Q6VC/7uUff9y7Yo3zK+dt8yxRMwoEKn0XQDli
Pz6hsFJ9MEZSwhtwt2v1LLKN2jmkDk7vrHjriXeauCpZ3KwllvDUP70Mm2z8TwWs
qlTqDTrjHLVRv9hgvmSYI9Yly5/5j1x1yKXUvGEvw8oGpKetci5xef9TuqnfXRS9
sA5/BARy5+7SNTYkuA8vj16AzciY/xcSkDOzwISltSYtiYoC1SIHXAQxMU4yPHqO
0sP7F5MOHaQ+HV9aLZfKQlBP6B3LGpUNUPtCzr8XIRPfqXzR9qWuTcsMdjohseGB
hG2QrIGTU7AGt8OifMci0rm3cVCnxzk0wL4XZWhYF80kQdftlWkRKxFsm44jXmqd
Ddlkh2mtXSlLkZJrFS3e/YfdUW0+g5zv4WD1F6aq8QETuJwJ3ew16kaxqP2buFb1
zx+MJ4f0AUsyB/JN3Wr/smSI98BwRPGxcqm7x1uv2Q5m6Bsd05PAGX1DLIxiXDbP
MDE6godGk4lLTvazV3R4SHT+twItkHubD6XTs80PXpMQwRZeGll6EXQ7UUOopYqL
rCY3p1QR/WPQ52jgjRsHZ47AFAhY53b1paDy3xpQn6en/d28wEBvVeRrTpxPpjrC
Kfcb0DyaLzZAAOLIXBtQrv3OpnONBF4iZySMfzQXHyUxzINvnEe4cDhyE/oaWVGC
AsHh1DS8Hs24OgKHe5ucxYmonh7s7Z2jFM+XSIdzMc+wPpSGdD1kOgusqsdPb5Qc
Ta1wI8F4LCVOXoqtnN6DLaTGTTpkijGheLOJz1bhQhIsEeBvbNCztIMZjmdSsw6U
eKnOQa6di5361r2NHM1SDrmD66+xQazoy8QQcezG3Tc65DIA8fVreXWAs+zrYcMw
8YOJ0H5p6ZVxK32zP8l1qVD89f/gGygEthfrf6rHabuq5RLFdBDsXtUfsWeZqA97
RRYLUUGhDA/y1NGwt56rjmPCzKG+xOGgCYSUhkTjJyWCs/mlxp8XMr6jZb8QXEt0
KA+vMyE1G2eGr+sgev/o07IYYkKOGsbbdXESqxPcc7YKEMeQzJI50NnyDrmz3Dw7
Wh4/VCZ8LxIjsXeqKVLLGgosyCmnQZS3IVXWN99ZfxJrZA1yEWrPsIisXwA9/1JU
DjYzeCPN9WshBRuAM5zo4hQAu6LJwzyySDj8V4LWIhRukXo7aXm13f182XcqG8B+
TIDj4aXUYvsOUADOgs/vXa2oWFH1AdABLTIO4iAOMTaxsqKZ5gOgdp0GD2Uy4Xrh
Ziv5RgRYMUZN+sj0GeRV1xBordkGcyiygZXYnh/YzGUWWp2dq8PBldJDpTogcKiT
3bcxT5CEQUgf/XCbDZxx042sgUqaPcZhqZQKXLiKaS2dQ8NKjZqP77BaCU16OBl5
+LQM7+KCEoz2sg8+PUkD6+EebFgh3u3/xAmqswRg/o4f3JqVJtzty5zP0oPCdc6e
TL0ZmQNvh2YW71xvS+w51MD5/3mf3BseiG8iCB2W2X3IAWzI3Vyhq9vqZjv+g9ML
tVcCtCa9gKAXUTRPpjJrk4NRJgu+sKBtkOCIuhfpy7y0mGLio7fyP1wJ19tu6Ozb
Wgl5T0RAnyNiewbZyHs14MacdBsz+pNP+3jOMiVQeIIYfZTCrK0baq5Yy0FIkUFz
wDj8wsIfI81XmkDXb1/FfTZP/hrXhBqrlTsKk38lE02rpRXu1b//hsnAA6GZsrr4
vU/mf5dSrdVn51utnpO83OspNxU2GJeTaA3veHV3n3ikskgL61Zgxfoqyr1e/pzz
ddiI3tqWN5w+BwmsQuOayAWDyPRDQN79jeib+0Tv2NmKF/51ajYKPn/7WAeT/zd1
S9kIzU69/NKVABZ1MhlqXNdE6ZIx6gS+zAdDirTzHcRbI0VA/J19Dr21HNJjGdHZ
H3Hb36YJzMrQ9gKH2EGoY0sjdZZkgoKS4UpkFvVHJuk33fLGAupog8CzpWx2z6yA
ptdwFE+qdwagmrUNfFIZjQXZi1TeD++orrjNCo4O6han7vzBTWlabWvIyutSIcnW
mjIAgGRjkx0OxduhGBzJ1k1/vShi74Vl63BpN6/I7a0rZKhS6mgzenjPR/dbqEaH
iWSOfaEiByDH1Uo/vBGiIxjb8LA5SBSZ5LaCQX9iVh2bsZXe84MxR36a0vvYuvqF
XxcDkARidhled1QnJEFQzfCp3CUL/Oa+0PxTCb4+1HyNBwTTo4PnKK9OUUnTyHeI
3tkD+K92mzOPbLy7eu3B8O4bxDrS+BwfIZfv5sWERMfNej9L9qXerZPbiYYM7CRi
YPuev8l1ODyt1rRF0UIhVWBNDPO96/ekE+FLf2H5GSF5lJ+cjL2uN91ecCZT4Qrw
bXPKboz0e5dZb1HUTPApwPorII+vzyt2Vo2grmHgMq66VpuzjcB3dyqtFAsEWhum
409NbQTULRvzyXNk4MkxrNOKTVn0Ra+JxunbcL+tff7NRaKOvxhd6yhrv5gYAQdy
HEmNFWDVu70GVlYf1hrgJL81ESaXtPrWsRurudvENzm8Gsm9KUduAQMLgTLBnkhD
Ls5LZS/fiCS6lB6hWaZ4D6IoJvsu7XUEeRFbRu0TXnxvBp8G2cwW/aI/ZQ51YZgN
Pgij64/MuVQIyHwZrMEdLT7+MnxcwKQcKuM2A8aTt6b5KFVdbTFmkhCmcVIjbI5F
JWS0d2FGKKLIkTCcMZUaY3PHbxvUPM0SolT13D1eL2JiJimVGmZIh7Ind20h6whX
EfIGJPh6yZXi+EQQ2B6BZH/D+POUEoEkTddpmWHegHhXJGqBUiI5bfromgWlMU9+
e7zK4bemN5vazlUz/ZYpwL5eLmN0L/xiKyNJpDG9Cu0ZML/hFAWcYXk85G70JpOc
T9BL+leGE16xBXyDE2db3M3+Aaad/8W9uaF+GmllTZR/xbhG9CdvrfqTQQuhhXy2
KlA5Nqwr5C2qQtZYTGgI5mmhvZUbtS1x1FoCpOAN1zR8xkIHdt3VUc0ifbx+IWO0
R0CLs0SMZRFD2i/3eArK0PDDixsh7wb3CPDFSFyGI8A2i0g7ZLSxKQhNqoD6cFLn
p64KFk65DtWp86y52FbM9SZ5b+TSOaizR3s2643p78rnXb8Au1IYZW2KuBf+HNqH
goRCgXWJBG66k5NxgXGInVAJ8VTbZcIIw4IwjlTwc2FYz5klsPzMkHmQ9OUrcGbW
RZrL8jNRvQuLYZUdWe+gjt7u5SGA6HuXFffQAh2pUwNd950hgPFbOL5VqCPHoW4E
d/SYfIuNkNUQUXjamiiwnLOOj94HAnMfTDCIP7it2cVZ1oRGkCpdix9DfjlH2Pdw
se5J74WxyhmTKEXZ6YkvYYvNczmQGPvPxN4L4GXCbuwZxhMRAGuckIgTk1izAu7O
rJdWnaOxv0b+oy+JinqOvWP2Fd52W75a2APSWnms/K8MsGafx4wTtvdXW2628BMp
h8v+rntN0Jtyunt1OwcCOMQMkw//xFI6l1pJNwEfR/11nqrMODZLoDo+mm4eeIU7
M3mxD4hSx7L3g4YNWh2WawkOgj9xPaVdwFbIW33fSswFt+CtmUZO8qpJG0KyO5Pu
xCcFxOiJiND1K83P0QqcU3EX5k/CiCV2Ig7s5KvdvbHfpyiN2Y83udGGUnbvtmsy
2ojQ1vX9v+P2DPhBWwgs8WOFO5wqPIOpXjt65lNexQpk/avgwsym49o0Ey+LUHtx
OEdBnXeLyisq/Ely5XzEMiYmRcbCkJvrCs/4IqZPhGnxiOcXspyp4oON/znGLnu1
2ClSlPu0yw3oq7X43jHlld6rtfYPdKb606McE8bVaQZL1GlxvNefJcYS4aEzeJMI
qasqxQf1zxkanS5JGDKfCF5FH+V+eDKfEVKKpdKjubosxd0bW+NTlRAbw3fWBAkg
NwkAjzpQYNB1iIXTY53b9ME+SKY3oyH0oynDr4FdQ44S2hOQsPRKjgF0cu6A9d6Y
BcKHjxxp4GjuoPEUITusvzGJLJTGca8n4TYTc6sKifee05Zjf6a+Akoy7fkEoZbP
YdJ9arB9W6z1kPWb7b/H/Nzci+xCqfgJ9BXLrpWLxu2AmDTEOL68/MUwoSSpoJ71
ML1RbxP6g3pAwtSqt9U24h67tCVRpNortOXKa8mJREoFHPaZXnYeXwvn4+g2QsnD
VKf3jP6B9omeGzPalxmC6P7KvApoojU3CPR9RKB9mMaHOQ0buaiMYOBycPlwmXGH
S/QS0Bhr69fwjRtQ7Zln3mBGGzU5pZH1zkS+Sg8yN85TxWQlpVdJ5+GmtxmeuBPJ
7lY4HopNO8DMdlbjoEro4UWzmXpCajxnt2QBXhoZZyCPNmn8l1IxwUVVn3r2UdEW
AeA+aO/mm/0wX0S/f+Qp6iDOq9A1i9Y/z9kintL3fwiASAZ8q8QKUxhqIfObWy6f
C9duFxQI5j2VfFKsZLRKB4WTtC92F/oBHCcblyQTwRqb57jfY+KO9QBLnJmHr6Sj
v9lphWECBvQ12bTyT9u1VQoHkewA4bf2BCVB/6QqPHguxTuX1IdWc0nfntDZPTcr
12cFzhtmRSMzVuA4jNFntysrLZVm780tMJraffCsorKDC6lOF6vY0PHvyWP349pQ
7RHUADx8MABeRNRs3Qn4alj2lkR3NhcHLf2R7fVdw+t4+YBEBr6SIB/fgpeChJZc
9AcOlKvdc64fPdBJSmAuRBPHxd1tUP+PuC1UuWZy1bVFNBHKbOkKsAG98lK7Su+T
6JHrCuKuNETBuZ87D3QvSZHj55jVs99LaB8XzhChccKI9vP3SdY2QZl4HvjEOeun
jvMpFlNRPlRysHkubqSZAu6QbBzxanhuW3GG2a3O2z7vQ7n2oUWX2TgV1O3vxfs/
2eE/2yB3IefZf9hZ15dkCmOcVGZrz10FhGYrvsOZtR861efwGiy+rHHy6rSZK7Ij
PuU72qcR00CVn5ccuglBMm9PnZe4FawmVpXuVDHw2xZzJ/Fn4KiqSyleVoSmR7DD
khB//3SoireRCT+faiILO+MvLUGP4tutkPiyYQQKMzF/P2cbmg4FzvC6aPB7uTPA
sHWjPQ2rzuYJ+Eml+6RmK2q40iqV5nxmuPC9RRDt/+d7LnbeDyqlcXHYSLaQqkMz
HVCNazaJm+gvbBunK2wfNdzLxGRr9uwMVmC2ITMYIRdMn3Q+JjqSPaXBBMMr3SqU
H6tUn2shBtOPu+BrQVypVjWrSrnO3z7MRxeiC96+tic8gl8M9gyLikeAmoFl5YHX
mVQrXO06d4y8cBoKvWUFivDDY6BmuiRSa+EFDeMCIduhRay4y7qhDO6mFoxeUrrD
GnAkA52DOnnBvCkHlpxeig2EfMZZ4YISxJUxg+1MBuBH+72xQCJFSWo8zrRJPdxF
4V6O2jJcHiHh+4QLS8hbIP1TEp7rDpIlL6vgeL/WkrE/Fgld4e50t54GmNwuGmwY
6OrTaPejVR7+VTI6MB3cQb/qwmHON3Js7WtlXj26xwzvflrbu2hd8dmAX9OBfdWc
d46jwE0KTFtSxdFgHew5dzHa6AREl/PoYvHYhSAlaSno56o4UMDTuRiQ0mcp3fy8
CcQOl74BLkVyU9R7ZS/b5cyoshq1U2zLd7aqG8vAzFfPbB4r76TJ9fda+X9AN4Wj
UoSqswCchQ2D8uIt9bC/9aFJjgiaEl2CUnPDlbo+zRJ3ruIoqRVNuuEvoNLDBmri
sM21QkKK5TSCUqEI0QCFzrWep12Xl6o1qXwUD79BwzwaP8XZSOzQRqF9Fcd5Flic
TwXqAlVIQwO+cvWCeh0tQFUGiK6b5uop1EGRtK3A1RVa3SPtx34g0Z63TSVUMFin
VjEbJy2llX7hjOGyWJfN7ELIs6Q+YjgWlf+vCoK7qjObjXHI8u7MpJqWAGLChi64
Tmaa+jhxdXp8QA0HsM/hYYf6O6u4rYFO0uPkogUdW3MOW0yr8rkGnwds2uhv/N1+
LqD0qf5xPDeBBvVT6LkIjzahR6mx5BZTZIH64jNGsEjY5c1OuKQgwhA5xU2KDimo
DdYxlZJpH61pC9qksihqDoahGZQyo/JpqdxW0YXhbuYNEo0tQoEneNRwSfWwqpbD
Z8rIueWO445q844/cqyeXAZJqr9T2kaO1uRhHwdcX7RrBvW3wSwUD9JS+ssBE8Uy
z575HRzgjoy+sfi16++IYHJNOLkoCizIK+82sp1XjIW8daZYCw/iXiWfHTkXq5r9
ZAKiod8vy8UbfBIjG/HU+/gfUTzSmAK8kJPmotRSDKohZvhmGwPD23bFulVomIYS
f3ptRpYQsKjnnMJAoy2oJmAstOFowdy9dOvxMzt6gsAgbVOIHiDc4Fn1dOeoFYdb
R50jAKxxPuWbOuYGsBgmqvhBSk/4SXiv3Cnu6e2+uRm1JIsXsSOBajb9lIa8Vx5+
EV/aYx/llHYwcQL0HW04c6izknchLgfxDU2BXaZE3wHKaDNwQfqk4E86FbioF+h8
AlJGnR/hoZCQeTkreklHezIB/npatRoEGPJ5/yYRj3ae83Vn/JSrnItx+g11M54N
jXd5evu0Zm9I2AdwwCkYNmHd1iOiRSYU6uMIKf0DM1gzc8WivxEi4UD46BxHhZHY
dZyH5ON9OVfoMK3jHlT+e8yim5R7RmrbLVaVYqzblX6R+l0p/tx5g4s1DKNGB58k
hWhjUFdguWUg3wkMx657njv/UmPPuiFPBgbF56ZmWPIkg+q5nzeKt5DpjEHdXyK8
d25tYyx267NFl5qSy9c14CXFdK8ajCMCmR2SDNrFwT5+9cb5PM71AlTUp28pG9RI
SeDr9YoSRd190Z5A0/WOi8et+nBM1KNUOoXfz86tdHC8gsaD+i+zL2zRGprDp8EZ
AX8ALB4nusRiNhVKbIPGkIJxXzeIvWBY5Xvl2oEU6giw/LmozO8wfbncSxeJsLFH
udktEfaLedefjWUcL4e9BIkiTlpNmokU+WgTbpJsiO0Dbj48CNQPQbUF4dU4gPI6
TzDTQBulKMhkQ8YnhCmGT0Yb8UoXHjG7EGu4tu7OV5ngOynn8yFg5xzeq2M4oJ7z
REgieujZVNylBbvX/RfEtWik+qqYRmY0IU0mzOEee5jcxTbqSFdDwZw1Fy/F+Pvg
CJBenLvGAbHIVFtvAPQUbaTDuYyKzUExvCdtOX7Lhsj+TUeEg3bMw5slj8WAww+d
Z8Ojzj64rqYGgrlgyfYKgcV0SZGFWHahOhynDkq5VxguEB7IXU6RXO3cujxT+r79
eB7o+EaES9M/8rLzdqDKKhn7mo5flNATCjCwHBiK9Raeq+saq4PwTuieUJZQnLFg
E959Tw0vA0SKfisUeScQ3SDo05roiSTeZnb5T2FbuKqBcvs8FvJy5onRNaVkJh8z
ztwDPqLP4WQpg9XQugOKDdOTbSTgs6tqq41Bn9fXVc86fV1NR4D9yNyhAKZLfJ+P
/P55ZxGR4COXB49+3OTcHyIf2YiKWk0oTeXXqVysX0biW14L8DAul1QfnNXQoXPO
jpBYbHOfZNOCGTQwF/CLRSJNL8fp6qQ2Ib3j5GzhnIvloJi01YZjFx6Tnc00DDeW
yJ47IhTDBLPFHxjzgK9zEsqh8zyzuc1He33fTxq6RCPVqvvQCpNmyJBb3s18oQgL
kXKbKhAgIyzWZUpIPuY0SWk6rdR2KWoJvenItrUIBWKvh3O6YQoZ91x63HmUQOyj
ar8kt+m/kTq3l8EbiwfY/qx/tnx50tI4d5VlOdXeF7s5FUekOLOwDu+wFPFqOhXr
ZgR1Wqb4mKjRkysuL95QU21ECTBaFLXReBOh5TAW+CJvhztvLrJTtgtKffl/OXUW
Op+u5nWzEjAHfqT28GU/1ld7803QM0pmSv5fVqfeEWSABHUSaWXPKYiPorKMtKBv
2uc6l0XWUhqoMf3EA4kkkrmH34jRWnLtp+WJAikxtWxFbHfL/rEbNbfswrHut4kW
IeQ8rKEdpClr8AVMEw40YLWp5Ws5815xl2hTNe043y1CshTQPYR03HuC0QQNj8x3
AXvcGpTyA1i0DmlhIq5GYxV4nqz5AgqRKG3/XvkKAOK+it2avlLXgeQ7dlAi8cvd
wLTo5Q84xIB1xkhCIhTy0/N8DVvjH0K/8p7YO+fbDYAHW77D31VUR26R9gyb/IdC
/g8huC1nvIRsrDByW16kt4LT7G04iIsAJxAzOupEPcZZ9O9UAWWAlF0F0hE2g+lZ
1K+rT8jcNSriMWbpgIXsBCLLKbhzFhHIUIErelO5QSyAp6hl/PtIfUroXopzboPz
Xv+JU9bV2DsxmHh0aLON6k9cIZv0t21kReRv12ulZAIavt7XMwxVZTGEDZvRXrLc
TMD2yn3dNsipwTRSsmy5PR4V9s3mj96hywYgRB6r42Oo8SpiLvvGb1ewoAY0u/av
Zg1irj5fqbT2j0y0puItggaCDByQbp7ujUHxQ2eBj16dAz1JOjDSSQEAyRayc+I8
DYgsn6VZ1jYr56iEIzo7J9QGI5behxDJDH6DAzI9G0lX0zxtTsljNTPqYL+RYxzQ
rNXpq2HmBunPJAluL5HV0OYTehSa+KjwmohQjTKckRQ417eKsGp3RPZ+CaFSzCnu
y1rTxvq79JR2HRpCkLfGfJSkvRoC6VNavuNQpB3ZF9gtwLYJ8GKAoyie2I2vmPSf
LCQKqTgV6dxpkN5q9osfDMY1G5yUuETRemhV1JXGEVrhDjdKil9d5HFG7XlgtbMj
Ie/X3Jymqy804XsN/KiYZLyz3IrARsx3+VHW00Tkem3MlpUWyWB7lVKGPfgW/40c
TuOndfguLmsuamX+aqdHIOXKaGKajzwkY8WW+xHb8g4O7g/wDOzZwLwpYNn2rlMf
qqpkuMAa9w7bf4Bv45KNjM5zrbvzv1Dpfm803orxdI6gls5UsUUEtyVE7kodzCE/
jKj19XGSsTf0SEgZJJzsjurFrsyEJbfRg0SizAA0EmTnujsgmPyKqceTTqqssSVO
wX8RiAMLvYUvxyjeMoqIrcGnhnLwgB6c0VdbNaLNSos5+RK1pxtBBeIv61FswzzC
NWSOEoYsB8cmyo3DJulPxK+mUSzRRs8B9HBFmD7oRB8Yp1n4Uz1P+UoRuePz3NWw
e83Eos7FRpayZH5Km3sfGv41rWOEQi5ra7Yud07tj/LJA9TRXy3AZgNARQS9/ggK
C+MFKXAqh0WsCqMMZIqnnogwTQuU10725fXueHLEq/9++x+7pNqS1NEsehlPSKKQ
XdNZ2SS7Y22dLj9XHON/Z7RiSDDY6lckjqe7IAybt8UoqDLRXHeTl/qAVgPESd8W
WXaQWp75PxnQpAgS/yI5CSL5I9Y0iBlxfzzNTuRuv1+23/XpME5qs+p2/pu/n5Rg
3kvw2KPwNam0S8I/44bi8l/SsckLx05RbV6TxtSA2GI5auhCHbakZ1j+SBZ4WDD8
kYFnoMjjyRsedOGsqNcOSh5Jt8LE+AFW4c2MQDqpk7sHGywc7rDIlErc8GDxQsuf
fDYqEFfvt7ynfokA6x0vlC0rmWk62JvmafNVUfcyCFTJkoQBlSWkpoMgaQANtcLn
EgBrC94fep8YnHFZuDS7KAqIykQ/G2/E3LsHewL4i58RXBQJR645qIFdDh6Rw64f
xQBu/DzbWKMqy9/Lot6kHYKKaUX+SbqCOMg8hjr4askhFXpY/+mVOYrGe69gCfFD
69f+Oar9BV1nhl13AMwvc8qrMpmKpxKx8rvLtVjfXZGNsWQ2XKQGSK9KJxQPSjBS
suoQ4zCP0RlkNj+Sc2RhHquPoDEBYp1xVdvjwQqnWDTBqkMaFZukd8e3E44k+Fml
H0lgAXunswTkVMMJUdoHy3Du6YEEvaT8c7qy9qtq3SRyYzLijtXPYdYAIH9+eDL/
K854THWqK5S1ht9UQM0iQ2M7U8Cvdd9p2Cf0Adv3p9gBCaEzPu42fr+sqjxMjb+E
FM2vjOAcE4VcgAZCN4oyTRy9Rts+f7wyWw9OxYbxN9A0P1yHnxP4gJpLcQq6yJx/
ublXylD789dhX+XWZt5011tHa9In9CHgC8/SMqrOJqU3P0puvXfDVdxTJetZ7IGO
uUQFjiBr/F3PotagZsh6Fi5Ij22xZ82nnjGaYMKGndsv1THOZiDHfF+I6w+ua3lh
aEuRdwnoDtrkI1USUj7lL9Crq/QSmoxkwNfEsMV50pT6jFYBNjK5lPuALbtePS1E
ly60sbeYgTxuHkszcYO/dVkVzkKIHxb5yVD6kp++tEbcOSH8PgeCGB7Uk/7Q6uii
Ie4cj0KC4Tpd+ZV6xSLqIMt8f4USyHuiGnE06YyiHYVS6k91srSmSCVX0lIwud71
xsxPzYCHnmV3L9QPz2OOoLh+B0MWEXILT7JtzaMFVdOsmGsACNDSY1ubzXxe9KtQ
sDBSMcgyciyhtTAkWzolj+jXR/JThXGjwYYF6o+hKJoahbQ7mscw7Vtc53CcnUiY
rbEgCaOsqX1VxOtFj5/HJsotT8RHnKdkUgfo8NWhs5uySHqENI7xM3E4lKC872Wb
FHx+V1ClCF6HSWuCl68AHmRQkzwWrJbkWlRB8VvSMsm9XHn0OE9V9fNux2sQwvDK
94zB6APkUODcp40ABimt/vwpB6IBsD0fyLmOdKwV2Ef0mRZ4Zr5ON5z7yZ5+/LUA
gZnK47FNZZbk2Y1061scgK4hsYG/Y97gSONTND+FZE823my0GW+UT1oT9/y6IdF3
fd7s6jDlfE+1h1Ul70TC61WFfZDiERcaWDmnKz2Jr+JUUjE/kPZ62MaU+wLh40O5
NTZAJYR0AETqKezkm0sVy8Bt3es3O70IjkJwDtQHKqCo1IUqHoX2ZSmd5YCku14x
uwwHMpz05JwaFM5IdMhN+MBApgSkJ6P3/19QcqLiItrxnYP7qBuRbg0R3tJaSUZE
w7p17tf9htFOSN68vZp7EzeuvRhxPSJ4STpS9j9EWy1Vq9MbrwpdGUJVfUdawwdI
v47NysNYdhEiBdVjMKNY4PNknu8pwk+RnUI/l+RhnuX7rfyXQg7W0zekv7iYnUuh
VxQGlcLWGgV80XngIyWmoKtu0hQNd+597jZqrEs7lHIoiX+xKT5FLCU+1IlNAHsK
DBXFAcYSKLGLop3g9AMkxg6qyJzFxnPnhDOgDhOPRUznAnr4XDJCLontnanxtFfH
wRoQX+copm3qM0wB+jED7uSn/RKEfOdgToBUcmCej1LIWqj1uMziOCaMgDzliumA
LUpX2eOmmtjc5Wb0aMckxPVYm86Bm8Gc0vCNsEPfhf/AdA039gOCxnEtUh3oq40I
t8OJneLWnXzymrXdX9vMIfWZDrlxvOisYDl1l6YILp7jTBN+zzqRn7h5emrt0K4K
O6W+zOYxxlgvvsBYOn4PEhfLaWUAZd8irB1UCwYNYhsRY7etqPb+oaevWorjAnEM
R3sEqs90TcteMhrrpnTyohnbIZkHseSIx0eoS5eiCYIRwwF6OJhmQtFLkFQI4lNL
1FKG6edOlbdDO+T2K16TopDfK/1BHfgCmnrZJa69WXy6rAZq2g3mGOgdX4iDmcPT
WBBuCJNhlPXGL4gZsdrXtczm6Ej+Q/kCn9c3ghnrTAol7udIxGQPrMXku+87QnA7
lkKSUWcy8/GFEE7sLkXH9EBpzgIYfPEWDpcu3HYB7kNKt0L1GftgZbHxeHs8HRlV
u4ExWnNamnFzIfXUTGtkuMd0nOowj3lYBdZGc+LjFvMMM66rQvFBF8FD94dtpKek
wWgIDkNZP2H/TNvjEAhKyLvYqs7BqlnYZf5aYAToIGF1GVBJy9eQkoluCBaX0MWe
JveHe6wMWFdNLlgDVWpqWPY9Qe59zkMVgySlH9I54uYKjB5cdW5sVqAe1iCcuFBf
s4OzACYz/HpmfeFd428A6SS0U6sBjtVckh5BPY+SiUzTT3sNr+4vq7JZ22TP89Z8
+EsgKoy9jRP8PLPIkqNGVtVDmN223blYw66MbclcjffVQyZDJ9kJWW5pvV/wlsg1
Bk4aRsqptlWLLEUMatczO8e8CLIkCYjqvCEcUWLdtFHzboWTxC/Y4yYNWmW3T1nY
kB+ZpXpZaTWdiF7is4l7S1wmqAQqfFR/hDbeq5v/MpVdo+gr7iKsY1oMvbdfqJip
aiJAGg9KqNjdZ/Zj40vCn+XOXC0TtIt3OkHJZkiL7yhvuDw3M+OYqD1piou9JSHB
OJL20f26CALJg/f4YAt9g2UYP3EeCIIx6WudqYxcdL1MHEB8gFyU/0+lJnV4petU
lwLyKbw0HMYbJsO+iNV6OHzhwysv+KNEVDpM6I6S3RYaGS6BiCUkbZc8cLS3Fewz
4QDjYGbUvgP2h1C9NkKp0STdmnbze5g1SPJlK726tVlXvsU1Zdu5PB7k7Qsfgq2E
2LFNFojritk0kr0K6ezPKyHEpWRxCImS+kxk8LWhnj36wwdbutvRQHuNdcsk5XPx
W8OIG1mFl1V6OQvzOHtPKEWu5ET411tGdPW2im39X2m6E1hokQmJczL6bRAS1I6S
O4FQST6xqH9wMxMBlSlTtUFocs2xtLxE9DiB319TRCy55lvEST+mYKiWDTm0vPCJ
Cq9+DvzCI6J3w0/2rUW/67Tb5bDZzin221keINtKHBzjiYbKTtvrrByg5/1oaS/7
8eE0XfwnyVDIxvP4KFkEwBdSH2m92UXFRgBwb1f4ZVscqz44i9uRCc9TkzWpBR3f
bTa4cH00EXvVjpgnr3OQR7vrPZiaOqn4Y6U3h63cBcndrd21HqBtMwDX2sbc2nsA
mIKXnHyCq8ZbaJatEO/L6tg3AYA4kssOWrrYlwVYxzGOjEC16Y7GXCxqiN7ol4rg
N76I1r3HaSlWbeQwv1zuUK7KwTylfUUCib0ERFb/DINVcZmfgza8oZkLDIz/G3EX
Y05919Gs2AaE4RHZhDXPQsmcwMR881ZibEi0U6SWW8G/x4RQRpvrBsJc9En7E/+o
J0NH83x1FKcjcuiL6vW9qsA8X1K3p1V4s96UC75tzquTWp2yKkKSG4McihcCV/2X
lujlpdZtg/v4QQj+PtljjOrRr+Zwi22Tr6v6Z6p65ubZ6ccvje8g3QO2SICHc88E
00/S5XQ6SoMx4zjqkBStwva34vSOo9t33mKj7DRry4i7qCWeomUE2WVeycdL+ynl
+cHXg8lmQWFIwkR8jzSLL9gG0eAK6OxQqHruEtADvEHDWHODElgQvljGOiSH8+ar
lAL9GePRsXVqKCmeutIuC6+hgSTxtYtINqoZecDxwoXEUppcrK3/QQf/VcEk3MB4
xW/XHk6GdtuyoSoBAuoUMtn5ELeUeCdCZ2bDFeb2NlJ4FNpqA8Ub08CJRWNXfY9o
UyyMqJuPy0w25vyz26n6KfAlGZ/dXE/gfSFWQgUzsIT11quTemZD1hgxYJ+B42SF
fJtaZDixQ8j3Gon4V4O18x/5w3fcVATJLZTzMRkFILs/ZVc/yU2zKNrLnkWr/uby
6WmJNXpcLmG1slyPh489ZGkSLs91Q1fKlRGcNKe+80yrgQZnu4/LU+d/bvCVrl40
+j0BLRcniHxXFiHd6F4mcehtMby5k79vsURmlibXJSIPqjKTHgDhq6LgGjtwfk8X
a5sxwEnykcl9VJ6DODGkaoQ6ihYO4+xzRmhtW3HI8QrGtp5t56CiBk93dhF830xu
6bG4Un0gXpVC2w1vL9B2uPDWIAm6TNyQaT289pFVsOvGL/T0rPjbuwe3qvxF1hRS
7L5E2ISkpPmhKA9L3HEsbNbbxsVq7Qf/JErDStJ8vsyRsJwQijY1TxWGj7N/FQMg
g2TPwaBzjjkHjDjWcXh78jHb+y+bvx2N1jCq9w8qwK0UCKW+g2xvEMEOU5XhUkic
kgdimV+f2fZzSq+rCpsPPPNTu+fdF9d6pSZB967BKPcSzTd0C/T3w1kzqI5jBzsa
DrifayofO0K7BDmh2mkgIpZdCJSz17rNkO6+k5Q9bGHeCpomQZDxasPmXe6tpyZu
Wgylj+3/9Q+WTG/uEFlWymBstXGp960GvJvDgfV1M1LhWEa8Wh1ifWKZ5C+5bY3N
XSi9KP83C71TnbL/XnvtFB6BjRzuG7Ah9ksu7Bjmz4ylgAgzJA8Vs4sfZeHS8D25
QYSJnrBDbba49g0PrshdBiVG8zeo0aZV4PmGRCPJmGOJ4vCvTM3rzDXM8GghtxTw
C2yKbdnz4LlBgEz4s3Z1xvBGtuhNheDuv6PMHNllxu6iUR4JqpOWRgKdHJ4Zj1qD
pp1PE5dCjPpCdrrDOfOtY5AedfbYq9iGu7VuB1XDxdZ2jmj14AmfquzgIstZuCRX
TtQkW3aRxhBYVGDKhOfvYnfhdmFhUBNVZW7+ozpDfHj8YR0NaR4sYHrzOydSvFpw
ki5vIlQ1BLYRjc8w2iDUFNO/bTC9AtxqyU76FBO9iFbAaenKWrjtg5fYbHz2m3Mf
KkCqN5qbBwp7E7lJPK2lYUAv8qBCp2yXNRv3juB2VGnw7EEbU8lvk96le7ng01ur
lAt4/0CGp7+aWAU9IR9PJqIo37goy5135ksG1jxCRtL30Ompcor585XHnlUja8uT
4ljK+xfGhrIP6tumsIaj4gnrrw+w6z5SBdAxMtlhInJzpruUBZvbkNXJpXYBzErt
wgfNOe8FxJ7mzjuuHlzFxKyCYVsvN22OV527gcu9eA1yps18Q0G3FJiFR2aLiDUV
e7jWPaxX3Yi2C0zph0EhVcVfc3M+OIC8bGckdLi/N+Pu2mc+VvC3bjPQrVuTp0DD
gi47Qy9r6jXSU+3G3a0dGS1zMYbeJlKnZIOfOXysOwyTaDDRxWura5xOGg1iiqtN
nsa5CJObDSZA1+umrGQAcj0tWttXOyiNGWD5WcqpwcbvTZ3df57rWuMPq9ADi0Hc
+aY9O845NRp9xQxoBLNPVXSbNlmGB00kOcjx0Z4pC/TowIceU/2/mcFrTGjbam39
i6uUAyMMpmL5WIVRjmIYbB50dGixsGvnMXXaCzdhg+V8ugYS5NUtWuoxu+upECas
UVguigx9lsY8nIkyuwThmnSpGoJ30/Ia4lCUxLCv2/GPYtUJdYPrRKClTVFy0061
eC9JrbeyqFxn1MGaARXc4mE5l+NBBOruIag56lYXSExWAInvkmiKXj7s3r/aABXX
tc7V2kbZIucr47zLL5ibpNAPPl2lgJ50uV52q3dXpGMcdiI6VAplgNbDrLbY8xnX
hYLRTqZdAFl3lX4hWH4b7MNSKCkymBpQ2B4Xp+kiJ0hpe13HCRqgs8cnrNU0ScNY
c7YppxFlAOIgljG7b9haqce2eGXuLwzWN3fk7sMGCcJrrUh7Zjw2d1MQMLTSZcH1
5sFgpF+3ZJJ3TlVqVlXaWcQT8sdt4gaOe2epxwFhc75jtWdYktiXSoiV1eL7oDZq
OnB9a1XW+UqBa4NDdWN/rQqjgRBCrPy8pBB2RyZnT9oHwd/aIXOJBVZ//lx1QpWj
/7VZaTbsuHRahMr7n6f1Ck7kjWtBn6JDH0dFCDGNhMoCpKrD+Yq82Mrve3LRrNMR
l/nLCKFesF0JnCh0FImE9VgFxCEeCWzzKjVJcMSRlVbXj1V685p0WG+EzgZRohhG
8Ls1poFcEk2WwItDrFsGftbwhWpt+BNOw3HJIvBLkzgmXSdRB5FoM/tf6ZR7F7aP
eApQZ/OTOu62wOrLs5opITNOd2moH9B/A8tsaHwi+IXY0cZEd9vc/zgzCwTzgNrG
h08azpQsE7+DZNDP96O/h23BxGnPhZPZLYocRwCgHf4P85ZvlH/pmC/WjhoJQ6Kd
cg8rFTOZ6/bpEOqeB//rY0nBqw5oqWch7KIPWF1wzY+kHdpQmNvQqCPpauTF8O5J
PiXJngHkZYqf4zih9S1OaxDBslCJo4keSWxQuAMY8xrO0nSE2TNSe+MXPQsEcQFw
27t8ykTMpnHkGRZvKGMkcsSugn683XQ0SBIIlpz5vrSG9HnHeL0m1ES5ZDvBSqKh
DhsOJB6NpRCgPFnYzaAV7nhEd5YVNLclc7CLfC0L04tu8IQIoqpDEOfb/DLLX9K2
scNg2uZVLm1bLhgclrgzdRw5OAgGTHQff+rmwcatlI+9PYf16U139J7P47AB5FJ8
I5Wbauzt/bJZESP2U1ApzJm0bSW1XQCzEmG+0kbejGIF85ion8yjOjNGKfpgKXBH
8VQ3zYc90Rn06KyKM8Wt62KckoNGrUoCMm6gyvOw52gz0PnrMbCsyoLDsSMWZOMf
HpkNlt8dA+sQEuZoWmE7GUDgSarewsSkZF83aD1S/if5G+noMaYhi47apOTfMeGw
eVItlk5PY261NzOoMQnT9RI4Xp07rVnAcIo32WpVOth7x8I4YKfNVrhWuNMoltLP
GFehKB+ZOEGn3o4S8J2blDLMqhZUCp35caH+lApcleJIvvhqSMtn4ic1U5AHn8pX
ioYAcOCVg4p0AA5n1kjdlslYWngEFLGiKbK+jSREN4127uhlOXE/5Sx8hLMCcmTh
tGPoPC8w4/VZzJ6aVIRvu6mRccB5BCBTrTWRvQe+5fVfEOgRCuGIlKFdJrS86oum
FXvqfDQTTwlfQ2/guthIrmzdbCNPN+YFlCv+vKchMeTIK0BrUNxfRsA0FvbZBDKf
jGek1LgotLgUEexk03av+uf8vmveAU4WLcZGJuSIWMWg0/FeTRGqBjD0qNh5xDmK
XjhjPMmkdAUuQrLTHv+K4sMCfmVukkFBSM1q3mWvktXfbAX0WZNLfEGrO4JCZSlE
XrjYVf6qiwbFkHrI6H3GtYAOcV0kAvEPZF3OkmfU9aVFPTUcbOLfElMMcHxVajVV
/UnWNRpPLlP5xcxtm1czHQhs+/hyAyKvJI5t2VBqzx0hp6H/5SuRyOR/Kt4knoaU
Guw8hhsezAKAnmVWUE2hG95s3/eGF/G0xXT8t8NWd54ai1WbvPZYlzkvIDj816bi
3KupOdSIJjWUNSKYU+caWLyMWOhaqXcoTF3ylU4rY1IhESUSOvyZwD9oR5y+Yx6L
VTwFy6+M2Pleln9/ut74lNSaa//emH8q6vTsrOe8BGGvhVavYPYL6q9AhfeW5Fzd
o0JdhV5fEUS0RuZkmok6FZAAJTBTyMZM1V20cfZCw1MdGzQRPMS3gog0WJ3KhtP/
ADju85FcB+RstGfwiqkUUnHb7A21SL48YmU3Y1uVe3zIjmpCnL3Ud2yIvbt2FMNw
nR11TfalmIP5UyrGIomylkA1kL898HF8mXQZX6rBX3wK6zvHebfdULHmkC3zVcDr
BtPTHewEKwrEP9y+BrJumMSDOhqZ71s9ItIMDWB0WEJ7JbPTtQzGy0nrvGxwSzxn
wvrlJYaadLQuShtN1UsESnf0viroZP7u3d3UsblmyXCpixCajzqBoiT/lbLArLfO
bCAL4n3wIguNufnq1MBrnt3tu4v9uMudxz6OlCgcmzbSCDoWfU4BEgm1RY3B5qkE
sqYIsFgLgJOjZGxeajSoCL/EPXIWui5w2JVPHqZY7m3Ig4fuWZQYx076YXorqBNP
ozkXxX+WO3GLBx2OHcMKDGGil1GKkpwn4kmBqwmDvKU3KqvtxsjYN5OrGAn5isDM
RvqE0yvd0OZgofsnuZhOqptxOt4MGhwmGrhahFuuHB1V7bnJxylk0/9kTG0Qq0rR
5mPctSIOSIzQeVbOqFCDVA3AwtGtGVLteL2/YBaaxPtWBVDDYKrvW1/bT5D5//ga
PGvjdivWbekW8UXsdSDfuBMHCM93w9Ecggwl0cF/6vscjQ/TRsTzOF1uYIlHPT/A
iJWhMuB2DI7rRPN7Q4GmEh81GLUlC8lIImN/xHrhqH6YBFn6k++iAEuc4lRjapwQ
etfOprwZ0Dp1rezQJp8HNgsSkH7sCoDl30bmQoM/p73UWPVIgjZuXvy04yeXWAz4
KpLGt7lI8sBgU/3T/JLiygQnVOxeSxfnO93lz+Co2yfPlhL4IBlmMDk6CV3T3rOL
OJqpzjob/fYi7fW2TNatPzAWiN5yjSWNr/qkzz5QEZIgnnsrzWfeM3zGsSZAZ18R
HL/aQ1GeAuRzXLB69zuzXQ6ouamKN+VRGNejafIp9LcCXCpxUSbBt5G8y2jJsuW+
j0WXZB+heZzlf00Ir0utgVt9IwIVyX/WAT3yYBcEBR13Obob3VpsajcgF72aKi+9
p6Ii4EeGcBCAw8yKXPN/2l1Expy198znVI8cyDArbFJUA/pUiTYKJFf/dVgOJ3Jt
XWVU/FrtuKLxoz4AjjgZaoCYlfMoR6UMj9Beh9eCU8FyX3Xk5T8XEEpf+jBgXha7
qSZUF6EBQPmbq8yHJ87KlTyktXz0bIloRoLA9LGnO4Yk8jmZViBoHdADFdNJrOil
npb450/yCTJ1PuLMjC80Uah/3YNbXvNqhgeKtfTCsCYz71WxN2VlRnViYaeGvbbX
dn4Np0lNA0Ofd5cIqOej/7Ot53CkByvcUYCIu9kOMNPro36cDTw4faqXO2Zqoo0E
qKCaXcCKIU7OiHxBSvxkExidcJDjRywzNYB/Dwej9Wqv9NlU+igCnYjNRU3LIfjp
UtwHewn5QugzbZlhHT3ds4b51Xa+Jy+q4O82pZ1guUv6TJOTxn9F43OdnNyeuRrg
mHI5ilI5Y3Im5NC22XqEZPglp1Pc3LGSSn6YLGznGUHmfl/TzabWaY6dDTI+gacA
zrLN/lk4STtwSK67dAm8+lz5p9bObyl2/yq549xhAkSbczNVcihPtRar57biCrcn
1PWxWrxmPfbpjqQlkDCiFfuT4pbOQj+b++sBHUQ4TY35Xs+SENbAfNXn7jBBH1wg
b6Kjs+xOsYQX8T3CxSe5Iw/Z1TMn7byHP0CEeN5Noc/R0MhpogfdT4AQBtOsZDeh
nAJhsdkz9XhOjjXhYddm6lJs25CcBf4hIrM391fQ35ITzQMrI7iYilwu42cVWV+D
oaWWHEWoqdXK23jRLoCP8ZOEiX5YI180qwcCHOL5xrYbmcWLE7lIOyUBa7+0ByS6
DYUuwTGI9Xfjqq2//oVUpHMrPiIV1FIGnGHZ8Ky3jw7ijCau9hFD66Zx+sKMmkn9
w3gtXYSSbLBlDuX6fGa3KyvXFKKrRm6NdEAf4L39gWcZotgKhMpPkbA06fZtw/0m
Jk7wc2y2YI0sG0QZAyL8PKgJkDZRZR4xkAaxSlmjy+seLwg+OpshMDGCV8SfaGoo
LXVCiJdtH2VC9bzeykYFok3xG6wRVsWXULArSK1xHIH9bMbDSDbkTfOE0nqVCVf2
VPh4Js8yyOeDzJS/xx6+EKhbvP6KVoS/PR0r7IhtGM9VA5G99o61hkvIGITgN182
7mJNJxZ/orQkrACKEv+ouhH0cDQ43tCO+OfUIN/mPUw0wmZmoYErHIRqX7Y/Pci+
HaLMV6cccJb1LFh2bKZVF/U6aLHR5OK3SaaoqPwOYxau70qlha5vNY149YQ1oN7A
nQy61bI6ZqB9J+m4SsqSGi3vXflj9P+trDJrVU9TYoonGV+Gjjcfa1jh6R5l9Qik
39ouYwzWaHQoqPQ7UuSBggE9oHdGJnz1ma4dWrMnvKXGzIzRHL2aYUbVe1MLZJJI
oNeLSfIfLtSlFgpjVNYV5qzj9Zv9QXUiKnK9WAY7QQUSsqPqaPyp72Hyayxgghc0
Cj+KEzJIRWPh3ohQhp4insJLZedm3/0l/l4vRgWFgtYgfL9rEVep/35w7YgWGuRj
QYWVdbdGsEyvkxsNjR5HDFSbEtGZV8tm0VevguGvjvmj7RO4tuEDF/e0N7fyONKc
Ci0RneqKnAjJHvMOF/N7b24DZ0BiVnuLUxnKDNuTIXVuGOrk8nqiW4WahHQRiXwO
GR1F4WeJt2r+TEparCJBQNLitCwGiCB92VqMDwAGvKDlT51F/JPDv+Gh61KDAHo4
AiPF2a1gNYWwt1CFd/69KHgs/PMNPus5SWw5jR5uXBJjV6nVBy2sc/uJ9OdKbHfT
FoSmMhNdv05J53Bc7+KKjRgcgXcLCL2ByfNxNuK5Z/4Jll3o4nn2sT3rBwfsDmwA
t5cXN9g82K8l2BA/crIE9g6xNSUhIaGgJsQFp+LDIqiEZU8HAEfH1gn8BxUj2hqO
CoC7v1cd7m4PHzarQJf1VxJJ8zTKTbqT5OzMaIrvnHSAePkL8gBofoB620tUw4A4
4G0zdlseTCIiEY+dmlq89CSST/zL++0P8zKwIIHJT5HPkQgSsqBsj3bXShfm70gT
Dgj+IB/DD/lHw58pWplsCbaDlTTbYDTrNuGZuA+sXVWNzhVpMG4kAlEBgv4UbKKL
MjwtH1SroscfZb2T7+X2EQys8vE1E/jDeoSMzG15R8gv3U3Bkuh7SblX5z6Ti3oc
GUu/lBsOlDYM42X40CE8CDPMb8Zi3NX7YVdxB78vL95/tstTaFO6bRljRA+fjZTc
5Wcqs/jLdSAOFGFDmV+/RPYor10ZFmqDb0bhxH1CrmnIRQKFjprqK+Zhgt9Yx6mR
hN/W1PdOTFomEG1zybXWrulU5yhnH4onZOHHkGRr4VVisaF8xX7xlp6WN5MxENS6
RhhQA8gk1wvvq7PnSK+XujuZ+R61rsEdAcNxNmtO1ouJurZfxlXBlNggc6arI9H1
TryQ6Vl4Q998yjE2FKi/VMNjVsmIdNFdLSX0cAT60ChAiE8OOizTc9zZEWvDCZ5g
biHq224wkdWZnkJLU4PPalTJqodsj286u+Omjn3IH8kbnsBSQwV4O8wi7GK+XKbE
sIpqbXBi4gpfw5UbMptBdtcXLEWp7zTj2azTCo6JppugZPq5Hjo1UxEjSEC4iX+q
brFOiTNOz03lAElE+cChJi90ZgbGYoqQIh/CVj9JhlxGFU0fRXZWyrPLcO5GStIR
TC3shNWqTS+ibGyHd/k7VfieSon2VcfwgMfqABk2lbf4YyDMHtmsABJVPpSIKuV8
J7FEfIW+ijWmtcare6zqmx7tJeQYX8EYMt8bHe19BbyT7DHz3XteW35P0eiWiKh0
Lk3wTxyGj7T1toqHB9F9Q/o99GhAi60a28mF/uZl4ybioWzmUNvsMHY5KUW7EE5J
xFy8oKpTFaP+TVu4xqW3pzMupM4Qw0d4zgpr8oYOSF5SlWM/vqRZGnREpHIKlnir
yk79DAYVkFSwC7ybjpUJ7Rg5NTmGgJA6lmxbSTaMU5+LKw0iK6Hf+06ZSF2f838f
G6pAUSO5pDe6qrNwAe4s2Ze4Y2ahLrb5Ul6k2Nl+rXcN4vACE9CX6HpW0KklsM2f
SjhFz79JWUct/TaADgtL7CPIWQS8LlrLAgvJ/jdN2R3H3XQzeOyW236Ke9wy//Iu
6POl2LaE5TXkAx0aZSMs3/mD8UrQGeufdq746aUZya3K9my1/Xe7m+YzLJlJyVbM
MWujC/r6qdxHovQmq1gjeVRniAluIOTUDLtCpkRDqelJk3SD1uc+uLGUXw+AcmbB
D/uPwgrVu1lsuzb/KMAOv+p6PtyMw9jeHJSe5c17B7QmJxAOpKA5UyxoWiE+9Dmt
o4mYrRiW91qzDPQn5eMxJxTvToZTnjt2OUPTzfTvW/NxYZ8LN3uk4Lgeaof5o6Vf
nePcZWOvkTJwZbBdfGglWGlyKFU4vX2OjVIXfxMw7wFtv0Itsq2mbI3KeAHLUwaK
gHDDMEuo4rY5qzRQ3WK650vUO6rOJd2bpIk1XZoRcH4FPhk1Cmw9reA4jAUq/sZq
eAYNcHeDElX7m8i6Z+/dlOy6fWR6T1tPHtGwedRqjanK5NCAzvIgXD2i4BXtC1lG
SjAWBpJcxHXUZAN9FJkPoAgIrbQYKG10GcG/efls32MGKXaaidRsxAfWmFofwSFf
anzACts6srx/TutJeeu/lxRj46Q4FulZEOGdlnb8xqN2G+LX6qKu3kupiKR9udYD
If/HpnD5XJiXUJGa2mZvP3Cw+SLppzl5XP97h6sc32asGL7MZzWYNhMf6DuNjdS/
Zngyn3TGntbcK+wwzP9gpIgFRXp6vHYeAk9UdkBI022G7e5DT0llcLXymB4w20Jg
XlbcxUGl9pEYicdeOxBccg6XRJXDjFqU5plwnXimF6csdpVj0x6YL7EcvZV0ciKK
kB8jYyhCVrDU363Ne/FxrHgBahOltQglP9XP+IrxK36Spu++PARjkUlPGSBZZ+Mf
g3mDQtZUJknHccL02OIOp63+rtrnNbjKoZbJoCe/RVyrEjI3IDPAckDLMx1cWfGo
9ap6uSN8ZrRdiZWqJixm3zOa8gC/Cjxq6qQJ3m1dQfncDP40XRZCTh5YqD+aUcLs
VD6QNbZspfcNZFId4csaCter5BzkYoNfneVHJc/HXaRXfH3oTiZYkt3zLCpgH4Bm
6ylC0jSsmIKD37CvmCP7uaTb4bcBBmCN/jeSAtOblFiTKKeaJCGfacRRtcyobncn
F7dOdXHEcTuprQRlS4YAWiTRGVl1V0RUMwudWsR46PMgVprw7QqSp7HC/izUv/3F
slzrH/l0yHc2lvM57hKzBfzQ0RqjOB6M7lP20iCIJkcW238dbaXPv3z5toBVb18f
Y8FpwZux8CpXxNbkzhzo/l43rfH0AUs43UTsYJCBmmJ7dMWONfnJfFYak3R8psby
GrKRN7wGVoccxjE92JPeDqrzxcB34mRAtNUmOAe+dWxPsak12rF2n3oYV1fDge4D
VpVK3x8zFCtGATXk0dqF60Rx2Tl2mELse+CzKrXNtCj5/rJ4GwcQoSjDeESlPT8r
wfCLy0XSGNfE72gFLvt6FV4a1AfU14Z9BIoRrmmGlvjV/OW2USs2UXaVUkCDaXeI
P8BaIiy+bkxPk4R2PQbmhTWAhww9zMsvvz3WxK/c+FEy69N7QkMPbUb7+rZx/noJ
MaumQVYosqv/guasRV6CPTQC4G4M9Dxx+8SkSBy77KZBvVim/SLbsHUsH4jbripq
8WvwqXPc4gNPBpmmRAegZEYYDB7olEON0MGOTZRNINze9BjNK5a+X8V9E2/R858q
ih24eJy60wjd+iM+KU97mLaRLLWv/gtPGNhoy1iZNhpvRgGOCXDX9mkooHXAFmKU
+8bMseIAKAbQR6xUY09Z5QpdiVOdsLmvcl2V0+juwpbxphJxU+qFcLlYMMTrJBZt
z2QH9Gp/yOiFGOdzz10Wc0Njr4ZgbOCK6fU3Mau2VKgzoivwnuQ4T6wRtgwp74zo
8fXvN3swci3nyKjFctSywk5XOFMmW8iJzUkg2pX3fjJAp2SZBiskwCabOjD1qOGo
YQCqmKvq4VWEPWNMwa0zF6VS7ElwY81rx0x3dzk5vHJ11uWWQXLQm2RDqB+uzZYZ
wCDHr4boUzTrWTUOh0IjgpiNtfcNyZp1aw7j64Nk5btvm6FSj+h6xKo1yIHYAn99
DTUZbDTzqtV99tljBoIa/OmxhR6VkGB8yrH5S94fNWg+Sj0wp+kvcgBLP9Cj7QlD
E543xWJEarGdLDEDAf8Wz4tOvE+DhR+3APYZTJCrTJnyM72ErRsHCg4uc67u6U71
G4nVggB9Os0FgFt0O4xwbWb1L4lRn2e8A9hoxvoPYoB4xTmHZ1f72yDOhf70biOq
OR2vCvNNpjOg7tk4oEzWK9s1jcESCJ7Wc8J7acqcGTh1tHrRgPYXumUoeOeU+GtL
hn8QeVvKyEMXXFFRXyR5AZLoMqEwUlmguwUMAQnhoZ1Xuwa4BVUDgJWse88OpqvU
klBaxzp3hKtl7KcpGzui6Pi8ii8gI9Hx6510lHxxEZ8RjCHQjZs86fqs2ArOi83b
juxTC6K+vEjdUoFdMi7w1zxIvVEHH/AlGqTo4kSnCvr7hKFiUY6Wzlmw162LI1lZ
Uoyl3lU7WYKQ9FV7t3g7N2pM+HjXUGBs+BvFj6I/+F5oicYvzPpWJgveSaJ9lvEj
NbRdbFOmz3gWCp4BlaVxwoxBYyBXsLTkUIJjLfw/UvlEOlSItz5mQlZ6nxVvAVUl
CLVQUT+/BSziZ7KqsR5QvvT/likT9GYMzNI4aP8H+25+kktyP2fMgrYbt/IqzCgR
O/FQhQG0pNHp/gAmIx8BqSvDgTcGdS4qWkAfgdiiXWvIsXTVvPNbDJwF9cG+YtyX
8wc/wDKF5S0BNeNvnTFLhn6YghiJ71gRhs2J7UARdM5hSZcw9wfR9W9+TbXo9aM+
hBr6U0DTv5UBrfUce316NagphG/hhlCGJhLKJGXI85O7USFxwWIztXp5/6LhFEcH
Nu1rwOSI5AYcootm1GHaufP0hSOEX6IFhYQSJr9xOCcCV+hDmhIAIWJc8QdNw3DA
1hvFpORksas6pY4uh/yEOcpJUoxYyVoHMmOzOjFjLb7GBiMNSH278dKSALUXqtx3
/4HWw1DOTzQaMZiD7yCJv2B2ShfZFiUmlO24nVy2PhfyiDJdp034/vXxwGe6WiU1
osWC84s7vb8XdghIGEh5PqOI/YiYcdjlBB+o9YTG8fprmP0nXF/bfX/HrB2sekFM
4IGaRBrV29AIODRsmg+grGQQaPXzQkRv1+GyC6qZ60Uvjm78xeRufgkJW33qiFa2
DXo8wanFDSmw2IZlnXVIeQkZntnA7YPCOlasQcKW4RULsw1uKCvZRQYZol5u5isX
UNY3hYmZIT/8joeLPZ2yep2/uS3UzNrMDEDVukAQHewQPkMLsaIR3JTnkwrxfcwK
5rKH9ytxvJwvGaPl6PhT2XgDSK2XkU/5dwAgN3CqNfWpFcU4OToF2lFBnayfF3Jy
jE2/HZPscavOE1y4g0ZLkXn3Dvl5HE+fWtlDcrJa24+Uvf1obBh5F3rfYTSx5esJ
iYXS3fIxwuQ/X8Upl5YfjD3mzXcXUigUs5d2zbH99Ra6as89YQ93scAi+POqnkh/
nK9qajz3FXA1mRbqLQgm8hh/XqIGxtQBxPdoi+0mqNVrXnw+KwdSTWUdGk0TMY5S
3uWPPqpgVmnpEWzuV9b9X0fO+qmlMOOBYvW0BHjW06kEsql0G244nSpM+7xakOO0
WFu3vJmA3eYhySQiYkRUcju06cA+r1WaB96d6Du10rgyPSUyqzvR9e8MamaUuPDN
x2bcIEDbZVhD+YWttzjB+MgfPUwvOxBqTTWris/EuXGHPBvfxZ0bMWViLzODqFjs
Ny5O0I2hBKLCwCFC2IrXR872DTgQkK+6UoftTX/WkCkynSlcqqk94TH+uQw9rzEE
J7PqsbG79Yv9qR+bOC0rDs89Hkisf+NyC5O3yuzdKT9wtS8i+o5r5+gCZuGe3EQc
r/uZ7Ld3AY/QqwtmdbtpGr5IuuslRdFYix7XLHKE0/LDKWdwE0zDHa3BMOoDb+8x
Swg8GbQLGGKmBImjx90rdXKI7J+hp/ahSvmDMpvEzQS+W/wYxwukgyC3Bku1fsOV
bA1mtW460qkACX3jrgPnEuD1zcbAPohVraJyGQpPDZhVcr3jf6Vp4e6fnu/AeeoI
Z9d8Yv6QKr+mnKU6aRDTZ0jvlbp/ekOtCVwtXq0JjW1cQYo7UvNzX2o8HQl7psat
blPeIyQCGbgWQlcebNac9DzYXi3YBU1hbIGpve9254PCK6CD3up6Ap2tQqH+raln
+3i/0KQwcyj7PfeDzbVTgKP7BunGXyqtcvR0cLdXwFAVHf4ub2NZohtOtsbDEHFg
VI3UXTHgwL2+gFmEieFg+Gl0OhjnhpY2YHhMDQac2G6qXYa6irfzgQ6Hk2fPnbAv
vPScIKv46gPQsm8ENQBrVKK66++CjnDUS29p/wTk/Vrkhi5YCYwWMAwjZjmGMag2
qRQC/cFrCdxPLuFU2sGIXCoSqaCuuGqD0yifxMboCaMPlETKT6j58jObLX9LpJSl
/CC+IqrcvSGQ/c5HOtRg+mJHB+kywNE+mSauprY2gs7pCU8QOddXYmdLDC/AS+TF
G6E12QUkrGEty/tQ/40jDRwJsTYqAz7a7YApzfK7uKVpaP5QboI38xM/4f2JMnf1
mB54OTPFreoi9Z5tXhYMOckKpFwlMzWp5nqH+HD8Cw1b1Oex+w1o/cmmkeG/tdjR
sjdy5b8q7wp3AXuwlExc27nL9iS5SBsMHc66fvaFuowiUNy3CxbGwWIqS5Z7/CpK
ELsdUkbWbrNy41oZiCZQ1DmrTxNzkPvvxoiAo6oqNTnly4eCmuoqxswr4SgmqunZ
cvbE/drMfCM5PCRvJ3ktq4mcVjkrgMqdI21r0h5Bn1lmrsKXamck3Y6jImBYDdkT
m319sCAZmc6uZqRv4d90D//D4d+8m/d+S5lcnbCon3ymZMMQChM4t1VOpryRuyrY
vy8qOVT0Bd878j+KqkqxbQv2XIPxrxqqGhhSGU6keOBZmiSfwMPRua7naT/PnJMd
SHgJVfKV7qiiMZ4gG2c2Ew16nH4WUprnPFwaja3fdEn7VfKIMC17iXwCLJf4VhxN
qPovBcztLAX8ThZnyz/UV4LGK3xtWFc4NnxxUjBoXB7rA962rBoZorLn1NexQ+M9
2i9/zaE9gY2Rbx0IJccc8w==
//pragma protect end_data_block
//pragma protect digest_block
4weJSQH2GYtCXUZXcjrrvtAb7io=
//pragma protect end_digest_block
//pragma protect end_protected
