// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ddbwliA88HhxRlB7rYO5hCuXAP9mi6JySeC4ZkVRuufK2biCDL/AyiSwHKDMKaPJ5GkkAwQYYlPZ
cN2gV6SZOnE0KzFnpf3l/tchZPkHzILnw0h6a2swGfQsnM3GliPDOPtS4DLiqAVX8h+MsWuwzDPy
pEi6tu23EWG1W7Sl6C1gOhzkdl52ZH9sCmrDsPq6oeIn219f/Mo6GNE+ZBcnTyffVjjkgobObggo
iYjnViU4d5kjXrkmn+VUU1OhEJHQA0lzShwycAltLiLC6yjFAN1poZFsjQvdtGZIh9B+P6oKdgh/
FA7/ZLo2p5rlsS71oU53IJqoHoKGpltMucjHsg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 54032)
a2D5jfh/zO1RVZZHZy+zqDUyvsjiAbbby9EIlHS6Ex/Mt6F7YdyViL51lG0/V+maywA6Ecz7uB6J
/0mekn+oScmlyxghKbmZqcJwfc9AU0v4JSBlc9e3tlvIjYVscncVistLEqiZIhRfWG/B11YdvGOl
v8+N7WUZMV/w/J8MWFnh5Tm/E+5kPa6FCLQ1DJ3k9+4XZutbmlHuFOGCSNjpHwnlR3DbOtiTJ+oA
94/B5CPIJTeVgLVitOWuUNSy9S6nlIrGMA0ETWajeG04ynXYdIQgB92V4iKmrOwnQbI2gAsrFqHD
rIdVQOnKLngPBiKMCzB5EbKAfh11uiAG78QG8+TMLq0r1dJD90zSeleFzZJ1O9Qy4q0DLCg0mjNX
E0ZQbKIC3YYgTak5/XD1LwBnqMFffZVFgE/I6Kt1kpELHb0r4c+o9EITM0fZKIQ/ShKJuzOaq8ok
njOTMn4HQIp3w/3I7qxXqq5wIaK89sddX5BEp9P+h3lBKp6rlKyXLcZWBn1roraHfdxyHf328moc
BrR6SIkOAV6bO7arMrv/boJRahMYUsmWO2NCeqEWiUUYbyde59Div4xVI4WG8cGJXxx7YJaIDnq1
I98d35uVdolZ/kaxbGNKZSQRha1siwf0bw4bWhNPEJ9F39jUfpvrc9qAbGekqDy5dy1oOJuJxRqy
yzIUfcDXJgK4NPs2qVZq/R756U34d1u6lXdI5yj26iX4x4JK+w+tEce9AqonvyAHDVB6GU9nXtCl
1xi/SikPhO6vmKW99DiAKu+Fyiv6c1M0BJYH9/s901DjmZeUv2flpTw1xvAxaLEPGFKmpxG6NQz4
/SEgkWtY0vZ+iNR9MlDjmTE28QNi/zec74wZ1c26rkO4pgyjLAButHVe6oAg2rGsb4MZX/Oe3XtH
V4JPfGn9LDTvG6NkJlDOWp8nr5fTuMEfiM8bmRiUEuVkX2G1Hh31/JqWKLjcu9JOdSZPTCiR+cfq
CqRGbzrVn+pre8aFkF4VOTCSogb0zJTHmvSRdsAfC0RBboKtxkRoR7ywtUABgh1XknEB1Scb3B57
TBrwXMc9BTVoc5jA2fKvE/lcehqhvcpIfX8FyUfU6YyzIOxaKF1u4uMun3i8xRqEJiQMCnwKoCWq
FWPml/49r6xIgMtK3DJAwQ0A1CPKFOLVOBeVkpAoVXnTYPnBEQ7Vgv9o+KoLbcfwOi1H2Bd5Gp5B
2SMca+2QzHWHrTA/lCljo8+lPL8KWThCIgDieIqS9La5d6nXO2OeMNNfWV7/woql82u4qcHAZlwe
D2Z6FRm6eW9vHCYReaT2tFLS27rBQMqDU3P3rosg58RFu/2H7F+HIw5hwLxHMem4kyFan92WZICu
vlhZc+Gda+99wAUb2clmF5Jz2+dQAr5vey8sm3YduXLaCbk8M8FB1S/HUgXo81eiPN3ZiH3qp/+3
ukQqvQdBa35garCZ/l4jqKxZEnQ02dsX8a19REjc6s813cJlTEuvnsIO8zEXfdrPSy0R69x3JAYF
taSjoUDjItgOBEyUAoL7pExbcZDq/x3B7tBIlrbKykLmifozPGFUhJi+DTC4cddo6J+UIkcqzR9A
jZKuhYfziD15KMk7l6jEJHVqnJCYsoO7sZq8W4NQbJy81No6NefEgXhS48ib4W2WRy1jmZvX2gvZ
yfwxJnflzsBmE17epuHh22EhEXpS+613dwS9DPKJqisi5G+BU9MWhv4Od5WRB3Qyz6ihSEGh2D8j
0SYltVa+9Bot/VEdXfKDZSvhb4pe9vykjHthG4/3DKSFViYDsjQmVVq6utX8WhxgdJ0cA9bYuRZj
jE9cMaCQt6ItpuSXnUQaOlwQdFh5kueYsvNvqZndwbjQabvjDIHju4vVAkymtsQdqxi37KoO7Kio
ePqmjjuKN24VfmqfB2JgO82xiAT/If53lhWU0CcC39LcNEpem51d6hlHpdMZapqhjiDyK5dN0b0a
rn/3MPm90I9ri/KjO9VP7zHTPh08gLD2yU1uOlQIsChJMGn4RASwC7kItZtiVctfRXN7RfXwvEgZ
M1FK+v1Q7pJj4hPtLGh3UpqTpT6pNVIfmGu/iQErZ9SlBCLVx2GXVKFGnDsXToqL31NCnb60AytN
lU71mBJSxXjvG5GpI4/L7+2aeYGIgwkRfhj/boFoK9CPO0AUFvHzl93Y/wg/wrnHv+wExH8BD1SO
xayX8hTTOAdmghJuUDouBcHs9NV24gO4tZLuEKK4aFzDd7h9WOo0kug3896yHMc6Agn8ZKuGpdGQ
nG7up+T2QZHlL8xUFGCNijrI6svXIPQkuDox/xX2EjsiKXZ/Gqxvlb2QHU8S99Jd07eV2kTRK+ol
hIsaMiILbBxdBGqFQ6uiSWe/fd3ztDh5Hfi6jYRaAz4upXWOMSHRdEGyGspfFmMGbXQv9wuotMHc
gfKqICgezACrmOwUtxZyHIn7MHEvS99VYrG/qg5Sx3+tE3X4kn78UWV/Z5Iy+tsaL1nd3kGqjXJx
h5/llqWw0i0d6v925P9xDXPOof3xzYOFedW7NH2PUdcqXiM0DydDwmatNyQ/bHzYdJLOQs+yiEkN
oS0yeQgcVRE7G8m5EQXtxWFmWHb5wjwiR9dNviWVelBEw9R1vL3Z1iyi/oFer5Fa/1nhJwVyIHux
HMnVA7ag9tZtCkEozXPPCRF526ypkHP122u4fdPtCcwmpmGHmB9zemZ6OmHwgJeHRUjwnilelzTR
ZyXc5b9YgjWjISHFAD8210CNsfLxL7C3gsZ6F/4A+GCWvpLLBfROz5RdZvNY3Jcg3KKp3gaWHiZk
X2JvKRCdootowB8JQgJfnWQ0n8v2VA64uC9UWjyM2kjWAgGKJ6VXFR55ruwhNqOxxiNJIUh3BXpV
3engLsWgToobmEBJD/HwpfODayIhf8OnAYBrwi6kLlylmhgueOrnCXQvD5CqIHW/EFFc+e+hsD4L
//WFngack2fR5sXIjkkLNeGgU9t3enAe9SoyLq4sPQnOx/xulhZgFEN223xhwe0DK90Upmh1dpOi
s1XfuggTuF4dRlN7V+qrueblV3TC50JWjOpYNSykPygNvx70eElhm9LgDNtG4KXaTRJJ55F+APPx
VbH69cmgEiJmtH50E9WESJUF11uqzd/D42Ii1chHyff4I/zWkUKM2zBt2wWQmz6GEPLmMCJfP6sA
DbEcjcO20XmEoRwBpbE7uVRhy//GNA2zF1pCoeEnGXZdOU02//bLzVGkOr/A5zr2EleSvm5FAUU+
gtya7jxQcwSfNvsJHd9oOSqPfJ3TuTLmaXGxCzrOyHAzQVfghM+WGNw1IK0IuK0Pctdag8Ucj0hy
wLDyMOSAiJBTCbVWOtz93viOSTGWXeVHiZWjLCJhUdtTxFJsRTaOAR2HDIlCZgQcaOb9AJ9EsFhM
wkru6OpbASKxqQC9Q5TKxTo6m0dV+wqCjSaMcHPCpiFVIPnocaKAUjMYUO/LWkr42Gqp2TngnsPI
JSg8MhWcfNM3RLNQOzhhvL8jAvkcBiF8Sc4K/Y7slHkYiow/XO1zUlCvAkTMwkGj/hlM72cbA0th
2ltjX2egFXx5IO5VGRkczedjJNMNz0zDbUTo4GnIFot7VSIigAe0ONvvHUeExYVizKZQUTo1wX1S
I8rRk8cv3AvlW0x7FVH8W2HiMpLrUCYqOJVGruNbghzl2aplLXtbFkd6zqREe6TqTJ4OEf3wuqbm
Ze0G+4tcpSMwsg+ZJAaDH9IcanUsf5KV5aAs+Dw2zaW2bR7frpDDdwjYVCbOJoL4SlPi3LNoQDLU
wyH7giKTK7DzVcQ+THAOwi79sxs5J2Qa5yv72VOxBlxKCPHu9IiKo+ZKQUrmvSR1iJhLarXyZC5V
/1xmmoXpQhnFAsozA+V8srTXbvBgVNKqd7zs3x5bCp+ZE3ONA8XJ0iqukQPGMPBoNU62QoIOsd9g
QOjM46v6smJxS5csFZc30qYNbAeiEXNck39W/AilSA4Qzd+ObORftS10p9ELNBDbZJxPmrbIni8F
txoPVUxmOSSFx4XyjNIK1qPytfmxr0M2PBALYBBouuxrJs7AfkH/i+j5ygBs14HEaLaso4hJJV9q
uQLuxJQeShTmHP6N1h30afix4Q0orD0WdP06YbnD2Shr0Joztay2j/lvd0+1aYVtlxuPTci4e6Ng
8yqaQZFlI94P24XWREoRgBAOdDHQ1zeauBw7aKebK8I1KWhR5KxMtbPfFlQNovmFUP/ilz/wzsSH
BYMojG4iPu5poyE5AZ/ZE6BpDRBaeKGq5CGdQo/h4yXEz9GrYQngB75uxPtcG2nQ05xngiYqpx2o
KmG9bDC2p1RHTxmlrN30UNoWIkA9Z49bIybz1zgGfJbb5kWSmu/1piTZUUxcg2sIRbvxY2lTaEOJ
IdXY/hD33gjemhWWqJZN3PNF0N/M93K2u7Dw4iXy4DvUuqZ4fDootfHFKK9MyQOgGFSMnVrhfVOy
9KGKDVpoIEtrd6L2lC0llvdoLhBydxNB5sqlGsNwLTq7N6TVsfovbLr3AHVsJayRcCJu0+FFiJ+3
AO+jI2d5o/1bx7GYfR8OP06TrdLsoWaT9bgc3v7fedbK02UaH6azhtXg+hZcYbGIx7pGQqgaiSsb
yj2WfTfG1xtig1O1IuWVI2uGebjBROtXgikxYkctJ51BuKmkefLDffByu9Sm5PDO8RRLWj7SO0KP
YbvBw0tBALWkPT5sVMH5IF5a+BSvNyDCXB1GkjaeW3nuLEddZEyhvYCYpQTQ5YAgJYWEJoE6X2N3
EYw4o0Z3BM0k/q7kqPHxtSAKOyE4qtGVIpxW9AB1BX8FiF11kHHva5IwWKycs/l+DjB7jtTo4m20
xpv1wXeqmCR6DTZ+bEDaPwq/NNIykihB321Jxpzs0BSXnjFWStJ5aJc+icRMJq4VAdt5FCWhKH1x
Mtsy6loBdjGcP3HJmlIoii/WO6otv43cUPrB1aLrmCRxK1mQ72hhbGUYqywCX0mXNgfCNADM/IlK
HUifPfScnAYZvEkK/fM/OXQVtGACWDi5rJwxxX0ri0+5HyiDAvjVrr9hcQe9FoN3Y4+eFwZuNz5k
2u69q34hJv3CSf0zTOPTeJ9il7qJrKbH42zgfRDKo5FRXdxneXvTrB+EBaEJjmkcSWP6H6nM+sO+
kI6pmUSdJ3OYxeDejxpRFnHXx1o9zJ7fB2sprjGZqI2Y9Spiy+ndirbtMnYPBLsOhzv7ZytLRbPl
vrYo46r+Je4spOQj6bdntmgN1eGFIQlvtZJ9xAuD3agzmQRPQdVSfRiNWA6S815kKg6xRoSqOzls
Fysj3/lbi9+oQIk4RYDz8BQFP3kmZgd0muFghZuXYdXgp5JTf62LjfA18bBeK0JAC1bPOmYnJ63t
oCFDMqlJ1J3X/E9TCCtsKpNVWETM7OEuP5wc+cTqSCzH1ola808Iyy64QDZF9FQRRNHVlzDkRceB
yKB4NRIViEtnOyGnWOZ7N3F1PZTu8/p4jcS7USlj9z01F+IsHSfn2QZbKcF/u5kHAG1igW85zLDL
EMPKyioMsZHSHC6eh09pYl7FNzJ74J/FsKbVru6CmJBr709A28dqyr1/fMSwQ0jvdKQ1GXC/qSHq
QgZZGDlgjbWeXyAobjNUkriXCK0ILPJvemXH3JSn5h+7QfY8+XSJg6zxi3JgpvmAk7wtNHqmVaEl
sz9JYr+GBq6oTPxKG4o413b0srSifrokr9qFDZT+vWL6/GhUV5mQEu83MyibdvlFRvXY9Qefhx3e
6y+m5FGUSfzhY1mg6brNXE/G5laJfhLMLl25yRnJ1tot+KKKrY9jVp8jkxhb4H1P5le3Nps1lP2Y
On4evtLEmuWNJHvspco7l180hadIy5Wr/NX8TOpSkRgvjm/b/kpDaMaQeAPOlk4GR7l04W0AAaom
rBgNv7sGKNgpelbBSate/g2zyQekQfBavg9aO7EAfOxCbUyrmfbOZCyD6sHrh5A1PrYoTNziTN0k
kcxX3WIsfBd6Wn46bHoXKx+SEmi1dsyDe4Me6Who5s0MonM0466LRiwX7ajFHdnyhwcKGdif4bjD
VmTmLUB117mTfDI60PVj5HGBPbTb5ZOxiTn185COYmp4dm84BnYYbna2leDhvEl7YaXGr9q38mN/
VCyDTDt5G/KHx3miOzcgF+WFIv8w63NWvg9qMjoZecnf4r/LxpveIpvVR2K3M1ypiR5U/6SOgKv2
vhpuScnZktCo62McpYMY9529eSgr8f9Q/kc1wYyNdPnHZutDPlb63zrnTlgKSXTX8C3qE/yB6Kiq
VxWA9Ggcuxss45i8e52jvqrXWaudxnk5Lf0HAu9m46yVh3634vWLNvh0FlySNJk19eAgSwYxEpv6
4ged2mJawLQje2ZCidcz/SpbZbaEv6ceWodUpUBISwcYzPHNQfzgFKdBa0y1S4SYMb5CwZVydAKD
GlOVZxxDxFxL1SJrpEHIf9jMfI0kWFSp6YG7ZfmZLT3otYAmmRfKpwgMSN3ZcHBoH2RU+a1oWtqM
dvL59rB4gPgeGYt+Ui83bQPOcItpf4CSS4V9/lOgCSMYXxnj6jjETe3t6cg+CqLiPBsFsxSaYv0u
MazTNYDzzFHyOVW2bLM9p6RL/CjS4cHs4sOGQ3yD+/AgcoKzwtHi6Wy3Ng1Cn30F5U2cqQ1EhE2G
RdUnGMb8oqPj28ZGWTik/+WjUhFuTI8rpYlKjQVeJNBcJOcxpNuDiT4Okgu07QfQ3eWaMBZNgkRI
encWK+9p5PM/+vmMW00VGPge/Tyt1Xzgn4ZVtBqgLh25z42IWAYJWNEDzIWCeZrug+kK40N00Wt3
0Gs/l46MUaOMX+OqhYtRxcIzrYZYsLduUzMk9KmXSggbzf1BZShb/m3guydV/ZTf9i/h4hL2eeFO
1ydWmxDFeCcPeJrpAXsMC+kXstQIxVSwrm0YondN4kblJXjI+j4s5EfkLkCNBm0qc47RTxh4VZ92
9bQTSHz3ymUYfwMgpCZDLfQIKXOyaX/j5QnXd/ALNQG9Ji7dSVvK22slAS6JYha4S67+Bnv7Q9jV
8onSaSMbyW79DAZo5FLPMsYOB4pjl1OemiV50iHdiejkrX+0MFZU8Bj7NJ4HowM+47sFEneXxNIS
OPum5qCHYrRKDq8AOZnTXLDFL2LzU+fJetndCBKy8MKDlwA5mNbazujkCn9nb8tGaRz7dKKvNyQy
Hz2+rZOj99//tCN7GGgc1bXF8FRmDoPRqjt9hqKNVDto4yeuA8g+PqZngLOIgb9oDBPXLtlOy/4x
pCsmPTeezKvSlyCs3Rf1JFN/Pd1xDckPr0dcqwrhwKcNRLy3AGgbggg4sm8jKa5JLu/XwMVZXqh6
bKdvpDM/joa03SILn3CpiaGxCqfzzR01AuLegkshhVMECn/1FsOp68WWcbCIa0wN9zi06AdU456n
a0n7Xa6rOCbGCqLtwQQ478SBncNM/MV/BY8nx7TTMPqsjKzoM7DISFoPDrchHl7oeLr9L/RK80YA
0OEkz2FdGIBbMUnS4/xf4Xq8iDmGAVXhbJ5Qr7NvRgPKoE2qxmeeJhx3QVjX/qfG/2Ejpydafnn6
37v9pI44M9Mq/F1mY9ie0eWIGcTxISvFjpiY9+dd0eX6QI36gQkp2Llh4VPiru084AIqAaXYZZ5F
+t7ykNe9uKx8nDXTD6gjLnFSOrLGcExb7vgadFn/ZFXKLMDyMSdmbXXm6vM5sW43iaqgcj0Mpyy6
Fnjqft0Rwjlafs8E7qT2KY5+qFhvqIwp3IKSDa9PBaHtXQ/etVTnPMZkM3xfmKhc3RwFerAmy8CA
Hf7TKwJnrl2nhg7id6zQD0Oy/e81GmARy508F976i4y4vJyWIp5tYsHQ+BCohmaBDiKMkdSkwiCr
tnQJmFjS/0WAJ1SBPqQPTCLuNvZgH7XQAfpm/7aBPo6SFAW1Fjw+9dtqn5Y4/V0CXt2yRxeDW6wo
u4xCQ3/cqyUrL3gOoIusuet6ISUfvaTZu/4Z3quvVOXba81zmaUQ6WZXe0AIZHJr0Mp38FMQCTG+
hVeJobeGJXweLzWWx+MLE2Qmmf6IC5Y/lB3RX9alNJ5dgOyWwG2AAifTMcCOSkdLA/Wj6iFTMTPJ
pFjqELinblzfL7s5nLkyHagiPTVP+a9iluAq9yj1y/nW+bJEvZ1beTSVNjQvauJOwDv1WDT3yacM
YJF8i5b7ZGeEK4Iiga88e3QRMqpf7wgbtjG9+2lIEv97oIPE08cdwEBh9Jca/WQuc0KTumYoP5Fl
dQR8vEI2gfBHwIwQm2jgDeFNZ6+Lj8t/fnYzgDH8sVebN9krRH23785sL39Dj3KbZdKqp+ed5dFH
g+25nhDZlkpEtbC0QyMpJuBvfj2R3ERP3XDFAeocgOYzaY8k4exUj/eRHfZZ/ZDcdct94Uz5uA1X
4K7lBDdsxXSB3kLHfcFtUcPcjOf1OikSD1x8pyRWTyWbM96MaoaC5hMnKp/NfH3QWWfqhJ4ZZ5rg
JjRozVa3cl5JbVRNz6OPZkae7INUoa8mBEQIaWSDt0KJ2HLl8VOsCVkRREvYg1XPA3Zelg+T1rR+
JdDA0L9j2jsiLGVoRs0Cz9QjCwDjrENUW4OU5BvgOVJ9zcu7ibrNKtCmsIvMchCAG5NSJf3p7NWz
MRTIzmiFB5KWxFomvFDjhRxrEwi/ykfQT6t/F7aGykeKDuY2MmHqgDkry4IGM0Wvy2J5DC3iQ4zJ
siEK7Ops0MlEXenZjCCQ6xhPF3LsJV3wewKMcwQyYSqX0CN6clJRGKJed1wf9+7ZkaQzKZRm1EXK
vQtIGfjWOSbWIJU+IGTJjyvaeTICzKpgNjffeJvqM/KLedDD6xex9UXN64ZlZErsPz3cWLPDjn0U
yPLpLMD+q1D1GUj6A8r3OZFaVuruGWy+eOdB+MTju5XbqNFb06nYmfYAuKDavhMK2s6dJj4WYwUj
T0mMgbk/INuOitScuMK5rYM3+ZrBQoaKmll+6qgf2ZpIVUB7gYnf2BeuATQTpXmSY3aWHMQHEgM5
y4whG8x5jFsWrvM258JAHMo2wpqQMk43JPO1JkelPHG2qfVWMxilPc7rcK6VB5dM6JS2dfjUnsBs
N7fvJbPT+cRlC+BrDlmOK956hP86flGdFVe2SxbCIhgx0JYYbcgbGC48ZcTjSzZuoUU0hBSzGFQk
74lgRZQGwNT2x3F5J+9ehFWStVp8t5AC96sO0jE5KsNQCIolWwlns4mj5u0KFsoeTNGPd0+YLWnR
3pQVTNaWe1/htOX03wvBT0MBEuFzFj1HybKiaRUDOWw3UiQhtEGze7LbcaNEc10z6q0zeWkspBWp
n+UykFFX9kE/0irXF5Cwc93nVa6GUT+cONRx9ljPsalTkzRMmzjxboW4wUMOPwnN3jbBP9kFeb2d
RkpP3bWNv0PY+YQ/w2mJjErCxSSNqdr++/aX6yYD/PyK9Wh69CF2Q6KxcnsW5KeI5a8ruunpgVMR
NrDm0BcfBVE3HRdXxuN+caOl2C2KtEFTKgW/nC7J7aS9r6R4U/SaS6aOvdprxVdFcT4ViT9daeTH
9Y80lkaweaewWDXF8/6N3+8j/5pSN8VNkSs3EKC7KDBwH9KbB5dF7SUuchfsZHYsnBmQv0rcXUj9
5NU1498YEgFuxd8omZB12Gyd3jyN8hxmeSbKrLk8lAdaNAhy1KylMgrH0jOBWJKazFboQQvUr/mJ
ifoUAEy324fhYqa/qffpYtME88ppHIf7WBdywqWj/S6yTtFtR8WCEzgKVVla+UcCqeMRFO+LbBHO
2x8y2MiQR6HXz4HDJaRYpHVVcVx2ylMe5+huaojHFlMt3KOTCC+7VTy9E34kgsSejDFQz9i4zFzm
4bR8OFJpdZ6AIBaiMV+TTmHaDKITUqxVv29upQXCranbIZvs6lrVA1+vzY4UhlWcQmfzXGdpt2qr
KAHvq9qzWdt/kHh+b4C1OgDpXOr9/8gOB4IECWiBi6i6nXNatXrbhkQomv7OC2VMCDe3zawENoiO
B3o35PGGJd6zO6E5ozyAfbYuogJpkJsdp6oYg4FVXZInWVaCi374nEdt0LtYUZGJIphYgn8KMqWT
JwMf0N3vmGmHJkK/MReeQ43r+tQ54gHdMEmob5hxtzP8FBN1yuOeHLrU0bpc/h/gUhnVpcFkeq6i
M2Jf5YXO34ha2cDg6AaKG8F4wSIErT9BcgYTSNXOxaH/3jWFmay9InnxEV/2vlirHUytCnWxJ2Zx
gSeA5jdX/1IX6IuBpDF8WEw/xXtjdAmT1VMTT0o4nP7UqZf9JzVAJWa0HR38a2sreNCyBwz/BeIJ
HwkNcIEODm5yukovcUaegXMVZxHXV880z6vOVSHnQiD8qvY61+UjL9A+RZkxImGphmNUdlN/gGJa
8AFSr7i1NDDlT2kgVNsvwDtllHH2DCrpfvwb3wgt+sD6DVOXNLYCsyG3YeXS5LfYmvYVekbDsWb8
lwJr3sJYDU0SOv3MQL50D82Ll+Kmx8TZiDW7gcrmozsh5fgPuLKm1n+WQTpGAftdlUSU9LEs5iZp
ENxjA5WVqvRYXsZA4ZOW3g0eVF+JZgMy+GBVcU8Y8N8MR6zb2f5xB64/nIXiKw6QrlNeUn5n36j8
qfgaxdh6JUqPpw3X9cFw2kjR+dRtAVqxSKSrG15RkqYL4JdGkwS6tJfVJAE0T4f3h/VGSu4mP/Kz
4WMgfjZYsH6N3zb3gcuxAN0yr0RYBU0gT2nEXv/QzovGfcTqJsfmSBYgwt53vz96d50IbU3H9T2x
iNXKqeL0GsB1eWZ98ikt1ii6FPbN8pnwKqWxcjO7Ia17SuQxsItJmQcBjz/4VeSqps2v6QZfMCrE
+qD3j3fpvFPZNJcamAD6HV8DEim6cnHohWwvyZ64wwjRDnvVaeyiA1/WymHPbgaAf4Ug4YEdUobt
CG/u8UhrQcntCsHIjjh3su1lGnmWoRXhucsaBRhu5vbKwL/hND7BpjYaGp06mi0/H7iOz3ez7LH4
speZ9w6KR1zrpMQHk1VwqYwYc80UJyoeJEwIJQJqHMpq04cIaY6sFty+7Rofd+TZE8q5py6F2ALc
NxQS7pelZb/RlGNl+Tm6VZ4V3vR1WixMhQlp+y8ykEBz54jPOiTy5pWnTQfANogyYh9Jx+4jfup7
Yuolrj1FCVkP5wZ02E4amRx/jzwvuP+eGI8v6ph0QwjMY4qBQjP18PfhiUIxNx7clDq4jA4yb4Ix
UGpN6WSyZgP04uvF/6HAE/wq19UoMs93r5PlmVZECo5GZsyVFnZyxlXD8g6FaeJ8kf227Al/AtRh
nP+QG8iSXddvGiLTyUccGhbV9rtbRYkZHtr37Kybnszh8fcAEn/cqzQ3SBO/6Yz0dD5G5/skuA8N
DgPwwiYNNFfnth3bJveD5u0yN2SLOq9INFaV9pBdXyh5vZCt6Z3BDJjdBxXVV4C1Q1/hRXdkdALM
UInEhG4TDQKp5trWKTmiC+hj3k8BrO+oecLtXNnrzNrYMFceaZPHx7zg1WEfwn6VDmydD0WVMAQb
CfDmAqudfBxeaxS02+x+oygnIEMFgpAPCioeb/j2jtrXx+f5rWbnqlgAQEpl2a53m3hRLwQ7wYgE
Du8oNq2aMDwZw7Aat9WJt8OHYI0X241obvoLjxpbDpzhKysfrIfLMmt/Gq2z3J2X5JYj8abwIvjq
0Dw6yJf4VyAE4ePT2J8uQctS/lJyV8hnN8O9AJ4YdC1IVDsmLbZsWOKIQMic1GM/WTsSWQPT1CBt
3nqzLgy9Sqahps4y8SDmYM6sTrXcnMA7gtVi8Fh7Wm+off5qGEX6M8UIDMa8D5kKr8bRXFz2Gqce
aghIWbEheKc1cKbnX2qM/5HlUwos3WGk138XjLj3oOFID5hXp8zO4acs3vJFYXqIVRFhINWvVN3d
LSGNoXxd6gDpax+uR1mbmFNHgyPVdanBdsEehuy5SBWFWXmMvtNmWMdXnRM/+++55koDNSnM55SX
ztdqjiR7PhDbW189M8rqF9WdXgijJ2OpF0w0bzV7vmQBwtWVgadZazQ8JlnRKh3pqzXh/ssIdQh8
EeM8Qos/rFykYTUmSAJqwCWw8h9L6F0jQjtUELbL6sywH9edhCjpH6CjJFnAeNlv2jDYapWI/4oT
qC5S9zKDsOt5anbjKHmDbedwZVqAUh0c7YW392EPY4sO+aoeHhw8O3rwRVm+wKh38B/T2qnA4sdS
uY/TMtRZoSykIfHV0Y5BxrNLoeCdUuJL/6Jom8Q9lrglgXlx6Tz1A4RHbCwtLZR9qG9MkBMiVTdj
gDg/W/XVsnfkJGeyeqCRiyEmyBuFna0ANjYini7Oa7QgH3nWkir/WxiV4ScNYgZur/62x3CnHKCf
G6DXup6kXfJ5prBk1U6keZx+s99AAqlfDjAIwEP+h7yVZcNIXNCkg2iy1nbxj/TLNI6maDKWC2FM
zsMvaIkxHPSwhGHruOz6cCw9U1ztXh9OGjczlsqq6bQb7g0QZwVGFGxJH4ivsHCyj4QWxLTv/Mc6
PE/h8c8Q0TwMu6prUju4eg5hZRi/EoW44wj3BZD3nkF+HdhZUEmVKULYNbKEcf2/R9e4foJhgEiP
A/rKbXpVcUCCsi7XSGaNK5O1TfOVU1/xgzp8uYw7TdjSecL1I3Cfri6FD1kHuoa9Pd0U/w62uAtB
hr4e3iHbj7JUEELMV+yeEF4rBhgaWL4wLr0r0QGh3mpKVi9YrhZD++t8lrAE8Cff/BowquYEPFfG
pIkKcjJxYw0JXQqCDBpTSi5ly2SLN1OfFfuSB0Yh/bYUkGrSKFlrSPDtHiacApA6fUXSUDc7XC/a
Uu9c5N/kHOggounQ3V7jamO3sPZmBbh4EV4mT20JLdX3+4KxGYSzjCnLQ1hXku26gBi6w8l6wICT
gydzstwD8O4OEfqOyFGU2zzpW9XvDQablWAjsuI6JDOSILX33C/B4JlHQ2JcFIdhE2+1D4Ok0Jsp
LDJs/XHtQsSs5turMB/b9zleAU47RJutdY+inSwQcZvtQ6YChn5paKyuiBZd8D2QViGNFZxxmsS9
sb29bCedvVu9Rg/ihJtj0WoGsP8DqB/fs7297aS9TOQBzbmbsr4yiid5xVQJKe2MSEGzleZlI8Xr
ozniKEeRd4tQjUaHC1Bizo+7KDI27TK8O78joj1CsxThAbyZ1yphwuVKJZPHIuB8NFp/VrPrBgBb
+Oil9R7VFbDiCoUb8gLdnUnDdCi6V0kXisoDJX6FPsnoyq/US6l/2wTRTxgTTHF2lyetHLFc+xfR
SFjvpg1EhK9AW40ldZ940AtFgr0f9d3pmlzeLrw6EytJzmETaYX9c7khdYXyK00JorhSdc6ooBxF
/53maWmRddS8qJVZIrMsi5UV2g7DcQLjkJkVRjsntkvSk7c0g6JmyDWg9BJ2HQ8pNgs4+7+kR1kp
xX24u19p47+suvRgZEMGXExsY39t2Tqx+5OulVgtqnBo0LNyHR/juXWHPYCU2IfZuIf4YX24WAVE
WEZ2jKsm5q1WD197Xck160Zocfj1rBIYIiJDuW22tkphdjxsYyZIwoVodUjjVWYcaU5h/fypuCsC
P0DL4gjUfRjrPrxqvMKs5zjh1+jTM0afItdZMnS/Z+UP/t2JdJ8fkv5IvKNLC1K004HgEatDv8Mg
eCWXIN+StywoKBtqX0IJgdzKRIhldNugEia8ppc7tr7c9nXyvkq/srHQPG083hEcK5T+5Z7FOq7N
AqU9bCyCdpDbnxbrVjBV0QHD4K/WO7ENikmMKjm2LBZWkwiHcoawRhaugEetUmHfXhZSU/RuD/xv
mxXiOcg48eRro7m5dW3LmL55qFqDsVu3Xg6nlBxs6QJXdKKrAIfX3OfjJXBXV7XA77VnZVVqRscF
TT8KPbHYUlYKuFx9Uyee+f6sovdrRA+MVhkhW7UZTp2FyRq1RVpiPJapEJWxxtgjKLXGdGYu6ncP
z6tupRNOxrAc2t9JsNyJS4F4WjeJBx49eXVsl3xvNdNm6dheO3uAHOuIyhsyBoMNHQaETw392NSB
PghZn9ko6i33DYzcw4eRsBGhk5z9uFN/On9/gr1nyqS/STlQOsH58Xno/n7xDuy88Rd6wYDBFYhv
u3FLnh2FQs2JFTMc2qwDMRv2ezjQtjzhvN7MZ91SKbL48Y4AEbz83+X33S1SU8mmYjL7W5mnxMSK
7iz3GtZmJzD5ZAOeHKtcJxhyZDxuRlkCIku7Ht84Eq3MQkE5Kmdxszmi1AWqJYPXwVnrcMe3Hg7O
SQUfhtMosdY9KSMPI22dG/Kt1ASEce8o6XQ+bUeyfj8i2KqmRvOfMqsFsfwXs3gzZbTt5Q4GULFn
qRK7DgwOmJ7GCsDpgj9bcCg1d8NX0ARB/dBsTFcpqPPy4c5HS+xbSYMvwUY9vawY4IREj4Ps/rDw
uTfEGxSzD0BFjIhHp/qw0JEPYp54a/89jbNgZH+uDh7nU0lNgPcPpmm9lbbmZ5dogbpP6GiofcCC
BchG4eEuzZGtj08nfZyNMUDjQFhZVHtfdg8Jcg2h1WTOKHNMFRCK2jZJFk2UYxdi5nRGxACLXJWK
GeTOD/DEX/NBippQaQ6XkXSAXIBFXniWfK0qfu9BaaFNkha5g4j7VWj14ASzycgW65NnsXejmncW
8EneQMfJAN1hOSjHDvg2yGb3HDQ47buELe7tw4aeyEN+tO8LJDPTQ3gK5CFNvtCK67uK1PfzKIKc
pZO+KCJf2p5srXT1GAJnjf+9nEPnKOdd7cpxz8m09lKJgtMI+XrfsePCAjS//mTNZYOH39nRlKOQ
deqMx1CvmqDTNMohgFAsz9u3gfksbD3mvGTpUtevAxEYniuZ8rZrSNtVmLDuHKGgM9yiePeJtQIL
Mo0xARq0xXQyEUVCQ6Zk8W4D8syDGU6pbApZCWkjR8nuPvRKEQXsUJh1S3dmR/Wy073oq3SAWthE
d+5ewAeJKFJttz2SG+4dSoTvkMlKcrzrMFgMZnFEJFxgdJHM3YK52W2X0DfYadTmfeMsXjcqXtoB
a0x9XfJ5CccGx/CjwpSICP9G8AOPAC8GIvNlB5qbxkh4XBVS9hvai75eYybl7xL5UZpUdI5ntLka
7ryYZTpvwUaRfegjIz9SkcdFk7AEoJccFUtQhCQt7U3clYLtC7OLOGsRkgEM+r+5yLBVTtR5FYSf
vPFgjRSr5uyx6eO3xVLV02fKBwKh0lsHCWoZ9Day/mZz74zMG6VyGmOPpcs8sJ+4yEN6KLVhGLLU
UBtVmZwTuNs1A1vldAWFIR60qSFp3G3NUGgbL8kf0In0sMTObyNRkTHELNWvYftqchSceBzaUcct
WA/ZRgIlxzJSDHUV9qddmq64dawyOOI1mE9bZUUb7jjoY4vy+FsYhRKPRsCDrjuEGoIuGloDrz6W
dw6hnTiwQuvkVWI8xw7CIP7B7vlejCn6YS5YHtPz968YFIWtBCPeJ5uvjHvtfgRvXN0Cd565ELb7
o+kd+MKQNX/T2MiOlykO6vpmMpp8zTaBja4UZXj7AHgoCD+eYgpbHsaIvC0pOOBtjxi1xDv4SeLK
k2k6QqFz/y/PrZFx/dou094/S4lUEzq4ntyCXDFhDB8qGJ+B2lmyyzmDwWZo8A3pbmRx3k8W3zxY
KiD4PWyVNZhz8C3dG1AMV7Ed1bs7B2qeTiCiBWJGyVFjv2ohbU+XB/Z5Gtz9yJp+lRtw4eqGa4Jc
el0OSrGnrBiWjle48G2vfb8mOgRosEggY6naawTA1Wr1jWwn7ZUwosSgbp6iELJittOz9D5yQ0kS
X2LIQapUO7a2kqN1r04i2WMOrUK0CnlyvGMOtMVEA/2E24LNcuuk3WflJxisNnsEFUeUD+RU42jf
elqmCEQ/Q7/s2T6AOOfT0/HCIwhrC/ar7859zKYqAlhlg8gh7rFS1HJoE5hd+8sSHRmtwWlvFitS
neRis9yhE/TWuKRqsRCMXRwoZ4nnq5669cZxTddq+LFa77DpReTh3xaqnMUSzW26HeuV2tFrJlLt
vQsX5D1yHC4T/BN9eJaP/4WoLUijtsi7VWCGw2QRM+BaJIKbu3AjZ/ydjWB81cNW3AsxZbdfZW4w
4LTiR6rrevMioj/1n8c2SYYRu4hCleZVGr9NMYOiQRoroCLUUJGZidxXEcAxKgFB4cFN+PtggnFF
HrdkJ9AG2G4ep4RI+dgOKVRyFR9akDDh/h/C7YcyuJEUJ8QbF+G9JfIGJK/7YIZlwq6OcGijzPpb
hAlqJXoRAFp9RP72ZaEg0XMBhUEYTHLIoZtPQO5rmtLeX6VtyJlaIWQwUH/sWDNVfR+ZlCDCZy/r
CypHmxQ5oAom2Q3jGRaTyEpbgIkSO9I/ZR0BTjxtUI/eN9So9Y7W3KCb9ipmRT0/RPKeUp5pTLq7
wgHNvZvkPPC3UYgcPf7LPauhulwu9Aq84RRJueJatpJUx7QkyITfzfU2qoXSDkmZmukA1jcDRQg5
5BnMFXiUMevQtVPfi1VY2NyTEWACJrFBN8/ZrI1/FQfQh1ewhg41igEsjGmKhrSzwJzE0ohg9W3C
o2jd7KZRzxD84XqYg53yDSKj2vEYZDHk7mRqfspx/uWwOYBNesPnA8Rw/N7L4I3AIz17JU9Ol6XK
IRC9TyIDyDZ8WRfenJHVIIVDh9NcCkV09rubdv36DrFGfF3bvEzk/79U8A6U0I2O5+Gvz4rVywC2
1HuMONg7aEmJ9i//YE3DiCdxc9MpOeTR7RU+p21KWEc+k+lm4DAi2SEfzKJv/PNpcoZk52W8vSJ+
O0YYepoSFb3fawpq8R9M0Ma5MYTofJ/r6UzARn3GOjJCFotY1fO6hpbZZcdCUMHZjK6cVTrtKw60
bqD0vk66RVTc1tdXwaVFzYzlJ6TBWR8YijZzB1INhtwH1Rc1iPtcfRPtL7CqjGL2RKPJh95tItkz
DCoU/ftOUxvmSvymYsKxNX4WmPEzWL+c2DlFewoZC89/FeizUG1mvGD7fYghWlZvjWoftffnC/IY
vy1yPnFCTnVbXFJCDn/ULiMudCM6hPPUcD+wCn9tRbsBnKzXJhfX/7n9A3UYUhmMbDGM/SSP4zKE
RuY6kf940YhvZkO0mjUmL0o7Jef6SQNz3aDlQdrHIhU6aL8RlFGI+y+/cg6tJkkm4hUjhEF88TP6
GlUqF7/QzLrMTuoZ48nUeWz2XBPjV1z1TqNaAJWaesOeEUOv6A2aN+dkI/w1yqvegoYe4Y9gRRxd
3HIYHBgbLjDtwyjeNTSodJVNauaxw5X2Pnip7nPNWhSFeCcv4fppSQygarSptu3roXtuVSFtafuQ
SnmgwMAcJkuSkWeHT/UZWK96a+4liHI5Bzs5VdkLygx7P4amHackvGTTJozcJ1xo5HMeQ3WTxkg/
8EnBRZPaaIeca3r5RQtn3JIjbID4JXmAFx5xZdnnUEsDcXYaJ/Cm9q9XzV1IHPv/S2fNabUHyLWQ
qcEk+lwtLRrrX374/AIDMeHmFfBkD1jgCDTN3+nI4/69TL6tjJo76IMtG2lE+YV98NhQF+9ufFnN
8p95OE1vu9JqNMe9tM6xDFSObNWiflbN2nZoX3na2OxL2blmaPUtnsF5rY61xE1b6Or1rNEJBGb+
EH08csaAzWjdqbG5l25BOwWNohGJySh6pQxlWt6XGFJrjzms7iMj//NPNQ3Rj34ZysruQZCHM5eA
kbqeqbz+CKfBXKkGP89JEjcsHhsOAblb2l04f199DQLSqZ/6y/4M1IV3e5NFevjAKDcdvjYJgtnI
hmR4vP6XDA6lXmpywBs1Jf6ZIkEo7ygkdJy6bQ/0C1gRDyjkung4Z6ZFpEt6doPoNMR/afTNcE1j
sgm6OmIW1Vsr6YM7XLVcVEbk2WjhqcuQZYrrtTxyLEoKeAgIe3WyKDzwpamRxIYs2LUppt2tBZjo
y5VHf5Rk1qIvBD+Lz1uh6Os2s6T35qtqPA1gqgJXc0ektZiZ3tj/AIryzs/CMLQc2a83o6Y6rukV
7XQ2h84qqqg/8lnLGLvQdxvqUM3+p/95qGDlM1Nh9RFUxdHSMEweImjG8J2t+PrUaalWD752Hjxt
pgFltBzSyOVZAXXCOlpgnJYXYCRN06yaBR/koix9EG07K2gFBuJjVDLWG/hcA89JLVdlxx2/VL0E
wIqKC9LIKQe0AeB5wBFcDbZc5cisD6aqGFk39RxlwVxQGgQAmWpBEx0guE0fi3y3RcZtuZEcEl5W
WEJ7s7DCWVJj5IL1xHrKwFyGojXu7udfPXKQW/+JyPKofbYgxIGH/x/p/HZYMmRRGzawVNrpkdm0
/siFQ7ivpnXWKYrkMV9ItuA7SO0nzWfdnN92Ntil9DHQwlpaLvdf9ropkIQx7w4Wl7hb6+h54g1W
9/xS0aXfWNDu32mFxdxFqRlqRFxT4TYlJyFnSiRy6xB/EhOf82ySV+0uG4/vZVjolRc47TNQP7h8
LNcO02N9h7sNofChfEDTUTC9TffQzk6ywUGGwvaohNV/z958Rq0A2wiwcR8bprjVkARon/Xs4Ovi
B5rkgNzcrt+8IUm7L/cn+ulmPOvn3eAsZJcS3m3cib7GqntxVORy9MJVsivk8c86LiTNay4Ckjgi
NDtQAXizrQxAWX5t/IuTePfwECSYbMW0mOjPSwHs/5iohHWJddyJptCkuc02rgit8/vGos6V/HVM
LdNED3yfzxjzv3YuMqYBnW3s+tS9qVsjEzZNTAdVvtScOpEyXMJyeC+J+b9LvJ8C7ty2CZ1oVo99
ti0KKIbT/U/Wqa6nzklxN3jbdP2KXYJTKJFOth2X5x6WZHFsxpAYrnZKr8jAXaRIZUbOmOy5uPtx
K4SOUE2BlTud73Ij+kJ4tPxsvgWicDbFap6BAQ9x5mp+pM2hD/ZrjQiJ0NBuKd836HwX2iobKLy7
ku4X/F09ybKPsSArxDZ9mtIua+R38YLhmlxN03S3jjt3g4SgSqH3wJh3CFCMkGipHDL2njbEdsKQ
iXXRiAcle52C166L6d/oWuzY757XZ/k5AlwtCy2GrB9M3AcU+3KKlk8h08nXJViz+AdXJZsSuDBN
JdrWvkkZjeAkm4vTUKKzo98/KsrFW1x3SYw3DNGoIoJcuru043S7MzaPg7hN7o30BKC6f2oCOv4q
SuHGoBnsVZYyo8m5vJlOsSqEI3MV4dquat+bBL2qaZjUfg2faQfLUjuLp1ChFGgAQ8exmnM3mIa9
UNUAH/RdJmShVl4EecQfVWfAh4LZTqgoTG6ihUm/ZLPns9hANHIm7jyzuaah08RtHeTmeNq8UOw0
jCg3yaG0WNQoH5OqWFVzmOnoc9kcr9Z3ViGs/3AAGk7C2i1DmXut3Syc2eHzAtxx2bSaKf/ZNHHS
DEASrxexQy5zWaqEP5ERSmiCqTrWZX1UhC8qFoK/3V/t4xIkCJj6xs3x6wzZwVEsjbtSQep//LhH
oIIlhn/Zx+bobTZCW52GjfKYSto0tLUqvHjudwnxOeqtq3OghmjakfAi1Rl+reWQSJzGjuJ8ygOi
G8EOu2BeCTud8cqzYqbxthFsfAZ5K+BrcNCb+Qejcn7+Diz3akqiizSYzKnMKj3rWm3rMYbiHRII
Vml0P7BNC99FkY2iAuoTNxf03jKOv+nBoi2ck1VTprC/jlEaj6Qz2Khnib1xnyrFPfjxYQm2RMoY
veuzZZTy51cXS/haxqbfLI1U4iZ1AXBwoVkWdYI4qpAVocAykbWX/KRY44U6FBywgrP638p97xug
9/QA5wSqMkcNvzBhuF/HcUDzeaZTIS58HeGU0xUGTc8dx00ZV/A1ZbaurP+oW7Gn8SWXvojVRg1x
qgpBEBLW8bYNjE+nJ23AtyC4TkSd55Nyi6UcPqdRKY6ElikQQhHNCRKjpbzUSVK9Fxq6kaIM8j2t
xaj18Do8Dc4UGRL1AEbT01EuqAKGuTawG34jLQcqHnLUClne1Grcv77PHPHUCe528QKNDfF11vxF
ritWpd9JtQxE5KNN3dqHhYV/2RcZBJwtQSV00ODGqMbSYk8UCD+HIDADOuyyAOy4ZPQig7NcUMaj
85HdXoLCkPk04MhlQC55mjO6vWGYz3N7GSMlyL8zvjzVJVggdQK6j0ay2LV1fmbFvWWVZ2kYdIN5
igH+CEFpGE47L3fjwI5L8JLweS3PT1H7FT8qAGb9hpzmgH9de/NS+/Db53v7ItXVcmGZJUe3blik
xEzdH+KW1dkp87Dort3KHY1aenlfkFQ0PZ8ExCWXJL6LVnt4iSIelhSb5BnNRt7koz+IHyOK9AYq
oAksTb0AsoMBsSQxkDA/oiAhUfeVw0T9mtmE91hoVcJ9xIqfGhvpfxKQWSZ8hdIEDQ+wGscmMYX4
5i1qh6p8239zSm31llrTvs/EuQnPcoYLzKZ9otwTbQEvnsnEwzzh2jb3zOaHjJBTV1fRrM7gNd1A
doan9UoJYQbyO6r8cgyFqAvf4//ztSaSUM7AgDD4Kv1QHKMyDz7qoXOF+UATgoXdqpZ+wYW7T/d/
26ioosieTIgKmme8aqCBNzHWRrhJK08mQelV2W1ThUeBl1IT9tCPl14V/gL7m7EipzRMC5JpJ1cf
+5Qq/RN/mk1SAuUSMs1kHh0msoHOeRN6niBS28Jlr/1u9bdWQ3YDdSAAe1NgYJ6778/Ih/BKG9MQ
F1/RMsJLV/hir8gbfqxb28fJrPD0sl8xB9LUKBgY6hTkrgPwA7h9Vkv/3jU6ky4Z3hvSyTvVuo8D
+FGPoVV6P3USlbxW9gxcLt/dlvDkdOp9aAv21sFzlWJXaokPxWwZGhDlH6TaDMcGewetEcVISi5W
5p948Xj90/2iVddSS6fQYdmVa1sS02Wx5d+vzOVrOdM1ZEbjG3gJeHbzefYgUs5pe2JDf7KE5yg1
+5Ol0GBLI0lLT/G+rQ2fYIo0M7f/ZWCoH5ucAbWDtxJYWAHrA0mGxYifgXdgv69XNV8GCSlgTLVP
9HQYs7kR0N/oEft9gmVERq0SGrDy6K9uALc80UmbGoeehGJJl3BPWpx005ubuj3bGw7JGhkashSJ
U+z19rGkRCvshHIhGER9yVUyjrVNfWtjL3GaSlVNfaixRNhzcjv/O6tqz72DDahmHocNPRZSAxdE
0zRoN1X32a2u0ARmH8evpyv74JrG1pyoriCAdXZyA+QkvqmZ6899/x4S9NoFIpU7wMvGQBPPtPQg
TJ+8suZdD6BCFkHBnPCKfYvJqexPLyrlXirGKdyjtoQwpjKO7Q6IrbbIDDTkpTQeMfRwuMVdbxcZ
OKufNKuxxRgNHc8InLWaHLyS2LKlmvCiU+RryrR5+/33tgMdq+2jh37HGMjK5ga80lLedtfspLgm
oJ8HLHUDCouPqk/ThHLmAu2zycAZamg05tIDLgOwkoledwj0Lcx9FX06zMcxBbpfDGAZvLbSjQts
JH3qv7EHrG5qgAa0vx0nIJU995q8ezavzkaViDhjLUtBd4syZulLGdjpkD0lAJBKzF1yHEw9hxmQ
490lN8IWuG1j233a3qbt+zP/KlyHNkbMuJwXjjKtSsO7c5RbK6VKZsHefNDrb6WMk4sJplenIHaa
jksHg/lyHgyjhNciehb1Zyz8glwSmLfbXM+7jig9OFF0wdZxyweoG4Wj/5v3hfYFvSLsf6+B2Ahu
hq7Wm2lHyMBr6lgeGqrzB5foS0FMlor2dTvZIxVQ01nw1ddMOXEw5ZvZ2+MQlDuVZwA1IeC98cSK
gEf1UBOvkz71E7s2f93VkHjdh4eNE23nslxDdsOqTxPbQqvPwzRYndy0ZDuMHnMwKxSbrIIaeG8s
dgVmJAinkr76uLEfwmx9C6c4Bxz7KbCswR6KyM28GJy42a0U+VT8YsCY/zEB6+tqE1HPOl1/Va3V
yTWdwx5myqxyWl5slnAi/d3HRxp8zBWzZUSzttnRa3JuhLZNMi976hLc8Q664ruLAE3HMJc1WF0S
ULEvpghDghSyY4LmOsh9imxdBl9VwsiY0RNf90NlHH51is//9kcFA8axhnzei9Q0/MAFi2sEPBgE
YGXHcRfDmfF9BXndq85/uTFSMGqZqVnvqXuh7srId9K9FwzterPUFVnr2RDr6luHr/V2wk3q7rNw
f7wx9nuH5RQBicd/GW2zzc7d1npDJLWyI9alFqnZFIo3nWJ+98M3vKBQarO5BkfM9HJGZvGjgV1C
FEiUqxQqHzF19RfD7Iv3BTeE9CdXj5boq9WAfWskSAuDWMzVTXBwuqLJdoJEBFzskPzTQcciLO1U
QKY+ua3421vNjj1+bIsPfVSlCxVUcfC4jWQtXMbrckDbdx8mLffk27ijouZr2UZCol/t6wWuTDMC
wWR3IVeyPLwcEetPV1uaVzt9OIIGHMMcvEtBGwJ38Hsfr+NHeUks2jWhgWsg6JAKYDiiDBN82Rto
DxOSlYlUWCSCETo2ezSXUHFaPwPgnThjA5ZEMetrFexVPA9cIPRhQ9DYsSYx+BatXEzua/A96ZED
/skS1liGpWA5ndKpmJy55dz6HlcJSv9PA7qrVOfdoSGHBSWkcadEwfozAPiOfIPGXe+HjCropTfu
9VUmgjLk47J3QKo4rffAK9ShxZZIVDru31qGVq9anTQjJLjevW0/62Zor1BzYru5jSjwFMhFbKzq
cZhIfiBwd/65zYCjzwlH1elMnNNqbSswEBJlX/HgncuUbWtVMcQX2YWGU86XTlZw+qlgumpaGZel
AISbsSlovZawI3KWG+940hMQVOXm81jasQUge9FlHSFogNUok5aFMAv5bYgXN8y30ELZgbSNJ/0H
bhvR6473c8DC7Jjbi+3IXx/gTWI/Sdukds7RSL8UrSClbh+Wd55xI+H1UznpTHEcDxvAqL72NgDQ
KunlNxen3WqfOM2A56CSLhGtayLRj9D01+cDVg0dRlWvHbMn3ChSMdsSKJxz5IsLuVVR0jzeyHY/
ivrvJ3PKBxf7YAVUsbmgAkFYwGB2/tCs4fUclCpYOVElsPzZzRL7BqSVnBTUjhAg/fVOte2RH9W3
QKvy1PxQ9pnMNtKjciwrnGJ6aHR60QTxSrGg04sDQ5lHVfJCP8Y6Ebk9AoH+VCErbmXMvXn77Xwy
0C13xEHcUbpOeOK7XXc85xiUzXH6UphyEqiYWX5vghgAye/DH8aOiVooUnGIWF+fWxnVqLT6pbqk
o41nemsqz7bLNimx8Y6hDlLVNLPESiR1Q2eeth2hIo/7w8nbel4DwGHCKR7U/pEY87D5T40xrN4Z
M4XcziHwfuaQ1Cs+Jqcl9+Vn50Y/cyyi5HzxxfFZGih9H93COa6oKSTz8jtiZzWus/tKBWpGoobf
WvWra0tLpqLtuQ5TkVztNjWvamRdf6zK8D1T8j5mjJIwLMz31GUkFg52wwuSFBKpemmsCPA8bfWA
gQlz/+rXUBetzGWXZoTK5opqWFcoYNPBmQz7R+5qPCRBPtRa2Z8ICEtq2BuxDjmLhGpVRhpTv4cn
/UMV51PNz5xUCnzfnJGr3mPbpl54th9iMMfgyCeB3/7BdDG5LG2cBo1LVhYQfHq173fDp0CCKW1t
cwr1CvV+izZvNjfP7eq1tH0abfhbwiYnQ6cm2FDKZz73MEPDzY2JJzDIhBr7Hl3cm9CxcWqOq4TX
3ScaGOkQtH2zz5QHTRlW7yqJp75Q9/YjGG659pHgjHGRm3hfDimOf5ZWInJUFOSWVAVlRo/5WKZc
1xwGw1ENPj7IO57V8AhwbamQuVg2glU4oGAJCiq6toztQ0oqRMvAoGqSTlxc0VVUUXpIMUolIjc3
97ExhT9F0ZQ0o7NcRWrly9QMeU+fqqC+FH+Zmq8xx5PJHXpLdh8apRl94RJLYglPgWtL6cRVUTIJ
VRGnxD1XJ7xrY5cwJaA+T0xaxayFYQJQFukuRRXNLeHotQ4VlbM8U2PaStnpnNX8oS1ldkBrXCuN
JGbq716NnooYC7kKycs9yJBAbBlMBRmDsheiLrCKotH6dFqAMFKTJLWAGTmAGj4QsT8pTcnLNzyF
EDOAtFHRns/sS7vb9NJ4cjL+bAeQZxEeI3psEEIS96wMJA7xN5jAWLQAPCOLXlKwbiLYV9blXUuE
8koOko6p2MUZ4+qrlA/4OXcB+ux/RZUJz8PCHFA+axeDkQvCbQU6gkXlEiKaRI1I+Mo24NC2DvPM
1tW+EIAUq84As3vklotpfq7WTx73OMQhSxaJEzmEXZLX0sbRmwmIG0GWUgmU0G6PsNlic2dlHBFK
oi1ohc43uL3QzYFd80BW6eI4TUgOxm+niHt9JMKj5AoEXxjyZsQvb3mJnv9xUP8/bYM0rDUIzofy
X3U/G9UGLAnk0G+pdymKAX0XewF7iuNToq+0zEuYR+Yibiu2U6VQRWx95I8CspZzBB+RlSx7oako
7cBmV8N4Wv6Xy/FwZQDszoP1SpatWY+3tSH30dIIEzamgbYhX2FK68WP2+ELHtUNAka+oiPjp9dy
7Zu4DkGi+pi/bcU70aLyPtt/Gk2DzDhCr3OI0Cen/v9oWdIsgwA9+wgUYA/zlEWpqSw9E8AGr1Xr
VvjUNMOKzNo0RHEe3FTrAS7cjUVGZdqQl2J0AhF2/aQsi7TeFkUlzAiRWc582IMNm03rytSvcKK7
u6h30ZOmd724EJqOPAhh4xok7c07Edb1/5zAMYTrpEaBQGpZT3p2/qJvajMTUB/8d+zG1iCz652e
91rQv+SmbRG4R/TG+HIWlFmt/DCWVB/wG+l5E6Ef8qa5bE9yGT3ybEOlWI8LJpdeUQV+NMI6Rm94
NCto2Icg+/571+jPuJH5+dE0LtjZNRRJindumb/y4S209Ic891l1GqoD3g4SZv/Z9xu21WpQyVCM
QeHDwjeNK02waRWs3pYwcre8sBk5TKHd85mRFrUqalkiF3dO7iCRSZwWFr7deMwMyfg1ALMGkiCh
AOfSNh6pkbmn241j+H+8LYPZ4RZ2HF2ZNBi8rce2ezncGoET7+uJBamTLU5ZCRg8GcfVaepH3Bcl
jcxF3TAKzs04PdbXMkodm1YJieSvOMEcFHnlGz4n0Eua7+czKxKLwTaXVOWzpQBLFTZzEhh9VLl0
EUmb7GiN5rJyUFwAghO7VlqEUM1AUwFskb5kwe5QpFhxK+NJdpMQN5wAX+XzFil/KeUmzAENUavu
z2mR8S67QTYVBmt0RYnKHGKI7uhChaM+U+Ku8il7pHCp+JJvAELaKnQ4WDpxiQiy9BA1ClTxghNz
5JrTsHxSubPdzp7xRZ2O2mS0ehhgLTTcsPHLg2wolPPCEO1JTN3wcScRysLR3ZuubOVVXXY7c5lk
ptCoApZGKiBAWxAxAsgX7zYHnxmk2HZoKe4/W2T4qa6aSztR+MpIhztu02oAVtH60gRQ9787Ubbk
EEkY5Qd4NYs/1Ip933GbCCiBEqjWDkg4ipOYZXjlAhz7sK8m3spUBLRllTKhZ/Hii+9jpGoOYg+/
IQ1S526rMXsHBEZtWExf3Sd+k6gsX81e6uO/pv73Iq3kjzcK/fE7JqeIGbCp0WQcSg02t+MYygFW
d1eUkNbd71SVi4EUfWHXjSa0Ij1nOkrFzEDVRcCMiUdXCjnl9pL0G72+B22ABGqVHfUrCx8GCfCE
9RDq63G8nI7OMByzH6ht/OJXw6qdOCortTSPnXQjSJJvRm+/MIpWTUG4gCJuqaEMGb7T2kUwpddW
DRgAk7JfPCrwJUyPGv40MIP0FmLmgkEhToDjx5CVWNG/xmqrs/DUEuLN2+EzPfhfAtiaMgNu0a2w
rYTVhASwAICwLv04C3LSopMZRu5QVA2VFZSJnVTsE2I4tlizLPOjyaTcol0yIycsHZshe1s41RA9
PNk960RO1rCCoEx8DCyYEQJLD/9vDCce5ig54N1NC+0NuSM/ytSmJaHEFcW07ojgLxsvwB133wu0
fn9nEqKEwBsnVPwiyA89lIHTyeARf6yY/NHU901KrUd7AE+rjeNCIwKNrz0C+sS56Qj3xHvUwOrX
Nl/Hy6eRoKB9eIsX01joZGOD1o0EI/7Gq466T+WQDIqOmX5vRuNEvuXwcGd6ajSf40MM5crICOeI
jIA14HS5C12bCfRQeJXILlOUTeuS8SlIjtkloKfH3zrQFNH6rUexLFGVa8w4MkuOEPPGl3R+73LM
8sfbzRdY13kL7ESB+Gh51LYpmEURbnqZMt/eh63iBzcu2hcElETqvE+lhxzLhiNbneo96EJgxkp2
gVzIVzv5qXfRlo/zSrEbj3VK71ZmsLk31JenldoIZDHu2iLGWLCFWiHaSPWAIYyxiH5JeV0O6qrD
CtQvlGTSDqyWBpNrFMjR40q01MBYXdEA44/sPaBh8/Ihk94gwR+MvM0F+OiefNlgmLNrno32pdph
Z2XEZeCAJDTPLHe9aVBFcOvUxpF3E6v1G/uMRXjpkDe6v9OXpMcLWBsmcAH6IPLMsaIZWzqhqCHm
K9g+P3/gzOXR/TEF39Be56ZjCqjlnQvv6KEoL3RvevVvDOizz43eegIh75jvFaIt0NmRhoJInV7Z
is7y/VYvLqZpxjki0KMUGDEtiKvem0oVxx6EXZmscjMLu7ntPZs7OfDZRtQeh9ajCMuxvUeLE+UI
llOLYNwn6YVhfVMgQhYK9m8H2bECVYUOKbxw6L8YBRqSMXMr2WCkGFzGROU9SJ5ynk00R7xVZOTH
XM5x3bSgLF5bPl5T800uzegE8OXSJHJgxXNWfJk4Pj4mrKlcHrV/i+gEqHwZrVYejf42mLZwPaAY
ji3kvr8Gikl22+WooyXl71nsXG2QHdA14rfVhZi3AEglsxH3PT8df3FfCkHh0d3QdgseudIoDpr3
MLI5JHpgHLiaeQUYAAn/MLrNVNF8uccezJ4IoiqhKC2IdMY6X9i3ymU8EVruJkjdGdqz4X+9amyq
mG15DN6iirOfZQyHT9fuIkU+t7goNuiUpZEBjWnhw6/rrNncRgKZ8nb0tDYAxN1R6B3VzkT78bWs
hsDKQ6DGxONK71NsM1GvNd4WQ0p3RG8qGxHhJmq+J9oAdDSZibb08pKe7Fj3/K9xLPKLw9AsPszB
wIGzco/qWvGHjZus3TbrFga0/5aBW4isStejqU+Mh2zvCk9zw1HRiy624xpXTMd99J+uc1CsueaH
kbFrakBSThGmv3irtxDA6pF/dNWy6bDT8vxbgWhtLmKk5VSVHaBhw/LVLrHR7AuAs9gdAM75dmU4
q5Yp8/24Clg4VyUBqmBzg1u9o6SiYxlG1YchXRKD35mni0ceRz88BqloKt+GPgBEjtkdApotSlb0
8akhXVsi4DRzRtpTiv/w4xW1k4ui+5wxhfQVQRTqNs9A1LxGp7RktuRwthgnwRsNM5HQuKD1gCho
Xjb4YLN288TYaBQAvWcO+CtW7Ye8Ul91NCv9Q+vc7+7NHTnQaybLPISt85D1/K3w3iUXHggsBPgD
fEJRcWZ6TWAciwTZKycR0PbpuGGhv4Kaf6DW3KZycSQShg/hH+DpKjG1yIcgQkS0KBwhsDmAomHg
/8kaHLDT8AHXU6hRBwxuc9pfzX2lqCgSEVq0sTVf/n8cPFrCwPKk7yuasBkM11Aj0+AfiIDcVn9Z
rxYtJMmeOPBoAV/yKwWBDvPWvI5kzF8H1mbFcT8+TBRGr8hIJ1wKqISo2xl704haUCHKwHjxqGyd
6DxE650VU8fz1oNsemt6+jreOlKjtBTefyuGItTpiS1cIZY9cGfBV4FnCxNqTCsRayww2nd8n7aq
WpweCKGqGisAadj2ukQRAL0pbSmd1u98bj+2b2HtE4+31rbtzb3A0udfL1gRRqsT718+m+UEi+EZ
zkHVxuwhXdGQQi3mqt3iJHDUcge2HDm+lFRtg+5KNx5FFZLDWZ9uhFySgurDQRX9NCPgjO1mJEQP
J7gCDJHUPDqiIJnpyExx3yRse374bnRJ8dKdnCmXkvff3Q50GUdr0I0SJbYNFeX+KAfNeNS4kT5Z
Xhg6lDgvo0kXKFpHBL8zL48GC7Nh1RJShC/+6lWXs6N/GvKdyeohszlDRwyTCjFQxs5z507fjSkH
SZGwtdEy5BpskK7YNpOC+6ABKYOFNXZbJWa/kiz6+YqsywDF/URRaV7m7zDnEM759m05jScG6OH/
ogL2RQ1nl7/jhPCiZh3tlDnyz01bJREU+GXL4JIHvJFygj9XmoC/b5xGB4yb1PFN5bWgB4vfy5mV
hZhKvj9IOHOGnXKksMCvH0Bc53Wv5U5mVoK7P5tDnDUIeqTN7SwsKXmMVgctVGyH0BMcBZDB5cDD
9Gsd8dfeP1Eg9uIj2qkic6iZQVxLhr7fx1KCvvp0iMryZWmT4YO6PqlXqSf2jsQpxJ30ZLwcixDM
ODHN/cV4A0uGo7X8+VMmF+yVEDysf+TzVTP83le1phqwQtA+xApqPxsK4/oroxddza08WpZLKJxl
VTrHQZvlma3LeQz/cTGLxCgTSrh4c+2Hoz0H8tT7Frlfn7RAZ1Az2b7YuCwu/DsBUANsghFIkwYk
qEt31JXVT7WX6xC/Hi7Tt8tQSWQZdkfmEI9fy7DCxxaiB5AeqPNr17ANIrOdVHaceinDPLt7ynFa
UZQAltlCfiD4iz+UvhZKeh+SrGgToR4sp+xxJyohOxzkqTsGuWyl8EnEdKGNgaDr5JrzE98sfurv
DyNI8v/KLmIy9jMS5aIRa1ONxWT9pF5mRAmahCkjZ7ND20YEmtBqnyW7aXoVVX3LgCseuZ/HlY9h
fm51p5eeuKX8SWA6xJYW70wWMK5jBezNUiA+NBlvhlSLit8WBu1+/iD9s/0bNZwphkWCHeBWTUSo
hmARod3PQUGHPju2TBUixr1G9RUcRTprrPJjhwnhYviWSBxlmNjgFbG4cSI6T2wWBRZadfKdcia/
MRAO5/tOFidJyQm8iJsN4sO1cIuRzF/MtLqXVVZYv1CgF8cF85I6EYjqrPFtcuR5lr6fmpKGDbkU
1KgtW25i4d20z183JdTG9oixK7IGvaENT6gxaVOxHDguYhgmui1oUsM4y06tFB2sXpsp0SCni9IT
HT8fUpjjHlkb5otRbMVv5yZ3z1tih+h6VeM5ktfEgGLn+afEerISWD1BwxyhgktauhdjkImse8KF
RqgLHOhRnZtkT++lr1rk87LOdzqbM7AAQsOq7i35Jp8zApSDEyrEPPekVyTI/Suy4L558XFK3c4A
jSKu/r+gcipHXqaHl55q0DqPb2J+Lc1FupBcsSC6mHcWodWYmKrELVlJ98jpQX5vYsZUW+FViqE1
IVO2qPu0F3I3o9K5FDEWHGV2pi/lESNQSRuRog9dbO+SIjmDSkcjL1rakQ6DprXrP4CmKHpw9M+0
aq1COSdQ4ee2SSmWrFzgVpBOlUc9pE5JGDp1pIlT1sXv7eTTgVDdKhgeTkIIs8fXvQFa7jH2aIoc
mbT6v8USYm3/2YnhO68HZ92ixF2LGULbP3j5YYc3gTZlPxE+5feYUpIeY2ZY3AxedMfDMA/bDIEn
I7h6a+uTYfn6PfOpXLIyvcJs1vFssfkRVcnnN+feOXCHgHON3eEfP1enz4Pbnf4kEn5sDPV7MvCX
6l3ejm/q87opDp9OHZl8jXGMqlb+I0voF9AaLlDhCLmOx5FIQ9IX/f8YjS/aTMo9goVV+udHjQL0
X5vrYCqqMo6AWPYFB2CTZN3bq1/a+EAm1aKbWZbEY/WqRYrgn3kG8MqQG8LduGst2Rc7djSFZu0/
6/UaEAsFQfMZtsnxMvgGY6uTLmQWr0NXZxVyh88AnIUVJchAtDZthPgj2nooAIjzv+WqPQISl8Fk
vVF8VdKUT3kKw6IL+YnMyakH+pWiwsD4mayShHahZzlgTOqEH3PEIr8q/KyF9OIhsn8+mo0BI7MW
4ijw5TJvySVL37YXFRkpCjjlQp1nuH4TBoF3d6Vx/hWP1kL9+rUVtlyiR2ZUjgSseBb81yh0ULkN
/C/yypDPQSMHu7SHKnVJwWt+5hpIfYKnKbZQqPot+ahlXrmqaS86/6Wx/MfDauEztfA9PmzeWgMh
Md+To7wBTiArnCxtEpxAdbVIAEJ3ZAo5J5TPhWi342siIVvJgfQm0+8at4GSTrhHNw2f0D1ovXcp
hSWRNJnVlL2xtZvUDvwwWAEzhyJ04ulmPBS4gDAAnppd2iqvT6ZkTGlJ+3c8nHLDFkXc9Xf9RjRy
JMAz0eALUwjusBJ9wdaCrLfgPtKV3eswKGLukZlGauh3Aeu/vAA+q9oyiuYeWp6t+oVRbrb0LB/i
EYqWCWasMeBJ3NpeQWn7Wz/qugbOCN+hw2TybI6/gTGbzdle5u9JoPFW+CocMcW00wBwH9xM+OF4
55/xK/qV1ipUOLo/mwuTvUUj8f6RgN6XbDglH2n0vdR17nwJgaewCrcrosihPvLsfVMltV7cOMt/
mVeFnXxTmIQ5yg/O3ArRsSaANpY7B2qiCqWRbL73hBPEuVph/OB8txPfCrqP6OT8V8IgIBiQLhRc
3npFPoioetNmEHdEf3gFdeCrSgX1vzTOf8VWB+OT5JCXU11BbfBlzb3Gmy3MD7cc2C1V3rCXs/Ha
c7iXLTb9tJOi++n5p6xp1U1zqXexXd4ZAzfU3aFN+6mZQT0zLgUFJU2XPoB+8sNDwpXu2D5GYyUb
vXlVa8jFI1s0KICOr/0UKttD2kvuOlW3C+Nr8oaH+zaaRhxMkHZtZ/j1NV8Qjl/cIngRvoPV6Que
ZWmXLtejZp8r7XLtPT0PlSTTLBdlj4ziwS0tcYBUqSA45Q/4+4SM5+U/bfx9JozzMst36ALtmiyS
lvkZ55vDDjaUD5y0i838I4uODSTtSs+Q7V7w92GHPGT49sBUq89/nkr/RifPVypNEJBcOjSto8LW
w3wH/LSvjssUI8SBpR46e7eSa01OY2mSAoJh3ELtTxC9t65vKoZZRSwdfqRrgOtC8pujAoNvPShp
+4KlVZesCq57vY1Vs0uVM13DsAVkQqNMaHzbHMa3aDQek2K/7MQEM7BOds0o6PFdjzSnxElZuIOW
i2wR/TnvBdPm/VF2DwrJ50fCRNPjTagawKQX6cLBNPkJxKXwLxxsOhO3pidMMiPicZ5D4BLZoqIp
Dn66upH5tI0l6DxxD5NqtFry4nU2rCtokZc6nPzyv2UCn7TUqQ3hp4/GD2bwTLx+R5r9/Ey0nqxy
FTs4pVJXa++efCTxbYtKInCtIniySJWJL6bAqHxp1hWImcEpj7c7qnM6xqJDAyHBR0ojZuf5tt6z
HiigETUm4trqe8zW/sbaI9etDfZVNV714e4SJxxQIsvFxEjK+mVXcgQu5hdD9DmjRGBRDfvJuM3Y
4ODoZsRostGirTQMq+DvirDR1g4+ZSDjCZu/WLbRDXvUCyTFkFYFfaGAWo+iLWzpx5WDXXZWSkQE
LhxFUpq31JstTYcAp/duceBusgjwxTAQGWBGqr3EJ3x3d9euZX2kw6riLjq3Dn+CLbW+4WDDOBbd
tFU1J+HNkQe+7GPJfxIf35xDCQOMe7TmEaxn8465ZL6O93aVW1fqVIg6PgvVypijoLnyY/QmeM9V
VOLqr1HWI53NxoGSahv8zL9iSnTYxWidB+g9BIrXKqZdvLVtTtUf8AkgJFILEkJA1uUfzyEeBKUb
XKG+7sOrrprDHM8jdO5gNRzmEcsAK548unCKPCQRy8uTqE7YrF6Q6SOUYcZoVsKPhHQ1FZzhdzVO
t6uokoI2M3vHNMTNYYTpr5AwnK6LleTQsnndhfS62iYlfw2KqwPFVj+ijdAikm8qP/eKzbu8DHXy
kPfS7Ic2V4RnGWvEblVBvpavYJTq595aYlVT0ogGu5lhN1RFVQovl1iTWu1/slv/JmWdWDUV8LT8
WzbVS49x8I0TPjhGmVCt1LVrxdkQ3fT1/7ZDihFBomZ4e8FyUNvI3w7fJXsMxUuUL5a34Dy2j6WX
4lzpgEmOel96xNQ/3LzkIzdFGzyazNBZc/oujoifacvYF8bc0+q6rRM2jwFwDNJxaxdqkg9G2WCk
x9ZxB1GMYyRG0isZkeU1Z/8xnVKwh0N/i+h0prvIdTau+Gf4PPW9izPTZQSQ9/Zese6CR1UMeQnV
Q5itxqMSLx6lyYYBcGMNDrV3yT3pbnDcUhuDMQZShl9OMu+PloOODDXrBQcxcK2K4gGmWLeVm73s
5OTgF6Hj2mxNo7zgROtYShU43bRVroqNl26hEFQjO50l7b9W5c1CNy7hjTJdtBrNIH8K0yUOB+hN
/7Tyk4d/7OkP0FHiU+cqjoFj4VKHONWwj8Dw9Nso2rMhQauQWMBWyesbJeg4fIxhdjzmstA6TKxf
+HYWjL5Akz1t74ffW3IgoNB0Q7Xq76v73drQ4d40msqYOIAtCEkox8wkf2tdb9kdIQkR1TCnjKpW
xEvO9THajrQPrboL1r+KAH/ChKpBzML4wnH3IsBiu2mybmawc7w7MCzXH1vdbMYC1L90KtB0Vywy
ShVYnn/a7/aFSRsNnOdn9FRTUkxuZjvruhZM1NAxb8D7inGqkSoZxE6MChPtEguCGmzhGsuVuzi2
ECNYKcY+y3Th5IYa+wn+PiSwWw7NXzoDCwqpHTVsqWJfEEtAYBteMSvA7oEtcf5zyrqqvdcj7sO4
vN2O/dnHCIGlBVFGYZfUTTpRV/8sSaSCJoO0ZN2c8zDBt8+ppoUfASk0UnNZORyla8x+g9eRfW1t
/KlEUUgl5GnOQSVzh2dZUKYrkMB5reLN5yTdFx6CLdHvidhEamSYAqCEBN5uula8+sLjJBxbZUXZ
/ggzJXnIbpqCyECtb8Qyz56bH0D5cftwRua0NEBA+llXX1pCU8KkX8Pg1PLRiMfkED8kH/qd9cY3
zzD1XXMfXwutaGWL0TFZHazNT5gYbLOPqipIUiuHSXlHxuxqy5PRh5x8tEUcOpX3mxHpnUkdBPfB
qTLUtfdV0imkSwldLqEKwwJO6DVXG4fDjhWQ9GK0Xu2keehbNzJD9u03Oq3+LG4T7wRKup60yeQG
g1LmWZ+EBb6KqKxni6tG6pqY97c0O/Sk71OfOIbxxMdEY/+B5WvYExrzEGhBa7nTNi5mqw1Oz+Pb
FQVYzMxgXYVxpnsknYTVPNH3WzM9Y8+JoxdqcUkjonlGsmlBpapQ8B4jkGMG4z7Ef2L9m+4eOvqC
2PJ1+HuucLEKS7xKpI2vebulevmQB7EPFerpts+wRbXb1QPtSLj7+ownPtjYn7zIbZfaEYH48JM2
kBDMofgm1lw3UUcPG9syz+6GlgfNkq2S62CrCwrnE400yid/4h0Mqz5DQq+aqkXJ8OAoDd5UIp0W
GCoYjzsL7EDP1rlzbEouO83a32BptzhW3HxSGiuyPJXO6tUCP7qfGUnrwmigAUXUne58KdfJ6vnI
1bwg4l5ubV36QR2zzGWEkPEk3aghnlvERVorlPyolXeiu993sbSlos/aTaAk+RtaT5mqLDQzBlOe
MJVEDJWy6D56vulQD+ZtbrcXWzF/Sdx4j7eO0b7oXBj9RSlw1gQNvwSTZsJV4PtLsb0ms10VW9TT
DRPIuTwFi9L8u8DMun0TCoYxvlyK3dmXTJpawg/XNitTCQTaeGWfAeYicNSUowTqUX5nzS3hSHXg
8CL0Nezu2TDfijWma3x01QGwiRAW3pRqRT+BMJyHYzgorrtR5VHZSZPoHPvm5tRurIzv3jhwnis8
ViHvGTOxQMj5iXEK5fPfRx6jE2tySUTPSb2C0VE7TfBsNxhYbKPz+n/MWfyNZxpMcPAsRsrwZR5v
QNEqVHk0QZ4tMYf+q6SOOauSH3MbQm2ND75wXlcLDGF6+n1dVcyypIjtUtieJmCTYyV8fXbIxErW
T24UOuXpomUO4/EGYfyPqzUf/kgViJ3t4xQp+Sh7wciXNx5rqGmzxQb8fWZ5J4cA+Yp39DXv+6+Q
l+HO9Fjrzisp/yJ1dSbbsjrtef5i9x12OaQ7aqr6jBlU2Wu56SCWEPcZSj8Xpt/U791dugDmYv35
IReDAHRlB2hoSRQ6bpYxrkGftD8GQlabRVPN1prlRPnDVMQyrD62KdTqjVQys84Q8XWvy5ieuY9q
iDafzd/ZVHrMBXuWy3UccPi5vOkiKV63IziMxDRBahRb4u/jnC/tCbxehIyKCUQLz6RF2GuWJfFl
RWXGdYQmHPJHk5b8swWHtSAvehIK2H0BNpg9WF+FDRUY3D0PGHkPWqvLLNO9L4muuprgEcUdaFZa
jHdxjCEG7meykfAmtJFnKUxSB8Ia6KfateLvj9bCXgLMRzqeRjCmpnBG70TwV8O2zGW/NKad+Git
UIOSQ4ersFHHwbciAT6C6FCfqSKXAC/T8OVyudP2+Rg11cMpnzsJjREAMEoNOW4ybRIe0Vjev+aE
aeY1Zga2xi/oXKoBK/i+9ArllETkspue8WyHADo/WHT8myOwAu8M94/azg2aSVme8uCxWdLPOtOk
Pw/gKYu0839+UQufsKgFg8RpsfVyxC9IQnplAcxjw1gX+8u8FtvySFag1hJ0LIesNKuwgM7dsoJW
N4hOBe91ng71OucDcyFAcxFqbo4ms04I5DdXjm0eSCtw7mkqxdsWSOu/hx4kUgfpQAmL5TMyx4nl
JlqbS0F9x6grK3anObCF88G8fheKxnr3JqQC3aZnm67Qz9fGtxRM95NHHSwUxQ90RYzxcdc9oxBV
npWysP0Io22+JtwUuIGpeBP1zCPKNCK3LmzrdYb2RdWs6F8GwJQ1/cHx5hn7kFLJs0fcAbkdeNIc
Mc/vz2BFdwK5D4HPP0qwJLblnhGtFBafijpq2aRphwcHpaZ2McWJUEuiDUXGeSwX9CdbY4jriXXr
zMNYYAwwKMyeg7BK5pVYdT5KH85wnsU5OMREL29k4Hj45Ixc0+mY3HS/3ZKAjvu91z4fFnCTjA5s
s1CAVh0+qMPPpnHXs63TF7JMUHRm0AmjPKtae4IeCriO+WMtcHaQJF1joaKWomLINdvwTwjZcT0F
OY6G7rXAWBXK2P7HpCA85La+03Hr+pbj8HbgMjERBh5cHAi9qFATpVgrvvz4o4nJ9pTvWRYaR3ve
9XwLgPXduUGHDXQmjjTR/RM2xK6c+6XYa1fycgEBSt04SliSoqrDHPFbTUTlRVNKQtZ9+zZD+sl2
JZR0FTajsd4/drszepLIn0T+ibm1av9rTaC3DN34lUd1sorsijjaaHqg3QPiE118I9enpZ1EwZ0s
qAYEYAMhCtnkZ+P6UH16Kz2iewPeGavHbeV8U92lT21Pt8fUNdJ4li6pMaAbxqDkoAk6YE7B8El6
TvoFjCtXZe28Qjt+XESn00qFVJW60Bl111fGEp7u77Ht2g47NssCmj7eDCinhtaRFFYJC729kOcC
yBuDwLXdJk9j15sI29a/jgmuVz+F+aRwTS2f8yxiIpIDlfR0f/lI2Fmy/v2vPOn6ktBDy62SyHDp
ni8WgT1QUgln/+gO18tXKPrMgnaRdmZvTCsimPhIPCw6QE1j3lyeyaN67lQcM/1ecdMZW89TBFQP
1b/Fnzeg4n42ygVuKWaQkRxMDyqpzQriYOw8wS/PA2VrLy71ovXkjGlkn2ZOZVHF6HCcfSLlQaEc
sk1AS2/EJsKzFTe/X03M4zxIwpBQ89d8Qt5fTBapeRhJRGYRDIsCvQH+u3LFWyr+ihFyZh2mj+md
+wOCfYlbCkkEyMVPKuHivTzh4MKq1JwuX/Fp/DvdP5QQwLGLGuJPQRJnwebp1buM8gG3j3IpgJBj
CUaSsXHoRGC9rdcmH6vMbqqbrOoUxrKNU/2w7gq86TlglyC7fH75QenqJVDtY4uZGNfWKy0lVpb7
xCE3IlPxaDZGBvw24SN3kGaLcfg7+glvHRrGkfJ7nGv7qNng4edm/g1B4g4bppdLI0NrE4o8gPOi
p6rp5NExSlKOTcneKuKV06g2S+h48IG0IvuTiXZLk1Yl9ADAxn/baA+3zs1VG2y4gnK7eYJ3unuf
DwffrCVl1Bult+w85yNz59MESKqkhNPKgIikDJQJX2byCqc46EWQB/E8kJEwX3Iq+m4zPp7yicCN
4x0dzIcloryCiJfakO2eZfSIXHJiXal7IKdfCCQBcTEJ4V4ojLPPhgopJ+5tvYVm57XuDKYJzVyu
0edqMrLAaq5oQF4n3L9TxLGcyYh51l6fYgSgiPY48R9WEb75AVbZcYkq8iRDDd8Z740NLu1qrgLa
wl5ieR6Ipqdr2w+cCfgfpnI/ZSUKF9gTYeNieaB9unIwvDbq3XLtHTHTVhkdYwNwqreiq7Wo8/mf
VxeKPYn6AAQ/UfailMy7xYjXA2PdWKf3dsVfzv/nFa53KiARkl40IHKah2gzBwIfH6iJwAWWMvH1
h389+Wehjnh1O4ivUTpwNhzOocV+V4UoiK5Q1ZqUFaj/erwaaQWH2DHJ+7SEZf52fsGxNpMehDZe
8yhtzCjzbI3Lr4fVUDborbyLCoc4feYoP4tRZIvgHFnyMX4pC5wDI9LWnOyNjxeGiUwY66NBoLlf
0X1Ugi+tEVoDHq793u7SqCS7PegmO6XT5KTbwQwk7+oMjK4vT5S6egz20Z8afcPasLBfImTYPDd2
7SFDxdvJMqg0QdhlcvpyAIlB4RwIcWCMshBDCBoBTa0OmA4mDXHZnM1s9y/yhJ7C2DfAlp/JT4cB
mCM1HewyyCLRiQ1HJchke0fzCz1BZFV87/9v8oBjqsqQn1Hk7toSiAcFPTEHAlDlWS3T+E+aV0iL
VibrGXBzarwncJACiRdEY3FDjDUJSVYOJB5/NVje8qdduPfydXtSMNNIc7sXQxykSNCJKI8T94bj
nQ3uDEtcGBNDBrWOSeEtHB6xZL0WPj5lQgGwQcVxh4D1ZNpkKrUMo/gSQCguvf/rodQN3fhdMu4M
p61mpR5uSMNaArkcEAYUgh1u+70XVl4Mry39cMJjBggKMtno3cQKDAdYmBquFTNlwubFlklyuLcr
B4qtKA9bZxrgzRI6S9cEenZVc1f65MphNfaPX4ehS0DhjKJe0QBpHiiQ2a7nyd2vgc8qnWH25JNQ
mzMsqeJBmhLhEY2yyP/yk+FG7XOe6xO8iTsbsv2swT+ZJF7FWGG+RlUWjv5KAA4ckeosZYow8iyi
+dp/xpH03b0Toz4V/olDDSD17NykG6I0StM0WT24cLbaSHxC4LAkwW8f+1ETNBKa6WzrpQd1LMN4
AR4i/ohI3Zz5EqmbPpBArGIG8ClxVJQmh8sI0zSmL9T58b8KcT0TGwa1xSIecj08eFUwgqlpJU6V
dcWxIQZgStPhVhoLNrHrJv8ahGYTEBNJVhrbGAKrtMvWl5UEvJOr052fDSB7AHWj9OHzF1SBXOGN
jjmQMlAQegM1PNkIlKcwKJd4Q3RGBF/tV5u77cPmnlXwphBHyYQio3ezPhMs5cZ14TCF44z5gEkU
qL8LV1Bap4yjyISJPr4DNCoYI6UfQgfW6R342xTvWyegL6Vhpn17ollEzSlREBgfqD0bzZ/WTuVw
NM7k+CF74RbkSteYg6A5cg0fWWVS/EKz1N2jsNy+v27xDN+S7xeRS5CsLVdpTfJj7KOoEnYYGfc4
YLImODiOBvisJg/CL4c1L5DTiNpbWBflIohkFinlh2H+137EXtctSwfK1JFI1wyf6WB1pkZ72ozn
kFg68Yn1aJrnqvvR3Fh2zo5e5DU3O2ccel1BDE0FP4TQ58z7ISh0vMQz1SRhXNAvQnBwIYUzuSUt
5J/kAlu2wfpK/cqISh5wD7f5CY5T5BWja6hqc+PiWWKD30eCmNL9lXYN+g+WSqr+jVMiPMw89TcJ
IQrWNm5eDdSr+qECytqK/8cGidses65GOVPmuQdZhHvUVzx8Stbp+fm+VSMFFrHSjKH7Inwrl9uG
3S//oxt0Do7x75VDq11CezI4wnKrb5PPuzyBs6WuyqGRG20YocLupeeIux9lzqWDXOPeu+znvwR8
QgEgufPyjdktRc7oAWRi4UwoxHTXtlkfAjVdFaUx0m3E4cBHLjzeL7jI2Bs9TWiD6CzYEX6YCLAC
6kdGAPHZffiKgMcInxzOWCD/CMl8nEto1rhc0rfdemDBz0oLavcbGGa4f3iCe0z/c98QSQ8Rf2d+
4D0DgBSTdVY2ooqM4ru+wM4+2wGkciLVuNjyoOnpP0mqVyVArLXYpvNTUiMafh379LPrD/+m+wPx
nBp7vVMVPLpUxo50yBZVov8cXp2FTsy2urrHBdECVPTDXNXGfTd3wzlL7KZb3r9H9CegNxnXIw19
9G1KdcFMvtbNQpj9/ObfDmg1Yq8VowczL1p0wkCPWIMoGACjBn/9T4XmppbLUSC84MG2qItbyzoY
JFrXlBUONfPrDM7DAPSZZ/qzuRE7smVOdJPbudrjk3wVMq0xHNirVAWusEgQ5mxAycHPoCaGEbjG
ykI97f9I46WBs9BNDlPvs9kwMVnd9yvijsZh+Ux0/10U7PAcb32kflXSCFBGQ/kSIzrhUOEGbgU5
42vX77IZN4F4gGaPhfA3UgMPKhzeAc2ammEzxqmZ+m0b3LVgwXyUHtOSvGqihcvNrgJrwASYbSoo
nLiQKiHNuDE3m1Zwr+qGsGHyDQAbnZARowh9JwaijBR4Mz1teNrmx/M4bJejjFKUVqFY8oFeHTRG
ThhRnkNzPZQd8rdMMozsoM2vWKbbc/q1VQEq0kYtNaYtIkZi+VqPGyaP8U31CIInc5FKjOe7YWsR
/5CMqWNmVDMJieV/I+M7hjM8xc+No7mdd3CYqOg0wrRg9MQ2p0GxS7IFQ6+mT/J2hxKv6tDCnzyu
E9/OMx9+VRfgeWah+Pj2EVHfEI+pkUmM+ipNbNPlLs1m+gLuhkns9BitoVmnyyIwccW2iIAQtMGt
UHasQsuKyrF6DbMkLPrpc4R81/Xw613tGIm+RvdnCtIiIdOnKHHGnYVV6VuSNje5Pj9Mxmiyg3SL
lThRlwweVgO+2/Jecec07DYCZdMydomWdpX3iUZj23/uXAei4hJc0ar18Yj5QFqkyOez20dkUX4a
JhJ/f5bnyutqH1b0sogl8pVNtiMWpf0+E5cjMUZQ1OZE1Zw5bd3DXEEQmc3BpOsbOyOVsz8XrGz9
ahQbht9RT2Z5bmPOekyytbrZ/OJhUyuZBZRragCGxibBIXOsXhmDc4qfoMzQ1KkfbXqMVgyioxp4
XzuX0N1aGQrVke1xlfsVJRLTsFQkV+WZR+VXQ5/W6idVz0kEiZ9QMRDI1EzYHpK3MlHxZtwsb1fb
m3dHPn6bInVvoREOpl5DLFRI9Y+MfipcNYHHq+xB93GeUq2go/prd9bYbIKkEDm+57tQcay5hyRz
16xtcuUly3aVbr7OjzGDx3xYTQuF9SjATh8UNg5SQQBEpDA2CI84NwstTQ77baoQPOEK24H4cvGO
vnF7JdlgtIgiy1A77OZL4gtd6qLcae29ZGyOyV3JS681/Y/TC9jQnZKedc6CDoEQdTYtyKIUs5vl
2l2FYO9eQUUFbuMTxmF0NyhIaJWU3Uwd1Rvg1DC4A8l1IueSBH8C9cuVf8CGFk/J9mEzSzOgorbY
eGeQ4Bw5+cFFz3mEvgsA4w6gqeEfb5lFHv0GECo4tqX6H9MRydkgclJyp9P5D1fZwrB+DihCzGuK
xibQfggfplgpwFbbmHT78gd2ozC44ZYuoFnSfi2lFF8vLutyZ6qapDjZeGucwjkTzHMctDZkMF1P
wC3wBD5afQXtKzzT+M4myBtxupsHjBkSEHf4kiJtpcGGjZAdd+9J8aVDfPKL9QTRE23ZfN3wmA9b
PY9qfyNuIn5IWjTmK4bjvLPwI/Qizkt8u2JLbP7dav2WPSYxMWDgo7+K5/3q9mP00Y/FTpsanXEa
QZhvM/NEix9KiCONwetauuMIUN4B0mPAg08liopwJz17W9Jt3Nqg64OnJfB6bXy/FOB21rm11Bvl
03hhjJi4xC8X0SKipJSsfV1ksUcTJrjdVKopQfnqeJdGuZhPZDakxkLEpneviJjkgHyvARuOF+2X
z400S16duaLizMqp1CmtAkLt0JhAZr1Zb2AdoyCHZS4zZwF4GurYO2Aha9M2rToLeco7SRHyjS+A
j8BOVIDdfR65ItvY2kdEcwE+CW8EFSbC8IqNHzg+hoed+iJnBto0cjBHzHFRMuhWsq5WjrrPwFgZ
f2YGW6e8+WSF3u5qNPXNtRDmSuavciCnP9oeBs5x4tN8L8W05WGPUSZGBxM6Xce7cZmpHXRQP6pi
iqJPZz3laLZkrqoX7+TuN5hyjgznDdbzbGjcnTXkR/Eb+8B7eMtsD5fG1Yj8G6bCm/zlrdRQif9I
gOIdJtx2A38C8F0JCAltKF3rWUnvtu9yrxyVHJ3MbMY8chGl7Oesnmu8Bv7yNc2v5vuFagmVUvOb
P1xda6hVxb806cS3voT3A0AoJ46GjxMRat+rKRZdIKRn7i1sE+on6a+J4y911r5UB6uIx5AoZWjf
PzJWG6FDUGQS4a5SMYM0kLPlyvfrF5tp/XRf8MsVk0F4njuCq0C94GumpNWZYVBFfijoWjbO1j0Y
kXDxyh/ac3IMUARh0Z5n0E1a35ubvodClcxbID1+U4T7S6JqDrOPVtaojZUYIZnaerEdGNMLEGNl
dimTy2EiY8uK1YHqYBgROgZ35X1EcYzzrwim8EJqtWbJT1TS1WTtdup2hLtTbKG5uYJ7VV0hcB2x
DPtH+hSZWSznJmjCitOBFmE3pDHSLTU3OXyTRAFuPXmEA2l1q2OlLp6SGzcBbW0bWFQxGPhS225n
xReEHTlRB5OL+2RpjdDNzOC67JWukgiLfD3umfzxp85hc6I/kPKil3Zqkn306TOdWLzr0Yb3or+J
v9gKV+MwjacW/KQSSrltwKnyrnBjx8yKH5BduoY0vTxP5E6i0Sr/OBmr+1jDJC7QVoq5BJBNJXjC
SEfR/tBGYlaaakaHNmq+32wxCSjcfgUQe2rm/YKTk5f6zaPqgun9xVlesdB50Kbe+X2RYer+P26A
R/YC1fDsaqZrttdtE3aWfMSI47lsGqOrQb5aSzNBL+2/H5MlAASlhKlADJtqs3u6dbcXOtwrTt3U
TSREskLbudzhE8vCqzLAiv0mWKqZadkGG1gBAgoHYLjmGjtd/tqzKfysIpETrAhohd737sNjJkX8
FsS4rm+WXwoWWE26onxK0kBN/YYa6rtNCr+ql8jxckw8JVjy3bHJysyUkRI0F+LlLv1XqwSk2yzN
YEcp+0C4U8hV4YXx2VQ8x3zqsSFOdw+3NywMIXcmreZakH4YLITz5Qu5rdTsPQJnZI4H+9RcbpcS
e12T5Fn07UmlitaQgLsjd2tKqgCksi75EutuSTfU3GzOuORA9H716rsAY6cKfnEfNmXAK+DOzdEQ
2kkD6+cj7mmodES2gHTCUOxnz+v9nGQ2UB1JWzFPP2//bYT1tI+iBRikARfPT65MoGfgm5LFBy5n
YmO9/QcPfTVSN0m8swLnbn/hXvJI64ePzeXl3Baw7E740Dm+Cwleayqh2HL+uP/KFv1ocBXXLEoP
4EHU9neb/7AscPmiMQN/G4ewE0WtENuK/k7UFpwxqLD5OSnwkqOB5566CmldWPCq94a1Tlpm974r
CnvMrowFjRQweMIei6e3v4RyoHAR235iPPFlM9TI40nHsf6IfXFJ/mv2qjD0QQSF/xbVfDwnHrHz
saQxg2CqISYcWtnqBRFZrZcDzlD2a1vTy9H6BcfM+q4zUJp1bZVKKEvinZ6haLy9cvKdc8UE//vR
+MoFEFXVM8T/7u1uvpRRyoh3ZEZyUsdFuAwogLMBqwr1Vjp9x4iMPq3qkNhDg+4/ZHpjIbQyWPSK
zRVcol5niRQqcSwqeAB76oAz0aaizHbMgyiD2v+xzZozGeasgrS6c3W9kFTF8/Q5pzG5VhIq3+sy
Xl4nzfq3+svegbYJeGs3WA5zhTaigVn/47gsc3VYJMkR0/ILszc4HRN8i2HTnwIIlSQ6AklxpK1m
JoWQK8uVtJGl44ADem60yy0y6ToVQmXI+ZKm1Uuo/mBZq5M9e5yS0//1lleCTSsru4MFvM3lqu1s
tOX2IpLhVgHEdfUWg4A0D1LN7rQ8SpR+nzKr8/5UggpBMFfT96y10HLLKS0tBfVds9ov4JJz+2uD
ldE4OEI7p7eTL15PCWalNi+dtMEUy4ph/3FNGZEF2VRr11ZcBt54JnHzqsgxHVS2at8Dw8/pzHFY
PMojTKpWTb5TTaDix1/Sfa2DnRHv/xPvohB63Jc/hQN2SL8mnPmQ+v/UhGcwZG9mSiS3ZTp+Blii
oKyxtBrNm+S91fRZkNBUmDYZaDh+ypqLzDQDeb5o8CPzG6yHfqIZoAokFQfIQM0NI+kG1d93R60s
rL39tfA+EHk3D11+rQjVarz+gQen/6+ckOGr3rLB/c1ho+PBCKXrFar4b8vpmxDh3tc4lL8qApjL
USk9vZMFIfLrflx9/AOTQoyXcbsadPwVXMts4EznW/kuWW3WlEJz2rc8yTXOwgSDzK3eObziIprx
KED9aWZMoswhdHXVHnw+b38J0zw/B3bklA9J0zRqNaSFqOWSiz4YAqz70PqdG4dC+LoRQkVzBvr8
sDBh+IsXnwNT9Q/3b17QbnnXA5drtmVUBnOujACp1tFscKYg7RodVHyOyOM93fPfbfk9dSl/g85q
1794hr4m/F0/6RkDmVBuuML+AS3GomcFm8eV8nUUShPGxqFURZdUYXruA6IewAFW/V0U4+AgdGsb
q36y6zNMuInOIVIvM6ZXPSmbjJKuaY+DJsG6C8aYR6Z50DNqcVZA+CEfkvtkC7FRUn4AKR81s/oD
z86Wec9WMj8gET3pKY46OXCHzKfg4tJ6Ot5+uUmtB76w1tK0jvVD3OZGhz6KtZ0ZqO63y70XFlUX
bhwOjFVah1dMfh+UpA2unj9M/5eixYENXY4h3EOX0DI+/jw7Q234P8NmnKDuC87UXNAnB3AK6Sm1
HzludtY75ifNXCC2XvTeg8rDQbHgzZ4zqJZw7B0zfzSnARHfOd0uiBfshJesZzi+szy3NdJAI9Cq
ZFBrKSaMhwP+0ZM6UdGiDzPNjxINaJhhwFYrLpof+rdSc9duueIPK17/7lYjEZUMCsxld2uUBVGI
xxUxxhUjW4GHRz0zoMbbVMbzptYykZXaPU6szkwhXRA8xR0b8ySBnnIBIsetSL/UKLnhGGP6VNEG
uLEiMP8SmOnuIXpSst3ZdGyPPhBSZZWEXTAfb9xzQyXMPvx56gFtRgxhqZ5+bjG012D1ZN5zQ+Oj
RHTwk2kj51tknwFCZhJpt3zO6UbAcDoP7pj0SV0a8VQz4CNDYfvUJVYJ9Mxg3DYKqAabrRoalGOE
F4mUV8GOX0t2w91PIRRxyaPjriZ8q4j/wPnQw8IRzOCWliU5JaxhUMa9uTBeWlsMd/3XglAJGTcd
MebEx7yQNn2V7x49qdC1wjvRkyyBbgECfm6LBao0cKIuLdaTIdL0HZEZzwpVcxBj8Avhju09IQZC
mkNlHG6/paAM+ZpOx1tA+Hxz8k8ZVlvE4b3dOj/j2YL8D0Eh/qVPmLD5VhIJBgmeCjh4tJRj+tas
i1mUP0MJd8lXBh7NsT0V5p3Yt5suFqSwgkAEudZanPZ60rnJWfEaZarA7ylxyago2MVncD07mvyn
vetDjI7xPOmP2oA0nHBtD9MEu3jVyO9zI27QfSlOCjRIEisPxL0x9+8Vhaxhc3lbnPfWp96JbTzW
D2JGLOSVNzt9y4mcJt1bmHYy1cBuytY1fVsKfcJ02QQWhCCc3blThsH/P56NZGxP/EipPTi4Ty1z
PSuDKLsPZH5z2nTuG2F4w/BmyVhhW9CWHF8M3S6hQBQl4TFM/05rCXKyuQjMwgEHkZAXb7A7Ouyq
YDg82Ou/Iqm/HlTCslWnoQtaf2aU3SFYtC8blgH/DXKMLhu1YJuyJZVoK3S6CoJLKmzg6F44naJV
TRzSXB+RL71w+l/nuNRb6IedLmYrk+WW/TW3qGZoZk6TKEZpdrLCGZzLmuHtvi1dOGDDjrG3yf2L
wTyVYEDLWYZ2DhvLnoOJILxvLv+te6JByVeC0zW1gp81xCnxkh9zeJ7QINZbHomEndg568bg2ycK
Ec2jZBcNuxygxvJPBcxdC30ySI4LPq9/4aneVEDHzq+n8mevKfWG2RSHYIcvtxlMuzakWA+U1qE5
v2dzTrOSToMJvjtISdkKx9BeKWE9Dz1LyfeA+eGWo2dd3XBNRV3BKDMnhhCNoGURmnBvJhzhT1rI
s4JixeQTuT1HzLiZTKxQHPs40lAefGX+BqAMmuuco+El4o6vzdPRIpWHq4wsjGeuoOVE6hYDjdds
E++Fs9njWW7wW/1uRte7iGdC5xGQcdSLG8XJmJN08pCZGZK33qWXAL+YjL7V74SQYMFWjv6AlMLi
Fz6sif/qSal+OI25QLJ55kbhLhwgs1pwbdXQiJYQ8hCl3l8dmzDrXCmNoTcaZEQayYYIx+/eohRE
hTKfxB+fKpPokzlJERuzAde+hCTO0t4SV5euE/7IcccVOD5rLqDaznvrUIekS5J9vkWWazHM/S0H
y83xuAFW+6Rmji/WSFnJRU4qWj0+4dWmN6y5YUVXKr3YHF39kl4OmI5fWbpPFhiA/yaJs9CILfFM
wgOk76N5V/rebbqIZTNK0PgkWPwdQEhUkjaYZGO0ZDkIlnYvoXM5RVO/WnWoVAgKrneabCZa4eNe
xBFIYnoopYa77gSuFBD2M6hGsP0Jlwsu+SDqslWoN8bCo6raiLThOBOdudtejCw+x+1QmSvS2ty0
p9zcLEn3FII6ZxSNizEh1QqGxTCpRT6ZDBvn0ryq8umpvnGFtDDBY6l/65zyoR7MGhnLZZaJauPD
O8gUGHYInD5zudwrKLE+OvglzA53jhaEBpPow4LpHek7H2X1R3PWKG8qy23vI/899jtbH0F0bEtl
cryNBxCl+VpAKTZUoioRddTqubXHEQYoPHhUvyLuot2rPEHU6c36L50cdFAAM4VcZEJc98GrpeJn
fk/IPXfmGUlJK/+YPBmvesLKq7TOFkp4iarADeu5rI8YV6GWNQmgv4dT0OUS6w06fdZweHnDVhwd
A8tH3Hw6KQaGqLX++BH30yxu5Wfo3gQsp0EWXK0ZdbMi93Yd2rqFmreaCzoYA1jbuq4PcIdFKCHq
Y/Jhcsyx7wMRO2JVny5sUoSCh+qzYH9+XhYI/xkzELzxgR17lfNloIgtFLaEPPbMzwp0ydvPYZyB
Vs15Yku0Zbuq/+CZivjrUV3y1WUWbsN7+WWNA6nOPoYNvrPXSo4vuIZUavTU7O1b1d/N9FiuTbPr
vE0ARvsthAJNUlMdL+465v2q0lK3bDit2p1GgNAYjmQ7OSMK8ow8ZZXPUpvJnpZC9HVrxPtC3I4Q
B2CgZKx4x/Zc2v7gMzSV1priRqJoH7eKavE9fHGOIdssPtL5kP5RQYOCW3LRL72de78cehrDJ2pM
8/TJpoglhrd+do3OSh9vEtw6d6SEqTwJ84AReNpY/2pE2jr0Q3aoQ5nruNkHca9jbq7clPCg5Wpb
kP5EfGX/e3OEDd0Gaolvy6jO1Y4UtkCZMjjBU4m4WtvBFSWI0dEo42ggxJQ2jI3lp9hnUnKz0XAq
Eijvnj/UgNcM8VD2LtKMLPnmp3q03hJ9SShYUZp1tgsIlOsfk8qGY6xqo8I5EYIseq/nuEZb3Wr3
+0PCTDD2vjCMVoJAvn1anfKOcUnysBOt2Jm9MmkSaGt/XME60L8Pkd1kh4Z9tB2Th0m+odKbX9FH
CIjVI8Hvr8KkZDmVHK8qM5LF+hyF+Jez/a8zjfYuejGce8VedgOWwIkW0l9bfzokuAf8PAH17bMC
2o92lbBxr/olZ2eAiAlkq37hFpV8tmmlGyImzvmaY/5Bbr+zMRkecQXtELGm6puNxH3P6N8dMuQX
ERtEBKzLLkVutiguZnLRVXiWPEx5Mij7kebJTZKs8M6qbgOJj4VLQrKCEAd6uSAQ3qGYudiOLGD5
ZhPzw3NailHXJ2cI+FUDhpSju6W/W8g6LFIPxTkZv+VwqCc1djgu2V5aMuAPuOBUvBHbrJ3zHVb2
q3E++DyZbG8uGGVTmzAPbjt/FzYCG9Ygr0xtxhrqN2b3mMavDA9pIhc/TbGFeTfG78FMATSkDRkU
uA/mdMNNX/MdF52/SMZiZU5fs5nAjEzVMLgjOZP0qR1TDA0/bkgnt2tvI46ZE0HE6vffiTDYhJjC
+IVbAH83tXpquVXrJd/DRR2eH4N8u45QRWmSRNFIXaPmmRcxVl6gFvSTC8C8A/093KpZvoSB2gpa
u9PJMcub+q3EfOsnakRsz3n8YliJXy0q3r3zFpzfaG2v77fwFlIUBovKEcnPxtkedNja6Tba9799
IbsWMaNtxBVY8NUqC0KYNJZY/xNJhCh25kwbO4OC/fAPqV07JuU0VjeA8QwiYKYDHUPIJw8E6yOv
yBjprDlgpSg/yegP0EaKBd5gIBpsngo/a0cwPd34n0LHu/2j3WOPcieOEtcrok7dClXfaJDWi9Rw
VXFj8sSUSJ+fOWCpXN+4Fj38A2w6T9s5Qsa2G7mh+EFiGrFKwZSYfiNp9Qw8bpvkgN6wugWeeLNb
BppYeA8O8TL166BKvsKFuEP+WU8qEaR9x9J+bXWjjS1HpEIj3qZvsCzlkqBKgUJlkMJl+UyHR0Nx
CDtVSpgPENVbc26rUxhBo6hJyWoi89G1AU4dSKNRC+JwFOC1SrFMyE6qg5ENej/IDJ0FB93tAxJi
Zvrb3tL5NmaA11q3G/WWfL25HiTf5moPPiH0JGT6E6OT6dIArz/XC/RNtSPDEXUnDVVy3CK27pyA
Kx/4zdPMs+FNmKpd+BogesVaAUlCznuRMHc3rUkO8I+rDO6mDA4tchMTw/y5pMNg1QRGqbyKOvGU
QE1NC8LaF5yAUQzNVl2eAFonThCzR4PD2+CmI9db9NnllF34fPKwU7Yw1DySpHJwvyTASkcWYbJ5
VwfUylgTB76iSEvfy0cp/3sHZ7D0a+7qemy+BeXYPhbUbFQW3yLy+ZlrNUVbS1ysSA6PdPunl+Cf
eNZsTuXNMUB1kin/MFS0d97bqYxjX/SVQQYJiXW0Eq77AzG8KeWhAU5ihrwMQvwvILhOwC37Scmk
xCWZtmhPOHOuR/Jj5yTwBmuMuETdhQa6Jfg2GAVAS8GKdPJgsSpnYhV+wzC88rCy5a1GM3itmeAS
QTAX9+PNzGyXo8o0KDEA6yDJ958gwiy9t0hFUeUlEdLbTiSwdN90QAhn75PJHXj2Ckw1yBbKCaWn
AEoQlCCDOVeZHxJ0aiK/Xgm40nBFlCCjAJtr+flo+92TDWLsuRU0lLSJsDZD6HlsWObmGUJAO5J8
nQKpkAeh4jOxGsehfjcZM1TOg9UtCr/FKrEnAv5jcZs+pxW3pQey8nbku5NWTCyrXqSq+nqqLyPA
Y/2oVRdXew+WGyW/TYfsbTdpT+ltYTUteVmxHnJ4CbzHh70xtcKWqihQIHhelCK8wdyjuodiy9Mh
rvPmAhwlG6iwuJWF2I3Qfn1AiORt5Gv3ml6u1icO3NfWM1hEpCVcoLndtobHu+yijf6hqIa6Ytyx
zwSRfnZOObzstwex38t5BsLqyW1vYjWHIs2tw+Hbt25ZgcsYs7a3DEQW2ohD/t84LPyzMWQ4c+nn
G+Hbq3vkbPCzPxrMYnNZkUMEY4AqYEgqZpz3MswWuN8WqJTwyES84VfGy7qiT5tBHZlvh7I1xzCz
NVVQ6Npog740KmpzOAeySOnCjspo6eU9QXWOptUTy6jInx2mA5jFXMESHsA+oelU4Q2iPCZSkB9B
WAtgikyJJPp5Esh7NCc8VLxOH13OoAtzLHrHvQ0g6CzM/H5QTzs6Wv/ewDfAslSbgq8hjTaiumdn
rf/WiZHidmpbvlZCJ53h4Xq5q6AbT5f2PlTcuU+MkA4MwbUgnCQO1z2DjOiXO/dRcDHDmW+H54YQ
lyJtttDKthQU0cN4tQuL5tQp/wI4RylX5Kq6ZgCWHtu7ZdvEGro2BpA+IEZisIZq+fAkOhLgHzgi
+f2C4Kpy520kqK1iNk9HdzfWo6S09l/NVrrjuNmHjt8jSnr61ErVQp5NnVspluarv9dJQ9R7uNf6
HjVrRGxMgmCjeBu5vzGcDRDkW82XRrEqvzY86sIvPleZMJi9V/+v4dX3OAMXvWzX4xEH49d+SJwY
HO3Of/Eqi112ATjSqXQqsK6rH5raVMbMT1mP/4qAjC3SKLAXLGDT6QL/xwhLY0BGX28FEmS4ntcG
Nujr17XSzGV32x1nWW5wLuMyAMPCqia+nMIkTu1u7jzqIuocDtXBRectV5EgffyaaEg4Xw8wsc2F
CibebSZBSIZub76cxyRN7iPB4g7dc9TWEm5DODvpLRqJh8xZBpjI4mh9gT6ZMo7l3Bkj+mvBQQLi
ax6QkxUM7i8rHbChhXeLZ37UXNV8ZF7uI7sOupimrY/EKEPO9lTG/kmC3OsmlAYz3Xj181gu9MQr
ZMcPo9zt8R1NVjR226HVHHW7bVdADlT+StPuXVqQZL4Mxh65Yr8503CfrVSWCfLCGnk+uJwD9Uuv
9eAxfs7a2Nfq4nmHXru/9Zhbex6luGQfFoM49mdU5eYfNkZalsmF1NIGasCygEv/GfuhUuiGf5KQ
65ZRIvdpy850nbVWZq4sWpE+21bUqSOGCy647SqF14z8n0vCgz3Uazi/VvbP8x+UHpGdg7+ThVfg
xmTYPkJl4MH1OSxPBcJIHIBnymBjyd+PZb6Es5s7LRZMymzhShHx0laaXv82nyqZPF7c7nEoNEXp
OgE/tJUKmkXyM5OHl34bcu/CpbW9JWR+c4V36Ly8oHuyGUR130r7v1iTqVxxAN0qFDRwxCmc2BAS
RHxdIwPxcfqagPwGIP2v/1G2LNzfI4KZm/frHcd5e6SuPuMlLvShjwgbtO7q0aQ5PVzG2KuquvgN
189qj3qEFaktNdKyT65neOGmPwxVvkZKNdiFAZyNwf92rIRwuQt6g/gNx3iMdTmpofmyk04tTpsQ
FyBmK7L8tHtFLlBgHoi+sAWRHrxeByKXTvqLaLznOldmECJrnR5KrujmQeLRSgD3+cSAtE61os99
jZXjv3moQRChaBgFvTtM1AV8toC36cNEcqC6OJa2nYLEwksbT+XQrimMESYja9HWdCmvjHYcknAx
yJA+ggSQhjm17p9ZrF8+oDARbskV5igHHhbGN+8vV+CNbmh6mTCNxnKx+921vuByoIYl0P06gBba
qBy604feY+UTQoKyIsCJqIf91OjRlb7MoX5Mm/JFcNKmsm9luzbsm+cPG35DYc9Nl81rJZgPL0EH
dPmbC7GhsehtGFEMeGZu16GhbUcSXtiUOujuHn+vjoZ1rhmETLRMVKEgC5vF3QVDB1urqTzQzKXd
SRP//tJSVVabUEQpPTLib6HcqjNwdl8nCdJ088MYg6/BrhqUgt2cY5uupbonDGg9bwLBBgUNhgSF
N70JboqTfDGiyBCQxPTk8LqoKAYUrNeRHYipOQHNplv4MTum0AB5z8uHlNMfq4Uz8E6tAl31n0u9
vsVM8ruSRlsgc9tKmGJouykUdth9TJgGSCkyidsHyIOWTBElUbStFj6PxLMUqPOiU8xEUJpzddQn
HeiVg9G2H5z5ubjzrBgg1migVd4FBFwL4HbZFuCmcx9zHGIMiaTVnGR/u+aBRvXdtjonM53eFe3Q
fW5Poma8dlq+dB2QhH9uOn2nWaqDprk8gUI0YNqkn7ZXj4YRf3cr/kO19MJilt6sJ/wPCWwaiMsV
h76YQAFWTxbA1DYWFzdha0OuqbgUYd95Yi4MqnodJIHYJ6XwH6uB+LoZT0ewIy47a0bJYezWmCXD
mt/wlHX62T9oaSe7DtZhxfYFkBmSOVZpjib6eEmPaAHejv0rQqgb4Pdi+BFcBlcF5UGT90gZ6Mzi
LOMpnkRfptxc5JgIxsT4fBebZPNPXLi+m3INIYUiF1Xu/84WpgiNPg44jgrvbLCw9ChnDS7YKWac
I/OM+QbWa+JpnK13OshY/XWVyL/m1txKVBCW2trve38dAxavbp2bq+8qBTUeJc06Th7KsY6cSxlH
AeL/lq3QBts/kb3m03ezvMmWN5sQGCAIEumvlFuLXjcqkRIKeJtqCJ7Apoymzk/+5QP1s7/D5ulI
Cr+Iuli8YFaq1CPr+PQzU8yRwpk4OZMSmkDEUEVR3lSCuC+Y4z6AZvqvpE/eeWXcBiYbQG+oXfOq
C8cFcxwW1TZn/VjoY7ptQuKPKpxt/HurEbffjQOLoMKrzVEEIIThc3Ehyh2noANWvB0RvQ2MkBth
ZAoZ/9eOw1+NxlQWjOTAp1wQZqTsbcUK6yDTsorzBjdkmcu/0ocCGsBTaCyvp4QhaAiWCNQ0RYnC
OUxpBzq3hNPccww/kdz1/HH09wF90shA3tj3qNC6/r6SJM3FsPp8XEZKRDvSaww+xa+sWceU7KM5
S15kJQZdboE4gYL8OVeyEZIA8m1GEmvp2Va+ysWbWFlOXTzsVEy4jJ0Uq0DKKfWqE4aSHd8L6S7l
wzUmdbtmq2ALwyZQsGCxmstKjT3+oulwuSv7ZjQx+2Zjolkzf2zI09yKR1RQEMLswQfIDrPNiwTe
SEBxmeKl8SXztREDI2B4EgHsC3Tdp9VkWGJckhuqWImyDRGY1QvjmR8YpY6gNoloJK5xNbaBa0pV
hMxHoV1cZqIoB90OK2z2BsUIy5a6ClHdaEcVqfI/zguoN7uGMg5lLA/RwLdTdpnJ2OgI33KKILJj
ukSkW8l3APow6ik6Z0KyKC6DgDdmNrwtwZZ3RZ6Jpm8KE/WxpWa1E6Z9vToZUZQTy7STFCBa1C82
0bFgciitAXgzxwSqFO0YMbVtOooVmDgRJ21U8ixDN8m4FTwB/SHPpG45jEXNvY6n/GVN4lnwIScr
dflWK+bhlHSdRd4IX27srwljMJ9mtJy65DELOtqQetioODxSZagfLR4YFzxBUldZ+Cre6zehENAN
M3VCA6XRWKA4z+18pT7AjjfaUtgohqT9yWpjBilPsHSsPS6f7b1gTJI1rkLdDbgZrn4Fh+IZduhS
zrCKsPgy6+l+atLq0OKcc7w7Kpsms6fuISZT1O+Fm25zn2vh1ARrHSLx9ZwgSBmWOfBo0EAoDXRH
k11/LTlXpgS3ufPxYr+8HwmQicq6oJFIdexGV7al1+KtTg6gbuFC4IhjJa5UKZqjcdx40uXEjqcm
fxGpL14BxvS2kwTeAXdV5NltZGMHFGAYvMieM2c75Sz2UrB7QgnIpGGC3igFlclrQivJLILuF8ZR
wstZG+3K1655pBil0LSD+II1S+GLmJbBb08Y2mEOU+UPTPZlSmJaKhgy546Xdaub1QTfg/XR4bi9
jlrS8vzDN4SavG8b1Lh2rtJUAt0vc//+gvAo3/Yo+ohT4tMmAMG43KHpV1+ueLS/xV6Hz/vBgaRu
FaFwFEf0I6bWjmGE1qM5vRK58z6ERL/oslY/SdY6Bsuzq3e20BmRyj0bqyk7O9MWuBPvvaFRLxqC
OtoaxDwpECpOh3iZMC0cs8+Xf6DwdmJESkBbCO2GZyRSR/jCcpbtTVPNm6FU9+MSPw973TzsZLtJ
aypWvdVJrBdQzhcA5sV1aPgX5MpPgs+H2IYwcLrLo4UpdlSo669Cd34npcOrTpe4RoxFh6Coc49F
cQ+InhcbHyVkJuwgaFM/z6m49trqQAMj3IAGdKMyYNoxz29SCIyMJYymmG95kSgCs7jdEoOmsrhc
Zybe0s+wIcWnlZuLUhJM7yqq1VtAelpfpe8t/0rCjhbEg7dV3F6nKow6vzE6W9l1ruO8K9elPQeL
5XvIjaJtetYQSXWUY6MzjT9mmsTNarIOkUbwKH/bRwSIIbRDGGNDItJVhKjq0h1LcHSQa4pH2HPS
O/ZcyIkmKcn4+q7rt4iKL4rHmMG9qby+04j7dD9AawU9+jS7FHgP8FaSHgE+Ci8ul551oJ0WBXtH
2imezzMfrIoPCMk/mDTx7Nd94CKOFgr/ccvTic+k1naKA+7MaM33d5PK09YBh3zZnpBUe+YFvUwl
orwoAny8BOR7Z7T6NqE0D/6tQ6Lh6Tca7BLedDoM2LRbJix+iTKfN6wPG0orMmzENZBlf/gT4MZt
4pOSueFQPFKhSNC8e1NSGW+RWD3ljLhvmQl18IyrYBZhnlo78m6a/ZhEf5C+jZycyVUWBaWmZ14s
o03ToYno9E1YUp1+Uokvp82xs6JAea0hOeW13r8QUXcL7QoSq/X9K0lJF8OgQogLXxmp0+jxmPQS
FptjVmFnLBN8Q7/+ZD1sJQyi0LjF7JH8SS8QclFnHIdSE28ffEgkzscMSEOV4LuykHmQiUhDowdr
so7vwopwlvc1wH/TNf+szT8DNzLAZSseAl1s5SgR8G80D9Jc4NGXuCNLilijQjdhGtooz5QV4JGQ
5hHEs06I4wvMr4aCebSa8tczfvpCIb4/JJO/8AED+PbvJ6zqzxgkHrgH+myPN0LR89hgmcJZQt7F
B21Wh/0zAYoUlOfWtlznkfv2Es9ydWgqKmkhh0OGHGvIHHuo9H3Gizuwc6o0Bx2YpAIZTPCQo/YV
D55WTzVe1r9hcx8pB0RuUS3lZhGAqH146YkSZEDf7n1lXUgj1xw3IIrNExBWx9h4yJKkgS3+gxmT
OzZjTzUb+0JIj1OyrgNuWczmAaqOSF2znmIw5E1oV43YcInZ3SOJtkmqzIqmIwnMKsGS+x6GxsTw
RTAS4RSYRp8As3x7E/3w+ObKpt23p0jiUwBD+tee761CAS0HmRKVy7viTpgyXXGnURy4mEOKwbQT
epK6lku9L15eXi90/YjUv//V70CIz+IFBYLrs+eGxawrEhbNo/AsJqLATR8xnlq9mGhVdccSBpoZ
Wz4PjZPmd3vNafkfUxquHTFfl3if1VClHlXQThUsSPs5WPzy3CvN/KFBeATawg0i7bCte7oQUtJd
GbTelJMk8CqRqSgaBgRxxj3/IYPrmF5BpFsH5sbfhdea12Dx2SOip40aicJzfEJ+DofKONP/3nrH
pyKyXT4+I71YdLJeMzow2LnjRfCivrtsY9QZlOOEe+HyM37xWQcubdFEX/GQhhny6jf2PJJ9yIlS
hcmI2QNfyHujLzCi2wM5dz8VyBh/SFrjf8HRUs0S1TF7arGiFhMLtzkLrzehNRLrBAkhQvSPMGdl
cv4/AJtRmY4+kJUlS8hKG3vfPjTcSO77Qck+g2TYKxYI547JuHgN4YRsL3Ve7CsYkJF1hwsL4t1f
C4MYp3pH4gabdKFZpNqM/kv8oXA3z/8iSFgbP+6iG1mkbNjW+5QIFwMJlkgotvyH7FnWywrQI4di
qcv6WJ5zMtwvdpwbZRKM0zv23FIm0+zx0YGYXw82KLFqEeu1e5OmKJPpjb24KJP4FSSYMCsXOfht
jHfGbhYTPi0wI0EworKIkDc+NG9gDIeeDFrfszng9oFdxEkNS/mrLuDFipaQQ0jCu1bheKymZAcw
DzrY5A4jMtp16hfRJTUz3zA/Cyl2RK/tgQvACVMSgDrfz6eh6vaYGpg5JAWk1M9XvvDPHCPF5waK
YajJHMNHTgQVC+5dOsSZdBEDqmvaFQzNZwzLQfbjudN1JfD5S7jkysJXmfCq7nvhOgD2liwnQCpN
FcBOF06ikHXjoHqRpQ/MHtZVcq+4j0Ku2a47Ekk/kwMAN9ehTOvP53hOW/zbA6kzU6uXCcloleko
QKBHvRXJH/qsA15cLSIcmgsVwiIi661QM+6o2uNeiUDkX7wzDxnWwH9INO4MS3mcj03Z9k1UaZal
afdjuqfmQTjDvrbYAUi31+Xpe+NaDS2T05m1zQbvV/QuHt/E86ViLjO4LrQ4BJzhgFE3yDmIYdUg
awtU/zOS4L/8K5r58SMlnizQa5Nrdsn5Fr+Fgcy+KPJ9plBZl3C2qKlUIlKrrTI7jbhzh0SnBUiW
C5+0GS0HzgLiBpP9wf4iiaykKmohaJd9lvKIGycOVUU+jICJXpRVYiEn1kbIWcdSWFETzBzmI5Jp
YvP914AcjYhQXnlT30GMdFtrzKZLSP4xcajFZf2BgFTzWsRr9U+AgN+M/jrnlqtD4eUUqkd7ppYf
V9glVCdmbbIeRo+QRn7Jmj2KQEmAg5TuR0ALkFp0ANbyD7uX58q6D6iNKImTo6JrQpEt2fg0XEuG
Oq5AZx7dI2UQ+seh8k0fYpgqqNtCJLHwgPGWTRCqpEygl71yFkni3w8qJ8KtHPgltoc4/Mgof/2d
TrL++Yc0k+czFLgwJGcEOEUy1+cd16B25+CBP/T25ZjCkeHW27KGo5vXP8cEzGjJpVjsZFuViG+9
zXZ0SwSrXOsR/zL4P62lCDR5l9lWyoNd9iY/TACST7lmipbJYKFeNRBecW8fq+/9xMwIMpKCf4d8
3gAEVzYD2FuqrNqoNT2SE27L7+tbAguBkNdvQ8x/S17zGml2kY4A2c7X2FC3tCXru96R1TdSDxKb
gdK2OUcl2rMQOFprAv20fbWfUmHlIQwaAGZabCADhtnrtUS5kznM8KeIfcm+CVI4Qcq2Sy0psD0c
RHf86iR5rSbvimf9KWDB80iJepISN/SuIgC/MKjk4Q6Api5Ck3QmtoDl0VC5p61QbJgh0iUW3Yv0
VXDheD8EYsXwRpdCnYvlSXpvDTJIcZXxW+1oVPCNwBum2oRwMSWk93tgy82p6CkdjPPP3wbjDRm7
3dsvfZjnc+urfGytbyHFkoUY4Hy73b8OriNiigGIkhHCfOlVjc1Nu4psmt4gp4o7TQrhQOmmoZNh
cxn4/7XWOPiplYBsN+1DVLsxew/UogEZQxu2q2bX/onzFusjxEMmTFNuodBKVXOFiPtQeaWlZnD8
5L15JOBoDfVOl65pKcMX0nk42loYyv5Rpn8+wa1Vo7wbkxomSunuiDGncBBp69YmYoEvTa8lToHb
L0N7ngjHjSMWW1x7CpU5rxKkpq4zMCBLpdisO5DiNP2QoRbGkednI5s+4fMHvzDqJWTyfWF+MU01
a1Dsl5c4pCVc+zeKoeIJvN5eqAE0SbptterMOhysDnv+Y7NnYPG2dMaVYQwjbVZf0G9pJzNQOxdT
5CV1PQgb3tOtCFNii/xFnxwBH2YLLu2xMbp302MQOi+2yhnDlQZtRgoDatSG8MpOCq1VOw/c+a6z
0YY8Wqv3tzJ0OZMfXHCfsj0OrU8nUQp0o7w3lm2Soc4suVmv2a3LTG41N5XZmDtxshwoB4i58KzW
5gm8PC36Qy74ZS6G7Z40863BcwARekBTosH+gWGm3co0McL7ulP9WzLoT7cgfnZXk4wlEKi1G7+y
ol5efDhFmX8BXSzVfOSO71lYBvPSnoXiXc24C3tPH/MXJtWgVn1EkKMFgxAYaBnqohVU5VzbvsnP
jXta5LFJEwyqA8fy6O9Fd1LOFa7KGHjfdN6jJrTib/Fa0Xw/3I+vmoQRvZkoOjjlipZlyNrKkM7v
7ZCNGgp+90FEAbNAPKTaB5eXq+SwMeHk08XwhUhYAdrVBGoa6TulBL/MD+ONg7I7Lcc/DkLrB1nk
LP3sjn0HKjonaeEyHUCqoKnFVS01Ynn70Pv7hBoI6YyXQ+JAbb0Hj8dUUEoZbcB7skpm1Ilfv5+X
Z7VR8LRrhW0MaHSndtv+WJ4ov1yv/hkng5vQFRwTFfQiUONsjl5AOGJTlwIK7Z2tYQv4MriJY8LX
bIdMvzzrb1LphZFWduIswnfr2aDONDSeDlC0vQbinUvvoYOkSK5mw9qO9m0zccxgq7CSMdXVvvHF
J8Qhri+VIL+XeZiWsjl5R88XoIXqCQL+bgjjrqeP3sNz5nke+O7IN7DEEojPooQGoRljOCV/k8RO
HYmjS5Y1EJAA3Mi4w3QtMAWTjjm9s/W9cOuu9iVer8Dhuf/YRTke2AejMvEn381GjGCSnZFEeyZn
riB0abVDZH3L9ObLeGPrlpS2rkbcBtAbl2AKkZpKAbropu8ZgFv3l/la6/+6IG7WVXgHPcKnXeIT
4x3egR9ezE6/EgDdw1lWUl6QJsNur41i/Arcfo3rHNiRRmj+cABaShybWtvB24rGvz2RNWBsmq+a
urjpenHm4ofyb21pXpdK5Rq/5Z73bnSK1UPBGHR6vYeQwCmAUJ9r7QTLpHbEJFlX3YCuWoHSFa3N
TJIOCzidMAqi8sY1YEXceoOCtoXuKBeQsf1pBDdBjIzi+zkQ8isbiRotWNKq27wHk5CWwBX1m6yU
fTDhVZY/2K15ouJiX/X8WocvWOclqydJF09AgQcOJHyasN8D2IveUlBhujp2DVhSMI8YoEajm1Ea
2J3rnwBavmUw0fiqrkQh5SDdhgmzf9QoSydAgWBotmWO0taI9LAezJyOyQXw1G3ylz9kz4S7MZkF
z7w5103GSZ4rdoCWGc17t0ZmpwDZIwIK/xz+e1re8q86Yd/ttLQqVkz5t34ziNyL+Kf0k6IIyJ4a
Acd/rTOYpKRIRveuHmXOHC9oYc4/AHfYTfB6+v6BRMFeX/dljusO7WnWFA0dSRRq+Z2TtRrPRHnv
eZjRevfPq2IwyvsvJ4UwxfCsNUUwXoGlTVxbgqskvjidzJ6foGnxI4muiCIV8DZAODSQ/WUj+Rum
1HxfmVA3XW43HNNDqx6TuCrY6g6ijcaPr+mZ9jC2w8YnBN3IZiuCuz5icZ4wAiE2tXWyD4AuCsxO
E0TDTEy7ETnLuWXaw7Kf1N9Tf1TW7JSTsLTuoDD6WhvmKG/+9fq3UrgCiM9V1JbFzRXjhw2yrJCE
ctMxUww6HqjHqs3oytrB0LuqUIEq8HwoxNs9Z9bEcL5l7CIDVqh7vb2F+wLi0QD1A60M087w7XSX
wALzZ7NxQoUNL40wAhxdbAuFL9yi0bxWEUXHMUKKCVGTlvwD3Kg/rRJmyq0C0kMKreIUgjUgLDkW
gEiZu7fSKq4y3ehyL3lD7JTFO6Xj3/uf5Gk8yrQFUud+I/emGDIC/16F8cA8+Qweg9pYdrhdTi3y
p6AELmlgwQwh+NsccQT5S+4eVwlmRbPM+9wKnxpV6kix+9Hp9WYBPWfr2WrjOZ5uja12lvodKgMZ
qhbJHqcVXn6TwLx7wbcG/I+AdPLMFWtBEodI+DdxNanPx2uRUyub9Cup+bPiIcGwXp3eX7uiEiWj
WShCPjfRiD7M6cmDiZivn23rFiJ1CsDIFiRQPXCEz2tkf1nG7JsMzh3u97wzWPd/BouFJWfKG8Bz
HD/jzo8nkc0YekDiSVa1LKF8BMcmsCKUgaSYqdf0kJ5lxh1Qum+UWcJS9RfHlITEPvZ7MX4fZgMm
HjBAcTQarrhgaDvSFmDzrkQ9o5hvniKNXUbTcqySqS5DuhbYQiIsbpqRBlgsd9igIRA/IOszmf8Y
UGBpCyODLEo20/z60bt9CICX6eXIThwqHEurzvU9X0SfdcNh8Vuu7RM21ul1+ssZzwGjwUMXMKRo
fP2ryTvrDNQOgUMNio+8Lj2HXZhi9cu0M4ucvkTW0MlsCr+eML8VP2G0GuzhR786O/npVyHGvYzm
ya6QK817AIFJGlOJtQHapfXf56eZoN64tATSzcQzWan5Wlm2Vw+63nsIYyWhU/sRThHTuenGO9xJ
n4sArVGxLc2sLss1Lc5QLBfVmkAv07TETq0hBlQqmun2fnsGgAe9etGmrXbXdveH1maxIcEsIS2X
w9JmeK5OpIQYBrjOJWBT7YzZgeZgw4131SX94UjocuhfIKXLVGxs3gDRuZ9FFafnBS1t5l07F+I4
/9ivigzPOPvDHWjsh7NeuvJxsy/JIjDCoueUhO5AXv0zRchtOvBpGOuuf3RWFg0YvK/658xAXi9J
KejSlPQlJIMf5Qq0rlLl/LATagW0XtI/xH1FALaxGA223LoqKl6R04cpvcZU3YyjceNVHGlqr8J2
UlUqKnSIX/XC6OzqBO4YQA7VbIaKEepD0lFyfGv5+zXywKH3gGWz3UsNDBS4TwW0hACqJ4M1Reac
jZmtKgn6MDxwuvh8/8JyJckxezMulrXNyNsqHHWOJXhH+arA6nki1/5lx2fCj3IJCuHHUByRN/Wc
+X1X+i0wQpUUB6KkgG2jx25qlSdMLf4Fx21g+YI7h1s2RxvahZjzd0UutjpNVIFD10f6g7XN/L2k
9hDNcNljDsZAQnIyW5DPjNjsHC/7K/HLr0HxdyrpiFUN4QptDYmGgNL2OLuLaBQYAdnoyQ7nCwXZ
EA6xznHK+KSeBGpk1w/HzAo8rXX0pGfVUOEkqzopNwpHChso4tbxB5I/aBXRxclCPUiQAnCpynYS
tCEYAc22YBRx6XeVKcjIomWjFz820TWpnP8FckcubZDUdd6Pe41hYkwaN7XMeK19ykMWNXChhBpj
fVv9xb+LzHRnCj1baM2w08kr23WZbgg9zoucFHa67fjGB72kCHy1hbKfeEre3RdHF7PQkxEjitU8
4CXDTvJIC9xEt2NuptRFUUZpe6ZUXI4oi8ww0FQCQgIMQfhDqGzhmcEPmX+EPi1TAUUNaEFNn4Il
AGozEsrQlBpZaqOTMnJ0DV6sE6sFRF4zfTDAAm9zJawEiVg8EbWU0oLotJhXeQ7jZZLCLeT2oX36
TK/BA9qBZwZ+T0N35VWMcwWEb4h5HCRHUv5v0ZAr7aGjAp2Nh9vFOzEpOez52RDzmdQO9hnowRI+
S3VnqpqwFC2N2464Cp1YorQlI31FGqavYxqCNPjcPBvZ3GjMQC9F1M/3KjTvSJRYQ41xh4g5W+4r
+pV9p4wCACMO9uxWOYLgUQdMrnJYwsb6K8RaYcSvYfaRFEIteG0x4rPKh+MW4yyDdzTayVj8iTce
CVWb/KV19L/3SUHDpV74Mce6F59svtXioSj7g17P8+hvNA/ypW98zDACJD94l9ooFSck47Hc+dn+
6pCLim0rA8cIoc/k/lMkjRfHnbegW9zzRIpTaGJwMO4C0X7mvkSBY1evIHt9YROLGw5eVSpVupRm
kd+blsfHPhBbjgUUEQ0ndi+QShTgDeKLrRuVczVoiyW0+lIMc73NOoIjBB25fnPeJgzsoAplqRjg
pcLcgpk7+++WKV+dikw1DQGwfqQo3x36BTC2uJ84zwR/wXlvF79XYHlO63zitzMBN3DsVaBVf/1K
IPdEDgr6OyxSUNzu3UVoQwo756YTczqvJlDVq6eSrJluMFdY1RJkeD+Ccfd+7jA8iMp95fJoV/tb
x6EPyP+AOikS5dO8llbzTexGby9iCCqmYxUGKlj8zzM6x8auwySVLWGvLybzi0FpJpDNAsTg4V6I
oppbcaan1f886wMTXqCwEzJ8kI9dd3dHIqyaUMY/oaAM3aRtlD/9fv9e3ZYeML8nbekNM1QoA7F7
d4BZJ+JbWHJzWPWFzBZJxH4xrjKWszdlJLWztfJVC0/VTEYILYbF38uVfHi4NHxmDgUzUoqgMeco
HV9v+cJdgCVDM42tBBlaC/5R11yBNkiSLNHfvFotOTb9egijx3kLCRAgpesxoq061/C5Q15RhDxI
gmJqz6l7SWfIZsWQdNuHXpHP9s3pPXngoEqjSz6wIteybg6G0x8BU+CDlDEScYYznJVMiAB11+n3
J4pSJ3NZCOS6NCtB9VNLkllV9z5w7jBb58QEpd/owunossdxNw5wP8HGHvyIj3kasSG1kZNVV2Jw
GlT9okZhvKr9yq7ahLsqndcDuo/FmAPhiM+sfPH1zgMiPbuCOJbJaLXq4rSBJZL7oOGUnP0dMh0X
hESCWrFcRRCLfhO/yt9k1k4Um+be3YARWXn5vahG33rdAg6YWeU7Vr54vPo4gnDQXzsyyxkw3E6a
zN7Rw0W+cfc3PQEsz4FlM7nWT0TiWeYZjLb9Khd+Sx8ky5chGvPfYvNciH0lTcjbWBuiNOFX6pP/
j7ZjRU4/DQKn38JlNggjqbYKfzXmj0IqX52L3P3z87Civ3fOK3aG6mLOhzL699qojns7k2QQGRui
HwSfHZ1fxgTQEWJY0OnXrYi/Bj7ox/hAtyNWX/XhwCb0MbDFFrOpzpAWsyWIfcv7WJknbG4NdyFz
FPVKpVP04IhH5b75RZu1s+X0zT+ootcmw4saeXSFP9R0+i5lrncwpMHWxvoXxObKUG589eDxQRuz
Z5Sn2jxo13bobE3eEaZqy/rV5ieVJAVK472VlAEO03CWmGMrGtb3rP2tgrvq0ewQGjYkQueAtQWm
zWLMTfngEW3s9v3Rnainaq1qL1tXW2wn50wFQiAj0p3oF3u1EdOh/tepJT01j1p9QnoMtWQvPnti
YVPCC20wUcl4T6brmwOm8yDG4MQS3vhR8NfRnLnfRAG2kbRmlvtEWlpu2gxox29+LZFNMxjA2RfS
wHGI8Z+7GJP3KxN/qlnm6jNizkfbjNMwY3FVXxJj5Jm8XFsTSf9RaaGgMH4ovLHUFr3E2vU24mLZ
cs6xp/28iWPUMSnuoW5S3J2CFMEsVe0l9X2/Erab2STtCKHpCOdP/T0Di/vCf9CxfoLalYm64LAx
6O+ggBETE7dP5Pmu54g97/SuiPHYJGdjuhLICWY3kKC1cJIH3AwtHMpUnt/V3V8egehWLNvLHFBV
e0p1oS8BI/fm81liCIc/ECqIshIaMeMrm8q3Rfp0APNa67EMgZi3I86o58ZYG8HDq+zUvnY5eYX0
L0qefG1ai69irOXt+Hjv68eccafXuGaBNMFslRCxSk4Fp/W4SyfQSLZMP235aQ8kC0XxYdOe+p5y
OHEVn8p+p+SHaM8GWUO3R33l6gqYX5/W5dFJ2idkGx4I0ZxTEEPN+b1NZnnTF4t7hw6xdORY4Q2f
H9gLgqe7Rr2OmV3O0q0+XSiRaY5Be7t71T2DJr1GJe9b2qZV0dNod+x+3EPXlmM1dsdjLJueTBwB
+KPLXqlnnscwXX8vQg/cFB7DG/kTkGYjWua5L6/w1Cvqni+BITWy/FiAkIM8VBsKRaghr9z2iAhi
yqOHgWYjELpeQdMTB3WEBJTTGtkmBdJpywzXpAOoZnXaGa8/YYcwEqi5PafNrH+1lJX5p+zWNpZq
Z5oMMtynkSfXef9Wfaq+tpRvlVaEJEiJt9Bb0+d+sRXtImBT49Lur5FtZBtfyOpBNU+eArEWNyWU
DP52+PkdhArP5nSQZOFqrwZ5NzHx7F+iX9qDyKr4rftYYFBxHKd/2b4uJZAm/5/KzJbR+SnL3BRp
bB3tG9LwbgwsYbcF8bQmmpuC5nzKJULJ1FdrB1iB+54kS8pLTBk1z+sn2xxbHbkshV/dWXmaKtne
wJOSc8RnjkjLZWPq1cE06xlfJIoY/Ri8cADv7OfmAGsjHMSuXotNlw8dR/UNHoTJmSMgYXDFb95E
S3vMAlzHtUWErOIZ+aiO9Afh1TMTP1bQ7j9tDRl8ZsDAFj/C6VMkh3UsECUgTr50mTgGN1r5WML4
SSJQecmLw/F0nr+PFp5FPLM6Kw5HiKOYiR0NrVKwvlFSlZcPfK9tuXgvtKtLnqr/RYHjoJ4oAPcL
blx4H8EWA4UYInFHkvWQkslZr9Sj+XljMcQrDhRcgp0NHBg0CTBRjMyA8Mb5znt0xRSRNGkMB48H
6ZTKgSpoVtMKh6iTGFu0SKDf26tHMeqTUyfFHJn0MefcYQS4Dxo1VqDbJp7Ib8QHiAf9/5xKQvXS
5ydqoyz/MPMbxSzGPHKQjIDXhCBXHXYodvg1RGw32MEuiMxmPiJQRNEsVPogC2VGMaDjVHUSh1DH
AKDZKK06F/kbyqixNCfxWZNtpiPg3BEEUckQJ1J9Fc7qjWoL7a57x1EdBDZdznUbN4RC0pFBCALv
6EEt7HdTDuAH8XesCs37F7jFXqnfKcs/ym29DHcHfLorJo5FS6D6u1PLsO6h5JcewbOuTMWf0FNh
WXnVYuWIoFjfuKYTeB8FCu8XyJyro5NZRURhaT7I+R3LmvWuzaieUCc1TZpMqtaELDLMvSZ1A55b
hsrcBZ+pp03NUZACsnceo1YPh4uCPu85ASgyWYbnjk/Yo6jsXVJluBe63VKeaHUMeIJA/m6i8knT
zuC88JSRGl3XWAxvBGvS0oiVwLm0agb50fB+KsZw9xEpjhwPHsa+oKOY1elyEBt2Pem8tMokWJXr
6RkO6NuxrZArutmEIAo9BBkiawJbkC2gdrca+/YZwzJOcQEYW+TkD/KG4J1Ka6LuQH3nckJgQFn7
n0RYqUuH4WMPIDPxFB3Berzb66SC9B4eibMr7c2FppvVaW2IaMklwjsWfn0AZM7SW2ajkIVLnzRW
ALucJyMYkka9jnMCr/SPx+t5TGXL2ihVgTLxsB5mhKCODSTJJ+0TPfn3QqQQnzzTPmjpbbELr5fm
yDll2NhTTvuLW8Kil9slmfHTKdwS3/jJYuzaWRh2aMFW9IxWtII0/zYNEpQ9Du9UckTWfAZD9xw9
hnkaYLbCG58bG8fNtYnCSGLEAl7eE5TFsErcsLWsheNkFCEU/LpUBbhRKaar0qYpRTVQR1eD6w/0
idfUzldHUM53L8gB2dm2IN013Yl2wzhdsOFAK5J4tffMyPordGmZr+y7zOwsE0fmENbrRPrRbN5Z
1EftSpriREO9haX0B6ubujPljMBxEOXRP8WOLIJ66d+igudiGOOUjtEi9pDn/S5YEFt3Hh3sKA6k
AdIF1HkqkCbcqeB8xJLTQNG643U9Ef5/q/2R7MMKVh6r38B2P3R2z6eHJVLEpSmKFRMexac9m6o/
a60zWb/a2PYunp7f7/2dh3AxZuuhGlAFOaxfUq++rUewiBq12dmko23mKzlgFLFnc0K2F5ESVS1B
CABb62ZYzIBJpGhCz5qRkKPRv5hbu9jnMEPWrAXmN204N13rL93Qe5oB0Flh9kRR4ePaeFdTuiRf
6HzglRoegFoV5NhqYwD0FPB/Iht32Zml0uYSmv7Q7YxlTpTRwG3M8zHuJgJ5rcyApZLMHXJJEegw
8kK8IHtj9cXkLyl4KVOshsxALAC3woYxA+fMxMMfRuWscs5i73wfsO8funPif06KtJfENEujEzq9
Y9DeMsafPGK6VWLmMzeUcsQlRhQO9x9U5Kh+WMg114UbHZRplKdGV/J2hIpfiruKWq9KPj8VHR8s
MUPpPrZOXJERMAHykO+OMmP0fcM/KAJR9iSzrWHYoCZqInGTLiWzICIbvBQ9VJL7klo61qjXDTNp
wd8JDwtB20ExqZZeCuHM4d/DKIE6oYIRzW30aHcvHjyOD2bEjGJOp533TOgShYmoGdpIHbRBZC9K
1WjLdI9CW0GiZ8gMpB3/r13rpmzlIWi8b+8LmwVsBY1LZ/zYEc1+22z8ABF3YT2yub9iJ8hP62EW
j4aoX0v1kPFXSERJWvtpjiZon7Lcx/oE4vicHihBGoFbfdR6/fq69svrwJjuB1mbHFXPE30sqQdh
ulATrpdQr3WervL4IWFcs1ppNtVqHUxcP/oyVtycoORgdMwNz83UUlSvEmzdUcYNBIAPatfbOdsM
wTUQF+HHQl350w64od56RODRGgYrxJKyjBCvYkg/7eE5ZqUp8zEY3uO6KzPwyLWQsOSSXsTzmoE1
/QX5/E7yHnHknwV8isR0Gp9VLvmDhO8dONs4WAmTZ45eENXed8R9RPewdErPGzzJBHnl8MT7r4ck
5DHPoipqFLhQMhvzUzs8hzMvU9uLaFOsDrkrYb4tmjv+4414K32XNn0TvqaJ2gwVb0VPPEFAVVkR
AMBBPvPmsVwCZq1AXUDWCU722q5mV2667t/c2ykrXcHiDqaIE7Wh5E7IhORYRdM6jRfM54fjfsKs
YOSuDKQtI0BUSQjv2yyDV71X9PqUguTBqiROoOPaWbDKcQ6jBpOHD5AaNXgeAbycwY40A+IpLMP7
ME9ogzyfLO0cXmz4F2KLjdEQTXY2+fLoPCfqmNYg8fblenkxLb/JBxEgTEoGU4K6wGtueNOP0LrX
fHt6CXsfsT5WvDm98ifbRpnMdb4HG5tjscfUPxmAIpGdv0fcsChsxR29LZ4of8ofSlHca7NS1Fk8
q3MgdbLV3ccwrroMZ6dNBJkP7PQl6HYnkqXyvX0/I2TUbf2jYfs7VHM2us1Um99tP+fquZ8tERdW
1xs4GZiAY2nj0B2a2VCeY9smQhZNZLJ7yp4A8r1sES+DJ14HDtihDC1aojPUU1d0cvdLgCo/O1IT
k4pTVYlYQ5W/bkOlaCkIuVVXGDIVb+nbCUg1z7+5qIY4CbT6FZHAQg6jqMo/Ro+D25/uP5BDBCZ/
53OKIAPedz5h78LfSTG+p3teT6ycpHMZPezXrVrIZPNF5C+MOCtFTNuHdDTXdnbUEq0GQJrswxml
qr2jbIAQx8f7Nv7qHctRhUbt2Wb0QHcLmG+2RDXK9rsF1Kp6z18K2HJUVaLwcNmR13GQuuyoJ00h
VMY9XdTicZP4HRlFdnv2BRvtM6t6egQshpYjRyXts1uE6UbA07DsizXMbDF0OvyietFYbdKcau3B
+XTLbebst92km3Vi3WmALWOpZOi7rn39oCY1EQ5SSwVY5dXQhty99bv0EG+9Swo742Pi1sYM8zHR
m9AjG9U/gGqZTHE6IwVeb9QKecOClAodcCyZ3q9LubWQ9ramIdaLfPwzyajuKUha0lUdbicYoG3e
D9hwK5v6sw8D+SC8SYfXCh1J982qnnJEKqvrcWSytcwWqxLgvR6Gt+zEUhUIRkr8JBc85nOabZCl
OSqT4/BRCzEWlDTeCupEwwe6sKhkZzbOabc1Wldvk0oIXZr444sswOv8ztlv0WbTG5y5lcCK5Clo
8utk4vkLEDvIJ0i7E04vI8N4TNK8W6RZZLU69QHMarvOKbRoThMeyuqFFcxWv2Y4quRO4a2AdLFI
AaycWKoE8ybIrhUAxQcnOK7FK7vMp0tk4KKJ3rI624m2W9EGvmRpLyN+d9YTdpzugV0YPWGX32cb
aGr+fvz+ofU64j6NEzEIryAwZhPjvwP0C16NIxFtvC9aEZBbUUvnoZqgwnZia7ZCKujRW9G7kex7
dUFM07b3GDEbh4V5jDmioCB5CtkaUm27sGzuV8TXLnP9wL7FO2DqCZIm/xjZoLOw6XhNqQBvMnFF
G1rP/LCz6MvixdrdezNLsIr7syfQsQ3ydcZSoVG791KtNn8NP/QQnhmF7uhC9xwkuGHhgiKoCAVj
4iksx6TeH/uHQjGfmMVP+o7SmkRFwKD6cIrIo3R/sG3ZdGjXtuvrQvFYEoHl+cAtk+am04p8ZtmU
X/g5x1tzHDMeR5qWnASGdlHu+ePrwLoD8cn/WWjIPKHYAfgg+w1q+IsxDkLePR+qeou3myAfMsst
TWLpNV1W03Qjcu5Sqw6hBgzqExnapIqiCcaMvXwRtD1LdTQXvw10v1dcMkIcZJZa0Ciiy9nZmn8l
QCJog1zIxPW05JOZiE5J5itNMNitNCY32dtutrgMmu1BTCu7bCTAuC00O0j5rOoUh6pNxE2fqinz
5X6S/dIszj5V4DWSkmCZ2cNfGODRdej0pY5xHjWQAynVctc7vwEzlGqMNplzz9X/jiJi/H5d7uIG
o72tXcyNIJNkszWKh9efr4cl6DfFvYEZ/ngFLww7KRTyP6xBagufyTVl4fbaxBl9/twuLcquUEoD
JCAHHo0Lo/b33H4Wnpqcwlsm91hhJuoi29xpM3Lm/Ihg6avtMv+yar8NEumfoR6SXzREZxJwnDV5
Fc0qd0xp7Bx9fmXPrM1xVaxLjfq5sywFebBJ6lzfvgQVGzGjSsGWUzVHPcbegc+dRAeXwKemGcpX
qjAV+OYCdU9cRZ1T4VM2FVqVXQHsjvWBZMrkf99rPYg/bhsL0DJjBU+hvw2FDqQqMrtiZC/uCLAV
VBBAO6Rb+QfM8ny9iAFcloYuWp2psVXqXZpLpBgM3NCIl9PtiUB6vZOMxa1qo14CmLvH6nTXp9rn
WRRuZFD/YKFuSCpSS0HewsCZOtRvh+lPL1ySwDFJLWoZ+ddpQvnKbXwUd9Im77/UL3gm0i0KSqln
E8BZLdE+NSbu82RsKa1RU81HXRVU7PCvuKsWvNkwTZ5DXmmI2wtD8ymKpFNM7wfBtvA+3ez79mZN
q9MIf+Cjwd7Pi8+e0cCaWZxbQtz8OJ1RFBga3oWMfQCjBlUpyjt7LiPCn6al5QZuFJpMVRUJQ3bg
eZf+ZUKzSLOXidqTU/Hd6sKdxkx/HKzDTrS6AoWdAu4Wn05C71oAjBxsb3xRkYVmT/yeF9UcZg9U
BC9QN/RZEOtlIGj0hbjzXQNBHJgDweaA1NDEOoaqkSWZBwHSbmnOVihhMr2t4+4ASwPmTC2yneSS
oDb86yXOS7fomdjaj+cQ3LL+gD/5g/V9CK/Up4gerpdB1JK6oIorIUG6nOR+PPAqRbaYkX1NZZ9b
MpoVomaGGENAi2mffGI1S3tXumfQk0494JefCv5Bry4F7mil1EmJIabpL2nhE3Rt4da1RhwaYvx8
9RT5vp/APUp76kK2S93XM/TMLz0chF2sKTCekCo9cvtJK58ZMy3O8RMEy+6B/D3YIKDXSfug5zbD
AaON2OS7qS8K6x3+1+MKfC+Hdljgf3DjeHt4fAIJ7OkM7AIEdqgVrzV/3WljiaNkriiBS9LC69fz
1+pcjz3GOWA27/9IeD8xTevrf6gaGNFk/n54W1sXQmBTn/WSli5IvIV8VvFwQE7HX0Et/RoQa8Lg
LZEGctyMSlSBSC38nrlzmr7uKM4IIVZU/R9aeYL5yhE/3eHpNABrpuU6rKV26D3nDl350uMYy+Oj
ndeH9fNe5AWHzMia5dwVsi5WJ4P1mLhwvsKDJTFDV1262T52QlMtN7qrGOi7VNd29PjDg4UiFXIg
dfQnNHRMug12sD9pjQ3SQoPHkl+SZYU/hdUT0KKQEeH7PDuSD28CU5fN65CQ+9Njai+d2f68px84
rmRQQ6Aj15qOWDhDBWEc7fk87BLApBo+i3pUnvGCwj+87N09EgMxYeV9yZTDJy9TY7TTT7SObUf8
mn3/J8nG4B1nq8iP7YZ6bpnECnPQz4YDgJp1HKO4AyzRRNew/MmlWVua3ffdriYcfvII5S2ZQOQs
1l3aVBHd9iUvQzcg4xMBcbb1tglW1/V9lFRsJjf/5k7vjwpurVgpJ10Z0VVue3TPAuRZIO8/iL81
VpXlrZL6mWA6y1ZWRTuKcGTWrovWWLvePeFAsw5bGKqOlY/hfOOyCtiWV6n7iiW9H7UJdwhF36pN
pqDMlycuhBDndjDIS3E+bHpSponhEaXk5sBTKfd+zJ9dfqPubBfb2EGgFWZG06I6SG9INon2iSiS
3P7G1D2NbjfOAfaaLiPsKY/LkOAQTqUqoIHMitm2lEMlAAT3dl5E4zvdBiho0nMwMKWL9SLTykJo
/Q7Jdl3qcnbbxaoPJ0C8NGv91Oj+QqTLlT009juBEh/tcZnvEOQYDEQ6gtHY/H2PSZJ9O9kwFr0V
PMYZ3UZzGyAoAAjUiFf3KMtBeUHYjqs2rKu5vVXVBdLZmFA/8zGILo0YHNq9VnjkBqxC1WgCLVxC
qioeusvuncH5PltJn1Nt+tF2SkhEzGInKHWG0MKd6tXe2s/RABHydTy7V3xMCpP3RHQVYFEc5mRs
ydXeFzRYV2pX26SWNHeauVMEyYRRLtYFBD8Mfex7OIljMt6vwby3Ib7Q+yQdskeHuSCkbvy3Ks9b
mBs6mr7F53IfziM8S0DpoolJ7+35Tc223yxFUxbYlyR9SYatWBaXhEpVIqBAp2leoE8cBsWW/F1I
EMji60WAICwu3ZI+RhwiDEdSyOfqk/1HetiL6NKvMOV6EmBxYy+zrZU5EdEB4J3pO5bgCzT6eNTb
qe4i4Lt4czFKf4GnIrS7ia204su/PoKneLbPBtX2/IOdfI4RWTaVEtnwiGiTwQuZArKrlQ5cLqpY
5hFlXW/8od3umn2BaZxflFTZ4fox68PDNNx3c4MZvovJIxCU63aJ/iHGPX1mdKLeJ2VzvnDwflzZ
U130LXDBsB4zbr1RbFvJI/Bux+32toEFoH8CQuGbs/fDTlTzH2jGrUTws7Xb9lf2UvqxV/wClngd
sOPm+dcFAhL9us6qPzP/AsbfUG7Hd9cWNNRGv8Af9+oBlNHk3rUz61/efoVsOb4rU+ni4ey2skzA
xpMQkYvmtvCeL1CmKsPRpawa30S3ubcK7Vi4CHhlWovzQ2Kl0+p6rtht/rQrzuuR5mv8HeH8+ZyH
gJIt+LLLDgybhTMcKOa1k20d1GOzUUi3FPgZ8HfVRXyJUQbWgw6ZdNRBiVuZNiCiNnIif0GeLtZj
pr0o0xldvFwE+g3iv9yasCMYDc0x6vSfAIYygoPLqBJTNw61ig7hMb7lkNc03ZkJNK7ar8DzVqy2
8Iy1kZHE6Q9PG0H4U5kGVYuNmq2P8+yPtNSGjXvtaKS50+mEG5MMVt4Vme/wLYJ6UR0CU/zoTsjN
yPOR8JbhkEGNNkiTZE2Ju+xMzLV6Gs3WSghOXrxoW1zsFlaoQNrwGHt4eXFA7YsT4IzHZd2fdgI4
SChcoPVwbxqKgghWe5SQ7hpqiBA91Fhqsn8f/ixiFBeKqdTVXEzLGh6K5MtvWU6Em9HHQQHlUi0i
ofsp3Bj7aUj846tLgmJhIImbsUj/4YOuo57vniblMTBS2FQ+/A1tElNzSlBQrSAHhXr/Q2RfiLBR
t8YvzWKQL6J4BBpCJnS9+NaIqgbxRbnsTiqB1pWeXjnfsNi3b7Xfo4mUhS0uR45/72qwQm+tUZgk
vhbE8pxaAt+xEZsm/j7JQ44hW1AxwAJ4vg0mqaIWP7Z64ZhL34NWrjlQfP2fUS1FScZGd13XeSX+
GN756+gqqB8ta2l5No7DngdSrLtGpPRk8YKTpWNngILUNsvHW6AilNeGxlFZjXFlGf+EAUOUQaS/
HkaVMITijl0ug+q2YJ3V7efdDMEnEJfM2XM2BWYFu5maRLukWpziwROTKJ10dhbDM2+8xMk8gpdx
8Jo0+qgsLLbMigtv+SlB7OeHDuWp1etk4nXTAw6NTGgsU58V6bXd5ZcBDqjdxKl3pKPAt7rrpb9Z
yFlPijfp3Dbl+hUOMEyoqoumqLXcJ+e+qV8bdm+B0TpgLXg7/MOvvtp7BDyyGCcDElBxrYc0FeIy
EUr/+LHaAqIn3cZVdrnDkygn0sY8HKoWApC6cjJSHgZuQwIvzjyrPwcOfYCL2I7rz3CNgxKI/7b4
5BqE6GxX1zAsnLyJOuJPd750jRkGV3LRBDet4FT5FgRyc1k2P4JRBLJ1bA5PvGm9IgZx+o4dgu0p
bk6WaeuyavX6zAT1wovsoEz9DEdJ9qCsJJtTs+7ynF8Rx6P0c7Qmh1R3KvN3v3TX1nNT/PiJEPTl
mw7rM67IZWTPgDAgnoSezgNitQlL8kv0qyx75q+UIWZtyR2fwjK3Q1IsvvR9DoqG0nn3JseP5ZIL
rCdYCDbP3Ga68X9oby+HUA9yJwnQaoaiY3bQBsKt/tfGLBiaqHx+0K8ws5AJv5uEVNI4DKLcONOE
0KCPMWbl0uy79LG++jDYcpvQiUSitfPVM+zl0g9CLwydpd67Vq730xx4DtzuUw8enLcA1FW+vqIv
TaywU91SJebH8JUrQClU0nZuxkCq2+lW6WAKbsu+0hhW9Wyaz7nI7eZAz+p4o1rXZbQyxU9qDzFZ
//t8tExI33I62wsVrI8/cCC8ZsB6rHUxGVM2wjFLh/33i92P180ggLy2PgNOcsnTAQn9Cv1WUlg2
o/sAlHStPk4s5EM703knNQYh4szWSJ8mM393omujTX5f2wDFjboK9NQS3Bhbozi7tUc25qZ9h+KH
99cQ2nmuyTZbttKb+HIrS2Uz3VZaFdZYUy4fLDE02+ZP/1+xivT3/5ktJEDv9g0eL5rId4Bcdzhr
fIxtlExyKkxKbPyfF7YjGQ5Ed9ihPzhV9zPzjKx7SiNRXbW9KxuIQdVth3Z/bq7F22rC4I5/CmgZ
15HkwxeKWegDespLOljyPCR2TjoBjLydL1f72PUt/AJS/DWMlzAHwM22J5SbZzCqwGiLtcdg/5VL
XYSBwtdP9O7yNSvYDnjwgEgSlV7bgRaT+Je1JSGQfQmRGt1lgCghBMvtKEqj+DFyARoi/YO3jzAu
tNhq79SFFRrZO4t3f4BTqXlrBarOXvOZKgfzFJkTnQMgRMMuGDkNdAVHXofvCzHfiaeRMArS3AF9
iVr1kueKefqr2PooL0zkUe3gFjXwPfczQpCqRf8Ktmk5hDjnI9ZbXClYEic7VDGjzCSb3MqJQITh
kolayqAtWumpJzBrupxFcPZXRf+ouun7SCOqNJE+afbP2nPfQg3Ejxm4LYqKaISTw3GDkDXaqErR
GtfjEIz/vzRXr5NoXXkKkaiZ81VDIEBy+V4h3ew22rj5bWipaE6yJvnUI9N0480mNc2Cz2Yq9C26
XLsZmf0R8lPMguUsHZYuQbG5cmHdHMDSVg3vzslIAIyEYgTuKk6qTg+JotlZFzMIPKF3MsrQaAMi
V7vDtNAoxlmd05ZpX24s0iBEpOjhHo93BjV/TgZm7YjQY1SI+1wheOylVwiG988wX3J3DbdUH+Rr
ixX+G8d8pXcwgXHEKN4aAo4oYufS9SmPGyi/DntV9BrrwJwm0O+QTaWWvdt+FHDGCq57MGHBmIbs
BQC8umsdl9mTalDBnztNwmBbunYaDgeYVE/laMaL3Y8uWHr4WhbBZ+U7jGZUHQ5ibIFnuI69l3o+
GoTpES3e/mJSudpm2CzT0S+AKetOsA/VbL8phdA5zNiVcBx53fuW+BseiyXilVWTNkBSLtW49TAN
l+4VMWWgS2J4fOMfBxDnD4U8NGtmLIq1+NsW3awnt+px1zMyRlFRL4tRFP5vf48ptUdDN13gCPcN
PzpYlyKypaAqKF6YmMpkkJifSoCsIzsdnh+h24PL42fTnCuWQbNiROhLQBfydPWvK/En/8+82o84
7FeHB0yVeiXtitdBtqxJfK9+h85OhT1UhZnwBP+q+dUBAgG4YkWmKXmYrHVU1m4W/XCwT1l+Wq1t
zMLwzsiihsXaxKXzVhDfXBbxly3H8NtllsCqxAlW0SdaWPRi2OrvF32ABAo953CSLTC0d1KzwnYA
70/6o80xxUEYz4bP/sSlsvQvgT2ADTByoe/n/w8faVNTy9IurcQ7RJOJNU0WiZGhoN+w7QdW8bHm
0xkZcCkP9SBIXMH2QxDT0wq4oeCo+HWLhiDizsK8ZX9tOcYMmpR8sU3smvZig3dPGn6EeULMfGmk
lwNlFEYZTPxrYDoYFCclYuWBpJO5eBPNOhO7t+2+1m4WRQaMdcbA2ai995VT7UjoIK23zptz2ihc
4LA3IHPVcVe+ZxYVocMMiWhghGkHidx3G9DkI+RC/FZl4CU2XqlFYoZ3HYEQzYz9ouKHrR/Hku1v
viNttwaI9/x4txNJ51pRsM1sWDH0x82RGaHdKAuYlsyPLdcqkq5elqCNzUuhH7+S5RQguRnspzL2
paHzxp+cm1qDl/ZI2E/m3wIujV9+GeS41tG1hND71kyQRqp5w/zF9N9LATH4hnZMOXojscCG4EhO
UQdtkIH+Vcwf21IdFQFD+IGEPDTPurpr+mob/DutaAu6Ei3VWQSssatsxe6W2fkgLnX1NMs8YNBI
O+VpTP2K13kmWOpVdyA2FUFPynUxzm8Bxgiog0gnQyyHzswEHRUEP1UG7rkbEqX3RERqWfbdGETl
7GAwq1IlSCuFRfTUG08RFyLKlVvF4Z+EZwq6iZHNCZOIHMq0QVLcOFwN7UYkC5WPecEsOL0ax//O
t5GZEL3H4Rzetk3cIlwvuujZtG++DnG2CbIYyXHacdRUqHmSA84AJTKexH8Gft9wIQCbOFZ45hZp
BEZ0GVor3SqfQFiqZqDm/uJeMfQYk1QVxznkuceMTN5auOwh3apx1qYTLrEstkP5sZhfhy3RFraj
+x5BguLBN7m39SCM9jA4oDcH0sAqxko5hlW9cknZUAM3P/r5SQOq3RY/5zUWJStPPP0Cv9GFhQ4Y
Rh3TZJfApG/iP9iTFuxxuCV5zRfOI5xMX4ENPEqi/+mGwuZA8GzON7Yb43wehYaOaBbTCAQ=
`pragma protect end_protected
