`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P0l4xS0N1ACznOIgwLeyPFeb7djSeIBePGsQK/C239Ng/ThQeWHdaj7Aqww56yCo
mV9+fpzH49lo7geZyt6H/72VhBtkZHij7cAq9rD9t2eTtDdxVV0G/440ez3q3/YV
I93tt0dByS36VEiy0eXb6ekEKO8AFoUQv3XLC2g47ts=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26736)
kKaSCL7v1ZaAZxUsvhQXd7/i6mMF62VGqDmzJo+MNlObLPdKHvwh4i29LNHPNyEM
72JC4UKvJwmh2NJtiHp3BGnJIu11gII/5Z2ZvbJKqpxWhDX5j8DQGiMLoPUraaH5
GbcZRoN/mQo5G0BHcp4Vn54v/d8FOZ0eYrZiPc8XupiYETjRufKp9qvnpFZfXFAL
HW+DIYxmoNnciAWiL6/MS26J4oRYH8go8VsaA/EnIKoVwbIeX69nk/mQKJ94suBh
dV8I144cayEeZfiI59ENBudHDvQtB2OUkSYnwN0xvD3gIzHPy1IZiLp7keakWCT9
CC0+mvf7A2nWB9qqbh+zWSsiq+pJ8Ppd/dUhwUicko2fDilgTYWCZxfilZ4R+wqe
qpNVpSFtOXobXdgwT0sXce9vPuJ8WKA+Bxd6BoZIxAH3IqCpdWCPQrISGeqpf51y
uy9iInLUPMEqU+/uQWBcKWOFONGCVKFyKhwgDa5AK2ckNqIBhi6HcSnEzcJFmDQh
6tPXFOIsw05hmWzIKHavb5MfmnKXP5G6JlDdwbCphT+o/k2ruCdiTIAAVFmyDf2u
wWGgzGqOvjcpl01cNWE7NArvCUKxcTNTFrC9oGhgRWGLAysYfj6ylANE9fz9YoJx
apYKd9azeHALTmh2AVuOJimaL9yWVcaMk3P2qjE68XtJa/jNEmmJjGpGQtuTZp9E
kXGrYFj+U9XkN53vPOJnPFlV+aKSfKWkgrexaLvdx0te9WxjrCtOogh8Sg7USNjD
ucLqAt8joE7Zsrs6F778u5sclgvQ5Zz2GP/pzbJ19COzK9iQBErhGFqsoEezl4em
7vl6utG61UCMaOUMVH3DQCx7dlZ99ZvyVlQfYnlyUCH3M8GYzJO3EAkY7eCDcfGl
4Ovn4uoRZ4WH69s7Wqr/9MjYzs89OrC1VenVfjfUjJksYO7VB2N7UZGvz9p9iUXB
4Jd/skDV0pV9ptGqd8NxxXgdV/CL0lyxKEcnDJ3wmMiPxpn4mEaTkW778NGdNPWt
1CHUnyH821Oozp0tK2efg9CQZN+BT3pLWXR3TkAutV9ooStega2pixvxGAeFMLXG
hd94XozIZoHq1a5yDvSuyUSEl5SrBEFwRHnI2F7Rjnj/c0wP0ur75LGrhQ5uwNMj
KadUEKMjaZMHU0O2vXI1i08FOMJx/RwkkEbUUx6rf+Ljt7PxPU65R5WTgswj8wUN
Lby2OnHj7GfCwcmWKzq0RRqDPQZtkGHdu7ZMAqT5StyY2YsejICkwmCXPg2uWhHW
iZfF9RE7CcDwgebYv6XUheEzOjsZS4ntozo1aNGsb9MN0h0Z5NX+pROy2nXneZ0s
LEPev7NqC0D123MvNPX2gngxVOHolnt5Tmlcv40XBe207kId3L3cWv3WDmIOmcF/
rpLWX3YJPcoMU3fookpPdKSHttJHNMPpcUTfn2QGkxJL8kcv4QsjyjozTtJuVXOb
3eLE0qvXR8T01PSi8wP3V/nEBPSmznI4yfC4nElM1YDzijI8dbfXDwYm0dqAbbyl
W+beJa9rD/6Mcarkc9SJYcuCClvvvlSJ7+eJac9lQouYWcMiPMfk7FVgJhhGvLSy
iN3j/y8wJ4XIi8NRnUUM5jzENn1wxbkbC/F1SeBO9TfqdClvz6ZGEJGXdfKG5uzU
Q2NvkMJo3DD3FRqVl4pXX5DLW0MZrkbNK/mBHxLkgucYmCNWC92F/QkESP0C3N2d
Hi70klXWC8Ag0IGlW2ThvJdUw6YaOqHub6rmiZbUDRDOjGGtSybG9/B7gC4FqYjR
kIerY7QdNXQSNcTEmyJwffOolVFqLz2sEIY2yYqpcTPQGQ/lDuV2hYCYci5OIVvY
ntx34rQDh8En9dTXXtYp4Je2tauxpPkaReY538Kf64gXPqLBagU5xOAltGdnTzKW
XseiuAS3Tg39x7DzS7Mm1QZFKRwReJVT2FCefkqvYMn/h3Vq36elZYMArTDUv/o7
VW5DH3aDtJLPaqb2EU9rFtyvLTFQKmZASctX7B8o7hdbaTKGIeqNTCLCWST4mtbt
+FeuuqFLKbljOOoJOdlS6eIhAlbSmz3AOo1ZNp3psoV7mqACsOuja3cjPZWoN+nA
kWjqFqR2z3vNYVbX0z/wQw7BS4ADsp9p/7EdvySkBOvjW01dEkUJltZXBDepZLP3
YuT7AaeBexfOy7p2dSLBJXv5b6Q7rrg0T+cr0D2DspPC43wpNaznNG0UgxRNljnR
22qmggkcQvjN24eWEp0d8TF2ZYMBjYIquyKWl0Cbt29vTGB01D9crsmD7aHNda5A
Xhz8YwQI9N4Xpr4/7TMuwFWB6Bvr0eHIB+e5C9feQ/SiYX07jCXZGtuBOL7aM/va
bXjQF3ZY6YWU4sl7OwMAmCxx6hlYaajK4V8wqPltMKcuEY4YzS/ZLNlNtF1CrAP0
LSWCZTlFGG2Z9U6QEBGlrtdo+RrIfUPP6eFz+W3jErBzEoxZr+xYOpAz+/42LGUR
myZr/ICbTdRFED6B/cFWGN/+J+esjaJaWgsghamteBDXMKeoYYIe3UUfVb+VPmtD
Ss0EOLzL9JJofz52go4ZoaMs8UoWszGJKGzAi1zueNjwRI6HOQa6gQGGAljP4/hR
wt6G7xsXGcxBSaBsG+IsxX1SZQeWN/G80/qGaRae5FCddOiMoRlioSij/nlCFE3C
nbV682EoUFxohmffOxPRw8kjCXJ6Raxyc7qd/p5cdD2PLquddlt88h5+Ml28pz4V
7mNi5SLDESuY9PTNH833sxoAEfYfn1+dLMgWOeXvl2mu8NDA02+NnJo6m71NRBYR
0C4AGKaVC105f3ROG6beUFvp74FKQkeUaCHPfZ25Tfq89/28ypudOlrDz9r4yLYB
L3Y0D5db/yyVoTVO0edqsLiLZCAEbEF9l5metVcmVKo9DVDluHsgXACjrq0D+Ihz
fC3LvlIyL/VuLNKoVawej5kgCFuKL5ajR1SqZjVeIPdyyVhBweC03DyVSPxtt2R0
2yDAxP+bQ2ehKa128VwXy7SV6p6Yq18xgdw0c4W9pjLN1kBz+rISyN2Xk/kUpsnp
Ma5h0iboD/bi4O4KRwBlBuK4AFsaYEBq0ZNF+O7Emqnt2Rb0r0yYHk0U9ppgxbU4
ftLFW44V2yMhqGdWgHLWT8YO2TTDiETwdxTmlX8dD5DM8OfsNwzmM5LRLty6q5Yo
h2Q6b2EBgqIF8aq697vId9WimAifBvB+Gfg3dgv6AefqNjUqWiwf89nRIQHGblCt
eFeN/+eCzr0sKI56pHSOwaRgC9rR7tUXI4ki+Km1CGoesIfpImzOb7DfiaLIRmjb
jKr2QxK01zxvO1XXkrMcT7mvp9HXBh7ZaSQlRHawcn9ZTQ0IsbNKix0uUGmb8XM+
KYbgkCFR+gZgRXAH8UNTSleFSC74vEeYeHCYNmsAzXNGOlSMA5xKm2QfsG60w7WT
nYNAowvgt8sKE+Yr76rjnOnaXI7vW+ydlzJpmjrHgo1Umy/DrrU/dVyjXAxmCQ31
TlvIyFkr+Z3rPwV+KqNkKMGliNLXe6K1cOrgxHBPrdQzFkiifsgqTZ0iCFYsSOqD
PAPMJ+zOwezGqD3yZPwA2/Kn3XWbV459Fo+lK7iCyJ7o9LSyP0Tj+udIL7RWX2Aw
nB0678AtSgcO1qOu2X2cjD2Vfa6g9rihcJcQOnGV8u23Ab0nd1QaSri81dF48RmL
2nAM1pzss6RRYom00UiGx3MN4HJtFzGAuTKMlZaSVGELeuyPuuOEEmZBlBzB6f8B
+7MYZsP+kLnyhQjKEDyk/108xkWbXR9Ipxw6PiNPuceBbaVbBzBi857Pelq4NfFn
C5t6xX/BTkRpnR8rR2g4ej5SKOoqt08xZjnh25GZ0JXvtwZcnc3SDLVeQwS6eMnt
JT97rDFBqM1tVO0uNOtNV8M6nw9BOfEUwpeQIdAJ+VQ+UZLAUr9SfG51sEuxOCAG
PNE+Qx4gvl0ddimOh1SQOkkOSm/aOK+RMAwQB8K+H6OCDre5YU/noEZ6tT7owxHA
068L8XHXgmDSpA0PUR6vXDugsHC9q7PausnDEyMlP/xUGfw5N+zbqzAUxXZnHMN4
hS/gyBC/Eer69zBY1Glm5RdxP5x3qqCkXOQtIbWmJ/SQN5HAYyL0Bs702gAjUfzG
HqPiYQquiJ6mOaIgy+JNf3K+g4DPGlyDJcmj2G6BdGtCgvO8vlgN7lyU4WYQdw/X
QSIXn56RahCQ+hMto9Nh/P98120XvHOGWTrSR9Qv7C5TUgnPkgNE5k6L0+Pksyfs
u6O4ORtPEeAr/PApZU1cMYv8x4VhULaJVEXY/evw7CvJ91ARj84Na/K8fGhxFexh
J/qeARCqhEW6sp9DmQw1UAAJjQdto2tKPwWu+kPjKNdRI2RENKeh/hsJyaQKRoaO
Xx+HIS+YKxwIvXwBi5qILcMVCl8pVMTzu0KOl8sNR7xKYyIiBhySg2V2ygrSEUls
TyFRvP0gTErQ466HewwZpQfC4u2iuGYMnHFBC+tLTWcdWa7sRG5wTaP+U1Y2ALUU
kRK9jCsGhuqIjUjNR79lbxDb/Nsf4mC5CY3ezSpwfP4POPI3Y55ylbN95hNxrfwO
UfcfpdH8qAsHXkWKK25QQvZBuObJ6Q0+vVTFQlbkpm2Swp0VQAE6INA1FshWz6aW
+wLhNUHscvbriwcrN1zX0j32E5aVftUxBvCiRZ5hRjFVg2Yg+sneESmA7Qo3ywM9
3UX3ylFimZyntrHxk/9QH+tTEOnXksN/2NQn9Q3L0NIe46qAJdacYdIc2LWo+kXf
wWuYgE6prAz79UPNwBGlREI757zxS+Y53JldoknJD3ZjpeUi6xG3Hct2Y8ni/6XS
Xb7dPl3iM+pOmUZlpJTN+tmXGH9SiHjraYsRxKrt2V0/QQuXMamjrfxpmWC5EG3z
g6p69C8ujs0mvV857IjtcZ3m4yLpdkUwp5ozD0/YRhZsB0rBxwh+XVU8OMzrxGkI
GbElzMdPxl+FMidXGONFD3MCxoEsImWBpw0Tb/CRlP8QoMzj8ipNUpjaeDLezMk2
xxPtPwKJSCqUZ1miwku+PIUk1iI3VfdB+8zAG2driJkT8F6Vlisu56G3tWgS+q0l
EnCl2sS4gr5KE04weNWuE77EabD2roO3CXKpFEw9Mobjy8CgKmKE6+P0aF1DpUym
iwYyCxlm4TjwX3BjKlt+y6qOKGtXd2QBM4VLkNDXyCRlOb/HF78yRoVRoIk8crrk
zXbx3qJelC6OtbBnK2MfDAtmteDL0uyrVHdCYyyf9D2prSqnJ1NUSY0h7Ahv6CmO
6mh+qmzqweL4in1TF8Fh1NLTqRwHgQcEWgXq+PwbwwJoDXQTwsMNEXGOLXbtKY3j
wNpx1wyHocp8uryMOafCTb8PmWU/oWJNWu8LrnzFrh2+8mT2QjYHaxKGUkbqfa0+
W5FRJF1ftmDeQvO90kSbdrLoTV3Kl2mvCqkihAeSknZWbtXEZnryWM9fxh6WyBKh
b28OOLDubD8GBx6o/vWeI135rUwTJcO+YHKacqn/7b6HWthxIAJrzb5R8VN7J0YC
LuV78DEzn5iLFSxeSS90F1/0K9HD/qKUCHOU/CwLg9uUzJvUCUg6vdre5zucLbww
eV+J9yU0etlT8pyFOP1OL2Rwpj19MCQCZO2eUVOVNYcmrbtMid9htiybsI5bPgDq
hCUNg9ak7JSi6/rbM41lFVIz+FQXnlthuRV98IsFcP9+Db2+RBkyXk3Euv37bQCD
v9Oj4d0Kh4EcHToidOXFk62frHDKEW07v3pw/OZgYKFcj4vFGgH9KY/cpWffWUfe
2QykVfirDxrleoPkHliUMIqR0Z31cMD/dZDJjRO1nYPkMe7MnfNZzWyCS7wx7pNC
FIevvLmDldSYG71BX05+fmfY9aOcjGsomvThSVHe+L9otc9tP4k0VS0sBp3Ni/Ox
CQuDD3nihjQi9Jl0aXIP5V/9QEFo4T9TjDlRT77lD/2nd+MerSNNLSUf+MA2oN5X
cP8t/6hBUajL+Gjp4ZPug6YgxpMi0lMtE/qwXXi1pztAHLkvKscD3Q/Tfwt2DnW7
vy2yyEp+icoq4RHTvFmG7Q+LjP0EtPha1S4MvPRByDnXtQc2sgsB0bbTGdrwxYZe
Z4Fu0TLlgWWyAt+UeXuI9SUaDkVM+lXn5Q2Nd93D4WOKzvy/RFJTkR8eOInNfbC8
CXTtPrEAC+osYqfxV7ti3D+aIecWb6r2Oxat8S+KF03pjfEiKj9mJ0cCpQOfeKby
b1HL++dbw7JKZaBUj26NpgGqWyPu/KVKEMMZAALIlDe+itget9fFy5BPZkj0FiU0
YsoRpM5ttBOCc/5XSNLct6RFy0fIsnp5An6wC/li7E9xstoA9fihXMxWK4lWP0sp
Cvd4ZCx6eJqqq9SwzRcUOCdOHi6dhq3MJax4D5AbH7YXlSSlIW54GPBiej/7F8A9
Qr1Dw68RFIjTWPLTPc2MZ+P4yF60rllo+nhUXfUFdkWZ9odSL7RlHQlrx5T2oYP8
Sw1HUU2Ea0eoqX7xGS1X55wtsd6YsFmBikHyH2NWbTF3FaoCe3pkknEq+pk7Z5yv
cGfFBqbqgbC2DOUxej1UBb1LkkRPxC/m9Le6CpoN4KTJOFoUMtePRZrCyVwHYreS
4/FnkeEEJ43T3+TY24MMTZPpPZcrXb4nYq0bExLDG75qWTB3iCjWKH1Y5UjcNDlK
0twabLnBcnz8gMZoZlRwFItVpGTF3fv5KsQcerbArrL5RYDVH+4cKEbuhej7JSxc
2oVpif4nIgYJQY1Sx3B97B+ex6qcNCB33+3eFjjS5e5Z6sidYtjPvaSqJJL6aHq4
0ZdZFY4N9ieEHSWOeltElsrLKniWSqONicGG3KpJcy9Ucpf0ZUOphGh7sToSQu42
g5pu3Df9DWl0oDGEoEcJtlPhcn7ceO1pCIOnWD9Pf1/y2jKe8J2wZP2SqaOloYVT
HSj4X+7JVm05xLUMQ9Pymwo4jC7OfpXfB8k1X2Fj0TnfrIc10lRQRYe767XxiyhR
9+XfPGlgJ4Fc1EmhBJe/0y2SQZ2D164FA0rIz48RHkWa5iTAuYY+9vtxKZrJaMt7
Y4ScMXiykayTuQ6d6WeLX04lf+KUWY+CdB2fAcBQUwmKvXdc7eQmV/0IVe18n6WW
Tm3kPkK/0EE+XvnYZD9MzsXIjjbpYTlHGnPeqXU/7dga4prLuqxBYbJ2Mp8IDMjm
BYDXZ1jKbyd3YtDInYjpJm2AEBcgFStDB5I6De4vDlOncAdtetp8KqcSlcUdpdeJ
FUMvNUe2bfiusChCeyjl2s0xH6FVGNSbAS/JqEx0q5swkZ86UZtvo+pgpIkFKWq4
Kv7p52ES13cuepgKNYFb9M7C548iNANASSUgOM3JTqT1LGTs7x+R9cFHpbfuE0np
nlkUwvRm/kaqRN2G3lx2g5hD/G8LAtyxc59/Uj9vxiCy2WeRLpXDqlF1Q21EbLwZ
Ide/jp3qe8LcwMlWmIBi121FdnOPZMpmaDJ7c2vlT3rFlcoM3IwMlT/AN2VRCicg
goWJ16X0C+/mdMAAEmjQ9OIkUp2eK2hkGcbZ+gZDNkZZR1DoLuigFEbKn9eghAYQ
Kl8tlbJ6NK7egz7SE2jMK/arwpi5b2L2kkHV/DEwfsDG6/2gpMcgTawtIcwQSikF
SJH7GJkFquvi6qpJI2obBS2eoCvG0KQP1FjkMpqO573IWL04BhXOxhH110thjGjL
ef3EbImTcEaSOawKfFkcwF3kr0zENiR305IVQC04piZej3Kxuc3gn2AthlkSRTcu
r2b4o953UUzlROVR3voiaCqJ25zgX3Oda8nss+fPE2cVDBYpY6MtsJo64HHvx34d
dA6xXUC2wGiNs/vcwWW7wS+sNBAuzQSIbGPzSezF9xXkeR5uEzqZ6HMdMkeVImY1
y1Vgo98z88Cya67TtHcFzi518tWDY+5pXA12Px87V5pVNf56cjlPYubLRH/nOGZl
gWa3YcpH9WN9SuntJJ6+Ui2eYxUl+hvUtl8uF+cOgWU2iI90BOpmhmIzBnIEvXQk
W2xhApreXfu4EEK6yb0gfBA14xJRx5XpGfzXAzIoT+Qn5yKT1cuSLHR1lTiwYdcK
PqjmM5lBJ8MgYU0JT+REImUOXkRRFBfA0TC5Zm9sISGr/jVT3WcP7UnUeohiScFQ
LMUWxUs1pKCmQl4eUlxcVvQ7NjqgUikF+xmGSa5mayc8nyjxH+8/p3HmEZWj9aZ2
+9pZKHMg8Z4Xz5dJr083eKB2lYGABL7n6uRh1S+7o0E0frzqVmOJWDCiSlzPg8Ps
B4lGJpS4EuwxFkzcE7qNCY17AKi9KDDCOPp1Znmq9t2eJYOVGDH22z4BbeutaNtm
TQsp/ZhWYi4znnKB8BGdJtr+Q8qMSi8Etul9jaXTwXCM/wykvdUcX3Fa960jIqad
xEvM1IO5WYQoZoJQE5L/tSAhcZJHg7gV+ovJcPaO2Ur5h+g3/+CAXMsy98gE6huQ
ILDuq4mvc9240VmnUPRF4un4qdpdbmB58DEWmibg5Gf72JzYE7nkPerxjL7qUeTx
x4r+0iwcE6xS320DRim4Bb5/zzXh0HLt0998wMxoo3kHI29+HsCxcSb/7+dpLtwH
hu5miro2jAfmuh3wJGHagc/nIUV2FxJXCMqlikxfIvq19kBSpurDEm/ZHYvWm/Uo
6SI+dpqGRugEPtVXF3BNwB8IbOF1GYD14Szf8i6H0DYuMReLrdLlqGfTpES7dDmj
3qKHP5G5EktUiU74miEvVs/QzZgm/Yg5LS8qqy5gywUUzhkcANO26lx9aEJf7COB
m4D8az7Sdw8HPabPb3lQiT3FdkW36WFlfEmFwS9wB98IASQOhJqmKitACHdaH8FL
vlYnfnvkiBmD81ZjCO0GOb/T0P9XgTjbF88fDIFeFsOJY1mmDdJWl9GBaW3C8yH8
2+YBG8HNh7i6hyRDirmZxLSyAgLEeIf2Wa7mhxoKCmn9bpqUNIq2Z8Vwo0zC5Q77
gDSjp8ukFaJzysxq6rc88FIEFDOcX4QO+AxocvIceT8+9cLFYMuseC6qZnsBATCg
wLsH5FvxVEtrsegwEesxmNNTvXBUmj2aiPhfQxCo7fAIXgtWydJ3msqLPX1aM6km
XI4HTgh689Uzif4PCEPyBhN2mxH7vR0RfyLdcvfMJ0b/LAeFuo7a3NNentEzY41C
3/3FZZBX337iTxeVbPIwQ/neaOnZEASYpPppXOtZ6BetiMherNKzskgSUk7YT9Zg
A9jdn8f5UkpO8Qtail5Q+N2uI/IsGi4RvmxtGPArb7/iTsboFWK1tW/46RKxUkij
n04AaZF+t60jUJXGe1G78RqoSBWMnBwD7c26DDwKC7REl/psrZAGZMU2F7FiM3FQ
XZT44Fr46XyH98ehjJ8L6VJSbOwb8HRqYzQ7s6i9sUmAawBaKfd4Q+TlBJjFPsiz
0baR/UkshuA2VyE75kq+bhsEdjIyGeZHj7OUyyTWIwR/7kjeV8z3vzoq/xNgddFW
sDmz2OiDZh63zce75tQLPCXV+tgtaeoRpBiHEGGZ62Jjs8fGOGB4NUwbV+c9e5iK
4gnqvr0n1b22cVJXaTpd5OlSjLwmV2dciSY/Em2ZkI81kD/tvJa9QWSXMq1dKINj
1j90VaQrXIsalJoThlgD0TE66szeyELQhcp5KQjBx5T7NonoOtjxd/C8zsn656tX
ZtPTvW2Xnxqb872i+vV4wpqQoHKZmz/GLqk336pQt0bVDcpNRoULGAsADgsBOa6r
Um2X+wJBxjfhZIZqBPPVhukeTg4rZrgeLu26P2RYFxbM5ErLO0Noh/YpFJe0eaIj
tM4x1I/k7umyEIVjd6LQhRgY7mk5RxP+b8fWj46vS3Zp5GKxJRS94waeJfyCn2E+
mOfq/L9ZROwkwC1kHOpvs7mLq4J6OYdV+8YXO9rDbVfpOAN25cCx44vZS6gDZS5+
DrQgf0hQZYxrHSNyyEa35xATQUaoqOOHc+gxzUe7//LR6ljlGX98nqJWUtIf5JU0
vPOfITrRhptp2Y7M1I9DOwjJ0cWj+zuw5LUAYq69SKGcIQ/fQPDUFSg45JjezmdY
Sq9G2MB3wC0SNhDfYPrzkC8DBr2KuhzCKo3Sr+76IGZ+G43xx2bH2sT3C9rhNiCI
0MhfwJ0iUMSOOjxRzvK6lkeCj4MGAkGne7QsX4+QPwDyrvssNEfebRri1ETarNrF
XwdREyzZjP/sKBafv/0+Twz/Nz45GaqWMS9dkJyFFu18VPvMdQtL82Qqa5cxl7IU
Q7xdV18A00ZPeU3zP7aNp1QBMZlX2yQ3zF1nrBOWwa5zDIs+Eycn14FLeQHXgKG/
RSE2uRkBK8XF1Tm+nRzWJufGTJal3pBvR+aU9S/iETTw9zrRBmF1lbs7u7TsjzRF
U7fFN1pbpToQ2EDJVcKbXGeT+vyDqVeuJ47CIsQYkYIPVH7BfJMr94PTwtoXfmWP
ppNqNr9yb1tcscDpBu6J/Lk7mL9xRzbvONvwRvANM3t4Qo80WvGVQY+6KcuJ2Unc
P3Xeke4aTsQWFV5cw1okeC8wjromJ+RmDOwMmXcMfnPAkVbtfdkF8HniTM3zMTZw
ISUA/Lreu8dyCyt34YM69MPc6B0OAp+4F2OLwfEpeVSs8qIpTpoacN6Zb0Jjjkam
lImgMXeocWFZI+ZO4l0XUOB6ZItP+rD6yRdrrVglAQ+6QCLaCRUGz1tK3Mzl1mcs
F+N/dIE0Tjq831mjKojOBC44sE2CYafQ74LgrnK1GdB885I4qKjIt2kRBFUcKYzo
gbd+y5tVKK7/vREOSNR3ZH3kXU3h8p9oNowXp/yn7FbXUCe7lpf58hAoVYeJ/8BA
R0bjKuvBdPiXC6SQ+BOxay3SggA6/3zi5Tl44LHH6KkgKzkLaA9mcg3OP0Z/dWjU
tyl57aEcp+evqhiOwoUTX58nJTPCRT2qMT1W30q83DeB8e8ASLtUjHZkfsrFzg/o
RImeOWoixcUenrWXz1Rc658cR68xxkebEJw3i6EwSVdAxcY2uLpMe7kORS0CzoIY
OAjbUYp9dft4+8wAU2OkI5DUHTLGdq9m9igI14uuo0V5iJ4+m1knK2RjsTRhTCqw
eBJ+GUK1UjUgdGh5cUpt6VPcearVyZf+PuM26QrjswmhQyaEQhlxsowwmwQjvABs
eApggcU0pDIMXkjSCw7DRHQzMW5in1f3R9/EL/jZvSkNr6+h3AGDpeY5I1hOVvy1
WKFBEL2cHITF4GX9VtQjWdy6xdyOFXZoITPxSE5V3m9zgTZA+HTVjcmx9384gk/C
+gQse/bbcR/urzFrU9N6AQmly6lDnFkKgxItB6YLO54EjPJ2I9IZWWDMVEKrQicQ
YNAXr0fj8UigSNMiCpYowqeVN5YGwtRmDftm9wBqceElnYbrCdx74b2cm+BKVzJr
VaPQ6QioR4ysQ9swPuOZOd0O7oamVKvrzATeznIFZlP8NTzRLizPB+AqAws2jC8J
IUUg24fnq9jLrkhGhxljrV0VzIJ29tWd2FOm+n8/3SYfdj1Khgewnmjhd3zDd2HO
fYnay6oWE/IW74v/indhh8jqeiVBX11O2flzgHCkjg4E358DU/DKwTRXnOsKwCeF
/KO1V49bQ+JsQfFQHGo6Qiz1WmPFCaah/nAVpGnFHLntY6wdvy7z6CgEngbQaOfZ
fVJ3/Iws3ttjd3CUw4voiqqwI6F3DTvxB8jXrB7k6u9zN21aKPwVHzErj6NfTmbS
DNrvLugnBV+mOT1cOmaNWLSNgIkYXi8Ht2EyGRDBaW9dkzzaHkmJ0pUWtG/ciYrB
rrBjzUQsg0rqT7bzcpmie3JY3PYKElYbvzHXCaZ/GjuUm0HB5GADPIz4JKPGbyY6
usyXYYj7Q/Wj++JCOtr7Zlb+7HeUDWJoNuGy6WfZy56ruQNr10eMRmLonr8y0V2x
2Xf+XlopimJ68Bii0PZbRXurXTrztHr6+9nFj3SjIulqQxSptQiCTG1C245j7jiu
YxIA42DnrpyxPBG0S5I4HddZir5p48e0RtMJwisJnQB4nRTO6Md06aRRtnX5OBIZ
X8gmW6D5j3qtLtkpHHW31qxEXT5pcaNQ+8tZ1emCkfg+/z5dtlaUnzYBjz95D4WN
Q1otfPU64p0XmUoHD/1cvleL63+cDz7lq5FUTA/j1y7aJZR7WkZfwLWxokj07FDm
CawxvGvTBMJ9+VaKdiCOv1VuizzlEGA0CelCJ7qxU5q7aULGSrGiz4dT3CyZoMJJ
fccA/uYuwqBGFNT8nmLyIwBcQMM0Nq8iCwYpZAeMILmwr8OvUmy8KYuUyLBr66Iq
kUKUYiP/3cffDAGvROm5uG1bZzqp3jjhn/YBC7nSCDfqgjqy+sNS4pgL7ix5qlVk
6MHCfuDm/d51WHC86/CqelezYyRehgtBXDRZxF/zh7Rf55oZsSL3iY51tIJNeTSp
ACYuF/6Uyd6+k3+0MVDwXsy63udR6QCw1hP82uaJ4uG5HIMl32NTNKnvb/HXrmUX
VGps5IxkglaK9jFw8AwQIK00PHMgeNSAwTgS1C7KyPrTBrOrrqa92Ie87ajM8iPO
/lbS8t4+FcZeKN+mO4fvc5Mhbo2OT2eRUte+szUkSF0a+7n3/pPKeQLr/377vkBE
YzmsZrDjPLHq3r4YZJt21/TxGLQ5fDzPxrHCXSuodPr2v8/pk9n8uZKy6IjZT4P+
bD1ImXoO1z7b7pYIdfFMKouFgMZ54OWiA8fp9g+0be3L0CBXE2XjA0WWITeR79yM
WVovV2D+nGrCD5vfbu0rlqwHdeae1KKyscod2kF+UVqwTDXxtsqc+jm16NWi8w54
fQGAiM2Omk7OFOoekt0VXAeCFHDQxSz7PvK8fF2o/ClaNhSdph51foomJE87SeKi
b9YRgI4cTtZuvERzIyRcVCwJajkIGSS2JALih02db6Zw2ylCC4Cflrjk1z8heiQN
2BPusQkU1dWNcgYwNJk7zYiekvhetz9ZwTGiEt/qPMFd5C//EKKb501GpNpk0q9u
iyqRSt35BRdGuGD/L0H4Kwev6AiE23MTLoujnAE35fi2LDp/7S5ryO+NM142QuxX
zWdLSr3ZhxvlAantu+Or3ePmvf+kHtUMvJjTami/hpFMxH2yHNWn0ActWthbwzdV
sGmQT1zT635vZ/2K8ZWbMTX9RvNBV2M/X8U3Oaoiv0P0jtah3p4En0zEURWLSyAY
ucWHtLDNjSJvjVbCxl5aPLOxqC8PEnCc4/sC46eGO3adsjLzz+sbJT0/ud5f/fkF
Fn8Eo0ACnHQAWPjQaquyuZb/kybR6u349jD4d9AP06k7GgLDcrHAcN+e3A4unwu1
kg6ez4nmRuxKnPrKVjUOrNTwFum7UdHp4FS4hOJEW0aOvnMjqxIewD//vOyiFPjE
zYJ/eFGlIzCnp2t+o/rqHzRkrR/BxIW7nVnYsJnqQivn06/KvklH2eRbJB6uWb6A
eMuIVtQU1W9L5e40QG3KXhx0jntNj5KX8ruWy2KLpfMjJGl1INe+yQcI4qbpTcpo
OnYdrZeYilm8vU6qaGUDTopyw4chR8TqtXtODugTLcLRMvhwpXEZg391HfwSvD60
jX7/DJ7XcV/UXbASM40kEKZJGWIFFeKyjYgFoAZ5L2+xlxNHEuQ9hCp7vED7ap2k
hiERgsSUMX/+0FrQZGXj2Nk60rsMCFlHU2XJ27UBrlldIYUPBnIvPJl5U59b2xsq
VxE7hNGHMJsuiBMzNBHQYCAg+wTMlHYGVq4Kb+vhojOVJwJYz/lFINUFEYi9AsjN
apih3Rs1lfa6T+niNVPLYs5GHJEZF6UJRZY6+3HP4QTyUAKWdsFD28fSj3kSs56k
Ae9bHQEqDu9oYgxc8Y3TPr1sLVAtLfoNE+yFwmZcc4w/tYz1tw7u7qJ0SRvX6cBm
eEd0+IVk/EnnW+bIiyVP/SnxFfzKTtRiFlar4y2e6fPgrugrlxeuBK97czqfytK8
dHlStsLPZnbh5x4DRcYcdh+N2cwycn/06kLnTstNBMP+lPp/UHi1MNnGLDdd8/Wf
idDcJ55yI3PNYGFExvPBFnWGba9qyIq7VD4U98yrDvCsYCf4ZzWXrWB9Gs0egSfo
tBhXm3cmJR9KTcr0tUrvYdfwF/rswDAJ/fZ6ayMu21VvaVr3kb6hXM8GNVytzhVT
6+OARQlF+P+NL7oNwb+veTrIe5TUn5gsedzgPjTnuepJghfQPDpQrFgzi8yBKHqq
+SNQ9r+Pu8750+UoK4EpR8psaCw+TVN1kWXnZajc5vMI0mCFC7tJ3mw6PLBFe/97
tHjxYIFJeedvApFeGFqLFX0W9rcQ6/VGF/Vp7X+vFQ68kgYhzffP9TFbwaEI304a
K19xqEEygL5q1vgRkXcCAXuFS1oDQ4/EHtqsR2Ipyn2mcLr3KJhq9fOdOZca7wfd
4BgCVNnakNej/U1elY8x0ZjdcG8ZyArksuBfTc7xSgxpH7rGVancn89gItXoRvoc
OmJhlZpi1TOO5cK0pgKZF6Cvh0sD/X1TnDC95c8RddZNxXTf2T4gitlGOQ/BVUiI
fTfeo90kau2qiz9OSLzPhPGh3yZNRfOMUxzQBj67mEJR9j+4Q79WhYq6b6Vktveh
myPDMclf6C1SrDy27SG87vcAQyxjngVnrAiXT5H61SkTT6eP36R1a81ny1luTBV1
lXLEQzLRtafDoXaC9uOU5OcHU7tmQ660u8zqgjheWVxlZjF24hlBXySrzI5EDpTy
V2at8pJHGVrGYsl0n0Y/O+levCDGcBpbZM8b5XW2zOAmGsZB9CAJQexJjAVnjSN3
RPds4SapU68anByuAoAedcqalxbuUs5i0dS3kAcz1f9ugW+WAqV8xF9rwdy6H0ae
CkISuuclqTV+0kliAA+bH//81aDv5p7QijkrSTyUJWaNC033+K0OT94BxN3ijRDP
Od3JSa1w1lnaLs0yDW9MEemym1mVOv1beO/wPfjYrBcXWKRtErycW/ngo5VQVkwG
MNGrUaMZsJFrixU6+It4gQAkfbOhgzcgMa+0UuJDuXZhesJnjM2r1PRe1q25DN9O
FiTIws2FJQTxkb+C6Zfaoxbw6l9fpfEcxmm8pvONSYiRfT4Vv90tNiSHPrn762Ln
TUy0PHBjuT454fM1+CZfzR+jQ5sdOFADqTBAnrt0h+Nd+nmohsOjejYpEiy6RBUH
1i+ChQBufZ2STKsPKPAcgmL6qDBKFI8ksV/IuFL5Mq6L1Uc1EEnWWReclh1byaqI
UHlqRCN8lHo2CqEMtjYOPGQ/mzPpyMYbm/T3sqxNrLR0GQbIhky4fcqH7vyLC8bf
cHdP2Yc6/FsCqSTiddT48+60np7XnyqayIzyol2f2hgHkeXsnRGhyZJvBdVASL/y
5RM4ldgPfrhr1WCwtr7R9ON+CbaXmW3yXxuADTmiDzSPoL04wFq5gIJAR4DIKTCh
UWF/tD//zekr0DKNIyBo9peUg0+1alsPudLUG/BpTwuxXiZ4TdKm4ISNJGA4nMEd
r9cPEymRBLWvzkeGvKiUwVjyOJaW1ofa62cIlEflT41Nz/LfdjDY1IOO7H2AkGsS
Tea84e6qW9VSp8PDHRxf9eNbUte+5TEhinQsRIKGAYP1CelIykECdAAliOlvHv6w
RIQEWXQX3SFxNpdvc7l7aXxQz/tMHq8W4YjaDRdstQS9qBkHvk5GRffvAxKTgyxl
BJ1/j5t8vkkDjV49hhGEyCkkIjgD9+RrWukIPIrZiZSAZz0VBm4/N42Dog9FLv/i
uOMlUhReHMl9PglFO+kgb3Ur5gvkk5eJwv/AHVtRuHU3g3H/YKyTOx7RwBfrlnAF
AzSTvBJaly4PRTV9bRSIO4mZQC+xACwrWNh9AI0QeKkMvvQ3K/9TK2jQ1Ofh2o+D
6XqGNTky6f2vQmV6VZGUEP4uPNsqcbOI/MjEV0w9QggT8TSkFmjAsyH8Yy2M3/iT
BSttr/lnDi0uzo4TNUSRsz0KHbENcjl//Sqq7RQQmF7EljOr/JCXR8dTHeuXaaFC
TrMnndeoO7ObmbkKJWgcF7OTazEOQlhUvXRWdZdVtUWhTd5B5EBy6EMWNXEwZDx9
BL89ly56GgbsCmuApJ2+xvjT5Rf1EdCnzZONOKma/tr9wXIJ68JtonHXxJHeh9zw
Ux0IOU4hYEWkkxmg/NyjGSJUYAt0Vs2NGjxthE/l679LNEI8fobzRA3NrRJo8siD
rgEN6hhopCA1uechAYX43qLrqrhN0lwmcKPM1frgc/LBWn4n5+JWk/+v/QfY5xrK
VWEBIapbhmFaMU1TOcOYLR0eLsVTriX0infpMQ/owzXbvQgnavquUXY4LMH8Qs/L
3NcELk3sbfW3Ug4gsoon54AiQ77xWipNDTlonGm1QzRjiaqV5qSC/k5B1E1FWRDT
gIhmOQ1XIIMnnZQA+2rtq2SxQuRivvUQI3swLybchURqmhG8NJEF8bL+IIiyR6NO
zzvV8Jroh2ZB1Es51jJUU9mR8tVV1mpsOPae4wPz2uk+1k8eTA6Wrsm/QBXES9A3
+hR/628LcbEFT8O0IWgVTjPdXEAqp/AsG0NmypR0zcX/mgoHVv3mdPI+kBd2wTc/
2kxrCH8q563YcH0gzaCmJ+NE+MpOCxZXk9XQRO4N3I/FqTIQkXj8vijcHlTEVsEq
56LH0kbnRqs1eJ4BAwD807wK5apKZGyfswhYglFA5X+m8JJKECqlwNX8Iz/e0eOH
QgKSK6YA4/D0l7HXd8eBXng9ilU3l7L4phHlFsFQENV/jhBbZ//+3LXIb+TqOHfe
rbZF18hDp6Ap9bP8IWU8be/5JeyYh4Y0/MTapo6x1u39Xq5bOKG2NgDsxTGg0/fO
vzPdEMpFBDa5yOH/ZR22kh6RyjfRH4Wf9B0BoJpzFRfXWhp67dHRPniaF1FgEfbj
LfEXVGP5aA6AqcU8mlX8uYYkI4MNtnn6Jh9Cm3IaWghyztLLXsk6BZgt6sJv003V
ddiFC1EHuKxMbMzwbggbfE1Qvi6KKKbNiv6S2oLP11yYtkgX6mLw2C/nO9IZ2JfO
EGGQg73zkr+jyPAA3JcH27daH8yiFHO+mQnJAiygbDkNjNtG7SOgV+cpzUqOPGhi
7xgUF8aKUmlrWoHnXEhaprt51Nd5cnyzrhAQdUE9t37Q1hlVJ06hFGR3N8qsKVQ/
0hhrOFlIqLOi+PECQ5B2k9sEb/yBhFvdEXKPx6B4ZL6N7a95GnUzDpJQUpXxxZ93
alRm3m39P/DeoKClGzqp7b7JKRd58i45uj143Saaz50RG/bSrlUtUcFcqFdzpPIR
1MPbfs8zl+PC5QW1Arv46hZ5NbAsuuAMvTRncOMYyPE3ZAEz06TKX6ct2YW342/c
nf/bjnKbvp1Q1XGF1wE32U2lRm5k4rAXBlww/dbMaMaw+i0zbNruJEtDf+k2Aicq
VVkzDCd+Sd0qeXe+gUKcexuZt4n3eR4fELnvVS36lezDrD1WIhfPduDymEDVemL1
n6/A4x9o7mJ+r4RC5Zy4mdmowMXtPiSV+XxREdYLp99ElGd+xNgru8+pp4DcGCuU
FShDQ64otl6hERE6YpjEttaJHfji+42zuYRkMtCfPKTwrC+67EBxBOyNizEUFxSB
0VxsXDPor247ueSzsBmNIiFEKyj0eANtGnRqWf0atBJjkb/aYPN74yXF0Tgo9Zu6
WPQX20yOQar5PYHMRoepqZ/uVHnIIU6alzzDrprQQzGC5JGKm/JTN2fJHSnPzFHu
IHNXx1Xnp4t9jVj1sn6grdPKP6OHWXV4hwYsDvpJfAUrstmzdzquCIR8FYP3gODu
Di5zwvhBj/jGb51tv+mMsvA/OKsHzlsSbmOBODhjQw17zLtFYl8kLcDYb0AErr4T
rReTofL2t63Zj5Zawb2cRrncFNYxlg2r/1tNY4CWU8hgkGEEXt0FllH+PXIfhv7v
4SpZUA9YPtjDjL1H+OmDnzpwVNd8B82FMJCkpXsCHUJNj0Xhnthbvgsy749UjHzI
OrB0c9veDuMILk0oOT7koBMLMtK6MXqSyEvMevyaRaqBDZqLelsHy51+ikl0DS2z
f3yFP+bchuWW4V6boPmL3MukNekZgaLkeLcVE9xO3yoCbx8b3WzhSF2yEFIV9F9b
B85PpC3AqdjIP2P6T3WS53t0+cHg2UMa8xmeMUR1esrzMG/BotM0WuxUoznU1CMh
7zkiXzmWtjt9twgbK2xccXVkNxALNoETdi+DX1kxSSDbQapoiuXDVIjiSoaTZGt6
3qNTB7AQeyGnmGmoV8yVpUDSGKRr/9OtmgkLo0JYMIaPF9se0d3z0ExKbVIyl9B0
V+nJ32pSJRpNVIPA1nbkdr5Uf3pDaUAt1m0Z8q6My0MCwhLkGjlAoXp9Jt0z6Rpg
oYdHvaSx6kYcSHfNiOuyzV5qMy5C4iZaTpNzIqbDJ8X0tkMkRekzZLcQiKtkF7AN
baKWrQiA1906Usbf/3bUjm3FugvMrieaYs6I8nFzH78CJhMqMdOlzujKyHNcCRGn
Xkr+0Ef4N3O5DH/7UsEt2xlOBLarXRR6DL201pbCUzJV2iX/HrgpGZ8p9OKPxB4N
gq4A1QZ3dH73Qdm46rIrf0YeuU9ysz1EDRAC9Z8itwxAMrgxDnQMZJ8CD0WDW5bz
0I4MGO1th0G8BXr3pSOOtfNQGuTkZohdUKRlO2prLuRsEXflePL3e1Fmkr3/nv9L
WPPqBJDTM9LQo991NnE60Z1Iql5Iai2VADBGEOy+bZ4UTPcUB/Yymyu1K+uVTdSu
7fPkTxqw+8vbMm0owRX3bvnwXWvEVRh6N8Cy5mCaRLsAdnSJ/ZorG4SdawhQpRQn
c9vNA+I5iGUMiEb8sKl6v3G1NX+qapzsD3SnRsvdi6v42VORvgppkOGNC19zFeIX
R7u1D7zSePUrxhvyTUeMUNpEey8lpje/+tKYOUpI2UWzQB9puIcMA5kX3sVRYi4O
EzGhjHVXBb1DSfHsjvk3m4CVxfw39B6ZbjHDZxk6yzhCuVoeIS506pthvuoYh7WV
8hz5xz0poXB6LB/Jou6pKLONsA7rlecrB0rvLepsE8mNgYGYDAfUoRLBhRAx+R2I
mG9fK4MU0KyQGvSQt7FE/DVqSvVCbfhD/mTjTrXimyBlfCrJ0VZxvHpxPqdesQkY
s8LtnGxNmujGjpUIJuCfBI20EaZLmnGmkJJszeUd4G++SRgCu2583Zs9rO9PIb4L
BZnBV6X3ds7hGEKZnSi0I4+Eq3MBVA047jpTXSEBbluc3EYqkOuz1CmPVt27OBTA
/n7FS9OQuAPNf/Vuz8e3MASOWkQ+u8qGQe60GJxQGhDmwrOZwCkwbMrdCfHK2/i0
hX2sMgf6FSdF2LKUIdEXhqnvvuEZr3psDziT+tw6s2XgM/ovdTxiFaopNcJJL2/q
5ocG2WxfJbewRBpn7oOA9uENSqtRZfI7VLL2tvBF3eNYXOgvbcqVWGywFBYFazU4
uiUZI2IusyA1AG0dVndJqIxHKCKtsmYidPUuf8LPWIHfpbWtEPKogScT1GWc40Xi
Z4ZoMJpcBliwFxzRooTn16sxTEZ0Mkx9bvubck16Aye3aPg4RkRMay+7m4MTO2BQ
KZMrY/LWkot6pLEvZsLmRid/ZRgTLCs1YTYvceivZxN9QWR8WC7EDNG9lXqmG18S
CYiiaX7DdM9xQksMmOV44Oi+XiPKoA8WzvzZh8nYzlgyiJo2VsLqDEdpDZSbm5EU
UT5XsS9edd1K70f7UmhRPvWFzkY/Nv3T7JP6RR9u9mRcpRNH6mPEs6MwlMyyKsEF
L9Tlt1Sa7QCRBtu6oQ3Ce9fJUmLAAVzgp6RNZhTY3NcN44wUJXQDkJ5Daxdeizb8
OWaRwjlOrJprs9AZhSki8AxwmknInnW3wVE8uVskGWEGMX2YSBedwx1TvkaPwEkP
Eo8QCbwb4OS2Cz/uk/7/aS+VWu1BvLvdAVVC+MOhQ+qT4doA3VkGoka4ME26b2Ry
YhEtNQXDY4t4XIRpfzA6K8BJwXlvfupVI+o5bqwKnGBnzzZ1IGn3y8rCDAEnY0C9
d9uavKYM4XZQi61J0vSdk/zSHbgt0Yl5sFaNl3GSnE9oDloDyaS2OP6i6YnthJqI
ovGfVq5ncCEogKQOD21Wbkzhd9tP+n5obv9WUqzm3q76XRup71JSE7pRDoI9Eu6s
t91+t68oW5u4n8xApp1QwhBUvD1XTuNk1FQ+uHdwtxb0aO74/u8vfa/YE43BIPuM
qYP72oWTa44WYQUHvnUEWsLUAO7+wSNc2WeoC76vzngAcGmmv4n892RxSOdsUwN6
QluYXJdATEVMMX8akfGC11yiyTI2OEcHsot0bNgD8o86cdhQ1fnWIJ3+g3giaMlX
MPm5dD7uCkXcW/MJJaDct/jIr9Oo3huQh3a1NwheXDBg7LDNGPoVTZEQ9QnLeB7K
+rl55PNd2idVD+9WcnnNARSaNlCmIOjOocWc4A/+u24iRBuVO5iRKtQ4/V0w/iYY
Wdc96Hu08tDAAS+yOjhOgCjEyqlEZB2DY5CWoHHPn6lX68gIuto5N5ClbXCQXOS5
8e9FXB+jgQfvSfgGZc/qzJsoe/ginAW7bj3blxWhue6WsadveXuPGdJCqdxaG1EE
U3NY/mJYspY6gNukACMw5H/eb5y2bzCs92TsDhBiC40/ds8oeoC2y99xzdAh9AQh
KZBzH3p24SqxzACff8xlgOvF5YHS+tS74noYiSpxkL7BE1U9C4lYopPE3yfoe8Mm
isoYR6zGPBwuo9DPrw2lVD/vxouOrAKQduM7m1grd5zs+CN1H9MATAykCqZ8Ds7i
jc/6YFbc6+SWydY3G+MROdPLX0mt8GBXyePV51MjulKdRxmGGBqWw15BBiStt0wE
LlZA//INW3G7m4yekfeaL8/VmuCgMMsC3eAKfjYR4bsGop010FBVK53EJE5vEn3a
mCNrPPpspl3D+aeBEuHfC9pjJm+cKLomUyjljnFg9lfrt38vPyZOhuY+PK/KxwcS
E6zLJKSyLErL8SELarDwWIhmydBO7LVpoiZCLwFOBGKiJviooePhtQfH1IS22ceP
a3eUGrvnueho4fzbHg+dNJ1idMyarPySV7UjOad9Zr99yO1SO3z6uuCsaJNzydLj
PIUoZfGfNnbwPOgiBGVelGShZaQf7YftuLpYgp+SjQ+ZC7dfxpldydeFep8ZDEgX
XeaQClbU/6/Lis/8s1J8PpKyP8QQyCS6nQDDNCD3eBwd4asjqYeYKeSV4/7b8E44
1FtnO0jIT7mV1BQ1r7ZxZtQLneGCZsrmtAbZPBCekqr6+6g6mxBbI00QHf8jD9ke
9a24X5e9v7Zprv+xNbJIrzpkQZay4L1mbq8nKFubKmrKfXzawaYzE1BtJV4qIF89
nZ+8SyGNaQXYNCYCm9hmV4pXPZ/F/K/NJ0YI2W0qbgeV0nWkKU08KAjbj3SAXyNj
58dSI3Qr+NupvhfMrgxkPAh4vmvudekSTuVpO520r+fMKUqZeMQ7HknlA1mbn6IM
zfRDveuHQT0r3FOI2XgGQgFw5568dasSp8xFtDh9ZWJiRlZjZ5WtyOXNn8tNt0pz
XfnVlpZvXmu4kPGCxlerTbyXdxHUthCm3NONHQFuxcVCscih3PL/xURTuYn6ICTR
206nfLgNDHfeUPVQcanf1LMcasNq9FqWwQZ5GHzrCYwPAFmmxhwGne4RvLDtzkm2
FQLmmtaDIl+gqLLxXPUOyapH7gPZaI2Z/qb6KliuXR8rFJpua5+5Ooy/87Yd8dRp
C0zqI4aJXuc9zPfPkFWytN7ly5elp/w6m+vf1TQi/No6MUtvtmurBMg2JA4sPN0V
rbMGjvgfjVNe6jUuXxhjl9PU8MO7rIq8eq7IpV0K7hCwMAFuLSvsjcRCJADtHlKI
9eZXvDO/V7nSncST9bBOzI096riPPsiR0GsyE9nNq6nzki3pKqnY5yo46NVsFpvU
cLpwWh+UzdpP7gWY4bBomrM21UWdTcKK1hw3e8Nhqqg/GkqdH+gL9A5UzsJcGNze
vOHg2GBlfeyARg/uCb0smD5x2vEyCPK/fWYvrWgVPhYQQXPsxpXlPH+sMbiybhJx
VtNzSnal25521SNXDt6z69PIjQlHP0g2y7x2Vj3TvMW+Vwvw+lKQ2PKa6SbNt9FY
eEyI8j0mCE73KRWEEopjVxZoa1ccqq263/yM0EkFhtMBYRiTqknvciBlXy5puL89
ZQNzM8gfnWQP8d3ckNbpje3s17Z1qcxfMhSWq3dgkg3CWWuKBDX+H1ISj+2xfb5U
pcdwrl6ZEtT2qAxkERd6v/inM27hVh4BK23/A/Mf7YJL9kzOcfynVQwktK0T5i0P
GkinmHsOVv/Vd3Ert3J0+/4cEFTWIpwPJRziQJWWFU9SOOio4kMboPw5bf//ISuN
gf3mEhEpQuCHz5gyJMRDEc9WtpGVv7MMrclPrrIF6sCee/sGUrM0QnJzvAqOfdxf
FEyTeG3EXeLVi0DTmgLfxCg8cE30NANxhIzStXBkX9YyQWAkUP38n3yNQ8N/QBcy
ircsFmNbmDA/wo9DLxQVDbTdT6+oBE+9tGiSDtMQLi001jcpu1zBrP/gBJC+97jx
ybbWKcUHNdZCQf8v9oVyAmdkyjZOB4fejngtEteesdG5jtP+8D5b1IRJGlxcTs6J
K8tX7o8PpqfkH0xHpGuIQCjtr6ZZNl1bkvrKM/NU4LS7JxiPcKwtBMwTJuO6CA8p
2T4oU8Y7oQHHNQaOPvEVgYifW5nGoql9HBorZX9VdV844In6nY2zTaa1XpO11j1S
DAw8Wq2AKJqxMFP4rhoJKydlW4XEa3Nthzc+oZGIuPrBRu2MxCQ9YmILDm6wgWQf
raaRLX6A6XYHZghl5jmIz0wZSn8yTW3mA8Uha8D/lYv54hvjrJDlyfsIIVu3gAbK
TY1iLYD0Kxe5aagadOTdTZwFU45DAXKb44jrjgo9C8epXKzHVthhuuD6jQWqfoUf
USMADYm0xnbuIVEfUnerv5kRk8P0MJEQvs5nZj3vuRcjCnQcG9g3xJbpFegF0VCU
LQQ6jg6VMaRLZl6MJo3A20BLlVENf8BW5/afKVgmLhysqnK3b5Gv1Keo81O4Wr5E
P9uMNfF4kl+0TXOZEc8e/TfDWy15ZliWdyGqOobPNDBkGVem9qqeZvPxF74iYKGZ
9DNb+CIsrZjkSXRwJM0E9VTlPbRW9D6vFkHT+Nk8/e84ZMC4UDUFh3GBL0iDghxn
yLMXQDRrqHwEjeWXhALM6tQz3ff7BVqgHBvNgMyg4wque+Xe9ZCrtYpQxm51fwIp
sEvS0QsKmelTFhDC47zUyEN1dkg8+JNbNWLhzeLmK5DOxEDnuUwhGdoVpNEQqMhS
2jiaWkbnOH7SVn6l1Bxk/BiitVh0iOU20N8ZUcDk8osq99fuchDmVgMR8iz15ZKs
b65HhNlbRJ1D4A0/5m8hosZY3Ru8yaYbuHfoW1FHMKSsUnk3txXza1T2e5k9fx8S
8wDl1j7EFAzkyv8zXvAYFjDAwrEJPScrtFKXLxiLmCq0uVmkrbvldxf+ebtJOr22
YG8zCJUgHMMCusYTC6vKI81LWNxEKvIWNmwCX7453za32EWkir2H4KavNsBfpVPE
TUGnaQDt3BUefZvJQ7iwahK7TP+cS0YuYGPmbiZka4p92NG59Gkg20hLTEQejsFJ
PYx53rY6ItPiKQg2i4R3d+8GN00Oh5vQPXlJoJ8S7BwSAjQtEJldIuaQWf0jX/lH
B5ZvCZG+6HyHj+ouL0sEW9EoOBF0z+UDEjfttNWYAlSeZ8OxQcAKjd6RplWVM0ql
/sx2WodJgZz9j1fJX1lmwAvwloThIx8I4QUY4IG9WzocrXV9xIeaDFnMRI4oZM2D
fTZEzrx6KjzVmqTQV3AODLSXuL1Rn4sw62F3+OPDcMpk7rXuScpLlirxdjBc6Ijs
zD1VPHGlYRxTzqw9klb5qfjF5wRbWyU2E8mD7fpMT200st7EYggH9pzJ9DXn/2h7
lYf/GFaARcRZCkHHYg9DucB3OzrDJcfIfq9+i8gRDu17NP+s9b1fKQSU3szIOHhF
eZtuK0B+v+/UM69uFC5pYOUOIHZeWymVk0isjCDt8IzvLoYzGzSHorO4VzMwCElS
Zh4M0CWbmynlOj7HnoCdp6R4npKz7gD/u9xmNlJtlV6ij7jVjvBJc+ZYKm4a8Set
uvWrVny0WRtPnRvJFJ3+Abv8Y7bE9UnZdy6eC4/WJ7Eb7TK8TCmiOqLaN3N27Rhu
8o3K/rniRNvN1XgSuoBdBTUqpi7QjbjU2I4bQehbwJhoBVc2/gaM3onUH1naRoxT
qg1b/LzF25yOHN2Ri+IZ52EH0w3bI88ahQMG73fFxT9B6qC4ODndRzNsj9tNIbu1
nFKtZHt16jwOZLYPIBEs6+5i/ouoXIe/hxuLtbdEWgi8cKHYS3YIVg/8tRpLFYXx
ZmS8YCSEWV/Ewz+V8Nyditu7Qqpf7sLNT8fvNWfcH1L69ndu2KFchr8FXm4XajzW
AWu0KTIFWi4esPkvqnWBvCMSJCLtylEaeqr4C/8NVF9IcVcYSVm46dfXh2ihvKtF
/5EtLXtmrtPqtLLdrpH0xtV6uEwjzcUNvU8y2Z5afiTtTstM0esyhgGB3UtS6x42
iDDepUMCZGJXvBebnqR8pdW6Pjqlgb4rsUnL9NPLxU0NKtEek8Avi58E7x5S8k1G
ekfMPw8WPpWgc3YN3+72sVhiq7QDd/ayQY476/Juu8FysfuBo+aMAKZOlNxxB/XF
IHaakl0dqPmMWFEz+tK7oPZiHJTqLjdNgdrWxEg5iB2j/Chdq4dADw1iCsuVwOuF
y6ldRXUyqcJ5D8iOmevnSnUHO1oSAA3kgnjki7c91yMsCK4dBAxAXD6ak/PtHUfX
HqbqfNYusqv3EosFb4VtFt3ots1CBK+tawoSEvRi/zWg8WRNAG9ZxFktzlHJ8Lhf
4OJR4sYJ68l1dvbhtdvzDcHCWVX+TcF2KEfreE+SKLHhcypzCLbivkXpafvPrqTA
UWbfA5TzKpgxPXZP5SEW5pXdh5pTbEc2dmuCimNYkBBWXq+MER3T3wxcRKWe48qm
eMugFGut/N9U1SqhLImpxqKEVWCA35Ga1wkUyJU4zXABCdvXxSAJzh7+/IxPjSE+
X56pFyak2XP31KSbN4t4OIpcVWd90NB1a/7E+A4RPZqLHD9M+vx048/468tbJBsC
bZjHYhtDYHnm5/s/GLK2cHlH5x1hbxOJBB8zfE267SldF0FMQXFWF889wpqJb11u
zMI4BW4QewWj4SBmYVMILieYbRCmP/9qML/8ZjvKQoDDvsFxMO1uYUU4DDGXXpNd
08k8Vw8+wQD/nYutNr71SxvjTrtiYnTIDLWU73v5TXYOlr3ADoWdFB39mrIjIted
3a3X/w9ZJ9aH80DEzbRQhzTI0Y2HSgVj9GsZBDSrmxyNKG082hyi8O8gvAxGchFl
MUYd/PTLxF1AotrFQRKLc+EapdeRQ+EIARigPlufXaYGUZZ+SIs+fEhDQ9ysT2w3
nB3IYYezsVpr2B7d20XwPM6kE9dNT2mSoFAncVj2FS1ot4+aN7rpOiww7sKso2ZO
jJlWR120aQf46dRszgO2LHxf0OCONPzQTq1bt8E2RQeSBvcke5DZx+1lEAbvtaqU
LzrxfqRAKcF1+Q16fjIwWXm2u8HHW++wxbrB7yLoqUJfI+EIkFAYWY6GCsWXS2Z5
zHvdNp4NjJbfFGrhGpXl/fKp1IJqZ/EA/sUr75ZUz6WS2VKhrfhlTU+5pWIEj2UQ
LMpb82ukLKpqPMNgR4WDL6E5CN5sS4slarzeESjrjUMNQOuQlnPpzV0HUjZbT6sQ
XbproWhId7En2yjC0eDSV0Yt3TKG3vSzA6N8h8o0dfgNsrI7qBlmLIPMtfsV2LKG
lyBYW7QsbBA96XYWNVHbDWNuNPsSyRkMP9F8oKHt4NMc8vMhh4M8K+OG6ELQB1Be
BnOnDMsQKi5Wb0BNURPBtPKVMiB3TJncbFosX8v690KAunjp9Dc6afMBQKIHOtM5
464kTfXGbLPf4PMa31Chh/+k0DQa+F95M0VQVTkc6q0P7wDjt8WwVmnAWTaOdN4/
21tQgBKD2k1gyZyStbmzYkamGsI47+df6f1td7IZajJwUFHts2O4UOT1TEDjz3T2
di1JxZthD6fxtwuk2YB4sj7Gs4pLDK1Ps6JnCRP1nKXg3/A84DKqOe04+JphNwoy
j0lEsEUN3RnnTuQzlweSGDiM4iVlYVFvMPvXGd4EHgXvJipbqRojI1vKqV9ql2GB
/Wd6dd5ki/wBFLh1OmVG2QHaIjmzgAhxXcOvxH5uZRMggC9G0E7b6YXr1GI9wf4v
f02G94PVo3/BSgTkwMN7WnEb6RliqukXZ6bbd/VSnZ1ZQ+Hs4qWRKTSAJBn/1BnW
W7FRB9f6UJsqEivTNe7oRglmj7Xu0VMSv3D6NPjSxOlXcHy9yIb0CopOFYTMNNq2
+rEaME3Oj0CcyLlS1sLKjqLnhFCxuXZbs0JMeA7Tdcf9meKJyVhrpbhHjTghAaZo
WbfS6giFkhCxBDpH5AZuV9Ku57qXmqEYiyRBCSxrKq9iVE62Pmr+saD2Z0UqfJMk
vMwY5ei9RPULfeO20V3ifIryQxmGIUGV8FUVkYz09og6hsdNIuGkXYSXGbeTTwkC
IjCUgD+s7mu1gatLwDQx/KzxvYrVeK/UIQn+FHESI/dcsQv+GXXcuBLrtVoCddG6
nKjGcp35mLIu2KK2mU/vbSQgm/TsCx8fbnNSTyoQdplt3C/SZ48Sa2KDrN3dQbl6
9vs3c6Ts/hGCa7q5KBc+/asVrNbK3/vaeX+FqMS18sG0cWrFE5kIYtmki0Q4vqUy
nfeYE9QdhgmLDWcBpaD2lkkpe0uhVvsA1S61MhLXeJR2jX5JjrgqZ4JUjngn5lro
P1re6DsOItI5b4S5dAGec4rZ6ETzOhGrcZjXjTkl69ttK0dKcuCfS+6MDf+PKeL+
q0xmi18wnfAD271LrGy9P4Qh1bOegtpFRtfKsVfTZS27GcsyedwgUPYY4DKDCNRg
l1y9Teila0j02Q5qpnCdw8Ej4ITN8NEbgIF3R4gUNTCreyh9hsKIfKxzgJx8vHFZ
9aX3FueYAWrM80ngNnsKN0fYTSFRPGYAlmi/KLRMCfvNrkzsFBB6IgTIeUzX7DCU
0xG+E66GZ0qAjGcheU1LWaCfgA5EfPhjvAvRU4UCPu0XuC/F4cHPi94dGM3brVAb
MMXchWGW2XPLO9e4WRE+jpMpfCBIf7C3S/DeWcRK8ROPYj+o+1/0zPNmDWFKvS9u
nu9a7oQfP+p6v+BzTKKXDHUUy+aB/9GQ0LFxIzqs/CxZ2zMogH48Az+tcjhwhlKo
uEyH6U/WtYgCd9z0jN9jMqikKv9KNA/c1BaG5GidnFiwUX1P8K6i9W/NshGrP/7T
KkJaHSHM/8cR/gbUG6+omW6ifpXlTv9ct+eKxAOKFjQVwTgu+h1vofQ2GvyFX70B
IGFjxOFApXXNFeKnec5EnuGPAdNyMe3zsC9Mpudg94/0KW//g8w1gmUjb60ypQvZ
WyyFSSzNSOxxQyh6dgZG8yJPBQP0XlZD0E/yDBltK7jvjyXVhl68HgQ3La1vAC6i
NwXeGsJmmDBksjJZfLmar6DTDApVs+Vkon0WaR31fz+cfeTDaBCE9KmgFF2ymkvD
8eT16Iltwq/CV0lKUoBP+E74afqdzokgrjE72iz1JXQSbHYKohIfHcuBhoZf/iug
j7ZazVw4/LJHrNBvAs5+BtPTQp2MPgS5T8yyKzS5BH6d1HvJKf8JVDSjSQiu3ujb
bCcJQQdlz697QDJ6Z/9qC27LSH8wvohlMirmGkLU7k9+Sf4xQ7HaMs6X9ueOf0HO
OOkVn+km6nOsl9rQ3PL52bUGwYZ5b2MX95aQBVMyExHtZ6jSD0eO28PtMdMUjxh3
fZ++ELPhcfesMcj/inCf8yIDuwleo2w2kxxqYWnsoYDMAC/c/Z1DHt1Uw5baK4kj
9EYLSJ418oH5adUfZQ3KCLQn4SyQttmIspJqDjUfg8izUwuOfqfgt2nqrPJ+OMmh
z1+kXLUySqxywGU9ZhvJyOib2lwE8xfadL4RB1OSuKNQCfVDY2z/feGtm0/dVizx
ouiGc403kY1gLNxcy/o4qDYk+P+/egKv+QHhSaUiOwGYpNYuVyvBgWyLsVMHv/qE
swBtx1bBRHtKlRzvhfdefeBsxDT+k91yRzbeUigfqLLVj1O4IB8iZZUh2krcidHc
8nNrG3n6WIDu8h73LbKh+WtbgAQsgGl5BNvy+Kih9oyyX0o10i8K6OdC3yw144eu
HCA/Iz3lTn6W4BRQtUde1U9rK8OL//xd36/ZHH123zfPceEAuXNiZ0gMCNLOIZVt
hMUicrAXl/tIhuCMCOrD1j2gYacD38Hy/8xAcyidyrCI/0slrxHEtN+FyqBkLN/T
jXDYqW6xXzFA1h6eSl/UYJ24CYRuXoS7WpvjqH7ToND1kgJP1aLrIOaJn45yqI33
46IwuXZdG48DjPik5gacVbZft6K+lacPSlTJC8tdN01sixaEhm5OzJASnjOZ4SeM
TbVFHr5JLZtp7o0rc+igVBMgiowCYFTG4u8HpV6wmvfCDw3HueR/F9Iudf4nXBM/
f057qFn/RpLHSXTUOdqMRNFoGCmDI7rOHpQhIejORufJzvVP5/rD1MiGRGwUBZu+
CVcqzD9cxoNbmU1QI4CY2n+bVirWiwoV0Wr9H37oEpX3odsk/ECvHcV7dPpzCABO
KO2SrhK7X9OD/cCotSdXS+ieAi416IbLUESWDuG6tMS1t44yjM4C8h2AHVfHiTSX
Q0mtolTJjRuD+8rYmBfeqgN3vL+EZle9BHAjbOBsZWSwCQ3As9y8ItS0isgrMghK
BOLtLL9+l8adK2+ZwMOVpsWk2wAu8L42ianYW0Cu7KRL0hhaxhrs+1N349Hm274P
TzBNoweLQZhCGuFgK9RbpY2RHSP8VwS9+JkEgWHJqwf4jQ3yo22qp5JDneOaBuRT
IZe5u1QDjVenHD/DMKivSlCWTT5aX3TfHo9b4Rgq/O0vJ/eqXj9jWurww6u964QT
1dHezqjgPhK86wAbLTCMh1SR1FcKGB2vFd/ebNwjF38RydId8Dq56d6IAvlLwvzH
UhKZFXte00cfclOd2RtdQVNkQyyxyfuXYvQXl1upxn/Rt6GW0V5SsZbXnTkV+/LF
eWYgw4NBorbLWY2pfU5oB2NqFdGJFipoFLYQnY5Uxck4QV+9DiBua68kGXw30nFe
kTaU0S8GQ73LbQkTO0MPSXI18VkwNgVvZiRN7ckvUwK5t40wPsxC6+MQxyBqbaaD
svexVbxSVLo69dkjBSwNf1sI/7/1utEZPNpKqfGBZozYMHotRNMYmYJ6pvm0XJcO
Win6uTzTDxfVMmai16HXQIQz5Qo+7tnhyaJdCMk6NziMoz+8i9wBC7CRwaEHaUl1
K9gHB4ycJdImooknNQSbBbOonEoyUbRWijbUwF7S5z7SLBj9RcKAjgufhkId2Bw9
0bOA8zPARytr3pnSvI45KRICjjRZmWySTTo5pIejyxS4cfr6CIqFYp1RU5ddPl7D
knqra9BijcY+DTqzk8nxGB019LqlhZmw06Kbswbe34T+IpTsLsSxSYJn5povTMix
SYgoyXwqUtpqBIR3l63UlssRhkG29G7opsuIIViNHUwE+wgYBQtU8zA4WAup/ZXi
E+xnAb79/MVUBXeyNaJ0RKh3KCBdK5EDE2apJsaCr6fHur1uvOaspBHa80IwNKgI
8s+/2oAeu1PLbvtzPDllJrc4GfhPPTJ74/f6CyuOSXItd2NkSKZhVhBA/XZ2KtTE
C/NmSnirfp3jyHgMUzgHEWA70At5rBSP4s+C2+0EbGhc3TFcsyVEFr7k8el+gG5C
BmCAaRF0qV1mHE6XIwmEnhCWyG+mHZ6Ux9pI0trh1b01F2luWk+dvf+H6YBPXHVm
hmF9HtC4EpjEd61pLwp17L/mhddPLeMAwZ+TouuP7mNzpcp0tH3TjgWbpmSmyX9+
Voj/27Z8cg6+bTKe6fWmNKQkzcPHZhxc4TJQ5ARmq5gCwq83J+5LCkvU5Ogk51j1
IETwdNHBrEueHmpjk/92GIKscWQzBLJ7To/lgBNwQ2wsUIIyE5mih9tQiT377DCq
C175IcTWs/cGVxkzoVGbTQIe58AZTue8X/LOgJ8qKQF8b0PYl5/GnLhNhrHO+VOZ
OS4C1fG7V8aauiFO+OhqQs2iqaPllfn9DQyZmLVGW6yDpbLbQA22Mz2dODPp1ocf
qDNUg3dwlmIqVkw6/Qby9xFw+YQ2FVDDR9y0HGPkBQsUSTCOyEy1zkENiPLIg0ED
LHLN+W7ajpa7zl7vzddzXURUjQL62mWN8Nr+7iEV6cHS1BfIOLVPM2inyq1yewSc
vks0tmL/CXArWWrc+4QeSKsxYXUx/Q1fHKkiSuQGDh7TZC0SuzI4yI4/KT8FgNNB
NSMaLjWo7ckQboTZarTX/AEKk7/jaNPk5LBRnxQaBC3r/JZX4F/uzmPVnj/EaQfS
6ZHphoHQtoNNVjTTleEBL+1nC7kzXsWXsWU8lC6FZHOVCXJgU93d7VOHw3SiHD/v
i3JKwq4fXR1CKvgMlF6eYEyXrMsdevJv7znWkrdxb7UI9/TceZBtwkekdoZJSF7U
M12VkAusuZ/3SY4CH4CZpywc+jyy1Wt8pUXS2Ow8HC42fkQwsBhnsMvq+4fSC9w0
YIDdfet8W3p8vHfEE7K0h4CF3Sf3gV/0idAS3HqXXukTu/+jZGhsA4obenIYH2mp
6MbIhi6N2QXck+uTwQizHuyhyRggWKqV7AAH32QETMpTBP800AcymZXa80+KjYgM
EPMdBksibrVd8Bqf2WdnzSVepvB/K69tKvVgFAqvtx+2TPq9jcJCIm4R4eK40b0A
cM4tvpg2k66YDHXwAuS4gCNbJX7me3v8cjcuuiegr4CkMfzPQFYOPs3A/0yhBPRM
Yvy1slB157M09BtDhMOE4aYSM2QMNTq/L6faQJ1mAeymjs0hy7xY+zgQa1FV6ZqN
UIGTMyHrbJj1XN8fJHtE6PSrn6/kGJJ2/y48WQMeGzBW+e1PHsFZsRoxQpiOsGzu
bLcboz0IqBxUoTokU2FeNGjJFS+TBylD3X4VexY7lDq3kbTxSRYzFo78Ie8SaO8s
KVZkJnSgLbn+SdYvW8kVu8Woh/TxjvtG66WixyrUxGUEnYaoTwYbhAZEfNxiLFRo
YVmtvceTOIocbrI7MC6zQDd90V2uJ3jgkC01AhbZc27rEilg/nn7rs5GL4ZhT6jZ
Ep9/TZIYVJiHV0rNScQ2TnJINKq/N7s6P4ga2Zbn6cHCZED0anHXHw+n/7GEdCsc
fdNoWMQ5CZum+ULZhVOSzOvEOW5UZXmHQibooJKqrfQ9mN2PzL6IpE4NB/8OuhQt
gWgv1ypENBC4g+vOzelGhH+VqwEnq2PSKzUcTPUo3+uyHGeGsZGDCnRdsxouXv3Q
D5DSljvlLl8TjGcPmCko4pkEGyQq6vJzMn+isJcYOvFeTxAWmNTfs7vl6a67vT41
gtkA15vTreXLaWclj6alvvb0flkmnx/kl8gMEErcvOrmJfKSoZk9o2zTRwWTcPfZ
3oqO9gtdSQnRSYy/R+XHAhgnf9S8U7iW8xWrujQ+4eEFch3msYMD7exj6zbIYxi0
cGckWUnnrMsteAgkoxBpj4ZuYIMdXMzsU3e4snQn+WEYaOL0tdrk02CdmoxLCJbQ
FTYORRLavQ2lrSRv5Q1B0QTEQySVma/4kARoiFmoGn4JMpxfdGRZlHJ2k36L6jAY
c2rwIL86IzVhaCSqY5ZFbfMKZUk7+/bUVo7GOmjLp/2EhpbLeTgWBeD3Wk2xXPGM
n/CyTP0F9eGmuz1RC4FAC6pg0aqN1oCmW+AiF7KHgS0vGa1RiZKQPPhAMXyi59Gv
MOoxIdlPPYO9ll53P9xZWg/hFiYSbqm+OhcqKRvg8sEtgVN0cvCzZdvFtht1V/5b
ocJRr0x9049pOS8c2tUBHqATpf+sGeV5qOd8sPaFQReSFN+/NlVvneHysyBfSb77
Afz6+gDkVqZf7xlWGI1EliYDbR2TtB2mV/C32I3K85J6/HxTa07Vq9GDXaEUUq+3
BEJdAJml1wGzZpXh06CHSu+WuworUjx1N77Ste5gpNegWRCNBRMDzAy8UABmHHhY
19gMJsTSrsBe/zXNQ20B2yQFJmDpqe991ATyktzYgMBqQthm+dOGyb6HnZU0Z8+V
WJF4B1MBeJXwtNipg9DamHz10nJb5zK04N0eJ1dSjHN4zQ06FiK7kBABNO4duYoK
ODg+wh/iSOFzdZpKbYpPLb77CvwwORGDDk78gHHJvci9Mg3gE1ZSQ8MRindJo2kz
zenYQGldZEHFDYNH42dBc6PsJ7aQvQ71hBsAoJ8XYEN3aeXA1hDLnyyqwl7pIndV
lpDa3Q3C763S5DKBmTwvWtpiQTrz/ay8lkfHiGWi5Rdl9ybhaxRw5w6D3QAVAaft
TJEHNWzcoU82Az66TeoPaqZjV26+d3us115N7i3UjGVG5N01M6ZGhSnhBMq+4ilJ
RkjUR3KYIyqA+RoK+jUdqzLuCf+w3yYVDl0HC26TQ3LA4G1SE7CRX3AjEu4W25wB
/eIZAMqKSNO1lQv6rkrKOm/XPAQIupAOTiEdNu+lTXHzAAi3KDpe5L6pXuSHMzkv
dtJL+/XpWcmibvEKBl1k2XZbWeNfE87gvtWecBcANDGjIMBZ3DupJst5KQo27s6m
QUuU7GppWtakxNGUROe0vtwjS9FsTPdg6DiJ84CN81yKmWxhrwyc/4SgaIg6S9tz
Of/xSzRmRs5ZgVV5yd20dny4Hsf46l4cDlY+YbbOAHTlQn6o5XJOTjW2zsZE2XQd
1+YPJpRaVqZBgKDBo3GiYP5uReMjq1afCpDdJ1a6xAIffA0Ic/IAuCpuoLG5zf0p
9gJfoj/ePmbktjcR4KCbUHH7mfqeMDqYmCGwAAB71eAMN8E0aTF4LCk2Ot+nLxia
hSAc2W4TyQhNilbxvd9N9xl00hJJBsH9tmtVFDVwuDBrqxy9anlG+vJDIwEmkvEz
pOsEIjKhMdwR5qu61/K5/UzgyI7K8pvnjnhqDZcNUjTAPjpeWDgWt2fCl97iAKnp
L/Ndj+X13QadGsbl1CeIs7H7VASaliy3IiEJiAr/QhQT8pGZQerWtLzHhHuvH+lI
sBrStT+LORJ2caQOBMO/N7PHQaO11HojIDDkJlWjAChWhlK1hbgZskmQkaTaUw6L
SQfijqftZSYHx52+HFwRDfJq7MHEEbIMelLB7lDzJDc7j9TReW35AIn5L8at+v+w
XrvKIief1knyZmdYnnLbR0NuO6dirDtlDlS7h2GWHG8GUwa8weA6aHlezLeo2T9H
qRbFzKHRfUuMWi43VikMd59VGpj9MuD0vKaBkkORYpKJ8cZkWZvges1ORmjWemEE
J4yAp+/QtCId9q2zgrK9rkkM4XDFwBHQTpjVGjPKjFsFcGpeLquVegSLWAoa4OME
0p1nRYN89hbreqiFtO0JWQmkZ45q3Y4x/RMQQiWuAmEc/VHC0T01/z4Q9TjcFb4e
GJLzFLRkkJwCBz6s+0pnA4BwWFF3K5/qMVx01Pdg5V5D3nGVTvNVnxsc31r/p8ci
LzQNC5/3K8WooZOarB5QhNMes9CXl2H/5/YaqOGSPQGv3pfSlGTcT+T3heQvqll3
CP5tLkAq1W3rE9WleejIwLIAjvUWC01WUMl2Ww2ik9RSxEX28sehm09pjfZG8lSG
KU0JANnXb6/srmHTsl1FE5YwbZkRhT8kaYoXHQZcbcZjQK8Sbh8KzHM2uWLtbVy6
puPyD1z6codg13W+VVM2Mrhq/Qe6U4Rs3bYMj2ubrO6UUwl3qNrbCyF/F98kMkuY
jll/I70q7Zx307MFDge1nqekk0gPdKxX/p645SxU24hN2XLNOjgqCfrASmlOzVhV
mlHWpe5c7J8WLaaorfkPZ3p/I8STKw+7FmQDLLtI2aJUr7XBisBaanSRkNDUfBt+
Q+qMw+kso8R/CtBP5ZDu01gMlcwrfThxtL3Pe1NaU2m1D8DHIJHL1yA7W5lMmFzD
bweEsLDBPEjK2/MYcR6OAwTEKyzIAfeXcAW4hBY/xnm2mFNimff2/pUYl/2FY3D1
0dfE1+/493ZDo7yITkyAGL0attuahlx8G7vFemtCCWCvNP6JtvTU5YietF0VMjF3
MmFJSGvUUcJlhNOvBW2iKbR9r5dpmMaYm1qo/lc3HtOluy8PLBKuUoqFzk2EPiov
/flKeWLVD2uiLRjpFoJ4yIUjRxWGJt7wmT2s0ewYe/4HQhvIaCtSJURu2pQ7rtxR
JYR/1Ne4dSdNl6RgcIty2CgBVtjMyrcEdqtPeb7Fv2Ho6yleb7oCiLjzQXeN9/TX
1wSrl0lAA1W05mKq6xbY4lUsxdq4vN5aoHNrh5GaZu++yDdxIcde9sChb83H6PWH
hKIuoPK1Hhq7VjOk6sZP7POIOMdz5OJpHTqzj7Z+GZWyMqDOQ5dW5yVmpTpCVo3W
LpoUmW7YNiLY3bxbfGY19E2f1aZ+sy0bLewKwnazsf3eWqFvXPQIbYtM+wgtmqyC
BYRU0mRa1t18Lzx0K3hmoqN3IwljBrrQ/W2wiM9u7sZ+nbLoEl25NrMs7L8xQ3Iz
NsnivcRifRhn9bv+rw/DSeg2Qfz7fMTbgZIvbqRumjYLCsJm6LjW1FZYY6sKQYdP
U3kSe9iaA9ngSoYU4hvj/qqvgRhKU8EdawV3fh/oJCWC5XAlTGsN2KlbzdN85dq6
7lZRlMnwqJgxZ7wWZnZfawGJ51ZhdbhEkN8ufw+ciBgtNJLg2j9v7Af/sZ2EaUfV
oUyc2+ReBCi6Z6N3b930vKiVFrvRlUHS9qcW3m121oxnZXw86MYfkeHKv0SwpBGC
oVel3yru278QT+Ch66Csm6wxTYKrT4U+R2P3IyGCVYWMItPtNcqoeEgeG1xfb1VP
D1mS7fb+IhoD9cwP4ifDpownwxqbUSKp2zcL63yDv8urjt0jWWQwRgZ0SsNDbXuz
ftLvOlHaU5HP8GREK8DGYhqyphydLdhcE8IcQHperpGx7ZXksM6iM/bMecZMNkvF
9bBJYyGz646hhwPUS8IaJe8uvJY8n9ZmitzqxRgCd5lW3ro7emZTOuMH8z8Kotxe
N25URqMr459J9ZGDOKQSQzUt/yiT4QiCiQ2bXpb+8DitbgSIuKNAJiWrGXLMKdLn
CRRabKR8fjH3+O4yIUPoy2MTzLrPLvQxm3mmyUBwT1fGfu49NSahLI2NVd4a1NWG
d2SGmyg5zn4qnYcrjKD4t6dHZgiZcLbMAXgIHQ0cuuEUSWLb2tTnGQah6KP6VOBA
uiC6B4OUFf6VmkYQo1RKED/03iXt1djx1e+PDuqSLGQ34X3t2OwFNhR4AmrMPc9b
qjm+IDayUwJkinrOcDI7dly7Cfwmr9VAd4anQ2dyxBW09svMN+6YIEIn6f3fJz2K
`pragma protect end_protected
