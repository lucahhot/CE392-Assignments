��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{j�X.;߅ţ3n�qJ�q�HŪ�/J�e�_,�cܗ�1��5ف���3��g�e��嘘T���a�^e��y�ϣ�޺�IH��XĦ~��j�h�lb�o@O/��`�d���P�c ���6���o��6���T&��ǿF�λ��KٍE�E.��c�'df�
"3���2��F�OR���0���N���A?�BDΜR��Gf�$�����n#~QۋA~t>��s&����\��5����q�@i� �N0z-p�$A�'���Yav�!����
�<�jl�AK��e�0-��q�%�G�^"�䉻i)������wL��Fi�?���=�I�#�&��i{��#��eS�t�Œ;v��L��X�'�v�y�kV�&�7�+�ѩ>u.�w-$�a��3}�-�da*5��k�g�}���%�y�b;Ү��4L�+�`Z�o"����Q]L��m�����g�b���(6��8~f	�CY�|�+14��I����4�yGp�#�?�Nbޔ������Ei�(z��M��Rk�gld�u�1�-f��%�4s���|� ᐜ˸�3<�E&`�@�lA-��	�,��A���M��y��:��o��Nz�Q���E��1���Tz�ʢ[��?\S��|��1r"m&z`��$"a8��g��!Z�5�)�r�"P�`Ì�����W���R�<�}�M�E��N���At�$?F�ٌ�n	�V�m�%	���+*:\7d�U.���x���W���3��T�?(�g��~!g���rM�Ҳ�,m2k�R��#o�m��?k>��U7�-}��`<A��UI�Z���p��l�j!:H�*p'������њm�q]~.�����9J���ϼ�������9��@	�c�Z�,̸�b�4�Z&���2�5Fsr�q��.S��F�Q��y��p��ё0����zY߸��~�����}������v[c�B��TԨ�4����H��0H����j���gUxg�&�q���\d�j�J�oǂj��m3�<%X��qQ4���^{)ۘ�yPg�wϝ�?O6)4U�|�Ւ���_��Wn��˽*�1�C���]=辙F�T���L_;�\�����ߓ�dO�Z2�gh��C��
�t�Ku�������T��j��Շ����E�9Px!�R���ɶ3��Hf�����jn���3���Bo�UG����ԋ=R�T�)���T���V��.�H666�ta<��y�|��k�jc�1�3o�*���:^KZ��m��mm�X��S��O)*�0��p��{MQ
y��>��7AHġ���M��8��(u��Az1�"^���F7*f=�̎�P��8#�&;�Mt:":�xv=tVxaJ���Z'���e ����R�	��j7�O�K�����`|��~��}*ܐ�������Y�v;��;Q/Y2\C?���4K��MU���V��e����T
m0�9o{�-R���l�ț�3h�$D�v�)��3���+�+!cE��
�[�?	N����c�l�F?��]s]_��DH�Pڛz�!W�M���h[xD���%[utX�1k54n��)�3��Y{�QB2�G~fr�J�@��^(���'����C0��?����j��?Ӱ��O�aM���B��bQ�X���)o� !�4L��gTg��_?%@Y�O���{L�F�^�����W�*��:��gH;��,��ZkT�P*������X�|NE��Fd���.�g}�]�2ǻ$E�n����4f˽)&�*�w�E���a����4ៈjS�l�����OP����z�@	���3�@_91)f��f�Fn�>߃��ď�N/����%�����%�f��*ڟY�k<�s�"iyXBS|��T���!��x@�(�!t�X,�^)-	�&�uN�4wkɷE�Q\T"}��>�-Bǟ��Z鮟	}L�3�_׀U�ѽ�'��o�� �G�솈:��^>b��%�祅�[���W��)�8a�_��9jUH��̘�wQ�v��}t\:i&����h�?F���Y�́��,q\9=ӳs�'�06;練�D� >�r֪ug�)
���լ��r���cr��ǽS���U��ɾ��cE��"���k�҅�spGX���R#���E����k�
��i�5_�k��9�fi�s��1ĮL�o�b����T��"=[fI�h�#^���i��r�*�e��VoA�KQEQ���!���ɄJ����$��=�|��+�G��HUwm��~G��� �J߲_I
[S�8��NK�'}��1��.{��rd�N�d�m��@��,L¯�}8{��);�4"" �nX_�CRw-�З�ΛT�؅"����/�#\XEha��H���c&��̵��1y�9��^#_Q�b�1�ߑ���?6��a�iSh�!Q��֦P�[!��w���8F��u�}~�J��;����uX����՞��\����Sܛ7=�$�w�+ħ�DQ�8��v��UU�!7���U'~/'����$�h�kr��W�تH�y��HA���{���d�������np�v�	���=/���9�����d�8�o��B����@��#�/�V=*�˗��@���ᩬ����&)V�
ъ�c��,�I2�� 2K���� �OZHd�imk��p��u{�sqN:L�~g�Ӯ�t��WN�w���=�D��;Ŗ��ϼEH`�tR�K����ӼD�<
K�'�͉���	?���
ˉ��1/ڐ���T�?8^�y��]@#2Â�1�$��E��cț�/�!P�������[�����Vr�z�v�C�p�;d�.ܥ�IU\��,V�U�<_�q1�"�knqńÓy�B�[a�ަ[ޅY�ڳ�nC�0�U��1�ӡ{������� �|�����c�B��T�J��[�Y3%{�:G�ez[}��l]w��	��E�7`6._K��)H�\y�P^)�W��P�p!;K�5��QYhȘ���Xه�G� ����F,�jmf�ƍw6�����Q�HX��bnc�V�����0�,Z�sv�K`��9<���5}|�c>�EOV*�?Lk�)jI�P�|
w�aL��Mx$�?U�]��z��nz��"I}� ��/���=��]�}X������$v�^��c9P�@�j�N= �B��5E����!��_�y����]S }n�E���3���H�x9f~'�C��y[��Yh�RC�\$疭�&jJ0&�л��C�v�B������L�|_��3�ǣݤO�ֹ�sݕ��b+�ڎ*�[�f'��\�{�d�Y�a�r���2;M��p({p�!j�[\��e��6�cr���=�cE��2<��8��d�V]J
����D*��=�:s�z.����R5Ɂ;��~G?����{�cz�!+�F���N���������������[���%�����x��(<}(��ٗ�4���/���D��I�Z�2yS��*^����R���Ù8����n���4�xa0�M)��-rT�"D�a"��8���<�F����B�h�BV���Z�5�ŕ�w4��QN� �"���E�����������8�n̠�����h�6��$��5�%ԋ=Kk�p�yme��o��M?AA�R{��z�uL���"��Q�� O_~o�q&X*5��WM�%�o��_�q��|O&��3�o*Sh);:���0=�mŹ^���g� `$�M693���p�s�C�i�
�Ku����h-N�G&.
;F"�xu�M���hG�h��Mb���cR�߹�q�x���lDE��9�4c�1�qn�{�{��=ȣԎ a"'��J�\��Y2�*��W��<$����U��	�H!r�U��,�,.��:m}~-<͘�Go����[5�./�/b�����
�þ� ����j��D�[x�� +'NxX�	o�{d0��*cic�j��Wo�m[�d�kF�QH��UW9Z���c��%��%X�TA�f�Wb���ӹɮ�D�n���@CkS�xW1���3���2���ؐUItYK�+�D� ��*�1�k\�G��l:w��6�|Xx�J06o� ��#x`Mbm��S+3��=��e��t4a!UY�!�x��Ԃ͜��@�����qXl�
/�K6~(�M�EOK�������jG)tT-c���kFF#/&A���+]Z^���C��o�DW�d�6�@=��Z<���䤭2;�fύ�{��t+��g�<��Za�yɰ����mC����Q�zf����+�d58G ��Dw�1\��ˊ�C ��-z��٠2l����q@�/w!�d��q��Xۊ�`(��vR�#��/�q`y��$�"!g�S�n�5ȊV��70By��Q�na��"��L�q޽[�ջ�����k�Ć���ys�����-�C���ޔ�h|��%�Đ��R}|@@�{���[_UA Q��Z:�akA,��$F��T�ò�����GT�.�1�Ls]xK���9An���R�����e!�]�hq�|�L~��!��$�Y��9&AI��D�5���P��{:�+$��jc���XZ��R�و���'Y�if$�U�>)&V�e�wk�� �Qy���5�:n#z�t�D��<���Z�<h��I��)|0����-�\X�3�z���FVo�By�/a�j딞N�P�J�be���W,���P��8�����Po�����[��ԙ�J��x�*��&�f/ɉ��`�Ee�Qd\��ZZW��,N$~%ZL"�{\�d 	�;�t^�*���"�MS�����W߯��ʑ�h �B�yr�X��_�y4 /�NHǰ�U�oNp���g3Ó�X���go���g2mB`��s�[����&o�g�$�$b��n ٩��=�@�@�8���A����d.0p#�[{�����ED�.��� �w�v׎�Ԧt;��h�O�V\�o�����DɡTy�����>�Es-��܆��u��H�1���L��#4�V�_$GC��`�[�%d+�%^!��N�)�ٺ�]�^�D��ͅ�8%��7�
�G�8"��D�������Y�w�G�����t/������T�Jp�R�2�<<�j��P,����Z�WA
qu�_��c�.�綳�`B�t1�����N_�Y衣�����rx�_�9��l���`�.����g���mϖZ��B�Ql�D_�#����L})��.�U\��r�]i�p]�����s5U�i��n:��!����-}y�J�#$~��ټ�O�����{�u)q<�<0n���jD@�1���NI,��a�tc�"��ۈ��i�X�.F�HJ��2�Q���$	k�; uoU�8m���i	ƍɥ3o9]��$��������=�����=��nC��;�H����K�}�B/�`Y�,\ô��y�C��;v� 1�5A�{0�7�����vnJ�3����R;KZ���2��T�e�FQ5��rs�<61v�pF
��Ο�U���A��h�\�.���b�YØ^��%T�V�U
���v�W�
� ��Y߀�w1z��=�'y썻�Y�&`���hY&�F3�!O՝�P�ilĿR����#�:�w8�;{78:�t�_ϯ�����\���)3b�j�V� ��&zQU�U��/�ن�;�I��ٞ�r���B�?�Y2Y� �R�����VC�2h��{Y�v*���yc�=~��'"c�����P�gf����������z�G�'�b &�]�&�$U��Hx �(q��q0*�ð�6)�M��4:��>�������X'���c��?l��J�o[��⹯Ľ�G�Q-f7�6��f�B������~m�#v �3��+#�����+�"H�J���U�#dp����t'���]|xa��,MpN��p!�b�F*U�"�7�\�>Ḩ���&��k��<5w�5vDV?ːqQ�k��\�H�Fp�s��m^���Ӧ=)Y�Oң�S#�N�H�bNy� v��Q ��r�"��ᚚl*%�Pe">�$�(-%*���� �2��|�p���;SG)�Z������^2�/�΋N[�� [�V�aF��&�F#	�$Y�b�T�j���6{�a�����@�;<UŰ��I2�V�D�ʴ���ϤF��;Z�BV3a�/�9#IގI�λ1��SгQ���#?tP�y4��#\������0{raO�����_�:ii��1�rP�ZF.�K���x�u^���k��^��KR0MI��

d#A͟�{,�E�e\���!�X)=���oN)��^���d��I&��o�ӐO��77c%=S�j��HVx8%e���e���H�Oݠ��C����Kߖa��8)Pᆭ3~��s�!.~��ފp��邾�w�?��`|���
:�"���a���s���Y�;�B&�~��`�j��b/!O�뺱0���X��a��,r>�~xDz00i�c(T�� B7\��.�¿��t�X#�2Z���l�t�+�v���+)a�+E�ӱ�fV��>5V|/T� p���� `c^�)�`�.n.�V�v��<�a�n�>Z����[��R��+���H	�ۓ���H<�΃T�	Hg��!�� �!1���_q{;{"3�a�
d�EI=@��
�of���#�{�5ZZ8Ɓ�2�*�E#�z1��I�O(h�]�z��^:���=^��'n����1ʪ��R���rX1�ݰ����Y��
;�*,>7����R��f�y\'#�/g�Aw������g2lD��=�tk����X�V|��`K�ŉ�6
�>5�bV;Ɏ��P��G�_�U9 ��lGl���ߡ�C�Uk:O���l���+P�����;M#q��e�-�B�S�̿�.1r��R��p�C�Q}т�0�6�����%k׮%N3�d-&�Qh�B����N�Hqn�[��.�#�h�|u�_�]��fp�7*rӊWmz;���YN���9G��䋆� ���8�9����6=������ӱc����whO��I�+s?	(x8�����?���R����kv�6>|&���~�������c���CG�Oi��C�&m� *A��HAF�.��a����ק���4-w^ ��Z�s8^K�)R
``�eOoQ�5U쵪��^wҠwG#�/~�oR����� ؄���<J��2�v�ѵ'{{�;�sh�p��
V�%�`b4;�x��&��7��u�@�i����A�a������:�Ue�imxZ�5�ze7�*�[c�1��ή@���E���X�/BB-x��qrN���֞�P.V6�G+�F����v��i���̓��+�1����~�i�!��n�.c#�Ȯ'K��*�=hX�����y�l_s�����`���<��6f�0MBy��Ӊ����}� Qb(���k� ���\�5�}��O�K��s>Q�4hs�̙�n`.���T%����8U����N�� ��ə�s�9���̖��h�x|�*�eݺ��*�"�ы��UW����hns*�|Fy�I[�ڻ¯.���	��\�������8B2��i�@�� ���"����I�]] )&�	����W[�'پ!�,���IbwsٸCj���s]Qp�.��s�U�����)>�W�%"���7Ry0)�y˶����C&�`3>o޹����j#�Q��`��l��N1@������V9��EPD�a)+���$��ע*��!7��<1��x|��u�d+��U�@�h�f�6��?��y�G���Wڙ��]=�u�bﰎ{de�ͼ�����rP��0{�����O�y�"{���Q�=��_�)"���S��-F�*��ٺ��XF���H츸Iz���������s�]4` ���V� ��8k|�_o����_��J%	E��9��o�W�iYZ�)\�&ֱ�[�P��c�<�M��T����|)�y�����aV#�(����p�{Oak����`*���*��H~�xf"���7f�&zD���AQ��vk#l�D�o����X���!P\ly��e�.o�e�ب��c����xOM��Eo�@����u�|���w��[8��Z�fZ���M-	y�4�N�Ŝ��ۼg���Ÿ�|��o]��>c�,�?�����f�2��:��u�'.f�f:�r��M�0'�1����	���A|���	��M[�qƩ��hyt���ؚ�]��ި�9J���
��0F��O̡H9�a��RB���iM9V'�jyS�V�O_�Xb�Ž��O����W����[��:1�}��ߙye�%@��� n,���тu�X�������:�y��~m����}鄆�IB�[15[I~K����l��eV�H�P{�̄����"
�ݠ�����* =CMx��xCϘ�?� ��p�j2�5�C�V����F�p@p��<�� �|��\���!8h�!��+�9I2�r2�y����*S!��8��k��r�v��R��I����?"�_�mZ����[��:�fr��Ȫ�F�u�K�X!�J�[U��XҞCV�v��1;`�dP�;bݐ�֯ཊNo��U�Z��M��\�A$R;p�#�K���S��+�K�Z����RSQ��{a	�Iư�;b�q��K��d��M�Xw0Y9C���;���H?��+A�\��2,�I�Y��)n�� X��4���1q�8x�Ϩr^=�~K����FR���5ݳ)83Rxn�ҳ�Q<٢�Gr��`��
�D����J&򃏨�O��a�m�" �	P���R��N[��<��pY��cz���(ѧgMa�ڰEd�i�yH�y�s���nK��b�~�m�H�������+"���Z̋@{̠QɍX�\U���ܩ�F|

�'p	�74�����BV��}����;+6\�,�;�Ƨ3kv=�e��W�M�N�����!)3������X��^\�ն%�d���{�9[��;�����ȵl��m�	�� <�e+fh����A ���O�WZ��f�;��`�L�q	��T<�����$�ou3����+�j�8Fk�H�����z	�5ϼ`�4r���{��v�+z���g��W��dlY���dD.�D�������X�s2��h�C���}����㿖���3�W�,Mv�L�M��tE��J���� ƫ��h�~�ҕ���;\N	MYl���E��-�(��y겜s�Qo��r�NUV��ՠ6���w����幤��EOƅv�=u���AR�^��
���{��r���H3�X[�R���+������l���Z�S��f��X������k e3c��c�|��N�<�#V�0��O��%]5)� ��{����aT�)�-�(�Kӑ? ���Փk>*APE?�X���A��F2��6�^��Xk�<���!�����S;�s2+��@�{��K6�'�(��������/�$]�P����A��˸��1�t�U{�P�,�J�d[v`%жԍ���o�4�H�2��np��fԆH�� b�_�ޤ��������^j�= »r���!��p�z�IS�b�"?�ܟ�����e��{?-�1L��Q�C�{�)�R�ȳ[�����Gf���ǽ� �R��_6_"�	w����l_6�:Й���|F\	ș���1�,�v���R�*˲?wѷ���c�ų�E�kR��Ie	y02��k\r���_�4�����N<&95Y��9����q�7���g&F�0�L�?���ڍ2������L[7ޜux�*1���FI��[4�˽��֓��b|�S�~��jvP�E������Qe<3t4&����R����ݹS�0@0|S����4���Ac��⚋�b����D/��i9��E6V0���& ,��,5�E���c��_H��˾��	1l7��1������P��^�%�]�Օ�.}E�gz�:���9�ګ�8�9��(W� ?F�^�)A������&�|�����1�T���>#0�������o�a�����;��jW�� �\�2<H�<D0�ܚ�������cu�
�Ns�_� ������5_�UF�>��U3�]g�Ԁ� ���˫���ӷ�@|�������>��Z�.!��5��2kn�e��[O9���Wp��D��=E�+>���Oji��`�ţ���@�)�7��4X��&���虤���8�	U�ͤ$�#:<@\�yc�]�����}(J��ϧd(1��'�{j\?�U�Y}ǲ�v�h�b�Y�I�s�f�~Q���,%=���p{X7rr� d	��N�Z�J�� :�#l��]�x�sں�(�q΃����	ɩw���-g@�:��OJ�cjsh:)�a*i_�s�'�[�HF��ҵ�	�����ü���<.�r��*v���|�Ǫ�c��Nd�Hľ��fDf�Eɪ��N��R��h��L�["����ln!��{t���?6����x��8 ��=�l̎2�Ϭ�L�:+����4S
�ay�M"�l�1����1�����s����*�]S�2ۀ���:��E�� ��������v؆�F�@RV(�3�����=Gq#����k#S��|5��a�����A��\�O�d"{��}d`�'ڬ�����}��ǫ��.FV���8Dm�r\l�{~	u�����;�!㚒R�r_�Qʟ�-���?�nR,�{����65�Cu����U`�!���`+��o�-�5ز5#Zr�����k�k�{�:\��G$J;뎰��ԓ/�S8�������;���l����� K@$��R�pk�F8�p!�-�����GɎ] �����Yu�N~(�����'��b����grz;!)��|�viW2)�)"&�Z�:D�i�)��d!�*b����c�pfV��c4Tr
��}mKِɏ�|�V]�m%����b&�-:Α�5��T�Ez��.8ET�u���QU��죳R����K"C��Z�zH�I�|�Kg-�g�T�	ۓ���j`�����v����UF��Ҏ�rw�|=�Nn��*�P���4��s<�X�a�c�1|Z�"�.c@�y�<mKm��8�Cf&�]K�����J=_giǤ���ó�A�xh"ٺX'#r.��Q�^�����`8֒N��"�-�^�'��K������s�}���Xtr��g�R��-G�+�	�:��L�� |ئw��������ۈ݈�$5�-�"@W?6˧Et�^�w�����MϳM}�j/5~0)xr����U��`��$�'�m���G&�>����,�c�W��vR��81�>Ӟ�Zmd,}t��s���%[9�_ޣ�,۵�C�Y���(?/qk����9��}c�ȫ�&ZM�O+Dx9}u���~N�x��n>?=����q��Q�������;����^8	@���'��0M<����.�����g�����hX��^���M`ۢ��Z�Iп1b" �z���lO�[��j ���W _�F���L�A�T�Mu�����F��sJ	-�I+��ݥcT0�;J:�٫噎�TϘ#2�_6�%	MBc���[&�j�%.��[X�P;��5�u�6���P���zFuۄl�xQ�!zxjM��Pv��� Ҽm.؜����0a�;���mB���(�8TЫ��\[bΖ�J�@��kf��H��R�Mcb�㛝a��Zx�
@�T�hwӨ�[{��_ʎ�+�g&�w҈�|V�Mz��U`unŞ�3?���,��v��`����`k����'�)Α�6sgz���![�r%�eB�����h�
�[J1���г]���0��%��
		$m$� �-k�m{&C��g�&IIK7�ⴇc�(Y �iT>fI�� w���LR{4X�'��*���`ϛj�\O52y[����Qt��ju�>�>��2-<i��jT	\pt�L���n�d/��7��Y�u��>H�N�w������ٺ�:R�=3��RרuЎl�H�ճ��.�v�	������w���w`��Cq;���Œ��r��_v�f�j�A��%��銶b�h`�E�f�~9ؼqC������a�:�}BYV�����6�}RO۰�����	��Q�=n]S{�'(�έ����Dź���qqb�⪸r>\���s�Ss0|ݩ�.\�~�9�@�:)r�ʥ5�[ғ-c�rQg�Zx��|�=د2}
8��Vs���@leй��(���g�}gP���.�������� T`�|���āg�����^�ԓ�}3�a`O	BYIS��1x(���uT�t�u�،(v ���n6��Q&:x���I�i�c�7�z9
Yo����������{'!��s���ufp�Ѐ�?:���u�ر�DO�h��_��R������\����ը���q[�]���];������D��|�*r�'ABm���`��i���;�K_S9�zUE5q!�c	�%,�[f�][o��m��y�2�0�BѫR|�R{�������d(;>�i�/�2잃��F�:��\�zS���:P�������Aet.x!�l�Пa{��jߣ�_%�TQ�[J='S�y�}�Ձ��n_�nw��sv	��ӈ���P��<��Y�S'?�(B�,+��0޽Y��FXu2�J?�� %q�#�i�!>���+��.����m��Xq�]����	hT�ќU�ı8����˸���q8�ٍ���vl�����҉��ՆCWK�[�2ٶpiyV�Ϯ�
�8���>D�Ҽ���Y�e���,�.�%���˅w<W�	�s�v��[�f*QN��U�ls�d��L��
읈�P)LE���v�����'�|ւ�b@ղ�_�N9�(X��ޚ ��W�D�_�▮�k����qHW����"�"4*��P�@���PuA`���"\�dXB�~MK�%��RS�z=	�.��8�=Vh��#pdR�=��ssК�t��:8�k�FwK��c��6�3d����-^9
;4=�����n:ւ�#`ڐ�v���?�y����	����nN��(�ʅP$�4|´k:����&���W/s$�d�7�&Ǎ�7�����ClV-T�]�?j3�=G�Nn4��e�����C���h�)��g�^�:��G��sY$��Jv��3��~?|�	Q��p?��n|��S��l��M'��.�!�c���� 7$��QY!6�F�Z�y:o���Onb��(^�1�@��XعF��Qr��Z`w���ڰc����{�������ST�m@��0�);p���kju9����I����b�|��
]^偄>Rc��1��y��\�Ԉ9�Y��/!��wn�����v���j�8^\&�x�K
{���]�cu
�Y\��N�G���A��w�:ћq����prU���(Cʧ�u3�"�c��n�j/�r����9>�𫗫kd��BVL������v�F�����k{:��O���fa6�C�'[�n_��2�(T��RP��&����'��¡��0��D�n�J��U.j�P�&�|Ywlg�]vO�f��]����V�h%*N8��wd~����%)8�|[O���q��ߧ�-��?U��Zn�.��߳�
��:ٟ�l�p��Ok����u�H��U��b�k�v�:�h2�y��CD�U�썜�E�~������������(-ǀ�F`�W9:pd?LZE��:�k���.�72��v&�e�`ɸ*��f�Qb����7�͟���!V�j��<V�_��IÇ?����Řv��]vb�(5qI����g*��\�;h��i�/]��=2��"���$�'�x���]^�@<��D����L�:M�N���d�'ء�v~x�{a��B�\A�-����%��9K��x�w�␅' @2�;xeJZf�7�J�l�5��Tw&=�� <�[�KH�xn�+遣�.Ll��5�5�*!���O��.�ղ� 뗲�q4���7�Z�'��㙞�{��F��g0�%=�&�g|�E4.8���]�l!	��g�~0��[�+�zYb�Eyw�Wu�z�=����;-Y�������Ԧ��ws2��K�Igw�fc \��c̢��mI��F��M?�Mߙ�Zu�M,<VɄ3p\g���',;3�)oE���b[�%���,x6u��p�s���{%Y��|�i��v^3��޺����������$! �w("���Q�jTԲn�vILD�����ǄJ�I7�ϙ���;@��T��q�����Yt:��Ր�8	�7xs(?���6%J�Z�7;7c/-�	'!�T��u�(!�*R�^3��B�'����%������漢Xz�%^����ٝEd6w���Q�Ӛ�e��������߶:��g�u���K�B�%��&0���Lt@�!5�&����e��N�;mR�'��Kp',t��d�^��B�[�=�.(!(�-�.������C��;�֠�lӋ���?Z�6@����4��}�u��c�1�v�o��������s���gk�E.6Y���h��U�1)�B�UHc%#�{���A��=��p��@n���X5sg{ ����1���9��>%r#9]m����س�x��:�w�����+�z��M��ƕ���(EFI��W��1$?;c20���~��ӄ�:��m�*
�mzή��<�Vc�_u�\N%%0k�j9�QKq������58��J���<�Cqy1�]{��NQj�$ n����v���<=�Ө��u�2����Q$�ʥ��`A��q�tTK3�%a��j��*Bu�9�f�'9�ԩ��vTZPۭ(�YL�@� �]P�����֘�}�h$*{8������Q���yͽ�����L�ىs�e§u��.�}%	L��ճ�i��Jv5 ۺ���n��\��T�����˿xB�����Mgo��	CC]l��G��U)"X�:��>t�cA^F��һC���L~Zl�Ll��iA�Z�e95nA�-6gѓ�9I
OЧ�
X�k���v��u,�E"��F�����Z��CZtR��x���f:���f��r��s�V�8%jI�T���5���4���V+�t>�)�l��6��k��@q)����ɑg�7p���e�V�����K���"�K6���B��Ҏ�Ze/�Gw����S��1�n��N�:�%�jQ:(�1�\d%�}5:��<��q����������z�<�i�1q	{v��HĻ
�y�6����2P����_��غ�/�H����J��~���~0��`�4��'�����m����Nצ .���/�5b�{3�n����l/��`,FY#��g�`�t�|�5�̗�w}j���MFZ�����#L�(!4A�,0��:ݡ�~ͺ���=[Ň���rFq\��	0u��o��n����;=�����]8(���~���_�1c�d�$�,۫XS�����i�:��G�O�{'M?��70O�m�ad�\`j��0@j�
��Ў�cB޽[��8��S��83�����4��H�r����̜�r I��=��x1�KD\_��m���G��[8�:�P�g�����"�m]`n�e���Jz�-Cf�{]'�r�U|���uE�u�A��Qd��aR������^�Ea��;�5�v�|��|�ۣQ�+K0�	�DV?���B��}�؛l�6���7���1c�b�c�j�uϔ2θ�t��c�=D5�����4�|a��j#��$���F����6'F�`�gݥ�n+�N��1�v�߶A����(v06H
�8|w�x߼�+Q�&����`�5�R�� z;W��Gvb�E��0R:`+C{+ww7XߚIK`���a{�5���Tl�(@�$�R�.���v�f�*^x���KZc���Ȣw+�h�|Ai��n�葫 ��n^��%���Y#�mI�)���lBh�0��q����M,�������Jo�>�/�Сp��&Z����c�)N8E��j��9��4���e�02�7�t� 9��j�w �:U�h�5[�����bM�q���┨�FW]��bt�`�� ��G��c����1˂>+�G �����a�����pщ��6��P�����HC$9�7�B�ĥi���G0T��Q�O����y8���"�T�ƹ�~Bs���8iR������\}�'�Qe&�)Y�0�/3�2�T��e�|;^\F�(P���:�:��е��� {f��'�_�+Ӹ�O�|]��e�G�kɵi����<N����y�`��W����+� ��^T�"~pC����}����E~Y�%��}z�cQ�����Um=�Ɔ��Fv��Jd=�B`�q�;��w�6\끉�ì��C�'���5k����	2�@s���HU:�je���H[]�����:����F"`1���鴶��g4��m8D��-K����7p��\��G�����SJR8`�N�K����rk3��ۿu���f���<�����U���ӝ�w΅Mcd9Q�R3��B�W�r|�(�c�w�4C�]�-@R���"��\�y?�Lڼ�ƈ����o�0�C���yZK)���/V�V��"Bw�G_a�����M��b�BǴ�߄�y��L�d�q�{"���R�`��/yv��(j.�[N��*K2!00�F�D�o��톝﯉h��qe�����{�fUӒ��i���C--�y��(�P���fǽ��b(���f.�֢ɞ�=�vuj�#�֖�77&�%��|�W$��UǍmx�����U=���X��J�@�W��2����R�P�Lw���A>>s�	��6𔙝�"��&�$?ޚ�(�!���b���"UNe�B����ArO�U�{,V��X�qǯ��懤ҦxJ>�)�n;������J� �J�A�w:'��R �g��-v���9��ek7u���rUM1C@��H�&�3�7�[2�.�q|�
x�u_���Zh��|���!�*t�o�߅Zl�	��W^����;Gxɯ{R׃����JEp�=����Wn`�;�!a����{�5����~��96��oj0{x<dk}��Ge
��~��σ��\�9d6Aì���4ژ�Lo��5M[��~.�3gQ��͎b��Ƕ������e �J"��p1ٴk�6� 9^�7r-E:�E�?�M8f�MJ�va��x�XxD�ʒئ����������,9]�
�]���rt��G(�
�q�����������${��+ԇ��,k�Y�]��U��t��m�WC� k
���k0���X5lD��#�K�խ��טl�d*qPŰ�s8�Az�j�)z5K��0
��] %%��g��U����3�y͙������O���A���� ��!<��Ys�bV���M-��$�)��f��������z�ߣ�Y����m��Ǣ���A�������;�>��/	>G��ElD[u�`�;_yV���-��"M�C��rN��
�ee�IW[+p�����(�A[��=�}>��!�Y���ր
�q�p�M:��hg�d�"lM�A\���:�;�#���.N��k�̻/�<@4�˚Us%$��),ѿ���c�eb�;�$|������FN=�l��rU�eu�JE��0@�&*^e-TI���J����'���z����-?0;���:>�g�����ԓ=:�F��������$����
`q+͗�C�8�>��x��Tcpf(
}�ցwd/��&),���V1$���F䋂��F�ݻǝ���[s
��6<�eA���>�;XӹM�.=�n�"vC�M� ��R�	8�!/l�������h�~���J�!<�R[u��uQ�s�1ד��|��#� @!��/"ǃF��3�o
V�=�9����H��^ShS�9h��I���.;T�a�x*��=dhG�5�oVS��Ҁz�"��d����e��1�J���+m\�D��	��z��V'H��>9U݅� ��>����%��D��]�� ���U};�^�::/x����E�X��8�;��rK	7��j�
�Rc�ߚ�.'0�~��b2&
3s��H�4?�a��k�xm�D������1�=`|�A\ɜRBF2�̊
�*Ȃ�&&���8{,�%����د�j)/Lc��t�n�`�(����']8ҹ?�6��_�O�H��U8Ņ �EXt�t��!Ŏ>Պ��g����m6K2�w��A"5��:ٶS��}���2��S���b)/�� ��\�s*ج�uy��� ��;�ؚ�8W_C0l����g�v��ù��u��bIi�K�N�Q��qm��l���Q�(��.LbJ�� ߗ.y���T����7��b�[�`�*��S���_*����:��s�}N`�AH�P�`���.G��fq�{[�_�A��7��é�7��c1�lGG/�wƶ<��Z�(UzM�U�l���e?�n`N�|�&��t��+����G#�:b����蝒6���ADo�!���M.X5�`Ocn tn~�G�5�oj;����b�Tq�7��bmg�#���4����1%����WB��3��@�-��Q�)���e�T���^9�@_u��[A!s�7�3�)�P���i��-��x�/�ϒ���.��\��3B�%N0~؀��p�)3=���$��I��H:��$�#=�14�$x�9c32)��Q�������e���j��a?5�M����?��"M*�>7��̓�������/��I\�s��>{J��*�u3�������c5y���IH��ЂG��3|�N�89Hf�p}'�q�nt�֣sPO��4��Ѱ���q��I�@���
���De.0��G͐��6��m�Ń������F�32ƕ[l�݇;vbW=�&'�a3��
�kՔ�в�E�G��ɟ��؍��S���W�x�����*)m�r��$j\@���KbN�g��)2T>DRE�~Fs�R�Aiy\�ѷb�+�^�W�~�Lm;p�;�p���|�x�A+Ї��E�~����e�����;Ȉ��������d%����|�:}���QD��W���tyl4rg�2�!�A��T���*�� �,��|��程�Ym&��������k�W�/� ��DZш������t�����X)Yx.z���W��o�eYjoD�P��&=kQ�2_����cۤ�}�v���.����|��)����~~�]��J?��k�uv����腋Z�$EW
�|Q /o &Z������(E�i+�J�?&��͵{SM��5J�͚p�st�^��0 s�n$o1�(%s3�@���r��/�↨�-��	�j�9��>ڊE>bY�X��x��$��0 �!���7�aytex3}	$p���s"MGK��l炫�ԃ��/\gv�sy�.��]t����ծ�I��#Q�يC�,�VC+-�U�V��R��cd�&�_�_��t�@���/�5o9cO��L1�>-�3�c9y=���EU�_����'��Q3�ek�M5C8��� ��u��}:��bt���u��J��|�.�X<~�����<;���:*���Fc1,H
5�Թ:"xSQ���;�ZmH�z��nS,�P�n,�vE�+h͖�u���y��]��k�)�ZV��2�S��~��\�x17�lw[7�\�}K�ښyB�%^�9�3h��^�ڡm�5~��"����D�C�qc�J����W���ƽ�{F�Q'=���T�/7KPĈ^;�U׽��	I;��#�!=��}���c�<�<�Y|tt�k��8� e���MZ�gbp9����*�\!5�̟^@��x��݉�Ӓ/sT�6�	�����P��J�98?����ɬ��U]�wTSZ�C�{���0Đ�5{� Y0A�j/��-����n�i�=��Oq �yG�9���Nςov��w�����ʒ��1v����SHζ�F�U�H\���D��'2��!�;��Ɵ�Qm�֬ ��u���A���-�3^�i�*�W,C}�]�+�h� S�UH +(!*�^Q�J$'���͇q�T�g}Hs�!A1 �Y�K��L��OR0S�;�9���)���aU%�� ���ئtkr�5j�m�ȟ�N��n��҄�▵dÃ1��a�#��ְ� ��1+�2 �2��I�c��#�����j�l8��i��6�'/���f�{C�u��>�V�����q62��mtc�v	Tڮ���fɽ٩��w�ܕ��2ƛ�~R�9���)ݯ��K����^��r}���{��s��/���"�Ԃ�E�Cj�G�Y9{�hk���ڠs�Fޝ��~ �/��=��}�a:]�D��(10��JP��ݡ";����rI�� (�	lU�Ϙ��癞��� �0XArWҏϺ"�n10��4�y�IE���hg7���t�g*�b!�W�<$�1�
d��U�	v���F��O���b�V>kzM�����0��#�>�|:�81f�]yة�Z��0\tu'��Q�z�F�8�eW��*�0Vf��7گ�zq��ӧ{ộ�'L@���_��a�s�����K��C{��>w����d����!<U���}�~R�d�3M���eN2̑�!#!/��z�W���k#�yZ��zR��*NZ�?�%Y������K�߳K�~ K��9*�(��i{2W`��x����7Q��LT��j�E4�M��}�4�~���a�L���\c:�Ϭ�Es��ȁ�ۢ+�����To�}�Mo�L�9�M	�	�|�,��������@G�m0�ǆ����	�����a����A�A�e2l875ۑ}@#ִ��z�?��qbD�#eiԝ��VVD��ר�h�E���wv3A�Ї��'0*1�Ъ���^�ږA^?i0G|�-�@y�.��#@�T�FX�puD���b�=��Z����'B�7):uȗo�]�^c����շV��_=�	��ez}��ǆ�S�$��:��˾��K!í��g��'�#Rտ�}�N��!x+O+]A�����No��/d�ևB%.���W�e�x`׈�]�N�?���Q���~�'��0�,)�5Nُ����-kv�m��B�_�Hh��1A���e̴�30�k�M��8��WUؔv�N����r���=`@�<��;w�Qt9��Z�`�>�f���Y� šy�h�Z��ma�l�C�J�q��\��NT1���������{
PAaה©��K�\�<B�T�U�G�w�5�?�u�QYφ���x�k������8J�n��ܐ�L��߆���֣��"
{�(n�)xSO	����UU�i�U�B�z�b)� ���HC��s�i����0R��wj	�b���p��x@���i.Z�#}L�3�
��dh�q꿓�W���z}Œl��R�C�M\f�m�z���m����Y�cW��2?+��sK,���B<w�P<�<>H#�����Y&a(O��;�em��6�i�4g��*P�Ŭ}�4���Ο�> � �0i1X���4���bJ��4n?vG
���,oOB��^�/h Y��B�6z��a)��0Z� ؞]�q�JT��[~-����/�q�*�L���G�.3�p�a��o2��y`p[b�ܠ�j���v-"!4Lc�
��ѿb����k"(婙���I�l�l��-})�b�ο�v�;���	s�2>�vб)��&\�I��g؇(*�e�G�xIHR�Z[��.s�)�ʋ0�d��!c�m~��k�u��� �v�~��h�1]D1A�TG�����B���S�n��0�2:���4cY��D��P�X��_��E��9Ue��`}õN_%D ~C�N����s1ை(�|N��UM`��^"C{^S���Tk��[%�����w�Q�׼ƍ
kFJ�����1̮&\�jīЏ�-�!g� g���i���a��-[�j�Rc��Y��:y
`�B�����+-f�$|!�3�rt�x�O��><D/�_�1�D�����}8�q���D�U��[����<����o�����x#l����T���o.BQ?`b;89�7����%>D��V��Vq�d��	�0�{sگ��=��Ձ�u�i}��'ou�[裡y]��r��`ɻ��,�"""�,1I�YKZ�~M��.Vy�<�$��X�m	��W.��O���f΢$���D��gȊ$CX��6z7b��7U�c��PUvC7b��|��������n+D�����W��d�B��_�W�V���,�w�|��Re}���n߽�|*$��+^�_�8��(7�z�'?�� ->;u4�;]�c!o�p��l��E�өWʲ��lZ�+B
���f�g���cixe�@���g����(�r��P����� �W�c_Z���tj8�@6=5*2-Xw�Gl�"������dkk�>��ww��M�b�oM0^H�&"a!�(��M�oP�~��f�ݱv���O$Z*3��b��g����K�[�jG*�auLGhǶ%�0��f�TÑO_0���-.n�_y7����\��ЇA��V�����ˍ�Mn�&g���ǌ`k+���u��C�:{h��>q�UxC<Z(�<�G���j���U�@U�*����-#ٶ��U��b��P�$5���|�h��)����8�n�B����P=����������9�QC��ŶE�~|<
p� ڱ�җ���M_Ѫك�D�W{Q7��4?Z�s=³j���l(ƙR@�-�I{Y���e:�ͯ�J��T�(���!/E�D�CN��r\�yE؉�>����T�ʅ��SD�l���çj>d��;O�d�bh�A��<ge�&�ݽCT���g�5p�7���?��h8�C��--�L��j=M�����n��rp�]a�Z����6q�ǆ@r`
�X��'#7�%�糥 �e�(�rV������H��ON�cL���o�JB:R
��z��޸��;�l�S¼��::%���ܟ���}@\�;�vy���=e2��!�@䶍\ZLP�\#���l��&�z���/*-w�M" �Y�qt�~Wņ,��c��1��W������gZ�ׁ�KL JZ�L,�diDZx���_Dk$D�Ӡ����@���{%y���F�YRK�^×��$!TF]��-M�lfq�=#�t���x��i��ܗ���� ���]<PQz����&�Db��2�fP9�vܝ󉹇nT�W����m�
NA܇����k>�K1�[ �ꆮB���h��@�y'����A�#��1.O"Uؓa�p��S]��YLo+���(ˊ�~y�f0�7�'��ֵ�i�t?G%��(+#�pҹ�4Q2�/��H���%#�/���ǵ����溽��z��P*Jf}���5�%
9/�0�#�)Tv�G�"�@�?E5�A������KA�Ibå�'��W���1�RO��*��j�.Gq�OuR�ir�U���^B�ضG�h�5Eȡh��Ku��{��)����|J� D�&���{�=���lKi/����]5�ް;�:��h���C�+U4�9?*����\�۷��yTN���q\��~�԰~t�q�Wo����^7�ٺ6&���B*⪭��c�0.�>�x��:W�G\�d�{'�b+ɓ�,�.�t����׽?H Yl����M0ƀ��]�T���@��H�R����8�QYO~b� �������.���XmI���Z�����DYUە�"��A�'S�{�]	��e&"+����v�� }0�AҗIu�Hn8̲��3�k^����&�{���F��S���]�<M���F-�qU��e�v�� @뺳�,��7�}#�qK^���.����K��}~�&�>�{�lr"�I�f�w���o!�Y.�*��̅@i��$w�/7���� D���u2sֲ�I���!k������J1�є~�MQ�����~���w{��Z��8�����B���u��X=�$;���\�܁ЎB�PC���u��ג�[�ߤ��=糢�xWv̫�g�1M�V1�_���C�eX�f��%_hӢ�ķCc��Dk$��F'��;���o�%�p�