// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
02tccjxi00OjdhnqjMyfxW1hM+CY8ySI9fi1fBkFuPw9PiEpaa5VHJzAGttQRbhW
q3IW96rKxMF+ODpqbt3G0DHd5RztGaeWECeBblPbeWrPl2SBvU3SnDR49eobwNbs
s7CE40eVDekHDHVBF+QAzvY3/3SWEmV6KSNeNVA4/6o=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 90288 )
`pragma protect data_block
o0OtOsHrPRK/w5w2c2r1yitsaFLN6AXTmgXrDS56RI2QQM2fgqJZO9fKfXNTRaOw
H9Dt3UH+VHzt6UjeK+boKcXMnNW6WaiZ1Apmp4YYN9Wo/a3ZZ3BO067jNkk4lNC5
xwtZvWVfT9M+MpISyKkog8bQpMYg909QUQ4JvWHSV1NJbEdh/DCRvFBRBgYjFGJZ
BzDQzNT2XuANOTDo9rVxxsFkycSq4cc+Bm1Z3rszy56KQlTXTxqv636qcfqDhm0M
vjk8STZUMtHyG8Igd0LmSLoI+XUjk3uA4tOFuuLsrm75TP+6m+f2hmvkuCQir0dy
JL8xDS8SlR9nNqykr+tGDOBbCLCCSGOJ4W+vRvQ1RQZnM/VnLmwkRpkZkrlElGqv
Ut+f4KeRYhyikbxXsmbeVsNkcA0nwLiL6rP9jlPmVb9YzynkBvoMQ8MlkCe5a6tg
yF/a6E1kV/IKSAe1+2Ss1IUBCY8C6Lv5o8HQqV771sFTUwDnTvfRNIVwno9+YOQs
kvi0LhJd5WdmLVi8KrcSlshBlqVuDaH/tTQT/LvRrE4yL3IQyzjsBgukJe8yHzTy
wq1rvh/zlEU3VP1aqJBNpbTA6CPZi3Am0afSzFLV1hJ3ItUxUHupDZktKBz3v4Mf
uxINrT1nbjzRm6wr+jkKg7OJzFVh2DueGnuMD0EFaBYeZar0tZ9OOx5VEh0Yv7r4
9w0MQ4mX0d4Q9zHpEV9BklQIPXGzg5DduijeBq2/H0fgJqATAVhaa3s9Akue4fmA
JM0gg7BWCEU4h+xD6ApCts72oRZlnGj+C5TdIgL6TEvfBOkFhHskxOQ04euCtI6V
o7JqbByVMooNJ7J9EAzsNXmbTQ02hcozFOqgOv1vVaEmfVQXogHXevW/AFogkolH
+fSn8QazvxuXjaD5E0aMmI5cM3Qt7r5iFBLVYf3gym8xMHKcKCV6Dhdoa3H5lRUA
chKa/BlV8XD4AL5ZYco5zeTSTm1TY7UbxvylkHAJmdwwtYt+0F04tjqb2OzqBixk
Sm8L2zJMmwatT1U4b/mJTokst602++lrjqaPDLvDuIRBASnEK2UZW/2Kv1DPd6R1
LshxyKWsRMru7SSV9lruRGsf0iigHcLDZ9ZcdGysgl1wQGnEKDTHXIgReF5OAtxp
AYQba98A4Cp1CFL9P89DWUHQ9CUbVkEN+usHhtzU4JXPln7yegx0uMYNh3/N6zQP
ZDmMDlIw6et9Xf/XHdLaHrODZtN7reNzeyu32UbS7nRbG7aRqwLM4zEbic6ZsDDc
EGABFj02ugn2aHDHSbdbgvI5846pywF7Q/ub8OB5lt0MYo1Nunm7B0FyOC2gHzRt
9Yso+bTBOvIL1u7msacX8SGi38Y9j4ArHTg3zZqO7YKkbenBeWRDuXrxQq5FASma
kbhiosP6NLySPJpIPvIguEnUxYPBnauRwyZW7Quh3fiGNKHcGAmM1X16O30bv2aN
iImspXyooQy5Hvzt2UPnWHCLVYcXcrCBcAYE1iyW+mL+w/T1tGviNTojA0gxwvCY
galsHlQXyqwr9MJGNchZvs9C7ozoO8wNHelWhLuHJ3ldc4sr0oM7opZMSGpSan4F
KvxG0CGa3enuhCzRtBsmhFhpxRrNmIgR2bJ3281blX/2X09IX043Zplm6gSMLqMW
XtWeWNmoqbhinuX9uQX7A5jLfd29XqBC5e9NAyjfW7v3HTrMh21+b14ehHrNluEZ
rRU8kG6d3tET1rtQTyYsCgo2xkJtkEX9dsMCFuq8YpRE48Nm5M+tL9yG3eEjuoUy
kXnJA0E9tfM5scLICnlWTF3VVLTtSB1bXxpIdKEi3qWtGuh3VxfLcbI8QRd2LeTR
HuGQy1d939SRAM/rGEjvYKiyul2ctNAOVDzGD7RdNPUCfJSpI+0b3T+o6GYEAKe1
zOwnj4M71riWpPnTwnluao/65i596/kQ4E1eARhVpWCxDzMmqGMTPFpKWsRh0NZM
bP6shgprlWEk1tfSn270jhovPRMYBtqEqHrVftcpoSBp/+aUR8pwAQUd93cae+ev
ZXVJLzLRD198jENMbqbGhd5Q8QTmI9qkA3X/1SH1IZfjJG4Ei4SFvdmWV8dipEgn
O/SQTOvdhhR4Pat7APFlypybs1u4xJpVZvSBvp6rkQvCllSF5bAPXDOGXBifQNfc
LjTCvPyYi4PWXdwIk6nXu3lyuEiGU+oZN2sOlXaJJYf3m8y3nLCnXvw9735g2Lz/
OJTKjL3grxMzqQw4wzFaaNdzfJYgRHBqmbTc/IRPAQtAMfi67qIr9MaXbfbqc7GC
5E6n4+bGY5mkcUh51E1poQIVDvLHif2WyFO0OJ9r47gIgxTapy2ynqFOyzPobQka
AG9sf+okSCeznvatUAEytHCgws7gZBgv4BrpwB9UDoTdGhuiKiGE5TY9o3CW9/79
KUcyXN3rREkf9HeLOua+px1/5kRF5LiOPi8fqaNNKPMsJzr6Q3eUUg6R42YPMIOl
bUcyIpaUtLlrNEgBl2Vl2Ab0WNa2yJAXDb60cSS0qDvP/FEcdnjHt69cXTNA/8nM
+poi5COOVJDTUzDZAhUem/xeBH43WUAU5788nR+KA6h1hPZW9G/I3zhSBu3km0Or
yy0OqLM+irvAbkBX+PYn6//zzZa0KWj7XUtX9IIrL+LmctFertDj1fGgHHZfMcm1
kHyyg0NyTrr1nFjB6NKiMT2hx1KNsoQu96SHRxLFrreZquegmQh9BRxrhRNEJcjF
75rp5H78mhiH7/sk8ImX5MdNkQ24A81Ejy2GG9Y4W1fip22o48gE5bIhKcrx8T7j
mc6RNcTjOMo7RoXqtBLJ4npmWyMoHacXunyGWWWL9jDBl4ao3eheBizOv7gtzpor
QRhc2GOZTWVbNXeXKDD9iGqwNVmMKxLn6tAQIZ3E6AasabySzi/5/vNRwfm3r5k+
SA+ppmMt1FYsyzRTfnrye+3J2x2/jFjuLDm2fpIg534FjFeFlGEPYkce0U85MG60
RZtv9BKnyfd+I6i6RSz/wo+Echh/BVEtHbzhSX+kdmCp0Huecw+oiJF7CANdUEx0
5HnKqdn4QR0OYjTGINz4wbTukDCntjKiwMtX/yXly5R8k8mcGZSqzu9BuMImjjVE
CWii2JSTEOCVtLJ/soCVkTkA4wtMfo8MDXDg4MNqRNyreJf3k9wCXgm2CO2odBkm
qjcM9WtWmXK9eeU/+OrtpqOO73IcbnNjFt7bEZDGmfSZg5mJqrgcBOYsnQR3A4Mk
Mj2jfiGTl/ZgR5X5JCKEErjYQiKPwO2zUl5EZYCvTLFlvfWuPlgZ+6hxuOmGeHKJ
C0rPR8fKYyjw7Rb6eJFEuQ4q/X3ZQ270CD0sbZ8VGRDvOn/asWqc7puch3Jk8auN
Y39kn5mW6WnViv7w6+ySESLS7SyyVoFm5amo8t+OhWu7RV3Gdq1br13w/LmBwCj0
OKI6wcWBwnS7e2c+fXHPkEEGLYCovC+8dWCUSz3YZ27LsFiBMhRQI+7it6OYP4Xr
rWuALOiZFu2KATgm5xB2prsVvDV8oH3iG8RzfIcH+M4bsL/Y3vc5cDS1IYbdVCOU
Xw8gOkFaASzNJjYhOLK88kHBFNTwBNpfp7hnGkCig+ZRLWKYbH3Ch6V8Ocfz4N9Y
HSh8sbxoe0eeWeFxvQIwLIfEWAC9YCtHMzE9xBlenh4L0TVMykGUb0qAWDafK8Od
PnLk14qIeXOdPZUkGE0z/F2jYhIGKGxYRlBFW/k6KI0FAQ3u3st2ls8pfGgUBj5E
t9B2u5y5HwAYk3+QU0GvMiBPzF9m8cqz/CS192Y5Y2FSuHm/MNf2mqwaEv3E4Ii4
5hbgrTlhlVRFe1hHp/BWFpWMsMSWJqbRFFmAcPO1KpnFGBSg00MQj5pid+zwaOq5
LK6Yr6CoF9Lo37PMjxyJVQPDLTjAIpNylQ9DTtXrr3N5sh8/N4/zvcrAq9aMxHgX
7ZxEjrMnmvj0sj2b9WjkbQWgdv37dG52hABiOiNk9Hpy6usOP2vl8muOJ1j5fzcQ
B0+qzmhi3viMxdttHddIlI1h9ya0Q9FVjyN78nClhroZUgtVAvg5avG/i/q+g94F
P06Fwn6P+nwdPqTebHaTrdbzxKVnOZ4i7fnlMZDB4CG6dbh/81HWJkWbJFwx4uel
s+UjhHsRYrdncN/MqlYO4AjfvYOvDpWZ7Ko+d9BeoWp5U9LVI1Ad12V//sV+AlWE
RQzGUrU9KW4OpKQMT8otekq4AsC2XAOPYokAz1mUuD6OQY1Z1TfG5Xe3ZB/mugkz
pA2iyIASp4CkhU+O67lrgLlAW4UWpAPfnlwgZB7db/cgavndqDG3W91/FaVUTv7i
q21pzlpBk4riOLITKJcG0uShu3OUWUAesB1MmrR5zeB8tDV2Mgc1xjEPUi7SGcFq
FEb4dlMZK1X572mh/U6tpaAwK22gaWNFs5WtAKnQ5W+UGFsUaGVXR0R+HoT7v23E
NioibMM9X6qBNStleaoOdYrzLv0dOWiMqhjoR9Xdf61TaivcMNZps9TxNE9bS/Z7
JZ6aZb5eqTnFwJs3Ay9zOf46CL0bCewVPxJ8Kq+qX/e2MTrgTOYqPXbRwaT1eEmG
kM4fUIAYnMlllvTV80EaM7iSmO39ZA9gZVFvPMVSHfpuEyUS5HkCFGUvtwiN+fW4
Et+9YaMs6Wm896n9tnaRVY3zexi+luh3bOqi7dlVspAeSghbLv6rjKD4LSsY7afZ
Cc6sBy19Imwa44AO9SLdysPeEEMH5Zz59TZNxLuiBs22shZWh3oth/3us+onLCya
5bfeUSxw7rZigMQxKkPpUWyJONlaa/gDomopv8GnAKT7yUg7nzwfyTHPABjxxpZi
f/qvIfmgLvddBp3YOxWIreWIS5UQVFBtlrYOG4TyT68+9kA+zzYONudGw59reXWO
CDw70/+ZgKVR38T+ktB4z5qy8PgBtNtG92GFT278+2iv1BSZzyyxXvmbadElZLEp
a9y8aH3EMHj4+54HqZrDX4x/dxROb7BoqU2uek38BsUsCzz413VQyWNlEjUCFIFR
LY3f5zjI7B3HUfSgEZ1H187fZyeftYsDXT5IM3V8Vp5MhgIsJ5m2rxqSj2A3DdD6
TwmUg3diWZfIq9DXcH7jngcCWe0e7WRwfqduAr1aKBTqt++HKFoio5kNjNy0cjuY
Uv0E2SUvwZTbUcjRvb7meLE/RmqeywOFaoNaBdt23L4cc36dGYp8Z4OUmwJOgap0
kH00qqhs7qB2Fv/7+lmooQY1MxNqMMnztZFiBFARAfTq/3ccxeQiFWlVWZIDxXpm
E4L5opLn1LaWSaMsM1I8S/QSUYdYMS1kXZjuvBI7TVDJQmF49T4G35zlfDs192iy
AwdUHT3He5WNDAgfFuGCOjs4ijHpkmn1aUUu5xG+4KqgfEhFF3pE1C1CHZOQgb1Q
8L+N9XSiU73gUWHN5J4MqhR0fTXiLZUGd3g3/43531sO7aPlfSUnG6WZ+rrGpk6V
lxuiGjMw1/cJf2SrIcvBdHd7c0JvSLiPaqmexIax2vtW0/kLoozHTJFuzSszn+28
2L1IHZhKwEXjKIqMi3JgWYPM06XCQ01PMKboT2BSuhrLuct1Y0zTtuEps70rHENU
omfK3Cb08io7WXPrZKm8Oiy0xYgzkuIBPAXeSp1h1ohb+djs1BZ7Sp/MDD2gBmrs
rz5X7/ZIhITMNSz9X1w27xEA0rhY51udUtrtmikxARCJJh1nCpfuPOJbG9yJ87z2
oUSNSdPTPUitiqzLRsqx46u2RqZd3Fpv/drfPN69IW1/B6rYrbLQjnrs+j4EtBKN
XPGpocVkwRfdLAS/czgJbHpMdfFUXOBjoZeHrqtJpY4nVyQVjcvamkOn5DDo7Xbr
0bX826E7o1WSqLTf64nu/3InLOFuatlM4aPaOBLQScSxQtM15L6qZbOzJ1JVtPNa
j6HKh2QlQy7UABFKgQz1XYUoqNQp4GRoBOPkEgvgJYBFcc2WbO3fDrpcZ2klk59D
FEWyDzcLCd4ex3MPB6A6+IY10M9lsgnPHfXK2QKrXznqDkYbhZQKbFx1wsJbgV0y
clhlq3C2qLXN4V91lknPHeRWnHBvkEwHVZNMtV05UuLpNGh+TsqTnGxGtvELWkFv
UECZPzV+oKbFnc4gAQ47QZynx2gXhGQ3EzYpz0ll8QOLqV1zcfs4f1Q5WCtwrt2H
UQQRA1mdjqWL6arrJ3pguflSbDjc+wOPVTXFJo1pBuZK03GdsrvHMuRs+F5R8erI
VixfwuPESpyir0b1/IuxlRsKHfBzxna7taYnDGcKtrMFy+DJJagdIVKE+dKCa3wo
WKvqa1lrgBKQcnhC/UW5XykesEEGnpzYZGJlqc2UmFGGkrVHosybMAL3XYsa2gLn
TFoUraW4nuZ2bq56MbEgym4jgCBPe4/ZN3o+r93atvlMUaY0TI2olvbmh1sVyZDz
vWvJt+nXMzYjDg8FRRrErAukUXLpf8X1dO4aMDpubKkPmznbQBm9QyfKO4HiLzii
QaU+Eu3lz8pLXvdfb+y86JatCCaR5T2jDWNEom9yOA8NgbSRFkXfGTyKySVUWh+A
vnpy2uMYxDr4sbO6dAg61lTywIA2TItIcJyrtEiLDW9ribVMw2MQpzWD8wgrbNMq
dScjVgDzZZyiRJ/qSeRA5ZW6QBDSENh1BZ4+U87n03AUe+qSsBLPBNW1GpZK/V5Q
C6r6zlk0jVTa6C+HHr2gBJnOArkTrR1g56QEJO6vjl0Gtnl4unQD/8eHiy7AXRrI
aucaSgp+pPVRCJtkRQtrdm1cwhw5CdJtnthV97DIUp05OCcl5A7lAtZqOpaXV9tP
eRAZj+wCTmVfxDhTAw5fcT57+UF+FjBRttDZ2mZmpdB7pcyvKcnrGD9HMsnAvKqp
RxORbpczrItBf0H9CUjEeeW7uU4HfNrGCQJ9RZP3inQqhwXTi9cBilw92cwdjF3/
yYgT5L2uwwTVU5pI8ujtJRNtL2+FearD1t/bx4mHfv62cCsq3ThPXoIkBrvxAnSE
YjeDxDZaKIfBSZUCbMdWr7kboH1KqpxHJXoxZrJ/2dbskMq4N30EydEZ9Wm2lWd3
RxbUIh7g7L5NSCFuaH9pOl1PvFgwHqWaG7knyCygjNPhtGqwbqwKe7N2lyIQ+rWQ
C1VPr3iOoJT2jzYAwMFEV3aON0Fq+neJ2GYYflQkXReRA1LmBysLltz4Pl/W8YDx
pvNKKjhWzkr1OZxUMUI8D9Gq32jxlJqXpMoZHs+gAfzAOJPsBbpePmTLCP+mc93C
fkAI/wCNOvXyH4w8x4FALw/QDQvMBM5p7onYrUmsjoc2q1IC2YRI99aTwPj1cV4g
hVGHWyb7T668k1LBOrU6TLmohh00awmWT+iuCAZhh6okMmqaySsHWJwCmniGv8D/
HmoBaKitpHmNkuCkzBm0nVqlbkPRU70Ww815GLoSUEmQCrzQ45lqMX2mOJVkRT6Q
VYRKSvQmirAjb/w5Gtq6yBB6gTS6IoP8P7npyOV7UexTXo7Y1pMRbOxC+O72R1UB
/3PfMO/I+ziR7rpbdNG64SVd+tmsr0IhVqnY+Bknu2b/AnDw9sz6lPwfm3ekp14s
tsFHt6XeCjM1FCDsNJAFF9VTQlQMDhW/ck9qJg/mJdnGM1pyou0SeSTqVwOfQ+iv
uOouWf3AYKsOxMKqg1USH1bIi01KyMKwqD0dlLaOTvauCObX1sO9xMKGmEv//djd
sbZw5h2kn4Qo2Yz5ZHLcCwWso9+f0i/5RnkeR3BRGoO2HoBnS5UBewyoM0wmX+rS
Q5KWO5DE1cD1AEeOCfvlsZ98iszG37xDdpAqGXxIPRNnkuGxVsVpYVwcbNZPOSst
g0SD67Sqva3bliHN4sC+4T98icou8N8wYpFxpCCVPzf0fqoiXujpcj87UCl0aVOK
uW0hp/3Bp6UleVNFPa5drqTcKg2c9A7hGnpxSfhLMiA6netDCA3LCsNp1wMqTMq8
kCebeWZjIZ7al7ymZ2P+lS7t1KsxeUzid+4umxdyIekfsyf5VVLT883IDpBgm8Ya
UIjqEwjOHMqItb9/i3OqpYkZzrfNhs5cAAXmsgbX5ZumKheB6noa5AeN23JQ6T2q
2Kh+se9ljIVFWJW4uTgYoNjVtkOzEyPeD1h3ZAhh+hCAn5NVysXwPClMbqBW4mOd
4SKEvJf+NEZrTIL4CxP0xsXvzrN+7r9PuhgR7sz9vLbtFK4rwDPcwMHoD2isIb+o
gSIwfvXqVWd0rCRtjqDbX6XW3TYdyN3sSs07/LOses0+VLQv61qfJf2OPwjDhfbx
ysqZThkScbhLcLaeTuS4sD7V666JCTAPAvHzH8YtdlbQVmQHQLJrW3k3hdQ0bXUp
cmZsKRPqHH6TJbFEsYX1TfO4ZWk1ovjg/fgjw2S7rUu11O8dYnLeQuQ9+w6sG2s4
p0YP8u/ZIH5hTJVg2R2Oy4tGvvGJwrutYRldHlF5QH30BmPdMRTD65QNIIkx766O
2wYXfzSFEOqjS1l5fkVkPjjdn5+BA/7umSGfPXewfGOIN4DUSlqTIONDroy1mWVs
V9fXm7DozQxeFJx2P86RkSEJ0NCLb1IsPsS7VAOkNV9pkhfUE+XaOFQ8LzI+J1j0
XH70Av+G7M+jqAiniLxbvRHhOurVO1y+XAMCIvRUIT1hY98Pojx6pHRrkMHBKXSI
r9/jGvu1gQVXSIarvHpb45ANFe4C+IgoQjdrpEcfRQpt9g0nEbpHQhr8/NssB9we
ba5XhnDhTiGSgNR3ET7qqDpcI/grsC3d1a7ICGksm/zD7BwcaBjyAoKMrHNuygFV
/azcdX87MoZQPJHSEHna84bDb5s3snsH2KSXfsu9fdqzy40GIzTSiJtRyR1pEGEY
GBrl3FUDI0pAZ2nvHzqJorZd6qsBqjUaEaI9sSTuvCP9TeHxYG6UFb9+URSE+4M3
SNCGG0WVbRrGAkAU8NQWxceqX0qb8uTpuVM1wn/wo9mXpe30XraB1DEb1IyGwqmt
AUHWqI2BBpcZpzszGkGPwI1TewRc9uzGeZHSJA3Xm4Sgt4CC7VPs1cwcddpl+DJr
d/cqRRfhueP8S6axEtgb1gyHrYhSTtEPr7G65xm/83moep/4fbyJF6Yt+L01QJjh
iClxLWj9zorxLzCM7s+fmdneLU5AHIsV2ENnwa8n4Rn1THEYDNCTMFoKwn9a8/dX
0p0pGtQTsZC9AjaS6oElG3QeWNowNchGeCKQx63sXH5HXOzvaxHwqMxWSweWEbcC
iuTz3zVQ+7UgyjtIPHqkrrAtH8Gx099WWrXCxKQrOdqhqol/0rvpewgpmgQUMqgQ
nJVcinfKfIeIlu43siFfj37Bue3LHdafGR8cyfmdo9je88I5RopCtzbupsEbMfEH
7rbfPDJkt+R6FYKY9+Ou2Q1EOEEBC/LdlB0IaAY1CfFce0KouQYL7lh5TnZMzBZG
RoSjbOFMkZwGf7hKmG6RE/YC/mHRXGJgfcyZQUp6TQb90mYYezVRRvZsKPtaShuK
YgxI8/RR83s6BQa/loT2RnLLIza9gfVo8Yf/zZ3/O2dVjwA3O+vlCxKB/xfXz0As
aZ+LPb26C8ypxe40qAwN6ERcORStqY6ML6EX2nPnFyas/EpZk4BSYcLNA41cXZ9x
ICh62mN6drn7H18fZlGzoyZgxEe1vB3L0/al6eVNxMOInSctW3lthk1eMXaTQdyq
BUG9sgheqnUOj7sXGuHmEUm8P6KusDxxjIgS3zpdjijdJK2MLMStedEceR61zSh4
sa90Ybk1csTm4/U61EG6junrcBDvp+sZVk9SsSraogOwEy1pPNxJ1kpBADEV0YBD
bhp3VbU3xFZRgCJiMspE+UOg4m3/E5wmfE1i+PUQeEMuS9GAl+4xKmt7xszLI4ma
BJI1HDyxME9t2hug1xRSOHcv0EmsFmOmw5YrpU5F8308URM5bn3AqmzwUCtm02x5
fwkn39vVIo4VtaeRhBzbQu+IeNBBTaUdaWS4VDXJewijwup92CQsDVACBHyegZPZ
HD43wsOWhIffhBshJoBu1h9rlBluC9CyIUpOYDrqOqN0hF871CWSNx2T36gja/P5
EdtOSkKUo/0Jtz81hrqRq2ACZBDlHLPrr0Rpo1KlQHp5MUCOcRTZSWB1yJ0T8z0R
lbJ9gktY/qKQgKi4zBKaETm3TV6zSqnDraGvZSMaomE85hngKBTBs3+gdEHpU4wB
zuYlsSToHMLLMNgm4yc7kC3Hh4L3cZ20QAxZcAzzK+aXbdt1x4+uGmy03tl6J6IG
RgY+evAmTcsAO5rLkpwh8APS5zWEC90qfFaXRaXeU4dqxkdTSKdhwE30VS+wlJi+
p7TW/JttmlWq1OQzXddnGaWDeebH0zm7V+f79pKrfKlfNTNqHkg2nQ67QPZjJn15
H+1IMj8yYoAIfcy99SiMrJ3xlylS/Jr6uNDTaKV6YFAFj5eU1ypDWuEwPScScvzR
p6bnPj2JgUZsAJL3fW48TXgZS7Pa9GIWIAWOje1rpygeTGzZaPVOa3VGi/rBczva
Wz+vAjmopUsmVxsh1qIbZcKxsOZz3LX8YUIuuU7Q3C9IYhQysQP51NfZK2R+wpl+
oc+0cZkMYnzvbrzIAc94CXymxaVWVmrutI6L4KQ30/OBsVZBC7UGLSXmpOJ9kp1d
WAzDKNKj8TQ22cwDF7JXrwkVHIlaYHAjl+TmzkgklJr9HMkwsAMUPRubzk5mzJ41
clkNx8pe7hhZTwFIfg2LpziigC+6WyxBxRwkz+236UB7MgZP+pUisg7eE7zQtkr7
LbZPGIxibbg78lKp+gAy872p83a1ng7/nTSPJ8mG9NjK0qzXUmdgAOw1MS3RZ/Y6
E9bhqKCzI/ZkylRSzRai7RG84mhR8JGHlVyhHurHHmAIeE1uLgPJHWHDD8GKOyIX
OTY6kKbICDxMpVa842MSoca8t8i0EdMye1TRqFAtNjXU0IypItmmLe99LJc9edOX
CLTV6tLzxv5g+jSmYlJBODAzfGjANPZqPKq/PuHyoM5BxxhkYIOUDWWLPM/ULqhB
Rt1LzYPvUr+iToxCHngC5QKoMcnYxizYiE0Sh/tmwny1vqiZsk+m5Y1vhyNKlUvB
51c7arRJ8wjzIjZHMoPXIOHoF/dE6QqM/RyqMfaqMqXUVEkrtNLmrjIQHJJqlpPq
luU14Wjo8gURPvPGcWX43eMqTIXz84z79vP69H8BOJ+UbyNC/jGd2kIGrhV1AfJk
WXp/ZY9FxZtoaSvjexZL/6ufLEv5Nv7L/ylKtO153G81kQkWoGVXfrYzqvD4erUQ
h0+VrTTfm5AbRygVB2dQZcDgEqC2h1CFdW+Hud9E1RFierjyu3jz59lywoT1jjMm
KqTi7ksBq59qFPMa6FR6PxOCXMxTcPYKcsq2cr3JRMxTTEwHyltbvy3u63OU6bNM
9AELJTx3gRN8Fh7lYMLtleULRfxjpYGZdprs73/87eNYDcBV/nWpOYCLBFleIO52
+HX+6GuR8wBai+ckUPH3KgMLayru4bns7CFQtzaew7OnGH4S7mYNzVEHby9pnBLL
qTqRaCED8+y58RqIpqWLxvXMosr5xsIxOuniPuMa4dQ6BWV8NfblUUfiRW+sSO5Z
LqzgLhZpwCR5jdoxRtULpQMCHzMbINKqBX2XDQtTe8YFUFGC6tXC2XHUysNW3tWR
J7mEbqjr6fhmkmk4PAT7KkNFDXsID6mBW9bco+gaqgO2LhBjAELV4sk1wLk4Zhs+
gcelvki7C+gGtYn49YvUiX2D5ewPVsJO77ds+TXiaDOHPcVgj7ftA0R/nw/rfr0N
OnPKvrX7EHmKNZUiJMoCtuzSXt5zIN8YQQzCD90FXjkQpiT+Q8PxHVeCMkok+//w
bE3KM/D1yLPsvCwYjMW8CjNBMjfDUA1tI2HTRBIfCicn+07BF9yVVFGsMOVbCkXK
E3GsOlg0aNx1JMyQ1KeFxHKWyQ2Ff1Zj4J5Xnb1bCCdRjynEz9XbzxidjfKCApYP
n6C+NfeTrWrXWCJINylrcqZ6DEtHpAWgvoUWc/+fbJ4eUGGgP8eB6EOvEdOZEkc/
zN030aAOwGGAFQ4Wq5XqBXym55BAPW0W2d5fY7M9LlQN0Ivt9S++Yw3qkBiqwYP3
b5SQgb5mGAC2UrlF8zN11Kf3a7Xlds4qq3Kjqut2B5ST7wayiSXd/9wDhaH8cW6M
xbq+nQuyvNpOXoApL3khV2tb8nYDLl2e3ZFCrkKFVGjB2vDt/jQXBdbYNCzepJmF
HFZFWTkmJOOtCBXADVAwNR/1Q+PUgcxwUKo7yr5dC6qqiZo1iKcJsaVUFDSMFmf+
oteRpOkroMc0pTyNmXmyKSM+t6M90iCc2pW+2o31O46NVXlzmJPTSMsXFSApoPml
pe4I2NW9/MPcOWw39xjNwBuL1z2l/V3m2rwSGWs6do0wex86Q2OENDEhPgmopXJQ
oKLEGKOOYx3pFbFaYNObqg5GDYf8g1is+g0d4KWLtD3/2F/vBvDgyvK0Ye+YPYI7
TtcujA94KNOOcDghiPw5rSgERR+GtAq6C8hKmE2ZRzwvZ9hPn33+adaxHkoOgZ1i
YdUsgQ70MctM2TARtjquBocdVqbCfZuWxDXrknsuMRnf28fp0J/pBFUNoObIIBvf
S430ejcrKn0Ii61hg106aAo+rW2DRSX2jGHUOcC8LrR2ELm7xQn5snsKuKduWrO5
pTs5D905cmTP3YEfaVAYLtJx67Wsr/aCgqxA7xFVhjb8AuhyK4fSYcN/yjzxYXsa
/z/tYXa2voT8PgCyHZKANvbIabUDT/P6R948CpBdv43Ymg5FzwMwiI+swK5WDrkW
vGHXxzLkYA6vZBmMcoe62EFj45ZQ5yYEoK8DfNwHmQDLriYzR7O3lNEhPT/8qZ1s
ozOCQn6J7dAoLeoHv+5e81WJrHnB8BUJooT/nCJQhxE6yywm+SAQKaHJLDwHzm14
2bIHDVf+24ZV8RKj9YiPKOdTGa7O9BrceTILMWjYylUbuTTX8tx280neIY8N8w59
CRFq//ukC+Xr2AIPY9burKmk7q4XkuOM0/LGvylJLxeGIx8+yFCHYeieYESSeDDJ
DFI7/BPcFRSp1xstsAcInhCMC8klYuczxrqY6ujTdoZF162Yi0PiK5EZQ4QByNNl
R8d5KwvE9OmTpgt4EBk8NALKGpZPvr3I2UgGrW2GDynewjA+BO2sAcABKBN0CRvm
94spdLidA+elv7UG4tyE6FAjO8VehHwDoLS+ydPAD0BUVgxt36PN+SfsWUr/ZW3L
GTECQPt0bqoWYEhZv2z4E67IgGs56K1C36UyCY4iiSd6wpvt0mKvUDhSbevxeZM1
i+hOPM0HcKm0fHPd2jcFoP6DvxBbRk57cvWON1i4WRvNoSYbidV6wbhN4zlK1NCk
L4cckYsAESbGwLU5WaTx0uOGIbWf3TNB/68arh6Dufa+5iGPQ+LRJXhRon3teted
Jf0GaL0Iz0GWfLtdVtDF4warmasID70oV60udtqc9KnDWSKH8MZ0X+P+ycIn5H/g
eYpdSoc7F5H6PiCgkVtJZ3TY+KFZreEmAIlB01l+kncmiGhEx14CxP6pRdrxYQne
SpKFs/1BYxqvbQpvArDfbfUzuOW0QlkiueTVgCiDCPAoqfsvBWhERLVq2w9F8cYS
33Wg+Mb93ExDXko0RCTrojhxSRzaapLc/o4anpOX0LzSqf23r2WYaKZHR6kYgj1Y
9wgqHdfhyIjX7aXUhxtdrK6Ou0TM310L1ZRDHX5/MbgAEJMIe9m2CQ3PToNP9EeN
qHNIH+wN9Ev+4tB80eR2acdKHg9daxszHDdqcVCGrz76DsSBx6gPmCxCGl918jTA
/pF5JkxHtEDr4M9K3UzoCo1XAhSgYMpr53draYMSBDCmvrY8t3zy+5N0LVlRSIaw
lc/GHNobGVs0Rdo+6whMJ68fcIRAlpYh5PPqeEdtKO9Q36ugWC7KIYEZNqTwNUZd
ZgGEf7pdAVgIt0n1VXv60dR79LK3KvSTx+Yjn9f7iUcJzWZKuhTmXc2yrURHtEZ2
31upw8mH0bWttw5Khmrkj1jPpc722RnDrxT3znZSLmqgpkkIRIsByMhsJm++WwTu
+cX6j/9SKpk4Kbl1PI8A8zzVOu9g18ZjxgQ0pb9h/7YdrVwSLPGd0fv9cUMInK8e
c//9rIaDfOtxVpbk6MgwbWuvXk9NCVSv8nwuFl7SgF3ReJQ2ahqYk/njodxKgLvX
3NZSGFUHy5gs2iYZxxTLUgwIrtouPBlULmnLw6JPHXoprje7U8WnbrtJ6Fh7TQ8W
HijobwcskC4jMVzlRKk+UZfZB1LagCElon0GO8w+IhFv+BJvQT1+ut1CqiUFxbs/
BWqVHAca7vDAbZfZCCDEqvXpprCQSmaS1fvqp87LXe2/HYGT2/BuFV0xzbdL3R8o
5oRjMhfEQP0OwTvC+gbdWogcCFds3MHdEUPG3+EvkVukLV4Fo1RJ0NVzWvedI9U8
fjQcb+A/aqypcugUomMV89Jj4QW2K1Hncv+BwiVC1qlb2/AxD8xUnNmebOw9UHTH
1Lp5LHVwjbKFYohkJij87zs5hgIkw2ztsIQTFfsEnuzOtU0FcEHOAqURDfNdLH3m
te8yfG67tSEPWKDwO5fcet6t0Xd9EiQUfu57DiKFd4X+8fDle6/wLL79EbucuCfs
GzzEgrf8vtipdFcSKjiVRH9rpUdq8nX41J/FN3rPvwMXYLm7PFPBUzzJV3PGLoiB
QrkzeYNowMycmvQTjLgbhiNthmBL1xx2C6Zc/dyUzAhDS5dtM3leWnBBXnZe6j07
98I5xeT1YqrPchnxnch6GWSGLNCbYu3RxdELjZbj5xiGVGB1EgEZyPIS+1IUU+07
oBUO6YM3HaIrIZQfB7cvpjx3s4zRfr83VPTJKOUzHUUHUVGcbJUehPNqkO9mKJfz
QMo5fkKX9E3X2gKz4lVQ7lAGkK8PGqnHrb8gUwTcJetcV6ZegAJkvndjkKh14AHY
y41kgvHwAGsu541Cu2XoWrby1Dlt7NiUU7JhbwLIzRMeqbn8k2lDilNltSbrys3e
6ClRdPR9MTr/YDXTVu5S4hzoGLmsz3WNDCjBE4Q3LVANy88nL5jLtmXOjI+/YFJk
fjnvQkZsqzjCyuHxPBM85Gzs1pz8sbEX0+GQyh14WaxAGP0Mv5ylzqxfWJXUMhv6
N4xwtCIFuDSE+2ATDqzGzd6iPTML4eZj2eRAKybIGNlm2E6s/TZMXhWNHmHpuviC
BUM02l6W5Iqp5SFO9V0PIvLS1uZHqtGU9oJCfQ+zTiwvCPjmhTFdIQGScMy/XhDb
iW87Rob2nBZ4+lNHKDGicmMZeGLQmLIuLhxBkIY7guLsV3JbsXOzAs1zNtNSau6b
PZgPMHzpsCSc2WXocKeLiVCXqaWcw4uF3qx3PSoFoWZQJoCcw6lD7DnbYIU/UjDn
OdFY1cVKTi8+fTryqh0Q/w/+IwRfmC+MnN9Kmzc/LXU50OjfxwyrA9f1EsxCTBBD
9T/epkmyAguTxji2uc63qz0GRkfK/mHqycXAsMBsSOmmkYOCW02Mzekxkq8eo2ae
oeHlNm+QOtAh3FVGaI3U69lB/pGjXF2riKPeizlCyMvFueffYdR2TWKjsDSsB5C1
YD1XCfL9Xy2RYYbg5E6BJ9F3M+QIkl/uM4/LWVbpv1yKfLpqqS6ofsx7b/KjZwBH
27yNRXPif18/V7o63j2g4RshzV2MBIFs5wZEXHACaI3+BhTvAyYBcMb4RnvM1n0Q
mbO0seInpBrCc7Vrz2Uf3yZluczI60UpR1TO05ug2uGOxxGOGrzu/j7lpmLJgQln
uWxwR+pt3H4fXCZhCz4TjjfOWLZAWQWSk/q9m+z1bhKczGSRz9fVtfwmwV1eywJU
ygrptv9zE1nV/E9HabMjkGtQyXX8R64LvjIKLIHOd5k6D4kjWdbYf/BRI056xDQ6
82UAaRAZUB3Gx8CdScQHduxg0Q95JnmDqbN2o7bnhCfpOEShpJFlJPXQF3TTjWQc
a3l7sKZWldnXbL3zr+pd+J1lXbentR8noSI8g4d3ADXeVjVhlHFinqeFCVSkQvjS
0d+EyGplA1LH8l18RrZtDHM9mUBlMxeB0Ay0m4UHxJA2y9ObvBSBPxk2ER/HXcE3
W+CTlxOEE8alSoA/abEyDHunRWgXJe0KTieWRTbJgawTSdLuYIlN2yKduVBou8Qm
5vlkDiPn4L47900V1YX2B1hwQ9ciq2Qiv6Fv0Zc4I3hOfdRFwUnr0Ecu4YA0VGGJ
ihRNX6xEoXY+3E3paKmTKayFeMYdriGdO8znU/K8o7zpK6+yISjyXnr+RmY8Z2jJ
MCpH+gI64LA8NiKm5nHAOKNP+XC3twR53tVQtfivc3NQH6Mhzsh/h7ZYXlheby1o
BSk39ayQ4fLnL8xtYrvFYnEUM1LcBM0jaw0mMhrVgzhmzZHow34VbwKc8hJ3VfXU
xDmqtx914QSmlymxwTsb+2REYx3KLbGLP3GkI6Bi8vWP8uxiE/5p4U2DuEJWY5mS
eb/Oy9MbmWvm99z7FnupKDfUiywpFiRMHqZkNx65vVQSUPls19JuCXjcNzXmYXuC
IMHegFuxN5LJXDKRn3HTdUIRu/TG6FtpEeeEWpSiCyGYHCsWIPIY1U8Vdm6qTXzn
GxkJE0fiJjwYOQIqDHB1c+ZynE0yff1ibv/gbmdq43LnkITZ+g3oeDU/Kp6CndCF
FcUIBsxkp1EnJX52+uwgHHSFoDcgkUKc0qKfvXZEslmjHlpETSuNl01u44LIPbd+
6tMCEOXNZQQieG4VxrmKUDKEzDyBEN601gOwFLCHV53jRU4xtK8ZI1mqtn+tsow/
Fr6lr3Ob278sjyyMOTmNODKdqFMvkv12RKwz/ZPaiZE9WkyRK6JCTQaHW41j1JXY
rF3/J+QG9C+RKDFe+awELSXd5IDhtrb86E1v2NAIyxPAdh3qzR3TWRvoRELnL+DB
StFVc5gxahvbzQC7jAWF/9rFceu19GLczbajm1bqb4Rqjb6upjlat2besihadM9a
1qutYjvS/GPh5HdZtsHt6sipNozNwg7PCy8fh6l80hEi0toUE7QWoBdmaRJTk3lO
XONCxejsq0pbYgYKGR7/oPGtvpOZBfbaVGQJ4+szyY1Ag/9DiuZ70ZTROysLq1ZI
qRZgBciFydYeyG0AYmW7NJyRdbnYHVkO5H/diAauIyukX+H923SnUORRVR+OZyeF
4WkA9IIH23JWgo19gAsy5soECCZo72nnRQlD07LRcqlcvv+rx7i8oGx3e2kuXGnA
hQyVgUhNWo0EjB6Q+zVO0keuM/5EMZ2BtmddrSHy3hpnAbzBpbVURY+QOFDFzCJ9
eACt+UPSvHrlEL26Iil6RqaFWtewn28MJwvIDAEhKXDGrTkK7xSDhpNBqbkV4IRV
OuiF0u2jXqx1ZbdQxaO26aARzxpNLq11obmx+KFGOcjpPYDQVrVxjR0tv+6NyDsw
gLsNMi5gMQy+6mg0x0CYnMnagheUifBIIqAN8pxFwzniFViR+maKrULZ/SNdI0lz
z22fjJv+rWhgPHppvWcmw0zul6TH4QW5CzswU6vlasZmiCqSLxAy5i4qEGFrP6d3
19TbCkmufgj0RuggEhASJlgmZ0Ln+bhWkJXhpozj6hN/HQgGsgvoj+vKin7AU+XU
jcJ0rPAOf8Pc6/iOIXxDmf79YACpPBr30ChreuWi3VZT4E5WzBOwSnObrbrPMOEQ
ul+43/8R2ybdkWBgmqRBGZQIV+px+DwpRCqHLvAPLaz1rmfT1Wvs5hl9sULSzRBt
dhHY3UPX20TlWsl7Kq29dbKscGKtHyEph/yOT4XpfFdDWMAb4zpFEl6aL0Ev54yW
RV+P8p7yB8gdFdS/EZAzYXo9YqqpdfgXe9G7KxvEVdNdeQ0cF23Mzr+/TQEywDPY
8dqZMM1O9xSnvIcHT43BVPzOOQD9DTIltfheOcPHc0Af8SOgHadd5Zqr8DZ15RQ2
vIOjohcQprkoOzQIQ8KnGgXw605+Mmkl19IvP/sW7aBc+YstTTYIVH1RPbJIDm6N
EVwrHJwldaW1s28RnqJrFnlWgrv/t2mR7YPc4s6HxPFCYYGXx2wEauPuzv5Ivhs2
2Dwlj1SNH3Lp3QXkG2Zbh6lPKy6g2hJscYgNQTds3rXJ0eabsC1ItA6WmLFBB5TB
bXDgYUGTIQmWGJwIv36nY3Oo5RU0oPWTFDwQGMW0/tL6jEB28N7AVjaBlzkg58mQ
Y4EGMl3nO7evouf8lyj47BdIon/uCJANYKdMlw15qsAfjT7EUg402e7vyddx8L2p
mpNwB/EaWYRt++wmiVG87KRVu3ySHl4Jx+byUoMZUKSV9PkDjZXXnh+rY+HSoip5
aYRtwv3Qnzk8GeDGgjRMrfImyxYQCHk5xd5DT8fD93O241w0/Hsa31snzd1EAn8q
OAwhTkr+nKw7PbW3K53762oQdRO/K/uBOYNCDQGg3y7IZLWRzbzAV4N3fW4W/tcv
IcqsxyKX13NdMyKdXj4Eujwj8UBfxFgdHzeXRksqafjH/kwZBtrcfG8Bz3DZEnAN
LZxb9K/kLjCBkGiXD+Gy678+OgxNZuH1Ogiac5Y62qINmPKFhdcUzdOJgtFYV++L
gMgMv3RYjhV5QbcVBShtbGXkE1iDxMRCG1MmHZ29yjBwLALmBcnB2DcZ/U5SMEkx
G3Y1xJ+Bb/1ch77MW8QH02an+tcShujyDnY19LVn8r61aQ0nWQ+U3fd2FjrUKjoy
sFXIC2AF40J1qpHstXajkuPLsfuVoOylgFr1KVYo5/in6ZeBUSAVFSm2ihoSD2G9
/7L4KXrMc+uGd62evf362nFLVKCPRi53YJzHENH/nxqaN61Ks1RvZ4X/09H4tLGV
Im6tnhvy5NvCHPn7rdny9GgEwhO8bucIh9T6ziADKA/E0/PBfySr03i5HeYDBaOG
V1g3ED2lDf5JgP+mFJOcIu6k976XoT/zbI8D/sHWZ7YoGytcOOKu/EW6ChMFvAOO
SOEOUOPxKZoYMYUnhqC4pertt66DCBpQ1DU62JfQxRPKaw3Ol6hAVP/5i1oJ0Iwd
Kq9yQ8sVAIckj+tUreWSvPxDkcnNEkMrymT61Jh5rxTLhfj/cYhvHZOeAVxGUfVB
5FsMuTDr81sSAeogEWIy1YIO1RjBRdJ0Ol4Rk3FUiA2qAYs5OjsH4CzLBxWy14VS
tvn0OBnk8do7niWUICxs1TscLurcjDusqGsG0W5/WhPPhIea7a/bnBQS1TKwxb+c
ECZiqjGblp9xsZoa57h7JIHGHrsmuDFROVFI1U9oxMwgORqH7x+qnileWJ7yhOdx
Nk3/AxN3F34GeMrjnSiFmCwwkBKYgORnFEgdtv9VEOdP0cnCtzUHEuXNtGxAza64
DdV8fkl2EdHZDg7XU+AznyD7IS90Nm0B3LcqNXdkxHBY6qJwNF3PJG2zafrGUD9S
RXch1ooBS6PFArGaj09GuXDeB0ucb5rHBjaVO/zVD5Wxr8CLbMCzeqQws+rzojs4
T3cuH/BdYA3cNGFU47AEc1n7LHXGzdQosgwWlUz4Vgwfz6qkH+7yERkSZGtm81/w
ngClczL2SjKaPihV7V5a7wfxLv7xwL9I0KMl++lrTEsQRhnv2dx5tbvqhUZijCsu
7cVm6+KUvX4/ln2grsuUvYTwy9wwI/gwGJalbjjtwg4wClp3jU1mz+JH0pFd2y0J
vxMtbKnVwoCZGWagSa83KCSQZ7G4FMXOtO1hlcSN96RxaNQezlJnet2h0DJ3Xo8r
AdD6X7PPrF5cnXb/QPgs5DSuym2B02XqDJnan8HDPdtJojCebRkWxRrDo0TY90vK
2H1UCrtEwAYJVETYdewxDU0BFlss5zxv3nlYIpHYnBGOT4PpD4a+QOqlMzDN0oXV
bLSQIkaURRY+8dp8ImbJ1j1hgOFxW73O5ciR+w0LW+TBBpUWfC/2A29CWopDOsGJ
xgDHCeNzEdpONzYkwgNmY7+P4HbVy447tjZHwgJ3x+ZpBQ7HJhBIdOEDJImXFzuZ
/OG+MW1EZIYauepFZpNKXpkz58/8gLNFNzlcMoDzNzzyKHP+W9DHnWUFAlqAbFRr
d1HeghEgwXO7aIXuHidx2b9X4m2d4Od7J2HbSnI3IHB3lXYr5o2ZyrUSkie4rOp8
xRuJU4pSArvBsRITQTZXSIMqjP+jTOyplcG7+CtA31Nx7RN6KQMBXLvRNwZ/F4AG
fdTey3DXy8jGGBeMX+jzIEMoJzPOhN7rZfRfchtmg+dkvwc5uILY6bhyphEUNE9a
1Bhkij6fTur6+7WG/1lOk6j2e2tGpgUF7OqFf+qJdhLjh1VGVSGTjGTyu8hAtrIl
xSfJqxCt/K33yTXMJFm3H/1y0za7JuxfDGp+CzpIINGMDJbuomdt8IPHQAdXeAh8
mQ6kv+F7k0g7H/GGAM5iJhyCzEfPsdxrGbY0MQxHyeQeDurwrRz1FlROmHmVyLYA
eY0yFYEuWpX/p2yqDdh7Dj5tviiGjalLTiwM/NVXjQEqjqmmCHOP2cuQXarHeaIX
AZkske4Din9R5PZKSZHk4W1hJ3Hla1dMbsHLgHCBUgxmvLhLrbYSgKjh9mRoA6iQ
G4TX/bWlnxdSCB/SEfSwqWK+UAcpv2Esc887+Ff8lM9GwAWNB+K/HNKIStFG02/L
5AimW3xrAhxU35WIoPCMdp6QdBY4dC4eVpz0EW1VmcgDjpIrAed+peYkkATh0h/c
oblukfm5XksdXajd51JIcZJbURN1tV1kJaC3imsWdoQ8p+ItvcRiKp6d8t49Juts
JdxT197oj+rZpWtkYvg8htUk/f1wWCVZbNw7GR2taOWNxgQln7o0l+2jaUOKVdE6
WJKH1asOfK0pKaDafnWm/cyyZkFJnS2KKKKpPcxhtspoKJpkHxiCr7+Mv0A2g4P6
Zh3/Plro7FOKpp6tBCbQYGXVnV40JMKwIQq7RQqHeW17NC1VHJScmys6XGbzxEkO
Y/5w+UHzb/Wpaw2C03P8Q4ThAw6sofaxyD0w62ULSlMUu/IfHlWa+OYnrlEKloqJ
iHq38NSmZC4IzYIMYAxFH7xj+EMGJrDNFQszMeSdR/bwHDRWLzdnBEdg8HC2GhSN
T+D0sMGxjAthqKi+V4wjC8UfsxbwAa81jHwEdfIlw3UNuZWwOVp70VKdLIYey+uN
6YaPbUe2P6XBQIxr/9iByipcqud8FjoVMRGg+RYVcS7CUzJNWE4mPfZWsFWIgXed
fAZE8bDTBg6ElD1+90g6Xr6hYRaTLW7QdjOsbib/9DOXCrfcCE5voHsr+RmnfTqB
EaO+mIp7KIjk/AcGcYFMlOUKMjyIGT0eoCO17fsjALFBsJhvahMpT1GeDpyQgwQS
Bs70fnak1CQuK2MNUtq1w95k6aXjOaPWEX3i1ncqrTf9mhVv+VUsfXKWj+T2Fi7A
0FA+jv3+IXSYAqSo+03psg6OyGZbANnzHT/lScZsqNA7YoIR+nhM7V05SSgU/86I
CgW3NoF7rQKemd3RqMNDL5F97T0n4i0csYLDKYP/iSyhyMSCu8DscVC+KvrwOcua
nTsMZe/RhTomsa/c88zpBm9aWdJ69QOxhAN5j5N4/O4YbG88UTt4XYzd098tfTsB
jEaM92QygW4h+FLbMgLNeyDsxE1EnnTnrxABE87P5gDReFJAdF2l/GMkUmWGcJPr
+LZlDE2GawOrr3ovmiZXm9625Bj6zbh/kWqjdXoLvUAMgEdFCsZCWGe3EP+PdnCW
5W8Gc8YoIGIIKz6ulyq9nO9ZiiX3q7oirnjybTaoJK1uvO6OPH/P8LzpMTbOVvCj
b0WkuZmlKqLy0mX+nTlMDjiIkKNrcLnFVanIy5G44e2IyM8tH+jdFJa4l/7UCtRI
ZChvZ1VuofUfSK0YWkGzYOBUFLNa6Se2qkP56G/qyjjWjdB/O952x82y5X6YzmTo
2g+kR18t/rHdDhZ2LpIKPd1WT7D7RPlNbhacYXhnWQr2LzB9EAYGWaQaENIwW5Pt
TkkuZZbXbL++0m4mDD7VA+ZShLTXtnEWIYyM8tJFGNY8tO777TcTPq+Ki+TG0vo3
NPM0N5yQ7I/jkpevOdU1CgbZTWWnOxh2GhPPH7YUPDW2ZYnYOsh7xbA3JhKU6Pd4
tUwWiN/mf6/WiDfSmuhS1rgdEPjKyLNrIlDPX2OZVtUYatWux29eacVbvD5Fdz8f
0OHZaj83qeSRHydIXYiuXeTBUPPhAmUx4t9zqZhrWwvC87pHxEr3taDWwFnO86/x
qX4Y9JsnlUshaW+6evbNTm6qM415wgbPDCHV+3/BOgrO2EY9XKJnA0SeoVrq6elp
NoU4xP+NoM2LzkYQ8SwaImEW+CzrPk3J2/Nnqm8M5L9chHk6H90EeLcsnWSjchsz
X3MGTt7crV1vAI6KdDR7+RZccuKgWpYQ0ycsnK2syn2Wip8j3GSXIjU3HbPlU0FN
GHkoeDlMQKH2zFpzlfqdPryDqG9sEANMRVPQsyDRGAydqEj7U/xecJzhB/6Rbfza
VNygX/+Zcr9Vm6bY6sVvA8e039a2FvAArk0w8m4x6GmGZXR2NYhR2JJFmh+Zw7WK
31mTGdt91YD8sBko/++m2jyBQyvCEK2S9QNwBxHH3uDE1tkajMyYrKFmffx+gssp
Q4W2V3EA5pP1zJ4UTT9TkyAP+etFXkii7q23xz69CjfwgIreXPnaSzKvy4V9ZTDe
BGJs531ecrT5Vtzck1T7/3rSM4k3S3tEq3aNn8NDyiyPHO1XXioqD/2EBjsnW/Iv
P3BmDxs3L88NwMp6bIDpEcYVeKuqJydsMOvRv2R6XkMsbTgKRd9BwD4tfr7KatiL
drYBa+PWFtSBLxZ5MWPd5ZA+vGPyHlvXwSBxg/46M8jC16Bv6Rkef+tQfdkurQG/
SdHg4+AFwVThlnF5nEX0hl//4xUGzcew5epEzb7AEhLkDqNRvkb0kAqkiuT6Ah05
PeOB5SkWjlPY8sznL7yWfF4PEo4LovGGnTGcHbvu7/T9gYKslffKdo1GynEmn7Zo
BgaNh8KXG8kHnzhCBQCGoHoICl0lEaI7pgUvLLnt1GlB4YtKNDQdaNKSyobWaJ0L
Pg241cV8nnGJDhfSy/0wFvWRiTYaPNQWsAzMRYR5pZo6h2+A84s/GDX8yF/JcvbY
jn7TvijjqgueDeAsqaE9NGC+1fkXfnbpxYtaHBwwcZNQJP03cDeatwGHJPw5HUmZ
iNJwn2l5AY+vsn5t+8MCFMv+9dT4OQdYo+UVduVPl6L5655nWRJUa1+s4Xhlo25M
zik5BqILlwL+CPzy+Y0A5nGWfEkhgKFGNvJV3jXC3X9OW7DyTybUnqspSeElqblD
OxbOZCfepDyPmek5ruHVCMnawYwwHaFdepRfXJGBLiRMPPUr1ABNGY4HBSpXoVtI
a3Mvuapzbnq5kSQRCCk/LALoUgGzGdnHj11//VVuo4DJkpwylR8fmAlTy7Ib/dWf
vpbkgI0AXfe9sKv9k1MwtwCcnRDemM48RNTVHBVmZy+QYSanq35FGOINItm8lJC2
RuWVdInUTxMCg+DRF09YIMgBcntVtfP9nzdcZ9rl1E4BquVbH0MC40o2ZTob8dn2
nb8hJU71FNeBcqPoGumO8v8hK0W/y7tgKaDOfutNcnf2qou/wUS9Ys9/4ordJOWp
LYKjEzm96NBuahqGv7f809SXPiGTl94qYAlMo7MmlW1ckkGmL4GcCuqYGYP1N3ct
aHD5LCIb08tqmAnACQCCWvL0MFhdaoygM+zUho/iUDUQDadEdvohTUBmdwC6KU2u
6KmKYvflij0gQW6g4Mnv2kFEjbgFHRloPxCxKpH3wMuicO2Tyvw9Xln9yrJztFEt
avUWZUXf4J+z/osvvJPzevnSvIr05BfcXlQymuwnWtp6KtDR1BcMLf0KR1eN0Npa
JUJZAnr7f08CRlQsPCfa6kNdCwy48VU9ewurmctjcGmavGwm9ZAZVOlG7SDFB8cV
hVlgm4P+zcQipCijvCF2PrL+2y0P8ds464uz4k4k5cOSzmWDoEIGQOdQb8IDtBkO
Vlmd5+WJwKpo4zh8TFd02LgWV1Vb594l3JXPd+VyZWF6/kKQR85AaJlC9ntsryfP
cXFavjkhyLq1yh7T0/g7RUCwauydIradTuhute6wlx1dddvXCyArS4G+4sMELczA
thE0OUU6d6VzfWkbls3DZwj+Dxsrnf769Tzk9HyC0RAzBa25ZELoxV0EqFtHmkMP
pm3nYjjL4HItXXJcbUlbYE/fQ/paYhAF0wDAtBJmvUA3/nGWkprjR239102805Jb
X5KAYyo9bjz/M4oEDZbf9xfFNuHfKfHMmqqf0yAlO/29OMgtod04hVoJUr1LPQZK
bpcR/4Y8nZ3soqjGzVeLx5ybjNuJhiuVJE+MhxS1vhbC9tGj6j1Ae+4M5HTri47n
ajpHzhZfeHwQobXwgqx03aiIKwBwtFDviaS7mZaRBbDaPEAIbWy8VI4sTEAUWVjM
tMF+4/7aAbuDSFPTZLJ2iYIbeOSH9hIlFnYqyrfy7ZqWr9PtUO7XkxCeDraE+kLJ
CnNKxxfGr1Rio1Wzpqfo7eeLtwz4AFsvt6uUKFpTw9etXeDuLbzuZH7sYFgNcPTU
lIpFUWCQemsRPs/IXEOmbdAbHy61fg9BJR33YqOsyFcrGzg2r7dZh8QkFqS3Lg0D
qsHAO4qNqRB2CqjNrWMLRsPxmmv13r0EBDT6e4sa3/iksvjadNn3gnhRwkUr6gcr
zyvjpdVWxiUfNPnN+q8TI7aup4o5FEZiaY6S5EjXWSJ03HOUrgRkj1PXqbmu7pUz
G8ZkRYZKIoLAd2dW2IzEysbZjmrWvXupA4oUaJrVwWK7QU6bVnMD6+9XuHKvVwKf
dVxEPJXR55UpoR8UWqmjcQ2tU5EZYhqK3/RGTDuuAAvXSLNnwPvU+FCwYJdg/nUo
FXKpLTNPM2AuX60YI6F/LLqiUVCoam3aKyC67yMLKRFS1oZCeGLV+oSr4YBHiUPx
rXMYaq2bAAYDOgM5N2Ec/Y82FQVIaU/i21czzf/7+Xy2pZOa4W4qO7678i1kG0Gy
dHQtsI24L5fOEL3OTNvfpQc6l1RusaOtugfnHQExDC3/479UtUcpJUHgNvoNbTuj
8VCYCwjA4QngkQaRmPhYsJ9c7pDtNEENcS5jrTpBiw4ZQs40iAbWzStFeVjfB/QS
iZWYK2DP6j4PvZ4ZB9bcKjoO84/GooVM+CQsmSqf8tqcJCLMNf2mjP1QB/EcXSOz
9DhZxMUbQhrgRSMyBa/PbehX+UOW40P4zqK8nlK2IL7DvMKdxFSS612iElWj/iJO
QrZ7EoTjp+bD7rhvI7S2DkQ3ktvtoWicq8ZLA5xX2lqR/CAOE6k1spZzO87sjijb
2Uo16JwVb9/ijgwOqQ8HTvUzrGeJ4LxYgWiSmTMQM4sf10B+6yfbrrRzaWJq0CmP
1xVnmq/1GPANPX8T3aZxBKQiKTQa4tbqLSAgE9zPR/Nh5PR9zci2YlSn7BdFUmX3
u7mJlHxQJkUmPmC4ed700oki3pae1BgCuc/I3m7EOMYSrJjpZJESkP989bvIpVnP
ldvI72zfrZvfYoMA4CUwkex2b758+czisXfJUuh5AI6gKKACSIXJi5QCFErbP2d+
uNCyVDOCxBihlclNDcsmJmsQapTC2hCsNV5kbKhraQJQ6TsIsdpcoFK9lRaMnT0A
NxX4EdbDvgYPyZBWzFttx2K9tcNryjr97DY7Rt1fEFluA8eROV9uS9N8zrVPlNr/
yDT2w2eoFLtSY+Llm824ZACd9bF45HlE/IuqaJhQV3BXA5FaZ42agxEBGcYwrRmI
IxLM42I8o+Nn0UBkvBY37dbJyoHzbbcEDf8zImhJCdVCRamp7vhiFRVTMu/jzKZL
l/f68sQDqJQIsXFDQ/RcMQFPQQUA7pTwS09EeXGX28r5JuNDgEGv89m0p979cpKd
OCRHjtiyULADOFp+agdC2QmDNhlt7REg/EuAMmUnu6UDjBZNo+A4aLmQVFbC/ZSV
JiGZLuntE48H117XqA3k7vyhlMglwEc3RhEK2VmssOkHzMa43cZfgNBOnHsbs9/M
vnV29B8Q0YIOAp0iDpvlSAFI3vCVdUzhDnd1HDlKCHseBuaugs6rUq6A+OJ7ECCs
fsmerW1V9APbbdfa8U/UMnZis68xixiCQdZsN+dcoOoKJhkegDj48ywkugSG+gtc
6jtMCU/NsaGLGW3hSM/EMIMu585Sd7BerzfGxlKSrNk8itUwwzfdHkpW0hIiWnLE
jq+DhUlT43UNZRDPp8e3BDDIAZTLxgVvoiruzX9f1yyMm80f5KJuEUEVdZ7Gkf/j
1WlFWSSdD/gX/Swf+C+tixarqbKrsFr37Skxwtipm/YlgJvE3kiwlbdLxIPj/Pyz
0a4CgTUgyGirH2cLhivNA3oKUCntkBiyPtxOK6VaiYMKPsV1MXs0y/FcUFXWPjyH
++HdbDFrCDvAk8jcC3noRLR0elEhU5gbAnx937gJA26bRTuivM5qNN0EMtqg34MT
bwRXAbY9yEjeZjwoMi7JJ6eCnmPYu2Tt8MiALewkyZeBjnfJLOqk8OVQSLdepcgx
ACMvf8kS/0GLqIr0cgIEjlhQl39+q42JA3jRfLk7N6blybP3U+jfZ/tPeihCEFeq
o/i0LPyO5+LWUfgeFJQi0s4+HBSrGzSoDt5uGNTArZ8lCTkhxu+SnMhfzvmPRrh6
/yfb/SefhMbdM+IEpUXdIoliXIcCZRDAPtcH54dVwB8/PdbMV3LdhHs0VVwuD0md
m7HPoRfIOhlTnciZQ14B5qZIY7ej5HqjK6RRSNpIwYdFpSoK1L3J2QbSqe/4utnK
KebJOY4v3jq3yRAm8yEC6JQ/bXJIkndv4n8rcID3Dnj7wgk2DZ2F5JYaasJqmO1/
G94wjvLwGGBrugDe7fY22Amc9MMgZ/dOdVY8EDhaTZquVBBwsDuR9oqpa2dn15eR
oHXXGQ5DmZ3/Z1rKMZPKOibYxxubO0aTxTUC3zhRocSgKL1K0xzMmchUiSXxMbNp
R+APs2E3CZgmtIlNGMDV/sFoZPxS5eARgzvdjzP9xRJggDWn2pj36bZSqUbm6krZ
L9lkX/PsUj4th3fHS/xYg6ss4uF9A+7fsTvttgauV3/nldoWglCglMUETLfLCqBI
HkoOR+Dbz+7OBaGpG5lVshoegrU6qQYXUTK4Ww0+DO6EAibH6zPJGFG0VQssJ6q1
NASHYjJlrzrBSGe+ySnplg3Czp+c8bbsRADDt1fBiJF62UYk7v3xbx0SEmAaRxI3
hNCF8kkJhmD3esjRnWNh0kxKfPKqOdP5VnJHgR2Ix9dObXw1HrU0kktoqHWnjshR
lukdz0VZzhtJESE+70cu6TOjqXgtCtfG3AeHUwq6WEq1RTxMwCSnEW5KxLFd7JJC
d+C6etrmHMBGXX8eAb8tnBzb3xmJiKJTDREq9LDGY9AzXw6teKYQFT1sBDBGwY3A
FZP7AWUk6yGHaO126LLp6/9zqCI+9ZRtzS7AASEhidSMN4V1oxv0amroC97QMnyP
9MoRbt4UOcdcJ24nDtoYJZIhMOM72vhqYBAmE9xasAzUBQcfMa91/nFcATbzDpxF
DfjJLDLXPR+uRWVDKW5PcoIYxj1hOG4KyfysLi7pHeJC+eP2lL0oBpY3nndp2e4E
wptZ0fqOPfduLJx+rcn7eaRXWUHAlrFyOuZ+6bPoWtlO8ap57Se+IWs9p56i4tTQ
dYBpCf4dMfIyOKEaB4CPbNc+AVBg8/5lRm10fRbNsduMm13cmv096iq5oxLXK8+5
eTidJz9aW1VpyPmBs6Ai8epSewfI/cx85l/rdxBGn9W79fk3nmP9n+nwLJ7H3tMO
cDS+rN7sYBjQzZ0WEoTwQh3txuxaKJNOMky4NUyNcweBo9OBWgAZCoHou8EsPm0+
szN8/FFbavJJWQy+ApqSG6VzvcycReHBnWRw8fHIKIRy1uckIfS1nzqYRkNGmnPC
9XrFG8gUEHd4a3Yc3Z5ku5QaRaWObzDma9cZtIdglGxjgkuiBut8VHdGLX8vW6zh
TFj+uTPhxT0yQoCXMV2dO1ZbDx0uX2cEp1XgcL65Fh8aMP9yPFNT0QKlFwABAK6h
SMm2H94ZssCbKmwp3Ip48SiqjQ9KpLncLlEE3TK2E8oeoXfFtSZkHNc/Z+2EYl/s
gPycGsKyW/0vq2mHvfTd4CtiHvxkdYSHbdlTSeQBbvZvRpvGuBKDdetrV+dA3KRV
yzQoGkkdHb+aOqZU1ol0XPRXRqVdvgNYfWAM141KQi6j6Lw1zQcE/N3dIUVfvKwA
tj6FKKgQ8FWI6/8RFofLniExdH9ZIvL+XlbnqKCfNyc5ohi2NJrzTZsDrLpI5fTM
ip/XFOdHQ4rxi6fE5Hk91bu8xgd61jgPx/sglMP+9uKX5nOV42kNF/WN7vs6uF8x
3e/m5b5CKN/SD9BKomY3AUIjt6ljL0RQ6GbFLr+H+Q/Nwg6rj089CQLwotUbFmWu
k6ykYWUm+4jGnD6AlOjsV59AsGlEXMX7aAE95qwD1AoGgRuWhawZ4+43ebOYPILr
NYdbZpkD3P1SirOo4plfzw2v0y8qO8l1ipw16uTcduEoYtI3zPOJTjQofT9kTyHi
i9ZucVWDGN31YyR2snX4pOWJh49G/FOZVBO4n2ziZCPQ3HVhEddM0WO6wM6uqYqD
A749R+C7cbkYrw5ipgYWVjOO1L2wgI6m3LylQp0UeI2AXc6HgommKonlNoyLy6JN
cITQiFJ3jq+lEH2MmULNd1rCZUv5qyXDVdrSudhw9EcAuwgfQaEgKBNLOeYiHJFa
H+rDwDnoN4TAPKfRSH9EMucZgcNg18EFpesmWT/Sv970XItaMROQ5Otk/sxWnXe3
tWOD4mdWJFMFdrWrNniCEm+yzcbFTElkz7SOvQtrNX7PVeGiHKFINxHrKlrTqHkd
cEI9G7OOQj9Ivsk/SJ/83/PGYkrp+IoVgQ3Hyhnkqv7s315TlQfKZWZoAOJLY+6K
6raZa3Qo5x1lsRW3InUPSfym9hOCQb//PjZO/xRMdEsmlUuFg75sd2tdJW0zMyC8
SH6Sind6Yo8ebdIrpkzIdejAGE5e1SdIFU/qpK7Oa1ik9Sw95jCATjRMFhohfraa
2ANkJXeZMdaMEO9Z2da8nsaRra4iUWiNTL4dbF3L3dBgqI1M0oycwNRul1RZ0dth
6Z540tuSYQE8hwskTTsOm3erVhu6GCqqckzofhIoNnj5b4FgrjCSUnrMsHCFyuHb
uWiJ5UejFBiPs4GhDxMSwDioCfWicxs4Gd0IH8w1neJXOp7RGqkWF3bKazdcpv45
tdLVoylzuj2QVBI8uPozOqXWfeloP+pH22k8HAjZF0zeJageaX7ABmJz80SjqVQ3
pox3gU43eJaRGhJDIBRtoC++g75sUp+JPvs5+NmGciNm/+N+hXMsGQ4OEH8vq8cP
zIkOK7FIm0AFTdpsFZftW+JcOugEBY1JneFv8STZOGK16Z82tJPVjDk/3yrSZ7Hf
JOLbyvn/lbLE6BsGF1mjBWSS6bgLRRPgSuG1cboIr1zDqWhTeO4pPnuVDwXHc0g9
hxmcDLzg54PetXntmu1A87SAIi81mUFYAuzvU4w4dxEV1BDSw3FXEKpxRgr1eDNJ
HEi+6gxTlFYA081gkdx3uYKoUhxga/SrVgR4yxxm7NiETfYJ2hsF15kzNBaSJgPW
FjqNoVFjYvmpTY2+67YMqwDmEyGVtI7x1brbtGPRN/QOCt7r2ZVoNXT6Cg/bPRDZ
MODAkURIvLCOW/lM5ovEhL+nTHkPD9cDw6g2DCkZC/lx4GC59YZcXaiHtIQbceeC
TFQ3CQfIuhQED9lsoBtKWMH8kNeWLJo8iP8NENmIr8Pl7B+bSd76nG2xtAgsGkZp
bwvn5/jzpHh9bDG+UdyaJoFp4o6oFRKpwRN25zVbwsmNtggajMSPK874QhrkA4/7
CKUOywYL5yKT27MNEarriwHCVGCqdnEQqI3PtEt022HQMSqYkJ/KsxrPpwfTJC0U
hEXutzCcPKiM0VvHxDX0DGaNUlbucT9QwXlrbD4J9QK6Dy8JNrznVXUsJCGcr+b3
R/SghdbkIkciQ4ejnkda4imFLYVcS6wU/7K4HGdOTXObgckToszpA+DW3BfLGNvf
YQD1Wd949jGMf9X0C5rW+AnKeymwLJVqfYle+Ag8eFausaNWstrUSyqmgpRKG19Z
p99mKW+ZOvowJTHBIiralYRjwTAPTDMiRHumqTCSIg/bvkmTPUe8lzhs5sIxAk1f
qP9IDWGtOug483DREQqifO6cJLmQPS7Gpe3Lm4f0K5kIkMcfhyacUsCVeQMVGisM
udvePgM16FHhmHLORaJTwYQdUckpMjRGqO3es9qVYNyE9jghHgKK1sEd9MiQsA5Q
UDB3/324MGIED6rN2ocBwSy9hmOpEhw5eUu9zLOATdS2brozjKqh9lbwGXtJEnlG
yjMJYevVof7kP81tt7+iKpsHIdOHHIeJbOWgxutgvLJEgTrsFVw99gpisDUCNS9S
DXDEN0iDvmapgL4kLcrY0czyWSKnj8RsQRa/rfWdWG4+bu8QFGXpMjvoPxuLBgyI
M8g877Hf2T+reiZWl7GD0FRdTVdKPvpq0jRvMqUZTGe30AC2ykdXjQSy0bUVW+Zz
A5URN1fmYNfLW44hAuZ2Y1nFaJ1dLwx2b26SFg8bDlieOxyoa8sVERz4f7/hocq6
qQWYq8ypiclUTYvpDFFVW5tev82p89uDktxlyvS5mCFwIJtowK8U+xAYBOM2onxe
Wl03gOxhQ3IfUq5RsOpRtYtXzRg11au7gyxfT0Z58ZqffFSaR1qEW0c0Zl0XE/DN
VBYZpRkqUAY5Uo2FkdRDXX+TffedTkIPZwqWh6JSy+kPAK6XaS5zB0nB+E0lPRXE
KodI5dZVVaGHxavZ5r+nNPM98gKSEl28hrA4oHWR5Uw1qhaX88NH3dGPFOZ/a5Ot
04oCV0+jUZBK+0Ky7+/lqWh5E0R/FZ2Bxjy7e3aLcOKtV112eepaYeEkNmN1Nva+
Dy6w7ARq+Htk2G6PsRwJYFPSj7+AUqLnCy7DTa2VjB51VRHk27lvvZ9VYJ5X+asC
QCxDyU32nDlnuG90dvJlzPlt9oAkrNhas6ObUgznELIeQWXjNCuzOnudSADZdEj9
QEBvYaYNsTuxbL7yq4KBvFxF72n6MnxJq7pm6kE659ErBlHG7DSiAo1xsOSrPyxk
a5Y0FV8j72BBXNpPngUX0cP5XrfqLd+RrPQ2tFnvuWTDy6bN9BMc1FZ1mq0hriBx
fWUKixdlj66/+4lmrp9TJ6hZHw78E/oqNGGkGRt91QlkbQtumlhQ9ZnCtMWl2ou6
gS/rh+jhghKVtU4QT9dqdEhXZkqaVDcexKEfJN0aGS/oYNzxBS7TT4uz4TjwX/1I
O/t8tE9azASDiWYOOWIoXVSIMaDGoilxA0wjNqMuzREHVeNAFXusEd46BWlOtDA1
lBuQ18bbwwqnENCd9e2mcHOJG51NWzh7KprJqMzm/hUouxro88w79dpbHRup7aJZ
R2UoThIk7Hg8dEGJTb1YHDqId3lo54BmEFukU3SZ931ADfPfF+TEQx+8zjnhYKWc
iJyQodlf+m4YEE7oeS4POsZluv4TNr/xqQEXZhU2G64ljm9/I9JsmuIApd1HaOTz
t9z9hbcXL/f9uWuhNbMF0ms0rk3U0KtL01K7j8evyVp1TQGqDtCpX9tBCcEO6YEq
3waYjZ+EKDa9e0/QDaCB8ecRre3f8GrDP5VYFG/WY2rwJwzA2LvXYYjqohOynRO+
tCKKvfgvGPdyfe7d3VQdHjTnmm0UI6i6j+zP3BAMCK2Z7T+8lE/Dw94jNLYW2DWq
O/UYQdUeVrh4pNxGqy3vPTcF8OHTese8EsG+NCesbg7/HAKDTUVys1O1sdMhXooI
XD0vKVsEk86+O/vfe0F9352uyxpfHtz2lq8EoapmhLgXduLg0l8kKRceeqCaLMG2
x/k6gyFMaO7aCRHjWIX8tgd8lkO2l0H6oGH/Yc+wRQirtDf9rjfMe6xvf/afjmzh
ih7zK9skZ1jITRpfF5gtPhtWeyBFwkpoaMu7WGBANUzkG2v6H22Z/OHmsJFoi/f7
1rNkUbt3PQKZX9LkfDCMNBZZ2GNAOJ9EiyezsBsAlIjK43lbVmSMQdE1HX99Ac3A
rSE2Ep09cqqXtlu/XfUT8qxvg+aZwTISXGHs9y6uh4mWZynsQy39/KcVhNzaTd7O
HLnQVOeRbf2acp81xjHw9GhCsd9QM1UThvCapmpOFMU6+cma6j6mgDIWwkoUqbbR
2ljOPsCZ76/QXl+XjJvS6+H4hiQaFx1axahNtCcGRoeh8cmv3c7q9/D0v59t641w
7ttIHF+TXKKO7UVMlJGPqBx5E4A0fnYO8aKenmz2IGFXUDvz4F79JbKXpW++5hG9
QmrT4oBfD8OhgE+nZAaDwC4jtCt7XGvoI2GiPUq/AKAmM2SScLdaJyzqeIO1Y99l
SdvAV4lmRP1OGYIdnvCW/RtRYRWk3j4W3mosoJYteeD7/HK6JemtwLYmuz7qjve/
Hx2xgQ3W8H8LWX1nv2XQ74ImMfNBZkoJ5kvSR4vPNf8r2zdq36TEjI0FRiNdkEs0
RrVqWhTRylvX/ptg2O0Kn1N5kyFW2kfHXmlM6ttkQLGOW7l72oGtlLT0M0n+0bER
BG4WO8iU3QkCMgWI74ym/g+kWfx9nQS5ojLmND1cICFZRwbiY+SlS5oZ1WPmjDP4
+jVOH8t+W5JUlXkQ68w9iKn95jQEv5+qwMWbC184hES9aKlt/uU3MhOlTxDQaS+a
AUiLFNgd8K0EWl40yEf6MSR+KbUucB5qPltYcoBeZFd8ygC8DnIwlTpglFmX13SE
gxLbDia78W5nh5baPhiD8sOwuAI+9rkE1xsG+LwQsYkzp7Ew/AREFl9w7V34Axb0
fkANpLwUD1Z9gP1eZBZaxHkQVOKaQ5sK8lPz4JJNRlluOxKLX9ZzzFDfvGPJ4I8x
CzqkCJ/FtKi+6E1+ExXWbgalxrDiGIakcY4hpnFVWTL3NOpoN+dr36cES84fx4GO
eyoXXz/vZCULQ+Jotsa5J58jjubORGEP66tW3X6zZgQ0CGTRFo/bNer5V2dk8QKh
Lmy/Ldid9rWXb4T+be3AbQIpgIkSt0iCqnfTf1nTpMod3fngXOh2xJQFuXLEHD/+
TkpB1J8J+FEdkXWlOk/fJ0r8l+eelCZjecZboRKaC3VCaEUt0FS2UTA0u/pnR1Dv
Gi10f9jlz+JCSqcsZ1HVzTQJqeVymZyvrIgZQZJqlsXUo7dlgcimJgJ2XmTPbutF
kX3qado5Coxc49LqEdmTLZq4FJmjX3AIxnqUk+7GvoMWZahFLyb8H7UiqfI0P7pZ
SpU+ojchTz07S/VWAHbzk5OLPayI5Oa2lkKbiizAqmxmIOroVpW3ii+h7G/CuNQN
2oeFHUxo/31NxKk6tL8zS/vIBI3EC37Dk7NBmtPW8jhbtOQzKiiPs+p73M9UIucW
RfrgZUOV4V/7J2JqF3e1OCKVo1qwUBe3ZoFfbC11WkRB/WYOsjITbBCuj6CJXhdj
hmCsH9uqVs60F2cUDhd9ZWtBsfdTTpZtEj43Qb3ghIX62JWZweHhjWfHzIXcTlwg
rRr5wTRldR0UhtWN93tYqQiiHtQf5dPrTT1zJzIXG/SetENrWxFycADkMON0XX+R
Y4kMstxFxqYGTQVvy3rRsbvtg9p+KyNixqCV4oQWEttqwQdovDPELKwieOO8Jfa2
FrfNQv+HWCE3z8OOKAuuuVgwMyc/UdBIo5ND5Ib9og8jiob6GYHCG8SHdif1KlQm
JhbtiIVwxvjP2s2gvHdv9COQc9guGWKwMT1PjITepqZ4dMbt/iZvG3QhCNFgDdRT
skes88AE3gebH6v4kx932LNv4/bLYde7kxNK/iHeIZ0V+nj+PfZs8K6ZRSC3Ahpj
pIjfnVflGKesLmNK/Al15+M1avOru7BTUs84CQy+cl3LuViu89DHcpwI4wsWZ0Jj
Qs35bp2t2dGDjZV92QAHtrH5b8R87U5AhRLl1mbBIpxlRKz9BQKRUO8xk55WpefF
oRmpTtkyo+ApHLZ9MF3VojK2ukYrEKZpIBZRWG5h3LZ2VW0NqLfnrQqMqWjbJs3g
rDxm9W48BN0rW6vLexuuznpAcc07C1rR72GXiNaa0kpub82JXI8WfuGz9dgcJUjl
50GvtSTEYoE/wvK/oGwMogcx0Ku7Mq0873AGU3E1WU9d5Aw00vNPGnsHgPt53rQ3
FIjdwausLYjekz53bwbp/8ybPMwtBelC4si80EsuKXY4AP59ymoi2QXPD5dVy0wv
fbOMWo+zhDExJ6WCj6sReBz5nEE8DaxaIKUsO262H0CAf/DYNf1ufQ1R8HvCl3Ck
L5n99fliMaOy8DtJ8wzt1j/3nBLWNgWx/vMKNr8+ru7wiEUaxaE+lYzqBAXuNK9V
rK3wgMgNtIiJQpJhIZuYW0VNZx/whwdxd7M0YEqNy+T1X7bsgl+wyg+goBhnk+KF
rk5ImxZh3Q5QNpMX2gmU21hacCWoPKRWoxDNK/J1tYPxCWzmI8DgSZuoNddzILgH
0TSOYCaRI8MWpQdsYCh3oj7F903RwaJbmnA82r+avi90mbOVRaHmQkbdXgPsDszo
O4N++EXrVXVr7ar9Ia/1t0oRmnV1DFck/cgZWss7Y6KCIRsDZSwcDJ60VVWgJr2y
nHLTTvQTPvs/WvbJRaPAbpVCGDGQc1VGSlc/zTlWqntuvBFMtX8Lqx/KMp7uahao
gIKJuR3fwdLPxXGThxDg7DLG37e+WQeL9YLpTea26QhymxCqh0BF48QAtywHgRqm
3KpHTYzuF8J+K0USNqjSxAd7iMFseivO5s1xmHsBfAsNiGCU4omAJZhOZ3qCp7LC
fobZIcspmxMLhNyDJcKXfdHFsHZLbr2sggf6mADNneEpXKPBhjp5TBwzurUumE0e
imnc+kIrg02cV/GWwAUSL+0ETG7Uj4aum3HC55/sEUaPgWH62cYHIGkAYjlPu6kw
FLejE7UPbECstJ0xZbeHENYTm5/8EtFsACJEY9qQZKSdbhcqkJXsKVRStnhARP6N
+/Xz9fk0kFfv1I8BnlQJZzghKpY2Nq5LPR+YUfw9BiYmCifa65fgQOCYrcRhNW5q
umL2GNk3oq8ALtDf6D8JGHyPuSESvp1QI4tKzTUfmaeU8Dfess1xoZa5EIOdQF+a
n/h6ni0bKSFT6lXNSZkDTYwOsReXjGP/9oEAe/GOghnj4CZ+FfahDE0dLV7KuXHT
nxDTnqCmVolLkEWZTRqeJlZ7A9E8VV6P8iH2oosvSNRb9nLVzi2UYxs0bAhAQIfk
368uB2FeNcZEPDR1pRIc10kE+sfhN7mTSnTauPhwKgZ/ktk6W4eXElOuzQ2dt1AP
Lop6FTXHZduTewxfznK3z93n307OghIxYYpadMw5Kl6L8G1A+i2HujT+m8L0Nbun
2jWvh1PF8vD3DeebWT8g1ErPtxhQVAjqT0zlfxsg+r6dLB6qwxxC+u7DtboY85Ev
uMKjJezC7VJlKkezXv1APWDCP7+ovMBD+1MdouigctKFY4gsQhfn92CsP1wS5Zwm
EjMMZFdVJPUN28qbC4lXC8mVeXOMhlDsFnQ+p4zrYCvff4kVd59HXOggY7Hjandu
ibKSVLtoeuoBFIQNCt8M0wkJL2f0xuLxdBsR+AV6Hrw5BSN1a/1uqsuK5bA7904/
Xd1tcTRR/F4Ygcptix2AkKdTYyYfnpdREfpIfqR9pwyGTnBf3qbWI8YfnllLN4nc
dNLDOk1jrKfCs1YE093VndBkD10sCOuPSspCDTbQkXYkbE9fC91RSZxzxBP1EHS8
xyNzyyHSdh0M0sfWUQsUqshmswm6s+dx+GRfjBPbPUdo6mWsTHIgBUDhSjmHI4fh
DRZujH4GE9yV+adp9Kb2KBNdq6CRhriT73eNAuftNnJ3lZJwBmtnHxb9qu/E00h2
E8DUWE5RT/PPX5LogAiO5nXHfUZq0PXneM5OXTjn8T3AyUmVWiZexei1JnSyoD9U
bizZKBIhaFbNs+v7+QsYmuJtXDzLRVaPBcnOI0sc0/KcjgpKSoGC0DjMzQm15uPD
vDrRCcf7wbJ0F7fKcMfUtmY6TAQ3Y372P4jSGiFQYw1qFm6OhL8JOGsMQAe0xAhl
P88kSqk3+hM6xWyjRDDr5A3DUmPQS0p+zbrznhIshYMIm69VtmAPEtv9zhr5sjpA
wHqpzZgk27kLmRnXjyU/qy3yy0dAQEVGwF+UrgwWBpSDm0PvEzf5k0N/KPqxjB+i
NB5rA48e1PJo8dLIpGStOapgQ6fEQYhlNLzix9j3a8Zl7Oh0INWGtpiC77m4nLaH
hoClqgzRQJn687Dpyl2QevIydbpcnrxUwhazgLJ3ic3NURm1VhSjpWT23oaqfVJL
6XPetkhbw82Tc/QUsuZNzHioE/uvLa1b6Ap5nTK8ywZ4ImbT6jjyQJHJQKWSfE8X
oRuk5eLnbUOgELbsGuGvBYnX4o5BKiv4DGRwu0MqCuBekSk2VAkxX3GTXt40B+rC
eJdNmBS1db5XcMD+GYnFbl2joaPzLzQH8h0ky99VOvDMXsNB5zLcwTdtyhBVj2Ss
FL1eXRdihmiOLuiI76FN2m3KyN8/cLa9JZy7vALSlkIiz/dd//Cce1m6Pc5zHtYR
vk5GlZHXFk1UJE6lHqj573T+OL8w4iY85uJ3A5jWBTRvJFpdhfm3i+mXtg0exUf3
MKQqpMmpTasCaY0qOnle2igfhlQju7d6oT6YOOehM09SyjPCDSjnICqdlY8/VQFL
wYiEBGClIWmypa9h8pymSndX2erReb8/fZebZScAqBS2CzDJIdw7+LA4EEdMZ2jE
DpF2JMYRwjQLyg/2EgzBZEnI7bA+e3tgsoV4Xs/2FpeoKWG3LRjF9UTNaA4QwPMa
/HsWEFnDfngBcarB3A9cGP3IO0vEnpsBd5sBgc9ukR9KQLWBlQIpPFK/5VCnkFLO
SEV820gQAWdDrB3njFhlFmv0XINAuga+xI8jwTt9/h6zWtISQP+5I7rdwNlHA6R2
osDIn+zzmjfiIXZB/fy0uwUQD6afcqTBNHZxiejQ+f27NhN+bulDwl+cTWObQLB6
QXO5eS/HBwwOSgyiMuapERV2HEk6bR63OPDL6oEdIFYPJVXOJ4H7hukzSSzCCqgl
rzBlXv2emLjWhebMBCsIsxhk83UpLofWoWo+cpn+TABM6/p3Vq2YzeE9VKj9U9Ap
y1dVjVSeG2kXhbCS7FeCKbkxW6qN8DH2l8rHSUBP3oJnicJsmK4knBYXt4NSNt2X
2ATSWGoaEzgaeFIRNueYuLRZQ3BjbFVRYSFhjLy6xFnddcjv2PmBW7oILqn58HA7
2CpwGoAExmKSNe4xCXWn3rJlXMCz6pdJp/EbFD/WOZBOKnhY/PfpO8vYRPt7rCr2
E8B4MVROLIgKPi85n6TPpJlaj6SUnky9zqFzSsEx9H+QJrJDYrcDP9wIEbtsMY2D
ucdm6wOuMf+3N9s4r7IZCeFF7rjPOWkwzckloUzqx+MeobJJwBWIYBOrOIHb8pqX
UcJkyjTNNkzKG41qdVe4fPd8bLpwtzXq0l8fsI+PQMUaat7qL0J7Qt4sjMjQwATE
Uf33noBIAywKeW6Q0ucA3l01KEauUu98i2/0bsHWFgHKHrVWIC7kg4+sOpr1AeyC
ZRwAfEpzQPPpd989ZXx1hfVB7U29x0qhn6lOEUvKxFQwtMv90cwdZvX9AV5/eCE+
EGaGQQnMXiR17kbE7/eizMFrIB3aAVzfTZ55ytBMavMPKdVn8Ww0688oi6dzft17
09fJX2jmTawpeJXAuDy/hAFR9AR3+uKVlKe3GqOpLsoQQ4GTf3dXEVRXbSYDRxxP
bPIfjCl0Y26l5k3SYtrrVPQCcRt1mP6vqMgUczNQGxrf3CsoX5YSaC2LWgUsn045
UXOzNxUO609EjOPsu9qr/STdzRo7tR9+Uk0PznqXv7duq3M7lHaUBrxhh3uNypO3
bwVbVuWgmDWkTe48Yiehb8RYU6gRYTQpYitcuw9rItevrSBOH/HFQmrRSr9rfhP/
pok0PiZgu+VwssGYHHnOWXIz9YYLyOdp/SHSbyi8SF46mGmiucw/k5Y+UbhN4h6z
bbj5d5f6nAw5kDI1mtWQqjdZcykzcCQYW3nOaWn70hL4uKIYRtsXrgMlD0d+Zw/P
Y70z8me0wWKLkjJbCkPiB0fYM75gFn3VPj0yLFHtnBPUnkBm2vmnGXe9reGa1mKK
aq67ekyT25rPelCu78vZ9WKFRJebuT7SsjKwHYudP8pvjbXHanLWQntKMd8nWguw
+SdI/3SAf/sFCIf5p8LifZfzSIRUPjtpysn1nJJU/9LYsj8TZsDVlvfxY2E4JKCy
8+JHM49K2k2NqCDkJWWiuG6hxqrPXBr/W++RFGQmHM+2lvua15xBTJiz4iX0/32l
fbW4u6ia1HaJG2UcKLPLF9ADHXHta1Xv38hqs0jvw1pWCUCWPvA1xZ8zZByKttkb
BfWYkDiutJdPcvJUMnakYqvUjlK6VesCyYH6ZyQM4jg5Qd1tcPKgHaANfhuzctXw
iYrl/XGH0fM140A9cnI58dEwMOGp1cLovpwML15H9YSuquNffixdxmZ3h3zSWTgM
R42QMhMbtcyVC5r/57XFPb9P/46YEjqknl9hSudhYV+JhdPvFHpwrmukBE/f/rj5
z6TjNO5SFgrQ9pjK/Y6OzG9Gj4rWOHpoS6gHVPRwbOFb6AD80GxOEWqD+o6Uz91+
PrhADiGu9IkQPiAWdcyHKt9NwfwdXxi46efFJ2NH4Eut4JATUUp8Tn7BXdpaKI7k
BZ8RhnaPhUZk8jg3sqqv1jiUabMsqKxaM9NWUe1QtzGKQ3e7y2utdrecsM2g7fvp
M+UtY6Vp71PojJ0BKq8HWdR0ZqzJtUw4p/sBw9SLj88jH/r9Bo73o8rQqsCbOE7y
GSPr/gNG4KtadERoEeZ+UZGIDWKybIAH7e2krf+LGyXV55tcGG+733ay3Vk9xv+e
73ZJYJR653I2YidITXXWPY/dKW7NYXPq8e4Y+ffOqNqRJ667J8IbFofK6QpCzUI1
fYdkPYIbAQ2KoPePO9l448tK8pnBBKnL/rKgxMjIdzuFJrETzAQR5TdQAgnd7GHT
2ZqxXtU6KM6XhG55zXEZWlPCB2giN2IaQSdlgcXcjZVuMwywd2pfu1P2JguiYqYD
7Kk8Sz4i1M7KeCnOe4wsz+Hrsz/jf6hTIw7dMdjiaonRWCyCLmFZlE16jjlLGke7
AdmgQ2aNsWqbrz0WJawTswluosOnKdHxEVB39njKHv31nwLEadNozWpHGjGWzXfh
xoEJES3Lso88Z5Fag4i1+WTqjUzWniT5z2Dn5n7cmz9DIbWsQv3IG4Oq9aphKrP7
CgYT1g2lDBXJYDOqj58tfPTw09elGqVFVrZU65pydUzVGZTzuLCTvO1Ywpcz0q+/
j/M3oMqPAhrMhCZAgSetygRfO5wkVUdnHR+Br834i1WFnum+AX8TcGSjh2hMy52f
epxBVZNGcuwSbDW1D94N+1aGPvU1ANGUoCyfXQroMq1uKQdPuTTxSP1KZPmuEIqZ
TWZM0fu/HSoFvC9OIksIbrvkxwZCwyhsEvCsya1Rhy94x9u4qAV32voXhBN/BqnU
IATq5GcvyVLQeoFd4wyqlhht6lviRy8neYo8/OZDvj33aPep33TXUidD2GCetT4S
9iiSqmvom2Ulo5Jjit0mom3wa2MlUTDHosuG5ijz7muKmSrYkVcTrUdAO3bb/5h8
PefoT0w6zgXk+YXQvGbotZTliTrigyjkJWq1BE3GawL+0n9JHW/sIjkY5Gm8UshA
zlI51o1CW6EuZyr7L9aDaUYd4di3egIT6WMf+CrEz4xOj4kgQ4SWimHqBClFod+6
vEQ+unk7ALSWRg86x6qof5/I41Zjo0JuzPNb1Y0qbQn8/ZLIGaIGYMA1i37ZsgfU
uU0+uFPWfBGv355m90EMgJbejcl25wSE17zORJn+R6PpXoYjcNaaZc7IfCKM+gvS
F49fVDYSoZb3zRX3aIdGRwmCVYxSaMN9jJC8DiyTrgKEi04RaUuJoUfLpJRxPpQY
aHVTZbFsd6h1B59gNmE2YAGtSHkSR4TEElJdx+MP7enQ46cxA9/I/vFl45LyoJ8s
xBZNPFSETV1U5THV/2yKO6iQBuUaTJuuayYFRlJo3q4XWlfBRsfNP6qy/a0YEl3M
qTQI04oV6oPXraVu5y5tTdRL2dlLpwCupmz4ovhzTRoqkHt7T3sdostFHNyOqAuC
xeLRtKT+Ik56A/+8fZyHHwe1ny+fkAgEnrfnq2Ucic/7qhskNwd5e/ZbURVkk2Qs
MsqOLCWIfWPsGjD+LEzseT6NuwEJqC3iOzlKAU9WmPe2ljHTEgq81PPxje34qJo4
RkVubQBIYliiSWKeVefSgnTd/ubYsL84WesPQhkCId1w0D4ZgE86HAHDLncnPv5Z
jf3i6BBACq83dG5xd9W/z8tBfk4JurEcZZwGjeYnb+zk56+dZSZLGOqeRq0e5Tmz
W4o62FWIumQYfASALetwcQCcmGD1teo/HJ8JbJU0PIwiMe4jpt/7kHv2hyf4hnqp
ds5k/Raxcf8Sa9DXFXTPfslPnUbeMOQBmZtgdWFhR9Fpk/5qapycruiJ858S0GYJ
hY7iWa4KoKiEeu7x6doWs1kBmMu+OZxGRDNzRgsMkuAaLuRxSYA64ga+WttKFn2k
BHfhgKA4bWO9cNFgxxaQRBjlxT0lmuCUtK3yShCHhPjuprmAlUGbJ0emPFCJByrN
ZeGVf8rIPSOVqfSjcnp4/rt+klbLvMWSb5DEjD2QqXIGQOIAar1Tkuv5NZ6i44el
E6MB3Eunymwg8TI777OzRxfNMNFe/m3T76sx0e1lf08sJtC3xxXO/byigL1aDsy2
4GJSJ2fNWhkJ1JH+JpQMmzvL7oyCMh6/BYCYvGZ8Hx6fwR7hsArhrKHruNF0Wgdu
5/MkTKSOCRvQvGfGpygEapCyINTHdu5EGrpKcNVONXfIAVCsszNA7XGlLxHZpk8W
OJfWQ2v1rzMCt+CFAzpYCTzlV6XO8xptKw1lCN5XQaGHlRas+gJXSeDQPO590ZeJ
PchGmnoylBGmAmsVh3P7kmbXaB7aWNB97HKaMBrJFv7JBvRn3TT8C1ridbANyM3l
3VzeI1dxsLdbeqJ35HD/Gd+ch7iBKmZeiV16T+PN6UgWCsGrljoAatJevLWBmKa5
Cz9K+4SN4mU7KnSRroHsGjJ4ZAlhhMaWwRo3pudGbECB5fkGQ0oqc/Shi3xWx8tt
jarSxNUSnQJwj1DTisqamPifvE2+d/UEt3ag1BeE0hqtdi81Kr3I0I2cejuUT53m
tKHXXec1593BTjtVL/RLI568UYV8f3n3MI4c6DjcaM11CgXaZj2ZlBCH0eTBAOAI
cbfatfedkH1FOYImAJ/VwwkS33w5u3lpaeWUXNmcEf5GstLkvYjZrcCMsDhIarCw
Nht+Y+bZmVU/I6GRMwiQ70kECQh6G/z8pqLqt4J6nSHzmLAN2AdpMHdkHsgSUXQW
UMPqv5a8ps9vFQTxZw0oTYsOD7hFB2DAnS97+7P+Hg2j6zhNvk+VNqpJUhERWsLx
rKXXTrt0aVTmFnmUeSZvwMacijzG/Izb4NGBX4M7mB8IxPAgIrN8oO+RY2DiiVsN
O0br4Pebl04wUlUtBs+O0tnWdKYmAJQ9i+d5dVWqgnUHbW+OVcy+bnM2VItcV481
2m8ZSfsSO5y4g8qbSVblx81NCfEJz9K7fNbY/tDxpgi+6Fcdg6rroVYF8siuzvey
FJ0p0nFmUaKP/tx/cqv8u165+xMZN/5cH4UGLl9rLZ3TC30uiPrsPe5rdA3vGtCn
mdX1AHX+6yQQkDATgEDJBT7wD3f/Y/NouBAVDH6zTpJoe8/gBawxj0ON8mecgZDo
oKs3/8pOw0rifY2ODAFX3z0JgVfei2f29XwDCMruQLAzqp15iYPfk3itPj2XhNYb
nIRXDC08TMnA2t/OLLQXVzryUoJ9TzZZFRueCWk6yydlfoeXZzkowXDKqC/kNr/G
Hu4F38fHMJxwkOi/NBVcyeA9KrTaU6+poPh19hWAT9JQ4/AF0If3Gvlu7i8c3k7A
XC76dQR3Twr9SjpeAZn3c8jv+YfyjAPI84kCGfoI2zkJL3bQ8T3A0W9OyQsd+Qzu
TM2wQl2+Hk3+LdyHiIR2fO9Y7XTiVqkca30v5HOomXe4I8geqFEm/WC6EDYOMY3j
WF/hu8YkbZkvPWhTk9kcsiiXirxvO7tylQCQZQpyyRPZcGlRhUer8kaH0ukvTOJr
T6Ql92TtU0P+3BpmZI0fE0CzjVgOdrn1QJsQ6rdzwT4GUl4mI+ULUacSA8DZPWKi
HYhyLTRrcM95VF4+p1MuFUaQJQ8cfxbZaCdw7denrMhG2E3Umqu7C6DEKX1xAWGM
Ptpric5nQC7MZlZM5cctHhweDNDdfG79FkTWqmP8bmw5TDCeyBlbvMFeSgIK/s8H
yhPZzcLNX4WG0MMz1AlO0UoT+z2y1Xl7S7lKd7WTizh1lTtEVYMMfjOIY1xSH8Lv
SQCMMbh4EdKH9UeUTIsCrSRmjXgm9NNW18sgn2snrsqdzT5GxNroAWOp2PJhPkr9
Hxws320dUI7p9ZQ3UiRrT1WzSC3nV5yF7kPim7lRiGJ8osiFMDCMnCI6rPZ/33IM
l96Vdz/mJfGHAYrf8ubYr8F9QLFj/mrw1CUrrguFG5v4d6AMS+g74CPPUqau2r1Q
jV2JtAerShJATaRQeIdNDnH2gI0y/jJ5GfjZO+PRu8dJkHuGGptbrS6AQ9HcWB5H
XAIfk2ux8bipJ28/rLFbm3DHoSppyXM9ByRzmVfNkblI02ZrfVsAaFnEdjKgq8EU
FJwK5TbmkeECGZhDjxFVeRtz5AMTaZ3dd3szGhTpkluQv6nGiQ6MqIwXezZ3JuNe
ZBrLjFrI9wN27O6KRMbu7wW/2Xlvof/lMc6CpErIjS3cOJf8wVJ1PeAnBzirnOpG
fZMQucZuE4RYL7fA7XxEfk8eJaroljCBkQts/c2qzBEFsE+v6/QwqjN4Rbyj96o9
gACSzyf0E0z2JOeJawqqHU1Scac+573lBvc1qSuODFcZFOiqlTSBLUS/sR/Atu2e
Lw9HHK/qIqU2jrcCPB7e+9OF/Oy1VMXy3A55dnxXASt+WD1Wx0d9aRj4IRDImo1X
aaSZYR9+RH9eqzCCr+FTYSP614NNFPg57jx1YGOITuW9KZxNKixPvLdOo4EL4ASl
WANXAGyxoF8aLY8/KbmZMBBjjp/MzPnJa4GMiZdP/03PBXFfodIheXX7EiFiNgQj
G+kX2MjBtRbanITjCAImPYOq90U8icBmyZEajBmyX6do6kIDHElS907PjZsdtlLj
FX0vbQnR2XbLJIYeXDWkBQEM9NT9/L7Z9mD9eEDG7JzgM1BtTrKDZJ0f0/58XlSt
6n3bwRbgFlwLJmbR71HPNIPMSr4jLVLgIDkIKWXsIif9TT/2pNQzZoY3t9nsLXVh
gIUHYZFtLxpILU6EiHzHKo0S+zx1Gx7RTO6LNyppN4TqkmkBZInWQPUGX2CLWIMs
7WsmmVrIshVb0dqmvcdZFoQM0rjZi6yH+nl8xDIjllgg6AmMTF/C3YptjiiPUvq1
QZDW3YSYSxdXmqZt5KAluCmPobt7bhf0bPgY/ibWO7vAEIiGslNQ4TkqjzI5jkvb
qKsTp0hZhCZWsixVJfC0A8Tvh+H0SdDnKZM/trWBA5xS0WwoPRiayPzfAM3Obcqd
AklyubzJHfDpN6L8I6KwAJqFbxYeQZqDE+lUkjhUfyo8EJGEKV9/d6KFE0B9z7xF
S3Ilv/OpgjUFhLtlcXYjQbnSKKzqc0++H9Y2Z1u4RGnssdVZOJ7IG1+uVhgxJLqa
YN7rxr52A93srfIaFVqBTyJxgrkKPsmZ85zd+mto979IL/w9s2emqoEHgTm/mhki
w7JqBUAe1tSvwy/1jiaRMBBE+b/c2EP2DSUFe/VNvYfvKB7o6f7C73tXNCYPHjt4
i6ba+WrYwQvyJtT7A8GBrJM9xxKAo252/L5r6Xnu5KKWCBpm0otnH6089/PH6TBd
Mc3W5/l1Gad1qO+7QUX15weliRKpI9o+HPkwSN7WkrXxxtX5F/c+IdeS16iDbeqk
JcEix/oED6gCP51hNiYdF/OCYcHc6941qHpxGMzKKfNNWvaey0LTBNt/RnBXu4iu
INYYnOrkJ0hSFGlN1uxOFLoYhmlg5CJwW9dO8QXfZpTH6oBPSJiKqJvHBtANMdxf
5Oo4AvJddHsfKRMdaDSw/r6zcgm30LiHWBr+lYv/y2pP6Tfw0oXnCcUCzt/9JLGz
cYeXqy/JTGHMUGnAnhZ+cHYfTa0mGNr9k9fB2vCYQk7mV4idz+80NZXyCcE3yOgD
KisiQjMB0Zfqas9Vntd02gqAvl0KV9i/G6QGNyL9OIraALlmndnAONrgxJD7MjA1
+LPPWAJYUAkgfYbUjMtfC2HhEgbVNy6V7MrvfO7zCMJIlDtxCQlZRjS7VRbM2UC0
VvK7sChotOD2TdXWRqWG7gbfIvyfr/qJby7AQlGK8KhK8gvkEl9hdhyMRHDKTM94
VOLcct2DOzQT1A7CzXXd+nQ8zDUur6MrBzKT0DdCGkdN1cjI7L4v8ftVT8l1xv2F
okM+vVV+NzNzGIW01rgqc5FUD0lM7t2vx4gMdY1k3e3vJ22aS/lfh5RR7NqKp2jV
MXQAwv1WPeHFiACA6OUib5QfO/O63l5qUftariAoDa2ypfAPl233FF1k10mJDtO1
Cw0s1K5R6itMCfSiqSZ8ohmCXRLKSiXJnHyHsvC51bdDqVsmU0S4yyDBV6flmEge
KtEfuUXIf9pT06FVrfIt6tWIbxKfbuF8wiFIpLipv9xJ7hrADOIn20gGZ5EhxoPn
yIBn4bzZF1fRzvgJ0iQH1MQTfTsHWyPPy23BEU+G320a85OT4ofhafAvkCdgORr3
CWyy/Ys/anjZRU+5OnBVhvh6hkpxtbmHgLHLolqPnwWg++pFRn/2wEKRwmxkrMF6
7k2qK+G0FlSWhbXcblmc/dlBD/JMuXgFhGFhj4Sm9PK0uPLiJvzoORl8i4hW8yxu
45vk7NQ+HEMLV7/hE259sQH+ClyywDSITHGeUeFIthJDgxdF3/kslBGox/qXYBf/
5rETe2pe1u9GJnuuM9BU/7wHSq4GgfTh80wDYYzEqtiE/hxZIr890fl6aTeDv8F/
bzADV18Pkk81S+ozJBZd52X9eFXL14ptxB+eSiUpTECiUV81gKFMMfvPbr9S53G9
U7Xij9fs//VC3b2HaV8F3UOB5DxSkb6/K/yxWLKZGytCfd2YNowJei8UrcRlPsVY
JotKToT/Wz1RwOI5HMs2FmYqI5Ba0bHyWSL0gqKGI4kUVMeSlvzS7yaj62gxPDDf
indF09R175+WuzUHKVg+He6FJdz1NQ8htKHFZisUsDlwaYt16NorIUUvRDfngF2X
YbE7OmahkzJKrLBLuCHT5P0OHmK8Asw8HVZhmxuYA0qZWArTH974u+zuv5+JS6gX
TRYzZ/fsuhuFMCfidu6YcJZlCw6DUewFaYXyicrCMfzMtnpSVKQSHojaq88IR4+k
6QbCkrMnovAOkCo7goaqbtJ7A5TNw0gbhMDPpwidnN+PDw2nRoFJMRRCqGnX9HXQ
Hhiyr/zHjIGCiOFo2HrbyYFXQg214zdQHR44vPk+S9+Ek8o++n0dHpPg0mzFla6u
5V7QDIA/RD2h9HfhHHeHkyDhlDhl8WxG++Ac7J4LITuc7W9TnOslIV3rvZq/xHaN
8WTOX/zwFEdywN6fy3a2d2VdCu32bht4xa5ojrNshnGKMkeVDkDw86zLc9u34Cxd
ChB0vdKAsmYXTYm/MqEIvWCpJIV+eqkFmqFBDBbxZ4MW+hwvbglw/LZWVO5R4Umk
BNKS7nlr7UzJFAF/MC9LHCT334C1D1mohI8vUjk98oi1i51S9PUQFfsXDXFc31mR
mbH56jT/ZfM87MQRzSK3d3OCKi7/O1R8SaFrwKka0KqcypIfXqfjqYneZ9x3MvGV
K1abwnwQQ2WydP0pHmhXHMt962VjzfHroqz7jAIWCRKqWweSmlJ42SBIvRel4lkM
tNEHjuOSAQ2kqa0ygedra4vSB2lpKPKAyCLN38n8qndsnTvZxYYucS4G6dlamNRd
WVWbWm+aDHvWxTT7SYo/w+j1vGYjxXU42QOl1n1KeKW6Hs+tL0acvg/ahkPjJ+bo
pxxnKZvDBWSLpj9v4m/at/oOYJcaZW58bN8hfU0AXDVlPlEKFO8nu1GIMIkAgF0x
Wu/4+VAMHoTZQvIUm5Z8X7xNT2i8uWsiFdmftYKqKDEiAGjFF8uGZfkDzT6cUxyk
ZAepH7KG8GlaUDJ2QsEH8GOOq9CwEXAVIqojkxZxPBmuInwyDkIyanpmGpf/9Glc
DVdd0SD1AiObh7YFC2YY1CDmIkdEGsruc15YbhAt4N8YtYF4PTkJDZ66Zs9zsTWt
YhMVp484XN9/k6Vg/OxVCoGK38fBSOJfNjJaLjGGR4W7gLz861NFTDHBpY00hSIO
Z8TvpMnBdgy1Vt9vZ/n5KaWOWCSI0bJXWYxo+zTL7mDjlDG5gjtPg8TJKOqWtQSg
WV2Vwl76DSrvWf3wnQ+r/SKJFaSRtdN2C1YR2n0u4ZdKS6wnBUAhET+3tumItv18
8X6qHabJf9R1/+90xM+I7U8R0ZhcGZfQ1thQykFCR6FJJkokIp0y6dg5i7T3R0xM
9kMSTAyNRwMAADZSQMwoJy+XIZRYKUMiRI3psg3iD95jhBjywngU79tSvF1EFdTl
paQeOgLYImzzjl+QFc4bq2aegP9gpBinZsaQAPcYCVSKE2QS4ir0eoGU9ooDbCg3
ugOq35J/nKyneMU/YDQj8Zh6SfmYLLFwjTur30XRT0XH/NPcjj3X6xRyaDsqUDIT
eYygpNg/oO5jXxQwun2oZ7uho3DEi4H4ug4q/pheAoByUbqARr6ZADwm/L1xpfRG
otfUjrppDLVDIvywNDtJ9Uo1FATsrI+JCEriO0wTFWqWWCaC4bfodOuPtjIisO/f
vIBR44OCNF1Uj5SKAZwn29KhKvEVhcjrC0/S+BMkcGYUmysGCC4GP6sZG3cXpD6S
S6on3PlyEFLPmLjVw8keiQoWni+Xg8TCOz025fxzWmzD0uqPyU4sm2FhB+LgLxtY
fGFuOT+HE19uiHDwOibiA0qvIhbcKsgYdc1h7JqrHsNOkea95ggX1qC6kINTW4Rp
ht4SeuHkwQfmYuAdZP4aDlr3RPc7xaROV+8Tu+8gJmADWTQ6txiy8AalYqFg55/U
dA3SL8oyaRh0+HIr/8a421TMgsuo12MaSdvWkI5S2KbTp9lsOpIQsvbla4jlSyN2
7foyXgwJHq6p7pDkv8LW0+RpB71hOke92bJ2yGNtk6+KTXtToUOGadymTEWbbb0c
Er1bJ+jBJ+HQwFN23CPJTnoj8cJDwZFFpuviRe/6BvTEw6aTFwcJKQJ5rvOpemte
+nttGCybn4cckkoxOTUjETo/cwIZnUAfsUpLziK46UmqLWYd0fdh8fx1DjYvQAes
wBx6lj0N47YZjEkyZvTa6zh9NwUkKzORftqUzxVUGEJa9jHTWKnGFMe9CdoFhNgz
RQz8RPL72/HCTvM9g+nDq7smxhe0j2S3S7EnrL+KcpkZZyxuUJ3kyt7vShrhp8UK
RW++pVkPyFkSM0g8KdpHKNofdOLfrowiQvGTtth/VJVxzsJ01nj3sQLS1+U62vKn
SLGdnu+9lnU207yncxXkjPHCAnRJfyQr8MbBbWoDqxlfoIFJ5+5jHKbOA0brz05x
kTLVl1zjhj1NUMdvVba376hTwpzPq7ZJCIHe8AYpb3gQFHY72NPviDdZBbvqevE4
BZjmLeYoixlES1bV0xhUG8rav+EOXFVidpeqIm+kz9mH51ZH6fr8lyoPCcNiGqnu
85JQAgPXaQtaysb+inI0og5iUXK6ZiStBa3MwOkGjoJvyPuG/aeSA5hOXBL1z1xx
RTJhrPD1rob5H6UBxxE+XsN2+aSEFqgeqoHGNaJbdBF4N7JpuidDl4edsSKsXMGF
SmIw/X5j/EZWQjGOm2n8ggw+YntWpLd9uuDQZV8ZHq2xsvIjG87W1mVIEk9rlW4c
c2woUzF5IoOud68Nw3P65fTlUHOvjreIFm5WaslK3NWRhCbUat5MX86S01nNYQXC
R8SocVPHZrKjuDxXZKS8Oc+0xrrUH6wBPNrfDG899rdxiBZq8eklO7RpSY7du3u3
Y8O0iGm2q7AVxswrVRT4XEhg9qoS/2UWqQPI7IYRU3g3fgc+nYmLU/yE3iejeza4
KmptcC+rpXVn7IqQ6hekl907Ray5mmIu8YvutPVoXD8pGneZM2MkyTO3t3r6m0NE
2YFvLrYTYhkTZG6naiqGkwgrV8jJe1joFMEvmXxwhnN8BrQz8+oSOqjn2IpsvsWj
+zVKNyKcHV5W9FM2hftsdng4mXV56+1GPlptvYUpSSbKdLqgk7m+3oZ4lQleBPnX
Xa7kyQinSCBrdbcCbqfyBPLve+AMp7chcFfv53KSP59YFm7ojJcwgQYluTF7yf0c
qPXeDpKelBLnJ0z0eQXU/QEt2qBK/75Thmu6UydNIbu6z0qXVjXcZZTSYig978Xo
cDdrmQg2gOIPOUtqcZfgmkqJNJU+LlULfkxHOnNe6BQqoofi9KvRrMZYNfLKfU5u
aQldDyvewd2UUFaBr5EjMzMnFyBQuds/uJ4tL59ImXc2yNgyZLjNmw/WcU5IT6eA
owWNguNxBgvR0irfwN3GipVaVakMWqXPWUKU3tbV5BWaDvArNuWL8WkRyE1mlvRx
zei8JyBrO78/7k1nki+bsRPWLYZjfH5OlXmDrcnjvHf2yfmdDoLfWuCEyJ/AjkSU
UjciJO7v7wY0AsvqGB15A8vjMcqXU8jPcli1ZDYZXZ/+XXaVHxAA3tYLQH6XFa47
ekC+nS3eCPo0mf0V99AQh+htoNgXvMDXAZk0E9vPYyo4VJSAVK1YOlnzd8944EVS
XDdC1yOv9yS151IUBqOXpTGU9rvVdmULbckIQQZ6CD3sGrGohNVD0Fgh1XkEl6eY
xU+54IdkYrP2UVKSIS1wWRxDKjmTymYR4fXqoSdDlQ+w/0t0cTAi5BIPSLwQcfJ5
4ws+pGjkApidtKj4M9bLvqav7m1QDmLJxQ/Hn5c+DMhOo1BOf5LLDaT74RR1HE7L
JOc3CVVS38u7y76iTUixk8Ke51N9aWxFH7rLCSU9gAjKShThRk3o6z4950zyh9X1
CbXuLPvMQPcGuI6dlRaH/h95UJV/FIcnEsSpr1I3ygLKQsCgRyjweViE3dnhlpDO
YmgLPQybS0ssOYHZt1X1kpNVrucz/7zOlzvNwUHO1X7QW2TyZO5BhQaG5+4R8fWl
/2Mu5OXhz+S5BftoGE1S+ACwoOBWjc+bMVyd5GKQDbzCeh4F0OlfPnbPYn3TOsMM
HzQFbQBNVfOHDA7ZQ2ihCqbA682CDallrjxt5CCsgKjB/4qx2CBQDV0HLCJW6Ms9
jyoMQTT8GdRla31IykX385+PhUlBkPqKy2ZaMjwIEUQwmlB99/QuobHE/7fP0irM
FWNt+fFQGWjfcKP0QmzcwdC+xf+asTOIdZSMenj7VPk6J1CwsajJlzBuxJjJ31Eh
PVjGzIrWAGlGe3M5TqeoJjJ6xXYrYlrm02QGI83RVK/RwSt4kC3BzWnmZuiXA+B2
Y9+glDLr3HznwGKJhZ931TVDouM4oQj85O7TppvgZzrwJ7iiZKlKELEfcxlFf+Mt
kMHS8p88m1SX9TwtiZnsUbvn018jySFRoaq2fuBfHZAR979pv5IWEfP/Bb/minvg
H6sEQ9x37IGrtmCuoj4mIu2O7rp/5MzX/9SoPwruiP152QZcZWiE9CuIDYZR2xb+
3FKKCizInBY6ZyuhsR642vTW697CBPFPWVQSBYkIDJfpqryI8dO+tguTqCBPmbZv
M9PIPHGPPVOlDh/uY5yuX90oP0jICtieP945w5OvnGuCTVGTPdxn/JPMHqqJmd6r
jtUUO5GomDcETH91DNd86C34t/Am7Z1qIbWGnggoX3ZJd5Ztvea+mTHIeQXz9NrM
HKMCEExjxhOBe0rOt+ED/rfFYwjBYOAB2f24XvvTPVjSVhb7+Gz2+ISgpLl1vSgo
ognRk9kP8FpJYUkNTDykFit++vDPfut8cr0SC4g1e6fAbDUcLANeVDCSBHtW7bxe
nw7B8CAqTlh+EtuZHJYPawh9zMy/UsVQxGO2q0NYMvD4cYdRFjlLiLcB5uqbKJl6
6sA+vw0whc3x/FU0XC27Yqos67/+cZYmioQJebYekot52ka/GSXqGr1xnzxRFRzy
CnA2cw50xAswiceK58h2myZuuHBUJh4k18UgCJxJYTRwQe7PpmSYBIiobTQnhM0S
hFXq7pD7vkPGBApOd54rhQf41aC4pqpVOuHDtiFxquwQU8FgCsOgWfhQIvsAIs9d
52RWoGoplv7lh4VGgW49aQwRSZ4214UoTdYe+c7uA/UKnFBJif9ykCz9wThMZyV6
ITWSGs3gGiuWBogbBh9twU6wQFjqEzkz62TkKT9+nStqn8hcewIKslaLXGq8LNvN
9L9qylvumBY7cPdgbcLFFpMUu2tHlTi6dzLGddpfLd+UpLpht55YtjWAeBu7vaag
kqItwc+Sg0aP07s/YQ8cN/MEbFn0JMpVfInGeaxuy5Kjm1fYYZJ2btJ9G7rAuU79
9lAdrCh2JM8gjxYaVRK4TdhvUUJTufrIUAwskzUo4rwYWR9nXjPBDHbKnXEc1/s+
tDd+7hzmyfQr4ADzK5m/M+YsiT9fDPdu8wnytA/B3t0YGKLNOhtFOxiRFNxNZyhh
nCbujcyED+kDzxkpUHazabR+nemL093Q8ozY27oMEfjoFUHRK5+cALQbr1JQj1zb
0gNP9/R26s2VQpgx53K8OAbSo1M5QBuBNWWT50X+VRnlwFCkY4CV0QhB4nXzSrSE
QnFGVKEtnsxvPyBqaHuPJxS9inaqx9HmWkO4mh+VHMv2QE/7q3k7/nEoWOiGQuIK
TQbMP76FTkrWV5hUHRHuwlL/W+ylhkmEsSdQnxDZTljMMAMSSneHlLZ53t8fxftM
U7vAD5t7xAcbIkf0Nle5h1cAMNghZVpR2uWPOKJ9gOP7nYVMG7ghGbvMXDiOZsLz
1kMQ7m1/w8w793ZKGwM6uWcroKT/EmS4OKGNrR1QDnkxbvSdSgDFsv/+eRKcI2xj
tjH6oTNekX9c4Kuxe3513Maj6L1qjwtqIXaD8cA2+Mb5rpiJSk3wqy/8JcLlKZSF
E31fW3efXSCquwBMY4WhZ2Bb2sRo4d4WdBI13ietSl/w7ZivmTNqja1sHer9JiNH
dFjcDubmi2m+vWitqRWomgFbuOFeQyU7upXW5+M3pZewpVGS9Ra8EKoWQFFzA9C9
l7fWhGwTi0Wa20PFIq8yXnTZAMofGB4H176lJSt0yppQWEhfvU/ZhdPiut3FkZ6w
OSnEOcgd1pmsZiEnSe6zV9FfnU4qZfBjTdRHZoRVAqvIwCIvtSnbU9wQ7bq+xqdm
o3gYrumNuTiGcd7ixYrnfOPVQTkzDlwVWD65mA7ka19WJxeeiXBZamndjPZssocf
iFxj6t4Nx4PuHe6bbitvV3Wpm1m+l/lWeP1ehSaf1QUHmCFizNGONgs3/z+VvHGt
3V9EY+SICjy05TT8qa9ehgs2KT6kIeljdEm197q44rq+kldCweaBDZ33m4YfOQUY
83W7iif877VUexPmmch8s375ZRdqs/0IomIGummLqWKB1M8Vn/CkvBSyx6rHfrNE
c+eoNXVkl671BuIKycSd8Chj3wkaFgx6NrJ8nhVOjMV5Tt4AGbBAkGkM4/8wEwZj
ryYB6nOydG1wL6yvxO6e479ky5KiVFrwiGQt1M9LBITxVnbc24VEp2NzD2GQOXyW
v03RqFLLZOqo2lPw84Q0pXJ8/oPpzh746pC80guUWSwhcTKrF4esDp8ZM3jgekIb
dEccQtATsZQQM2/+O1IWN8HFQSfgtKgyl6WslpoZj1TgTxSbFUY+EhXkJck7jiFP
LapVzhgm/RnO7Hp2eXRAlfBePfHX911dEvLEupLG1+ed0INNyaC03YNUCcjN1/+k
8knIqBAkzcRjUy6JxhiEr7VacVSkxVHHDI2NZmXAoUblWfSDtWAs3/A+cMlaAavD
BPWzZIR6GYtlDvr3kg/6CK9ay/Rcqh9C59W5IFhmO+Y3BpmEyVH0GnSsgZeXjWyZ
jg26faaiNfmEBR5lH6TatNTbdiP1vNXtaKQsgT8wgGZaiCG52gejSgkVrGw7HSgf
M2W1Z3PzEcX8eY56z88kssLeWz22mHPXET0/qrWm/mMo9tx7EECY0lCPVbpTEsum
Jr34EsMOaM613Z4HJuuuIvtXlyTHLsJM6GzMLjB8GgkuNjSWLAbGiPrbNIEntBSL
pL7hN6ow4zXmxIYaj3sRup0tUt10UzI3syzPBUax8Lq1toiw87vjl/yESTGpTfQS
coaJ1fhGhjjj8aY4zZNX5wn/skdBhMYbHcmCI/X9Gf4tSPL1wnaMlx1PUcJuSEB0
M5QIUWZEYy+/AMbAxcCxoO0HpIS+5e6pOggBPixLMZFCYecFrPtZnZ1P0Wm1qQ5u
NJF1jUvKFdYGPE43npk4Hx98WXDDNnCEeXFPj8yoCtT1BHJmDY3kz7nsf7tMWBBC
mHAyTXQuU6TELCw+1EauXuObycxqK4fYPNJTqXyC6hoB6eyEZUK9araPVQrvd5E7
1YFwIeNktvKOdQFiF1JiJxo0Qatv6O2J4eeR41uZVR0IhSZ565DmqBO/FkvpOXes
aNTXwmhcCxHn2QaQ1iweLgcIFBZpE0cQ2WwHI3tTnvQT0HCxvMvcjkfn4Lm3HPwm
Dg7DBmj4cy1aWfGNCRcZrRYVSMmOfoL9RqPVadzuRGzyvST73SVXZdEZKzfmzH2T
ksWUfzGFpuodwfV8Bes57ibyTpjyTZ2drLMOI46criOTZZA8b5E7pxDpnMfjXg9f
KIeT/Ux4QLXy65V8jhb9mRuSD/Qm0ck7dHcdFT/EQHInRKmCHSGmRP75n2tkPM+I
9aef9fl4Z2Io/1ywTfIKboVRrGsa57N/e5QkbzBQpnujAsFg0YX/bWK5P8tLMKdu
K4GPhAdrTPmNBZIdQKJvNtsF6WQ3ebLhpzO3V9FOYNdCuuf7tbbhU25+MV3/WjVc
k3nY61vBlxPB+Mp2hvtMqA2f5IO126I7rRdHPJLO7GCMp0swPLRzC8Kef52Ux1y2
LQzBYDZdSTpDfe01Wt06dGY0W8DLaiARKQVohz47c8UI//G1Fm8tYIv1hx45EIHa
UzBPqkFKFzFnDBsg5jZUungNBhBmkL1u7ieVD6XgIVg2gnl09zz3a33WJonYxnpI
XI14o3zDwACZZ/67MZMdJhisTYoOKi80zEYzFJYMJrv02FNh2npG1z+zczNtvbC9
FXK+5a6gku/E3+8ZzxFeBYGENKicPrMITQHVbuAORAcyt28kgJ9HqicPHYRh4aes
AbwwRzG0H3PkQqGvq8mz3LGPQk1BiXChdOLNhm+Ff4rUwqTmhSdmt/w/2dD0UcZi
l2x+5nO6PjJPTxpOeMUdVXVkMRU2xBx0QE8uEysba22FpIaUZaSFIOQ3wny5O9Ar
6gdaR4M/F3ifnxROofOg5cY3256DHbHTHMrlWCTcLCLPSC0tAfgK+WzmHkfPgpZC
yNiyGGxXl7vi1DPGsulVp0+dgmTeruwbHmWXcdNNhGjPj2eidmLp6fROI2zSMQ7Z
uVboZ/4vu4nCZaS7wb4SkleZXZE4ihEqMx08L1ncj9Wf95uKI/Q89d6eSv53JCYj
I8VXYxR3r3PhkxAq6Wsb/VwqV+Doirge58G1vtmfGg4O9SDio04OsQuo2XLO1Ywf
ne0im8PGjSO+svcB3jGsK8D+ijtTlTAEdmOjYBFB7lcuKgQJ0QiOyvcHkmNL8Fgc
dJTn3Am4dwW+0mYK+226/o3uVsyseI5Amfe8Y8/pDhxd3nnuvNmHklAy/9QXqqSX
aHbudbmngVgh+ZepqG7a37CrML65IMbJYZ31y7fCHtkZAIUgpQJAeUkYSVesJ/52
+fnaC+9WMk3bW6EjF3uzzeim0zOPSkYul1kbDpQ5B4CVFVFm37wlJEvgswwWf1sO
h1W4xi5dnysAkVp0FJ6MLWw5rMVfAnGMMHAeJruruR0EWt7ePnIi2qc6Q4yfBmE5
QhB6CCDuUaaOSJBx0LJ5jmJHnmDTr3NUZVa5CfRQfJSHAEo5Rnxp/Ui6t06nA94Z
X9nCqh5+ReYDKUX5b3RQe/GpjjJzsOLjB+llUNvDH3tP73BFejDgaj4L2aD4J0CY
dL83K5lGKKO3E5aDbxPGHMQOdW91TXj0FCZjqA3xOraYE0OcbKvfzrek5GuoYSXX
KSfqT9SJ1gwdTT4bxaNmSMooa865f4hHCR7tpsHqrLedrWIZWrYz7Dev/HWOQ94l
Tyu9AHIKNiRBGc81hjSsFwlNb2201lLQtZ5bhKTx3Eqp1uU6vcvx4jc/+j/c+3Ru
MxCYihySmN3QPeauuqaNkcALBdBgYuyPnc80WbMLFZY5npV+AthSfgsrZeQv+GoP
qyIbaEfnuPR7hL9EfylAapiQ/YvXMJk1kNpIGUUssmCVKIn/pECuKE9Evx8UgNfe
kj9Rg7edqMLgmkE9hwTY3OEq80+krTJl+Qbin/oqdVbNdBT1SELdt2IcfRcS3OZ7
hLA/m4o4BznaJaz0hhn1HqNAgk7KaacFatpncRT00btlGFq2dv5YtBp4yPRL4pV9
sS07R6qbPPwT0j9f3BygTb+QJd6NJgljtT37n7hBc2DJPdwKciiS4r12K+aie6Iw
SAycvARbWfpqK1V2xdTMofjmLE4+d7nQSNWYXwLkKdCFUGoc45VVfWr6CQ0KiZAS
Po/EVRjtDZLPvBJStC6QAx/amVIJ7ciwM5IbSM1Kj+zg0FMA5ZmC3CsXNAo87drt
o0B3h1MAQmab8dY4kiiO6NqRXBkFtd0BLVm4W/osWUsT4Kdnl07fQpp4la766gGW
d++PkUisgvjIBzyu/Lza2XJsg7W3MDEdyW4H/Jmt3dpOIczuFgEFZK78pCQaaNpH
wOPr3SKllKMrXwJSKFmsCqa8W/qvVEMKtJnG3AjIHSgsQsYc78PaBlUc/9bHNOvj
RSbyfgJyu+eTrlQTkEpK8mpf9/SZJbeqgqHNnC0TgwVIO7tUjbIJJdDt7b20KqmM
cBvqfNlpOzsKK87RUkvuHDzzjbqgCfAjQcRQZ+XDNfQ8lTBp+54EpEN5jzk/MH8n
L4wIeEBJzJq2uHGYPfHy7hP8P93Zxmz1MaHXji+WWxrJTyK2kAr7yevuTKqqa5eS
DuxlSXBcouZeTH4R5WdJPjc8V8Aj2/8M4UMbvP3NSmFHajkN32CYC9qjzuEZ5d2T
HDrvfyJ9QLhSBSqsSg+oKWCneDxtPPj7Iq+Lh8GxIi1Am877kysN3L4ww9GpU0Ki
3fW67/xdLrrDOCgxY6C9uZoLYX6rxt2XFalrJU9UrbtEQiJTqUFvKDIsRGPteQ1N
Y8YaELZzSBLJj/w3gHxaBEEbXBoq7cOk46GI+UBlNlJxYc5FubyzV65gvlIo1OgT
jx/GSFHdE7aYjV0gsGmG3kOWQKC8HmkJcSAT+RidQVk/iQd4pr6ds0mEIl6cdF0M
j5wYZKgtaBMg143zigqon9DAKPoOSRGXnGXaCzjfYTr2AN3ZwOBIhmbO7wFls8s/
vr5hLZfANuj4wOiv47xK+RtFkA8fWjV1XKzpu5uA4wJZJBIjeviuW+VAwK8LXp1W
dP/X1aNX6HSn4TS6mNsRgEqH+GLhEeE6lx+fAbpeuHggGZRbH/qMbXYzjoUOx0JN
j8ZzrYj4rF1kbCzoBXOjNUf/JDxQ+vev8dtx2hs/bhMBCr7W9Jtwjb+rFfWt3DQp
Xg7gkGiibBjTnG+IubJGnAlpew0u9ZROPYvvIgt2DNluA2nQpSpSnx1q5dvhPFWX
nFDTwl70AWJKBhu4w19iCs4sL9yplouIvK4dzOguwoqdBFtWIiFB9TlioDE+f0WD
PegE8KmQ4DgPGrZmlJEvc6RU/nE2uWMK2PRUmwJxHruPum5OkTN5w2b716qMtu0a
pzgjHL8cD7E2v6LD01Jx6PObyZdW0qNh4KG3LI/RKlp3wtIqs3BKvG6Tl1JP8HCv
bR1ddpnk/L8PuhFFcwE78bvQQzpwVrp7xgeMODku4ZKDeMKACtbyaXxFKaJwCvK8
ZpKpCw489X9J1upyRguHAZntnzA3kqRp3T7v3Lv7F0yWtpsGUGTzOmj57QY6OJul
4HdEdjAwyFI+rgqX0Zk/E+8gFu52nYKJfw8lUQKM+k0jztT/1vKQcbtCPCJQwZ2/
YSZpCog2kn5pIOSIYSz69qf8uFzI50x6LwebGs1q25/0tGnOIx5nIR2zly2o0JeO
uCH1ys6yrMUZxCWhNb9VomwHJs7kCgPgwJsk4UgivctBcqWeArvgPP4h1O6zjuse
XtwTs+FLIPvCmyC2NchkMzPbwGMR6VxsSJimT7XBBOs5ts9id/BTMM9HDeX5hmYc
+HeRZ/qeRQ1plKVRAnrcYF51OBMcY4tfKkj6SrswH2ajhvAW3WU/j6fg812zeZta
qffXddNFVLZOPGvv5M1Ij5AynWtzJjTKiDuaQwTPnI4Q0M0xI3A7NoqHvfyHoBO5
M6mYR/SC2G5+YzFFV/xfW4dv+PyosXPwvXe9xHK/60tp6ewNWVQnwAgIkg7LBCTb
lVzcLekxqKyqGLUaDH9r1g1b7D10e/9DP29ukbay9nCnQG6U8dG8twZNEjfL9OD/
2Pbehfn8yOAM+J9e4Q+t6VriRg5HaI0Cl/1/jHkdT3tbTQLymKZ/QNZaG/njXdll
+mTz8rFRQxyu5pI7HxXbViQlq0q0GSCTRIn2hFq9h1S+KXnCXEDl91eaK6raKxds
aYsgdW1zauZh8Fq+/XOyuunVJEh32jnc3Jhnho6pP9ctCrUS+W2XfxaGzvvUAf3R
IMbXdy9fjE+pozmQBUc3VCbPJrH/GBRh6KKlOtFmrP8P/U1TV6l87us7kX+if4hE
UKc8JarldvtWwTApylixYV8BAC/xCB+k1r1lZlQJleDMGSDJ+DSj1Ve4SaF50ZtR
emt+FSy+O9+Je1g5XCteGjCgCzdkMGPuxiwQAitBDUxyL6mTzs9wK8KzJ1wR3th2
rPZ6LI6Xww88kqn4TpK9qc6YUWy8sicvWcwam7f3i3tKZlAKUJlkr7MP8lcbj7gc
Am5XMNNTIx+adDYhGenZzpAH5PJFjlbVVpSVZUm7800ShWWqwQCYrm0ixhU2k2lT
7O71Gm7t2iWFPZJMQ1MjaPRYSdgkHSOuf1LFhOMDqLZI+53TNTpVmbyjuj//vGNY
BEUs2jhIRiPTM/OQhsPj/bGb+mBsxvmb74toF6aIPq+Dp156qsBHX625stRtSgFN
bI+DYFvn2bc6OaqRXR3MFDskhrhcbwHE43OqPKw18aHBrp1BkocvjR+4oG0HBba5
eO6r7FT4CxukED0YxB7c7IscpVvrFjfoMmPC/Qh8EBwtvxIhwfOY34i6c/WK3HoO
5Q5qFsKdieAfDUmah8rFQp50ACt2BspPnc39ZsxtwhVH6lU1BQELJot/LTVbHNxW
fhfZgGEOl8xo4CpPFy7HUIJ2gfgY7O1C4kYkOrz8jNFfqKqLypIAQvx18FikNA3T
Ovm5BRwvzWarFo6pepoeIss5fZx0M6RFR/+xMlB1oLc6k1u4YXnYg7gpI9kjWvxD
YaZK3Q7OmJFpDc8oe/kPqUQfLq2tAH1tITiYRnVw4DLybBJPJPOIzKsGc8bv0Xd6
VvgY7oos3Aaqh82AJq2QF3inv1+QDxQUTWyfWnc6QNfaNJgrAoRxeBn9XPZsNaQ3
vBZPsq7hIc8uZXvZ8Jh5WpweXrisDyeYVzlIlYJ6y0QtatamQdmB6M52ClKD9dlC
5+RtFid5EZaEi1jGajSWHs0ZI+S7Up5v8Hub/fTO0nynElYZ9amNi8oJqjRiEGOw
CAN3xdducaAPiYXeOYElSS/VcbZjse5lePrVNBeYZp1OOKM6HgsmRXi19GWx8yZ5
c1RT2i4LXLzhM7xbgdG9gpaANJR3EotZsyf18Lt03FwdQyCsCp51Hb1/1VpuqhfI
Wxx1pkP0IDhwwWl2UzLVqdAUKo1VQjlbsxDWt3u0Wzxi0RCK+FnL/4pax8fOOg3K
zPvELaIBI4tncQNWjzULNRQtsPfhtMSNPm4C5XiQmSu1O+R6A3kufV0NJBK5aHrN
LJVFl499otJ0Lkx71fhjVbJcoJFt9zutskQFj8iAwlZoaOdNUPRjSM2zp01oSDM8
saZg3N+1Nfu6CrtR92dIsWEPAVgWb15oFar6rq/BMTVYNUI/PStAKW1hun9nuEXD
g9UvSxTAg+lba2wxt8pl6Y+1PijjxW8bbAXtuWLNJKxyVtHLpl2b+olblzUP3WUM
fI40GRVW3uro3zns6ttbSurecfXDzkZKrBtsNPdX9yhSYwsg56sTnfTnWtvfUmYo
/l7DE4pjru38mXft14XutjVuBeZyxjNW1/GAcJJf3IyC+YvfTbVA3sdBcd3VSfFW
ngXlLRAyi3HRP5PCFZ6EpLtquPv33B73YWY3UWXcZRuWnPsIVby8TeWRDROCkGTW
cv6upijvPR/LN9yVxXkFOxUn39obEDXydiB6ZOwC3Bvufp727X4633bORxw3ejhh
xY/e6/AfHQI3bOHeyWgGeIT5GP4Eyxz9CfZKl/uXv2IkwIdaphgDRj+aCykEa926
rHR4/o5sgXwbRah/yxIF8OhQvu0hfID5l+VZXTlFG1hDWs+FEZwR68890lrdmz+c
snty+qJcQoIHYKWGaKw24TpzCYzGiJW50qKXkVC0h5Zmu+1VY/T24XIEPUM8ix5B
YZfXQKVJiuOmvSNH1I1Q9dkW32w/RvyJZcN8QHA/e9/06TD37Phyarqxa215J0Y2
o5WSfizkTl90ityhvftaWIwmKJFBwf1TCcJpQ1yap3IbRJXdtR52gWg8C3WToddO
AgQC0SQ7eAASxq7kw+qD1QKh3tXZU+HAoUmysa/BwXuYlBMoX3IgPuYIuy7i3de0
7P+lTI+15Yju+rbbbgiyn9g78KBnAuwOkcjZWMrqH4oKvVb1kjm2W83FvOoIT8ex
+m6GazVSkP2+FWrSyk1Tv+O7RP/TpM89Teqkpx/2/ggG9igKh+SKfA7t5FSVf8JY
QJ8oEKo3g3N5ibsvKD9jqJuCNFebw+ikEefMGGdq9sLaa0Hdx7vH1/0k+X4pgzkq
u1cgl3EM+8Lu4zUTjoyDrkHf6aEEXdIAlNPDnn0uQxDMHI8Y4YRPn/cbq8GjkfCp
rPoCugu4XfnTcgmXrg7tNmYQg5HK7p04df8001YKcJSYNay3lierY+uLdbFfepAn
qGsU+j0ZPeBJL7eo/lsMxqnVlPy01GQXxYGmJ665sgNSZbN5LdCZHhddq9mib1ID
o/OqhbN4+EsQ78+jG6hMq0pM5BFdQigjLBD5lBYBfwZyej3zp9wbiE4u7hOojXkc
KTfyP2vrlG9ZYVOe5w27K4bASxwqK3gB0DZxC4nQmcRKcBvFhW8ts24R2N3Yjk3r
cuEJDLSl4Fh1Xc1nSHdUBqSqh37oviQEWRk3Shbmnq44Z9FJnM0KgLiYMFw1bVv4
PJPG9s917HAxw4iPt4rT25Sxpofvrv8Hk7OBgxnzTP1uqN6OTi1rdLfvxlUEXs8k
itJvUqMpR2R1jI6bRVzwYi+S45PRjegKuEAVVGjuhaKaXouy9E1ZSZqVQ4fvlKcE
W5JoCTQUOj4E1eGu+ClUWl8A60Qc8X1mCujYtfHEhkJkWm834zDsANPWSUuE3eo2
PlBEIS2YMVUIvDbFiet4dczECgZvInGlpeFy+yxDAbdQh6r6hOFTzK4xfvluIXdJ
v0Edb29O31X3t9hee+v2PdUKGLtuMCfhKlQzcF0g/89fer1U5aFjVAMJWRd04sWT
4ujIceyIsG/AOqvfnZlmbjGg1Yn/aPeIQhXBgjw3WLNSA5L2uInvlLwBzP8c3+KW
e0h9mYDxc4GBY+lvfwyD+dbrN/gPwOq1sb5RTVFLhvwxcUspVKyEuwWDYfgMq6Ju
gjbPb6e4iKa46cihV+NwLS/FhEWsNJgeDr75PKaaTXeLjs/bmGBJ4vgV8hsHve8D
AgmS6pDtMxuVOU0ptiiOW63+AGNuelnZNhAzkhcUXFo1Rtz2p1+V7gF8Z9BI2N+r
Yx7oROTQ7kdgcXPgH1cbHpRLmVKYO3CGjSjSKBED1G5CjnrBbPtmk1bJQ9HClRR8
l35KpERWjYiM9frtnKQcMLnBT/PWvQIQk+Gzy+V+EZbZhkGFjiuGbGCqfisv3L2/
MlskUQx4br++uF2RlfjVXGBRoY5EzsGs5jwsFMY7bVBqV1ZNHTBIX1txiiA6r73S
VPFGmXSmLCPjUxTuQbdd1zVBSfvwBRj7mHy2h5i8mymRJShVcDyVsaO//9BucLHy
NY4V9EFJfJDh4XZwvDtPxP9tgYTqqnCiojnyOYqADcyFKErh1GbYyh9+xEoNjMU5
1gU0JhRg/yoHYXrzsTCOYaWJclNUEWsYwDkCut8CcPWwLvkO9wHu25sG1x7m2Ola
g2SE/l/STgyojrKGdOrR51A4TFZAON7YW/snzJVjThClmWUED65mVJmWWvKh8pTD
aGDbnvpN31qelvDnf3hf+M4CCODGqrrIiellAJJBgGhHan4fqoVOsfw0TMd9jhXF
1g/vnIuHHZOBNq3b2hid6ovXLmsH5tUNotNaNCZzsqJtQAwDqIW/mnXjctwD8EfT
UC3/Zz24anE7YFaSf0o0CCnQQvcZwKaE9qJ+gbHRkJ/Zuv3r1W8BxL8a8O85XuOo
leAi8Upkk8C9uvDuookFZnHAAnuFZWCWzBmCC0vV1ySe3d/UfeKU2o/GvwlF3gyy
UdbwYuft2K1+V3fKOYJplQ4H8GcJ0xoN9sdvtamJ49Z/oCISDlwu/FPN6bq6nfyU
8/43/JG+wD5S3WQMU+l4xKVRoUNHgjR/ogfXafvY/nCQDCtez5J0zxZVnlFUx/E8
I9s3JWxbtaphYFimgnVxzgK4tfClhu1GnOhowbBlWkzjtXmidCQ5nw7JiuFkjpKw
rFrV2pXqiHJuSQ1Nnl0J8le4l01l967IDMxByw6e2X7abA+3uN9kDTAlYKpWz7F+
CgONgXIxTGGKyXXoRvsXfLdOMh63Qbo3dM+5oW9vZ3H6IsXAkez+bV35EzUv5/to
4SRFhbRvMMi3mDJf7Gz9o4yosYwrWs4xTJVaXcdCgR3kszPeEVGA88dcDmHxbD8U
RLkubHJRovg32QG5l61zrUnyyz0QV7uK/q8r+AYbEq+bnnZxunUfvyIwt0Z1aQoM
AphIaxi9gIDvAmxAOWFuHOBhKR/7H7g45CNnEEhQCwV9BC49pA0Fs+domxHfyI+o
7mUqNZtFRZfRe0Nyc74d2Rh2ESPMPzzNQgwwRYhyuV53eR9ph0t11lHNrdlhW550
Fkp1yH2ZHhLiOjZ+dcrFlgFto+uivP7XLiGgd+SUvBjpxCfShChPaImOnL2Xv42d
7qH7tTi2oomwwm+AhE6Br9nxhmSnLaWviMpP3HOAWqASu0MHr88rc/6+Z2Q63pog
tj+0MJydtY5ka4kckGeoTq/1qfmajl1m/gEiApyttNwwYDxWFOWfP2VkzcibRtJX
2f0VEEesDfLdJEe0jWGV/PxpTmemwnlomixAUh7U/S8MD6P1wHMAK8ApqUwp1WrK
MtOOBv9kmjUrHC1pkFOmq3ibDGtEj3LfEjntMXZ305RS4OW1/w9f0wzvLUKlKHE9
DOxwVt7W6kJT8gOyfxxY51igZP0Y7P9/QeLjUy5uP/htg5J6DUkpSgt96HL3PqF6
feWEO8DT2a5tYAIA1J+Hb8abULrmavqvz9f9+53zZvQ6sPuIL02w3Pt10DBqYjjC
T49I3W/omGovpxd6p/9MjXV1WrRkIUC+UEvf6KXDz1JQ5E4wDXnYbDWbXMSjOvER
zjiISF8Kjy7VyTSwCPKhYELg0hdiIx7HhP8B9PK1brmIsGBzE+q6Sl4xZ+Sj1hg7
1lre//hldbo6UTCCFwaI5/Srz0hQzwukMc7KwoGB5UEyTVwtvl630RWS/EhEDG0m
fIWBPc+/IT9tZCOV+h9dq1KLXu7bOU1Sk5yrE3icLJDltlRfSUKyVDwPet+tTMpU
rtX2fX24abjpNkNcJ7p5U3B8D9x2p0PZmIBaTP0sg8sTUqgZm+rKO/l2XysIjDjq
CLzGaB0BY5jr0a/L4+DR713VdSQMIwz4o13lrIHSe/39Do6IGRTPW505K3QWzZI8
M9mCM5XCj3tJW/xCsKlGCD+hijxcWcbwhTuyI4i347lQW/8qpXLB0XKtwkw7ifmp
jUsCpDVEeoE3GOQUZK9E5jbIDSokeEASc4D21YeeFVXE2ZZWYOHBX3MTZB4MIslT
QCZTioUkK4yvPZT3eGGVPK+gn4eiUiSqToUE1i4jvbDEl8CCQFx4v020R9uo+n0y
PTgH17ohiw6xwpl0Xe5pmSbWE4AUfzfz6YgzfBhjChAyEbwkpO2isaeYrQpmwPoY
66bUBq7Q6AcajVFWdilXc7gRrWpYRropp1muAROwt3G9hvhcF1S3rCT8yyhQKE4X
Jgij1KJHNgEec8+dcJslum4ImOZUmOLDcw1Nsp/bCDYiujONraxbfuuEtF0BkT6b
L5maTgYQ36kk0aC345hiFib51tYysqp0uexuIMkR5J7qH2skegVhYav8K2iTh8Jk
eRMbEIDo5H2PBI7Pjv3KRWNynzhMpQJDJD3AsM4hC5uFZ/g3ky6MYjZVUiNOBicx
7aiGtfRmJ3DGRpNq0TmAUgd99zs6eJVY4tYBV2zPUTNqorzKGgBzMY98jD8BB1lR
ub+P7Y0Q5/zgcDK9n9ZeUanu2FMoIEPdvsx1Cgv8692o53F6FhPhNNbQ3NWggySC
7CDq4Apw833y8eebBJTTobhHSF0DuQb7pOBiyAZXlXqezFsVt+eXXG4EI0FIiand
cpJkbQEE+va4j+kEbsjv9ZmvpYX0Tm4DnNKoWxN1aBNN3wSERuWmKlCsqQ/lJEHG
s6o4ealHJNqj8reLVD/4fKNhT1UZ1UTPnhI4d0htnea97eHtQ7p/6wtfsUHjmuuT
niWXtc2Vu9AyIMK9vPQ1xBrBFWed1FUVhwZg+JzegQy5W99S+S2tycg3rd5IkqCX
9BPukT3STpRR4A7qAkVYU7dA7PfQIWYDGuTFgGCvLlm7JIzOev7sW2WwIVLEEzb9
Fnosm9aTVwlhMhAlbR6PcOqF0BDiZoObHfBYU2P/Ss/J35aJDkCe3vqpeS5bMQxZ
kAXlis9YbMs2jzt+UsgCZSIpnDF9hScUHk9qKbxEsxOyAPQVnbUW0ZyWKXg4oyrm
IHWjp4Mg4zEy5VbNQbmeW66LT9VPq9GQPT67uJ2J0klKDaaePmfuz5ccn+0PMsdT
0juT11FGcJZG9N/4UZeJ6vhnEdpnsJfH2jHCaxiAhOCerTW0qm5Q17ODgo5TVzK6
3m76Q1yRUHrhYYNkNVtq2ECYiSZFv0sMwzI9pyD4hjmT/c/YHDxj68uXxCJPUv+r
3vy0Ug12EAI+We9vDCXSHe5KYgbXD/JpwqY8C4mW1VyMo5Sa2kinB1Xh6i18iIvJ
ZzYomhVnz8S/SutxP63DAoejrcb5RTKETwLyW9u0jHDwgCoJpMPQw6U3JiHskrI2
HpeAwvnLbi7U35kEA31iu76g+TZHqxyKEyGg3izAiouFtqJk5B2K0B7ucdfwbX21
JBp5uF0yavuOSitFy1NohUmMuIRl8KGdN/2n4QG7UtOKqzFEPdBlb3hEJg/SgyQc
EqqRsTsq9cRv2Fcp2bstXdfvk//99gC32K5tPSOdmOX3wyrDK/4fmkXqPH5ZPZ4Y
jRAzIOiyzyx6WJXiWuMO6OysyT3npGEIddSW3FV2ZOYZ/5zQTxcYvzMAmWUntZPz
szbRhJVIRFJJoDu7s4/AzRpwvnTm+tAVpCcFJIyg7FpFDBRjfuiPwugmP1ZdDVGM
OMDRx7egAGrbQJNLngAKiUPryR+3e9n7qgC/t9YSxJMS+zLTElA1x45ohz8O5o2T
zab6ZT7i2FYlexxOqa0fEbDvA7DkHyM2TzAH+O9UxyIehJ0A3pnE3QkWkF4CwLwu
KWwTHxRJgzuPBMEkop0bD26wkRR5Uj9cr3l0AqMUdkzifVErkK+fOigumbCHXj+b
uxaWSuUyus0QEd+pYeqYUzrQRKBS8W4JzfnWp8WCjseRyG2kdvsYAzY3vcH4gT7N
brixlVI6GpKI5E5gBxbzvqQjU/GiWhHQ+cXt8HCZWTKwibgkDv03X7Z8YLWA5cFG
lWJxbTxf2bzTplLjH+N/O36C3Rt9lFh5jmmQB0p1skWCaOoM+2ceV1ZESKKyWxCZ
Ntet2LZzSfPefxXttrjZtUogTPMGivKyPfyA4gcR9xsEkfbs+Yvj94mKdkczeLJA
pnK9PVRZlXodgSjOf/oGWcKf0ZCodwvhMkazS+8Ud0ZFKIo8ZocmwIysq+gQNDtb
L3QuWGCbJMxYQ7VCkpZEDXLyvW6zAFY/UKM/dXfx3NBkaGtoqsWjXRTDhhqAIzaM
dRon4QwksTt/fKM5S6xWdmhzKvebSoTISjZnYxFb15ErbQZGPE4tgGQ37DbK0kh1
bmGMLgKSH77/QkniWsDKlS39ehPuFXQwTS0LzwBIcCBORfFGpyThtg1qkWSGqXiH
Kd58K6AssG+fvI8lCWRCvtf/tW3iXp1OCKFxRfbOqSNfgB0Yiyqz2da6ukI3xRst
6wiWq+Mvnw846DovrcfewgF6d435Pkis1IafTGwA13isnlgVi4NX3pKMhHcs9ON9
vpf8+fcBSGmWwm9IRa+J9ljNQSpbPkU4o+xwkyJ9daqZyKL67/AnUaL/+XmfI3eX
wHrcI9VpVSGudyv+25SnmAiULrY+fxBd4w1+xacCGfFG8+hNP1lB/WtDul1a0ZAg
dh9LtJg4Hhd9aZl3qv+O5ix3ZugQ26LWAYlYHYaYQo4g3e4V/zKVZMPjVLKoVNXN
0O0QL39D/nSczCshS4WVIaRaaUslfxHgO40aOT1TIxsTolsCfWjahyNkvQANpi5b
Z3BboW++GcmeQBCS7K5wueYd2jjR4C0Bg9oc4agiLQJhVzke5fjAjhSiZdsWTC/S
jSFNrbmOMOtSoFKwiepVw02Xpc0iRjbfuWtfJWtDLRMtlbmY9hfQcIiwEUa/M0Gq
zfXONZQZCa0v5lHeDfqVXeBugrzGfP3/KS8BJ6Q/hvwJVEdvImxKsWXlnphtDiT2
JEMax5sX4NMpox268l5f9ZyhQqmnuqpv525ZDPtRxT7GMbixdTvmwC0j5DvMqryQ
/m5OML8pKKTsXSzJhAOwesnpym6bDa5wmxCrntZOo4SSuao7DGHUDcgoTrWY55ML
k3mR+g/l0IPTE38Rwcuvy4Zu0VYYfFOCDrd3ViLXZbpzramnBPXDtvGLVWwHGKcg
/4tX8GVpZfAnf/Xh3LOUG4GsGBbyEql0njQLWrN1fD4ZVkKQYZEZQTe08IcEyAvY
pRApNxVwQZrdDqdo2OX56Pw9ldlR1czhvL1SsucrS+7ZwoLDJvYZsG1/myMRzazZ
P0jAgsYrJSLg9PZyvIPDy81vunHYHysCGnsL2M8ewNYD2WGPOOHaoWfYIEvc+thR
mTABaX7O9u4cyzjlbwC8o4QRwTP6W0ta8vB+BxDN7KRUBKauxnL9E54pf+ZId8rn
pQiT8ZeD6rXpofUizWnqoh7H74Nb5tFiUHVwZwzO62gS+G4jAClidre6aZjEVnUG
6I6Sbc+g4oU4s9QeXJLk5J9h+71TfFrZQhjVTfK/h8KGAZNJ+rUyPnAxN3SNxJu8
juEO4mhqZ18KtAtZd1wGTG5+ZB/Bmyu8Kw/u6YkCaPze7FJdyjep++zONvF3l6iz
nCoun7WP24H5Z3BGelUUNLkg03G4kqezLTIalD23rtWn4bF9IWfZpW4DO0j+z1kq
pyb9Vqbb9LghoNUL1OsLH/OhaeHasxc+75sTlEterOzWQ7O/3P70rSdtX2IoVgZm
rV/3bzqn4VZ0nRRwU3Go6kcawPTKuDfcKHGWikwDieGOd94FAX7P1X2HWPwN+sjL
URHJYlPwP/QGug+zpcHfdmU0HJa++NIFcaPrTmGHg5nTd7D4C89BwpUVYvxnPIVU
MAGisdvgkXb9BwRxjoF0BZScSw71Ur3BSaptFlnfVst4TcC2J9VysYo09bXPCEBy
5mfVLbUP0nKH/Jvl6kzgbMpWVUQ3CEKeZfspIPGQmPp0kllssweJjPds10f9itWA
Sf9B9JVq8GVQ842w06/EmxSJRL+M8Nl9A2grzphPOorjZJjVMMo5m/VaDEoh5mVo
ZyEV4JpmEWMV8kca9KxrSZdQEIwwV77I2tTmfr+rgjw8V0k7Kwrtvk9n0N86nbi4
jt4c22G3PXdxTtn7y1mmNadOqm+dUxXexlvCgF4Ana4yn1cY0S+mEpsBUNuXG2di
Z5h/ea6TPcZe0a3RH4M57qC3n/XORHMAMUW6UOrtA6vjkqz4DsZVGKzzMsbkAam5
P16/T3O9RJ3UNgQD1Dc3m6C/IE4EVjp4KlEAGk1ixK6orle/xtPf49jid9pzRnEn
Gug+pSgn808B1rTjmylRHaGMz7FXEAir3GCcZCgrrEEtEER29oRil8Xpo8QsbkMq
cxcTBJAhdnMC8YM4hA7+3j3iLAe8hz8enD2tpZ2ejbbhsv0oAiLtJQcDkYHfeWv3
YI8K3QnGW0Z71VvF0AsPVaTDA8RNMgWuzNS/4gE82DrsitrcK++XCdaBUeYieEsE
nQcK3djeDdk/r2LQ/vcjMm38CmDdt5UEQTPem2mgnHUDzPYXyQVRJz4yy6RvZDH+
1shohhF8pj/Cv5+rdsRo+wcwGgqaMW94zDh8uL/ahDqM2mXsBHtHfcM1oqqiog6R
/BKkvPZF6hD570Wh2229WuGJsI0IJxePniIqLWgb/e70T7Df7kneKgE/gSPEXEyh
6aVK90fCHVUmI8L5SWB6Wa46ujiX99T2pJ8gfN3yyXhYdEXVUVVNPFvIE708LT5S
k+PpZv9QLXQ6vHBe4DVhJkz1or2sQqkuqGYlgBTQOxgIFJWMurOFddIzoyKsn95l
z8x3+QkA1FJumGl7VnzrmL7i7VS11tfqj0qvrTU1iN+J8oUIBCJWMq3Vch6YW+Fu
ThOluiVYYbu7ngixIdSxDXC5fl9z6EsFUSAVA28huqb9FBL06DEsMsh+JsUgFviQ
98XZ847+Ex1DMcgAzM9RorrwPAoWTqIDV1rNrzSiM7aWJ5/Tcuc8Qd672+cUNxJY
Ug/evb4xMKXW82p2m+wWuB5QknfnyUDYxl/hzUvU/KoK5+5J9Cw+xSsG7jsWaJPb
CzsR3zmkWQb6SfygNwezyF5Bg3lAikcm8xFxtrZfihnM/sFl+WKJxPHuBqiPDgF6
l3a5d62iC5xqylr3XjfxoDNcydnpo78s+0noAkgcyf2+N3mqjKZHm+ylbHOvi+pi
tQTK5eR7UFrb0obty+3I6uVpA45ff9ZUjLyUxY3EXbmPaC1OceLFuO2Ag7Uxds9+
HjTb7agw3L6gAmq7FxEBYnuptqRiCe2kXWB2/iecZ9v4v2gi7ptsUwPuAmh+Poki
AAEUdMNDkqEdtqzMHtK1itqNNdSAqUaK9U/khR4V29CNSqRIMN/vYuEYDKPGsCXo
q1lcTJAA+ddNQ5BIHmB+Ibm1OUkxa06hJD9A+DEdGeZIRt1hJATGYND/zOd0fTpI
x4wgeK5kFt0qGRn5eHe7JCnqEFTxjZuhhdHsKAygVp6K1JnNv7JpKbfMydCpAG3N
LZ0iXI4QklEt8zESJunxta6oIttWL8UVfv+BOinD2uQz9x8T9jUH9wz86WLiIyu9
lanT/0Mx3vAenbBuTHzhKWusXIoEg8xQ5mDuM4pif4N//LUB75ANwh23KNMFqv8Y
6GjBl3NHWAZer13lSM7HlhhnTYjPbWFS2aoxHCVNLv2eQhQaK/qYmyv5+Toud4PK
TS8wdtbtyeK5eRMDIha+vxiD9zg0oKRqGZrzeiojszIqq4t2J0jH/R2261mPXKQa
7sskqRzSbACExC6Uw0my20vfFeTAG9ZxEcIhG6bFAv9JbX7pGJoW2ZMkKBqNmvWW
qg6mPK5YPhFC3ZqLaVJpK2+xf3WCNi3PdOrKeeICOmsxjUoSvQYBnvYyBXt+Ypjc
YVWn8no4wBQZOEVCtrR839BBiXdU7ndFH9h8t/rty5qWBMhAJqvrWhldeyXp57eG
GqoZSnRXHsV54y43gDcQvuoTlPpvZI26YZ2D24lv5kMxIYpqE5Xxir/a54KjgEKc
xnilMraeVxcQC73cQ6g1PIa67zak7QjbdNGehuBd5zIaWV0Em2V4zrUctkH6dfOC
++JvT9tQART//+J2ZAZX7jDt1djA4g9iasCPrDUg7vh2Yz3YRz2J+gPsBHPoRH+S
7krgW8CcHuzNtp+WPUJYXC8Nqu8rDcOMOXbST5Y25qD6UC7Ew1b9vpjfhXrL+Q3p
sjn6NwCC7m82tqE+h3rQ4qX7zyiWH60bC9e2+/FqwE040NNIquOUORTp+5qbbc0+
cCJD2VayuEKvXIAnYVapXS1GlJHgnibaunMFkv/vyHjyje2Hb9j8oNq99+gMuWfP
JtejiumwTGl3L8vfh8ONZNFkMSwVALrr4Bj7xLWZAP36C+fSI7D65xWSeoMo10Pb
jYfqRK+MOAs+4iueVNLpIJoH1x1CKFFzTgM8nO/w2HDaaVb31y8S93MG0nP3BiCf
xdnaj3/ZLkw6ltZoywLp5oCxDxR/3NbnaTE9ukrk3lM0rKxIEDgFmwHfU0LsJy4p
4oCf57c9WWOHiL3TQKVZA/aN9o7OJ6z9Kb5F2wqAOQZHXRzXiHe0cwAKdJ2ZkYMU
hvK171+NlpL4JDPf28cpB5O/vP8BueGxNmTAqrXhW9q5FP7h4l0fW+6GjPSQYsMh
DzNIXCMXP0P3iPWqXAGcZ+hrVqLle/LZeeS+kvUqUautjmoSnKdfmCyvmruTxVH9
5JfpiTZWciVxVKDdo5F1+0hBeAJu4InZ2HGxL/vGxzVDYFBySGmEYQW1k4n6LfgU
hNftpPumVva+23CO2dkAZTqppPFACaiZjlgfTnwxBF+FIHrDRRrxz0kE54DZpZqp
567Fz4sXDrXhmsCv7PXxZGH4zI5RL3b1s22bCFQs7w3UbCGIKAVHinkGhhEf/d/E
rkYsn8ZKWsoTPuha+pDiEYyHKxFexQZVL5x0FpvD+z7ZZUiHxIxp1SmUzzBfdIJg
3EJhFht4vaagJUP+KHKhJo53B3z+UhZEyfJfFPHy2ujA0vYvScU2dc74sQL0Yk00
lsUvJmk0sqy9mw4ibBZ37M+Qjhmdm1pCMMVRNeVIYGelzUUYo2SZGYY+nOP883zl
HtjiQ+1tFK/vuavfRNbrT0daA22P8Aeg9raIfVSG29vj6LQXWVxs/q5PTpA6VTFg
zjsqkTR+21uQqUUitXHG0yQ4gy8OXsthacPIBH1JSVMwStaWYixZfHSt5NdyBqBb
jOjcmHR9p1uhxvc++fM/EQImvr2nbMHF2jG0BQcXiKqgBXAftGUl/b+G+8mgSKlC
8AAf1fC17mUz6Chuxt700UhtuYkj1pvaC/Chugkl1K32jomlV3pkIx83q7qZ3Dog
59BI5SQzCvSw6O9AtXsKTUMerVhw0nb2/YUkcBipatihSWfiPG1xzh3vJQa/rjGS
lf87FLu8gGn7oWbfOcerCs4lT26asKILD/+1yrEtI8cwbP8hLADlL49917Wkv8dd
4ypEfv3k2BkSrxsb9Io37bcOYVBQcV4RNqguSg6VFsCKjTp95boXT4NdNtuiOnZx
SQtpQQfx2sA1OWX96dq3zYmflg/lMZPr2yEzna0JuqoXLjWW8ggVHkzIjqvYgRYf
FBWn3811knqNhKqIu6xrPKyWog9z1zjvFqmTuvIanJtwBrfDQjG7W/bk5lja8l+P
QY+vWFH1aZeGPaG6GLlSeX7z2tdhY3+jO1dTrYl1O60yKTfXkNy6+vbSkOX9t7cc
wPY7x7+URhV7XuteRPTvuv3JBAPStbCbIeUAl1A60phyWadxNwXVpWiGCEcDa7Cn
KNhfWlF/FF0PLQkop3JC5dhcCxcWVX0Zt+3cNlUrUg2Vwka+i/OJwemawxTnN0Yi
pojR42CcGYEXv2Bm6A6iByajcKDlyf4ZLdbz7q+gvvffwgosB4kegF/YAGFJNu6D
NkcNoETXa/byIYCB/xAdAXvdschz85MiJNb0ncpWwMZhE3NXYA6ooJ8DlPYjLW/r
WF0vDkjw4xFQlsZ4wMzVc4LepkV/Nmp73xjvBAEV6Wiv0fyNPqOp/q0x0t73uvvH
fmr/egm4jtBFd3sbr9wmMrfwmmy9w9n1VFiFtgWur8EX4xrVdX3MDwhk26aY6UJ0
b/HCKwqnOuhGbyZYDrC4fspOGpw0uw9thWFH3o9M82DLgwz22d1wa7m7zHVIgfY+
JAQTDcKFlg4UbJgukxT45p/Ix3nr0pevjA6p4p8PDvz8XBXC8R+WHDDvMfFnn95E
KHhMDddpL+xdq0oQDv+MiZfNp0B456gC9wZnNyqp+75+awLTiwc/lC5y+H+zLTWD
YHcxio00pZ2qs8dPasYhtFpDMuWfMmEIHAzusBgSQZlTz8fkexO9WuyUXs5pU2BS
cI+zD/kEZpNLxI1NF536Z3bl8GbOXF1iE5y60mfZX8lf8T4xV8FNsQqqCfTUgNnz
/0ARiiBdRJSePrDeLCA9rI9uZKFnkeYOGriglUxHmqEKZnJU6uP+ffqQLiE3DjW7
tvliNqB6EOYpUmVsQS4/gPtdd2yGHcEBgnHMu/E3PKIr6GhmoXoYXqP1z3rNeC97
qT07LM0YKBWIG8h1w7NMCIfGUgWr0rcdX9L67FrJB3AfD7wGRHOMeWTr+iiJwRAR
IVuACx69xnreV90Ixb99ZkMOn//qaO4zHLeQqCb4v9oSGbAzvu1XySwifJNqlAMC
Vi2TDhKYWzyG4OQ7qmlOZ0WtrOIfjuOhijFoGFMD25OTyHUcJv3gz4t8BOF215OC
NMHS5lz8CQBt8MCgQehsNiB8umhWyniQRCgXkROGIuneaQrrKAV/pz0F21JzcHhI
pn7+LrQSHbZ5UaJ9lMAS6pwJ27W04bS2grzXhH/at7cjw1S037stPOj4cpk/D1Q/
0uTLw/LMx4/5+Hq10RfdY83PmC7VXyFg7GDW9bl23c5xagVAG9tqxIJb6KiBl96T
zf9CRXYhYeEgNcX8VVVOa09pEDeFt2/LHatRL6UkZnOTwLDT4EiJqakgvgMqk+Qd
wDG+jEWTNe8srC7nE6L8TSED3OgqkeNkwW3KtUVXXZiy6s9UtG3iO9BhDFYa2RUC
wOEUrgOJCY7LGH1K3dglU/3Nh0yAReBy+63XnBersBzhlZlxqHvwvhoilACJjogX
EKEFaTU5y3nVkgLQ3W7Dp8Cp55RjZPu1+PyxV2851rTpBROngXP+ZmyICYO24JuT
0H3Uvzvsh/ZT4Ahmnx7OThPYZ8YQFyEi72Yj4lIWONg2CzXP6bXAU1B0d2LcEnnL
HHQ0KtpUz8kONVic3eNZyff9z24bkGYFNAbXwic0lT9YmbHjOaHyeolDxvzrdY85
wPJAsvJG6UKypLn6HFPDAivNzudf8dkmnaKPBCl39YhS4pxN0VqSm8pfN6e2ggq+
en/qcrDilJ13qL1/uW60J+Rp7KRG/XnK8w3KWBgE1e3X0SYoI1Lnc4A5472GumvQ
iLzmomfl+NZpjkPhLCtMDtVw6wJkVhw4Zpok1ZuUxlULJpZ/wHqBb2ASBJadyeFF
WERs7czfN9FGxM4AmvD6ZB82oic1+odfGqK6SOmOURpXRck13YKSxD50Q6vFKyWu
nJ1RBrK8DD7q03RzmIB/HEJIsgB7YFlCRGZ3W2shlrQqDPvDrjDlwK0HZzEiSJFK
tTOZNn6GuRsmiQhFJN/sOeAwwxeBG6PVoz/jEMeKMt/oECV0/BbSVPl7cuqzWWEJ
waVcF7OSio5Q4diU2wvHzqO+4QyrjKiEELVMDCzDC4yttAzI565sCC32LcvOS1Kl
y5UJXjHGqFJ236InpiqW3zvkQdoQR/3wNKAC9L7PkAkxj6JC8IB6m58CYVR1DlPh
W7YpQrlhLmtwsMntLk+K9q7fwGGicIod8lHhkaPwqdBgZRvhhB7FpfOQk4fLL+gs
ZvCmdNh4oLEHk/uTRXYZNZdTHnbImmRgawanwoQC458eHEoyXe9v/FZWnveAyhkK
05Js2VaJ6DtqomtLci+sijwfWc4DaABUVP98rotaHLzG4YczaWup1gNb0UjofOdO
MvDTzexv4woFvG9HX0SwhGmTPaEEx0jumJPIWoDXfyjg5jB1yXaG22qjF214D06A
JUNW6/vc35NAJp/ydhfyDByots3oRAEpXWYDbw64wtJZNkWjakxwppZKm2d2TF6F
sE0lSOvLKiU++zvFh8zYQ6m8I9vzU6f6LSJrJURXirCrgdf06wI/14WjQRmmiaPq
xfYSMAFvjLXverpNQoa1n1+qYScXVNu3T2yA8okKtOoN9xN2sqB0CYtciydyvlBz
NYah1ImDFJGrpF83qFE0tetzxYrt8+VBMb04+JYKHcHu0euoQU6WprNb2m4iTnBL
EgPMCTfVI/skDkC7cGLVqeqpPIqAozGvO3SwIAxP85Bm023bUACAFAXQ24G09/mR
nkuk/cahVYvJmaBWRx4uZmP+D3IR2g8yyfImnYnLy2YZZRRsh/NvWoel2IjI0tr1
Hgu7G3EqY8/LT0mZo3HWCaUxvvCi/EspGggdNjQTEKjCWU/y/S8qOYJGrzEPKHpL
TG6nRuSlaLXWqf7WgMZCshFgf7uQICwJJff2odItBsV3jOntXDOCaGwpyZhAgP5V
DQmlMPy++XgI1yU5GZuOLmyqVecO8iixEH3qCyekIDAnUrtOfGZtDFKxB+G+JUug
Pit64JpjPOh74ufuaZpGG2qxiEaCsq4g6k8NIMyo8/UK8yD4BugkgZjMrTzLvCw7
1JEYQPvmeYpWRZNugdoKsGuPDETF5FchxKPZYgkJpMTY8Hj5fTJ0gtfAa+8tysA4
nWBRwcvqDLhjOZWBdkDjAq+FXkYLEofBp684Pr51IEUpTnLgFugKpoiJ0/umIQQW
iqKKmlz7y9/cYEH/L/ObK6oCIGEGd/2HfXpIzskrfIy+S0Gzts+f7o4eaXCeAMD0
++TbSeq/Cn8LSmv0sG32MeVPMBV1nAoumsl/EVCO6cDn38+Edr0ewxW+Q+iW5KVE
i8J+TXt0IB4ISuuoegfn2+l15qL4Su/P1lX87R2/M/phzYBb8mPNiyFpTnWvKd+Z
XYGYRsBjETH7e41VzPMwtRyq4AQRB2C8SIWYFBcHNa6DIFl7e1RHrrJ08zbJiASC
7CFPvwPrbOn1gVYkEiE5gGTIsMcot5SCxo1YMpzZf7vG0UkqriSzodxiEX1XHCFa
61k5VR4XgritpNyiqyXGzRn0rbssnZI8NFF7Q0fRMqNfpOIG0SU7IA98a5vWZt6Y
Os0MlDEFjGsRkLP+jFn6D9jNd4SZ8Q7gH0QR0VyiJv0HHPu2cAZ3+x8sv1mOybNv
nxn/KxDQeNawVAIOMYvN/inqOAy7xjb4PQQ4o9e3f+nMnlOKgh10mx/iXW5BtD0L
5WclysNc7DBSJmDdN3WNg/rG58cPFHuIbzAX24f5fiuIT9+dQWJ/YHKO0/F/P/QU
s8P+VmtLOytDik3r+HI94fQV2MTdYpgAQMHP66WVG/74FfzweQFbIIMymbbcHef1
HOyLGRWIRZgvVcLjXTcbnrDXXtHqfBmAYW0XXbyP1GIINTLZO6pOJEvau9PJuZY7
Kw3bDhKkfREB4lyXN1DOtI48R9WZaRl/dephbBrszAwLlrB4jH+Vjm4rX8EyjBVT
HRZGV0Bp5IappfF0FthBMt7sfqHk2M6ACoxVUWIG9ODkX1zqAZI3DFoH4heXMaUV
Iy0G8NUqHWFNZQgRnfKUobIkYKz2kCHj2t/k3nMaPOzOnl4P4c7i4+VI8GazV1Oy
nBjHkQCifx/Lsh0Nl2bbpxyPVcXKsm3IJTcjejMeN2j/8/2kCmVRWE2SbLxz1AwV
XrDl73kpO62FTR27h0msiSv8ecTBgqkMgOooB8nOSWxJKR/PH+iveQbpMHzQiFmN
G+9XwDCaz1ZUmUFKcVKwmyF2ft7Jh2k53fJ5BcGRr0EkSSRhAjxXWOq3wjXZXSM3
gaX3+p9cbsApLFzY553ip2HE39fs08vBF0o0n6+AOvpv0tvDzvlUlXCuZzxpbKzP
3XUlj9klPRGb3YFm2aNx01d/BjYDm/9HrSYXx7XNUSJv1HKvL0EuEK6pfIadLyJH
gBB9J6ml/fNBsB+ZiSgsY+ByuWhsaITgmQc0iSlkKB/Mebywxy/XCAmz70paIOOw
uiYVn8gKTaUF4dE0x7ZmMlLtVNVVlqD5VVXKC9ceFJC+P+srSdKf0M/Pyyove8/p
S5L8bv4Dmz75+jV4OW3Lpo8ZtJ8MFzKEZa/MlygyzDapnJQiOTo7UOa7/GmmN7+0
Q4SNX9w3VfUgajLGMcjSLdRtgUCmCYouBAWrEguAA1w+Tr378GeDGpiaJHolUIDn
ZmgS20gAP2cY1OQ93BJRF7F5YEwvsjJU8znTRs0AHShtvvhb22QB4vroZ+p16VQq
yRNz7rwAt+b/6p+idjMrQ6yBD+dUN8nO1YJ4X3hkAYPXFLoghgIPZUPgiTG6p3uF
hKTDJ3fnlbUpqOreHCtuziRjbM+/mCVahAHsAsk33gA4UHd7/TvnTGaU6/Yk4zxv
BxY8ekb4WDfvSQOseGfdYZMQG605l5KAZ+iTy5rRTC3mmfceYNznKMs3F+cubPcR
L4LbXR36IhV3Y+RjS8vgrPOplNDSb3rRbXkzeI5Xx909VT4JRWMvOEraC10Haf+1
tAjTfF1pqGaouz5T3tuyOWrOwjI3xC6nozEyq8Evz/El6hiyONHkVYS70LwaUvHc
vPrDYd81apNFcnNM/4RbMtGzIHVcWdEjrGjSrkzod+6BBJ0n4x/GIzv5k/S0/1Nf
067dzvuRoaOnQ0nHs94bKiR9TKjgIb4NhVYovgjetXu+zB198EQuX4vxwrY4QkH0
2IfGvV/Qmzg7OfBvaLGWn4/E/F09BxWazjQKIpaYn2uVFCrFWJjXXwoXNmkKsXJk
IJ3Tps9kbvOoW1S7dxhdHLz1T0pegJOOyUG4afT0vNztcMHkUuyiH/ud1tkt7jqe
GjsW73IA2QmDFXg6gaTl8F7nDusOB8m6i+go7t8AXzAHFoMXkFvPnDQgZuKXCyRu
q7+/m3vBsFVbjZg0fXIJtiWcSPddb+JVs59ogz6U+e9o1slaLXlPjZZHaPYzD2ZW
IaPLLDsy+bcNImRjqJuFMWhKpbNfDOIiDEFKu10p5gDrL4RbaICNk/AQP5JYTcQI
WdQIl1rlOYDfExqwMvItk+ymGIPaF3Pzu+M8DCARNu/kSZaiOnDGtF6FTw9WKgE3
9YqlqvXItFGkVNi+fmBPB7EcuGuPZOLBxPkK9GFQFlZsHcNYbtpaMRysRqhft9+Y
ynq1cHrdtF2Fkuhki4FXfXqHTYkdJt3y8YyhWXgQl1/D1zmUBXHZEZdBPHT+Ki9r
sPGEKkUSNxOhYXDFNs6vzafE8jz2hQimlmWCVbEphXJFiejJ2iK6/EiKTHgN8zlt
FeQZ+59O/TtZ38vqH7ofXIjY9bLy2F97POJQJUSzrbdsl9WVrReoNmo49NkI3ykv
kFD+31mVRmeZFYzkDu2mU3W35K5SdvUVfm/GWuII6/MiHEehWDCzPDnVWLPQVI8d
OESHunrP/UnXwkpqhT8OyclIUbC5NBsnCk67OcwRWjJoWQGi/6f8VAv47UyiGUoX
MJ5ModHvV5Nyzph4DlNaarOYxEEkCfC5Ii7iierVQbSjpWoGrcYfkXegvnFgHeOm
g9Uq83DQxywGs3jwpfMOBpAvy4ZaBoAzj4JHGWT4exXVmxPV5ybVeBaEu2/pNhch
TsQMuUFmI5beuB8+CvbVmhTGi97vwRz9nidORqjHaVU9jhmbv17eEWFGxkVHL28+
x3PR0tRr1JAplS5H/C1fJ5vZVd4bX8HObHUkdfkMg7LxwTsytHQoqnJIPCOoRvek
QgTIX+31Kw3yhQw1WHiJACiKShV4aoTQY/Ay6u9IUAIWt0V5NepdrsGI/UmndexU
sMImoAgqODLPayxuNVlxa6E+uJfAaWeINDll12dpE5oRvfEDLf151C9SUwGGE4m2
MnOwu5wJTzQRvZbLOS5BZsXi4/NtPCcJMm30h5mH/0KQahpdASnIr+R3V/WTCCSX
HBc/noUslUAjxLYwt2vPKtGSOrQUn9Bs6U9UAkYxtyo63ycOSgLlvhTdv548T+hV
9WZaFNzRctHinlwJ3J1KHeuVxA7l9SR9AZYQcE98zuwuOeOMGkK9wzkAc4LJU/nT
iz0V3du/BHBHqMc/m4l6JZEAqWqL3TvKYwAeqfdNiVfwEH3hMEjnUdIR13k8pahS
BMOZTgP63AQzRTT+AoKWFvQYXAVB5lw6pUbLlCRtdUJAISJV5mefGwU3AwUKYHjL
Jm2oCThl2mJN8CHOeivWG7yIfwcbZnUYVlHIuOnwvwekG6sj5AplZYIIm58TDSbj
dPdzh4aTR94ojq+0FbaPBvkt+H6zw+k+Bt5AprQTBw1vKFDPsnxaOZUZLf9FqcW7
R+vng9MJwCpfl2W5jSOlZEE4RVIu21oZhI7FT8btVJZ6DRitOEuFJZiqLo3s0Tw8
tnOtDOSPvX3y9aU47nGvR0vJhqIeaoxYwMJLJq8Ajvg1UdNBA3D2RLVNZl8ojxot
Zw09998sWTQALLHwnxYhFPZNkXKyltjQVr+Xt4+r/NX7WrZE6ImZoSpFt0tCNjn9
bhjXHbuXFSeHq/qv5bC2eGpo3wyuS7V/e9lmULb/M3DZc1pqOkYcP/qdivsqG708
9tDJk+r9hkBf7OGUcEvKgtwQjCaWqqQJccCzWv9u35hwt0I3dLqZwr+7et0/EoDA
V8G3+lZwbZV6GirgSWVle4QXbI0uQiDPadQAj51R7PjTf7EdA6ZuwV+Fr/ZALT82
21RAjFV5jus8OnvyxHeypDmLUTd71k7/Vn1F+ryLsQd3hOY644oE877EG9CAL/yi
dph4wkp/M6FYEwNaQ0n2zZ37mfvLLidl3eyn9qXEw1E6dAr9FasMKSXzUvWC/JGh
9FiUsvUU6E3/CsOUpY6tYzbrTYaUknYFMBap4iI9hQvj4C+u5U8wLcypEXomy6Ry
rmGAB4Wp0gcksYjkJVFNg+2aOEm37DaTn8j6robRMZv0cT/FIxvJoE0LKUgD5pE3
v3MhDu5EH2UYeUhaGC0awsinlxlpSQndtSad5BL8l9cOGU8LPUMcULzd93eo+UMQ
lWoqiahlGav3eGQSF5/pTX4LEJUo9Gi3jfQaXB38BH4/7I6k6lxnJGRQPF+W02V0
MP9xAIoReBUO13/sN8Jv/SKn+W+7gWshviBRJzVrkMwjL4eWWXgaeQnjw0q5g8/U
6PwaVmSgU1b+TCaLQBExWjYW5n0jObsFXwMVh4wSIqn3kqZ7CkjcSHkTAUkRWJEA
bmH/uU0HH5Th9b40ToR1+IH7NdbYtWEmgh9lTQhzoqRxgbhROxPw1Dx/GFM2cd5d
oF5V031mLgU78CIWArf6MXDWv9nMXLiVBA2SPh3bkEInJhaJCY3Tae2sRgwbVTBq
L8iiEmsxvzNQywCyBfZ9ri7U6p3WyTtZE2zbcRHW08paguZt6X5p0FzutAC+rH7D
DhmzlaacA43YseKNu4aT9C9tsNIFZ8Tj/aMd8LghznuD1Y+WS8qiKtx/voOG0bi6
dbYAuaPHNs1yL7kBM1n2hABHhwxrzn/qNxgXjDA55bJ8qkkNAhwe5M+S/phk1lv4
Nqji0ir+Gv13OFmn2RDZSGrDazfEN/9fpUjhs+3VlzsCzb0tzt4g7RuEV6DcHTzA
b1H4z/gVCg3of6rzGaYgr4yi1YQxK5ISvvFYD7Q+hnEba+OxQruw2y3b0tCnIwZ4
R7qtKfJPvMxQ4/oxzfMPkGIWUr9lGDLZRCNv1U4okbwkR0Y0gNpO8j/hLdXZui20
CO7dbpOoj/XJ+vTf6d0Bhlw61uOyfdzTSZ7NSDBKFCIgv3+g9yMnblqX+lwtC29+
PuKZN1ssv/aOhIUKC4C9pQzPjVI119drgiqAbwZ1QL4uUgGwhRy3yunnQumQTSYO
7ynSqZACUCvT+D56SOTZaehb1kqf+urC8vJ0ScUndNxuDJ14gIH5N0hdaHALJpCZ
nMFhG82JqSrthmEV2yP7xjHgB4EYgYlKba8y5TqspThCqcdHVR66a0MAZGIY1pQA
tE1aWrQhZOCzGG1MN0GXMRzPSbZji0rGgG/qp2zpeSBmJnyEbM7TTcD69R3D5JGy
3kiTJAmoYNVmNjBDCiIj899FYtzLjfFoCDTEJcWaWT0Ni9vPPmgSW+MW9ed8n8+T
WRlBCEfsb3OMkX9uKazUMl4GN5mvo5HUtIKWOqmimWaxUY1vP5VDgS+YYHlWw+Na
6BghYk3dopZDZPLwSV/t6DgUfh6uSkDnF0T6xvFFfbpltoHkZ1ID0vhhiVm4yfB4
l/Xi+hWIp1fd7iYCBM9MOIDYCYH7z9EJWjrudrnERveT+KJGlIUHCnft075TJjmD
5xwb2dzbLBOh0Qov9yh/w9088dGqniaeUA8oNPOm1RNLQnQ6TFlrKDexWmplTNPs
zS0xYh7OVuOS4X+rEnpjPl+cCelrPYus4w1lWhY/ZOjlhidTRgfj7vji9npKilAo
yzsc2xk7u86BTV/YvrWVlY8UyPNQW/1nI7ZWt8ui2D/RQzNTnxnOFNTYHmRwiOsO
lhU6U0wdrVolZ3cyY9UUG5tnz1vAa2BIGFMIoPjGK1wHqigyxQNdl7jx71gzPj3w
mAqae9jDvfE8JchFjz9w8dJdrkStNYDkbLTwfLkXe2dyCF1woeRYTORWocNjH12V
u/AzUUmSyFhuxtgToC2VfRCsJkuV/UhvzPLVzJgwXjNVFpU8uYZk0Fp0LTKsajc6
2WxKT0KFOYMa7TDX9WbuH70zUBWKjNPhmFvmJvcvjMeI2pKlB7n3Z0aYxSzg2mYa
H51nuIn+4oXekFWlkyAr96LdGZFPI/B2rIlrSyTOR5UxU+HTcvCT7OFMfQU4lTvU
1yYK3s1MfVmqY9BRPXSLZMRvCwdjWPjs+jUuiPJ0Jex4Z1mWZEs+GOS4Stll6BqL
Hv18gd8QuWcngXuAY7mVnj5+W0ixp24f1AdibgHPcmnYPW2vCqVQWKESOV4Q6WTO
c/uYYcljEmVxo+JM0AKONBoVCkJ5CU2W3ricbQO4zvrjj4RZZf+81/NzE68eOEv+
yp/XnNjt7KdC7cxBOW+9GVPzNZzh2qDTkNYH6PbmgSHC7HI1uI3T0nlEXTxXb+Bj
BZvYQt1EzZQbTSGQzQ0AmCb7HL09ZRtQCmHSTm0mhGmW66MqqEYVNf5ppW0cNBvM
3Zn3NwcCdYQpjxL675sKJvoszyA8konsnAARJe49gIbmdOm6rbW9Af5zIepRj3+A
tF7xP+A+bMdaMnZ2s4BtWMNhTiEAjRiv7pWpLEFAbVZtbnm/6R0nPW2YNewImvWk
H5O/PbOnj4Bb4ir+mTD3DI+C1eKnZyhevDV1Zlduv47SxmvDMnF0RNiRUuCFKEhr
xuu8OhvVEFGJMc5GcDMtwujX6ejDAd2eWEnS9tvOH6K9pIy/ZepeuiHwTiqV1ql4
4NcqptqXeG6jTthLktZi3jqQ6kxIhz9WzVUBMNBudqaJfNQRqm1LXvJysaWdfbY2
YiVz+iQZhH5VlKqCkm8jDPEkgqX5QrGN0Z6cuJd2Fxf/nk/xuJt4Zt04Y7e8guW3
omfkucWUKgOw70NbzSAud+fyfoUtJW1Q3BhBU9SwrQqc7sPPRPLejsC2c9+z6lou
BnqFWB4+q6fs/InKoBasXcMwGocNJCAG3nfDG0XtiTv2MEPerFGNvlZVhTk/gD63
l/AailkjrupdorQHT4rXI+puBmzOtN9i4BJSgJDUa5T405mih4tPaFGs7tzRlUYC
X2hcGYxMUg/tY6u7b4VnDeLTqONMH9l282JyS+Aq/hV7/5h1PJawlQu7kYTtgC4F
FGWZyOgxK65JA3GUrsVLrZh+3qy1Z8lSr3sHKx9IuXeiK+m4sxhlQnpsDb63sAvx
pTU0Xc6YcLbtw3x9dI5ZU7iECjwaGt5K0IOXoJvieIdNRvxv+pX5NuvHPamrQ+bd
S4K+cA1hx/1fafpGgRZIAkvwGnYF0Iebab03F7pM27aDAwo5lLxGkF1J8bXvRYxb
gFMHHBySMwijtxC/W7j1Hh+xB+16staPt6wY0w3COYMSiMzqoqQNztFhs97vGjYf
anUT6jQiUfhIJij4Xnn5IL36Htxo48RlqvqSjbZKl8LOB6AIpEfheMPf5aS3ZdGx
zN4aCgmJxWGZ+ifP2CHVnuhh8+elUIx1aO2qk/epzHQjDWNeKrrRHC4okMT+lCUK
ugzStw6z2sFMpnV3FXK5HFfNPCZGrcFIZIGVaNEzXIwP4NkavOFyATxwQFTBTr4m
dvbY7da5r2FiKmN1DTzGNgkm9gGCIZA+4u+2wSfXZ1iDS+e+yGr5kgPzqeZQQEwk
GHXNtCDWaiuTnhdz9u5LoNOfchCg1TPHcaxFhypV5OEV4HrpMJ+VKlvOMHVvLhmy
+ksBJoTbBT0Mi4mqKmJjbMOT1ksnJbJp23pFXA0dTWXf1r5Qt1UtmkEQxRrM9nmL
LtgksKSSUrc+JT+1+sGDU/LhhaCTX1i0xWnFHnUhvyJUEImBZTNOeo9W5ZnRILg5
rrzdWCfSNKJBG+4YD0jLbOiuckFAHp5rzWWEl/t/duMTrije57WHMagiH/KA5j69
uN0Q4ns3n4JW0JyXMXBupA6El+jTtCAy07W5YG5OtVXlchnG0POxXdCfoW+yrXiL
KEEqFA6+3JGZ5q2CeCFlnbZWydS938bWN/5I5td8/Aex9A7Z9lVLFdbqprqiLWDK
pmbBbS818HnQwqeZvX4694fU3GPxoy7nySuNX6bod6uUr2xaAjtqSc1S/dsebXRf
pQCadGok3/eEcf3g0+kN7pxBpTlo6dTGWwriAHINbsIRUJIRupEWvKdj+6VuIR2L
uwmp04LZN3PK5vDCa35wLktMA7rh8FptaqHPNJ+ADNOIeZwElP/V5wdsYQl+v2Sq
qPhj/2gPy6d4EcU4M/BSs5997PeZJfjYoVgWYeKcGOW2hMkC69h3PAY1onUC14XU
UcZoREkzpIqI1+um2G/T0objypgl7pqUti70ab+kJgrqScwtO9BsDJ1Wt3jsUH7r
yZCj8GqH8ZQmB1Y/HqfCykiF2GFGIq+kPhS5IP4XVuSYcIB8V7UOKnzERRY52LTV
7f2bSryAAfBLhwj3/dzmJrclQQ+RnAX2NlIwgDEnG30/WKrTNUaLQdcJNbJgDKbJ
g+WNDWhQcZX+8RnVZGXbmaFdiVhgYtaPg999aVHeAsfs/egOoan2VRdv27i9Vpye
ClT2YBIKuxUs7WYJjbyJzKQg59bpdnuO5akoutOhr7LvYpK4JqCymw9Qm+2O71hy
Hzny28tYY0w2FvnbpqdcsUSrezTvg8Sh+eHHSQ/PV3P+CyUNneG24e8hZID8bNKF
5NsAEycdXZnEySAEQ14Sfm9t1QLMmssEFjxCeylUV2rbkniB7VelMzDhdXu9JyTd
U9t1IoPj0RG2fojxzJmaGaiejOJngRuXZy8P49J1gKfDxPr9xBfbpl8SOW7qxl9u
zRJMW/s/B8h1w9NVhz0msSXDbiHleUCBiKFr9tsiVpPU24GEd/swdiWZexGU6MI8
GWwouNutOZZ8PYHXDenDi/6dbJm05O85hndG78c8U0jTNLVhkStEGBLHRz86gtng
ujUrYTCbf5QHiub1th8PFyPjyclYJLkDBQuCIyyllYcJbYfk+orzV0y2KrAcBgW2
Mv5ERVgb+L69esmFNduicIm5Swn8ssIlbfoMyQAs6wvPl19D8GiH9ZAytEV4sizL
WUYQmxljAoyPlNilSl6pcgzBM79X0e0pLNn8nGPsqHjKJ5yIFzbTRW+nH8RTUQdI
pYOQo0+kpDTeknjjLpGejWvx/NvwJ/4/SUNOXvEEjgrnIIlWPipxW7F+1jaWkl9L
7olBL76BBz46OEHDRmd+35mfCX4HAiYgkXBop1uNuJm8H1+vlk82ZUa+cEfVisX5
sxiZuqYPCJcrXJ5/KxKmdpAL53YY3+U5VHeEwmsL3UphE1ntfgmms+D83H+4RzcB
2+KcCBqLSBD49JrbEi35QBV3Ym+Ufy6/H21qHEeVxU2r7022FbnutzBkik9xw7ze
7N3rFpr/1VL1+tODqCowbBdggetDkUOj55kfiXC/x5/SztHYBrXy07YyqUo3C86c
DG5dWVTF4G8nfFUx+uguAd7+x16zI09TYWJqM0TYPrPo8hAXiGyoNouKxW2GL17j
XiIwzbATnQwmhRwE6c8G8paV2K9RJ4CxFffU0XsTyvBSXiMsGD5ucRgL6qadChzP
yMmUTUC2zsk/o+Sn2AAyiObDqUzfEqBoh9JMCk8XrewsyBiGpwv80yR9MvDtg5V8
KJogitxWn2uiukoqTwawpJpxvqTG+FGl2HFedU3ziPRv1xdaKO5TqUWQ8BVvUIUP
HhdToMEnKLOzl3BE9WexES1vdnVx/7WGzPHDrH/grXVBzYssA2agM508nE8oihj0
EQjPcEywFuy6B20NzJ4iv6ty3lSfnQVXRFGeFxcG1RynHDp5bXX4Jlg5gB6AX7RC
MjSMBxqC9jTuUTxZx59hFC90EF98mKE+WFIO2/Jy+G3vTaIASKiZ6beBvrFp2KZk
ZmLGJFInuOyZLQf87mdHHGLi//cRRaEV3JcJogxQJEu8VJCGhWlPFLLJmexhuZ9A
YMYi+6wC6Gvjw5Hc+Ho/TtzAYkUTyuI+CXItMCWcx2rpM/4w2qcSJ1QtkV1ngTVJ
/z7+c9Iel2mGVmrqQqtf2HWN2a3EDHEJuyKsBP+GxQlaaplzXpUED7g+3c38Ga4b
mfwmPWUrwC/0MJOFeTFqRCV7tgT0XFNCTEged8TZS6HrIgWBli7cRH+uxldJbCVB
b08PUirwZIKGpVd1OckOCJ71Da3OsCwE/1urDjxbPK/xmfMFN6Nx/SMWc+HPYEA0
yrjKCRoA83/V5tpeYD4ju5XQjqsxQ09OFgNOllN7WHVQt7mF73KBPjc6fdUhIF+v
+UlSAu+fCWak+EOtlVg7+LjdI669QSDqgmX5r5J6u8Z0ieC4l9XO/G5oplQQpP4F
3pmnMD+AQZnuhxQKfR9sPgtQsSamoaGThJQQX7xoVp7KKGVMLcQfitS0iXSuFbBH
uJb5gf7LOxMJngvcQPh8of/DDQLp/88BsP2yFNe5yYwzu+xhi5QAkS5C+f4iHpZ/
Cu5YhCKquxwxgDe7C4nHxgAp2zAzETFHSvceF4vHVwOYucPx5Hr1Ce2ymM3NqxDJ
GR0qbV53OAB/hK0zS638cbQI5RU367Uv2fEqpIAEYttQ/SU28a36CsyH4oi5k13b
f7SmNXylkbu6ZbIaEzApLaq6mbM9LbA/iggfuiDZqZPG+GDUxO1gQ+eKVJGz4vtr
xGis0T9JnatDRJDkPuMEIwLr1RPQYqCmJEsG2iBsjje6eEyRdZc8toLfwJ9IrTMB
3C7hwnTEZX4a/Vh0p76XgT707ReXRf0z1V5TRbSBMp5LFkM86GbIh+XB6JMi7yfw
ySaW5SYD8R/ddd8jky9MSs7hU0i65A/vGNV9bsrgcN8ZAU7504EedaIMHfYWdmkN
DW7p4ZcXpOAQ7vaib3JAJGDM3MIWbhCFvuVOCLHbn2Rkgbm3atxw8TY2VX4uFuhw
DRDL+rg+uJQveNOnWXAJOoGeyYLmmQy9obF5BwhufOcwCupQBRA5LP4Y9wZyiKh8
QIQWhFpQZW17oqm0R9VQ17spBD4DloxmLOrTEEmUJIuuLFBOkg1PD219RNQ0juvX
8DWz3cO4rbbFCcLaZYCx9K9WdKhopRFSWwEsScyIBBuiPC99r3PrBN2ljNZ7LUl9
OCx59F7ZGoeRHI+FmGuQggpeSslV3z1vj7uPCSYiC84s5z7dwWPQ9/PQJ2TSKtQ2
whBvr8M/I1aMEaVPCTiyCc55f/+HYxk1W/IUatpw1olMiYSXJHSZFJB6Pvyf7FI/
Fa0ZtLtF5ndt/3FU+b/N5hUBJSqXNHZuI9irYTdCEK6jTRLiXORz1AvZW+a+u2kE
fDhfGknETKRbr7Vp+V+uklDxhvDX6ldTIQCTK2+BhXQGHwiZtJ+lrCQbwf+z4lYw
MMVkW0fU/6T+L/+GMwWLyoEePkGY4CicoLYQMIMvR5q3zpbjXxm/blX+J0g1/3KK
wAUAhj52ffmLk7KLjXmO4QtR4zCpIwImcWcFrVNF5e0bMm/lAwkUNnm+vR0C04EO
Py8kTf3AeZ2FS8OmLHQUi3OsU1WWn8M6I9ctG3sXiHRtMpBPbFl4QBfMX5Gmpauk
P2SArX9qa38om1UA4kAv317VLWsBRTKBV0DtkoX/t9nAIvwpgGpYlioPjOCM7taF
KgjwDqVVBroZjqJugeuJrU58DTYlGAhQetlZ08VcO3ReTLiSsLtri9LENZodDm+Q
Q8UZFRAwEWpa2y52e4RzC6kMlUShmV8mco/G7czzjDkjwgJMUGnGjgVQEuaV4WiG
Sdfe3+wUaEvzMs8KWjPVqA75BGpzjF1lMnLTBn65rP5RfCuTkSwxK3r95DdbiIvU
+kz12YT0qUjWq5nm6ec4X5p54BhhM/Y9pv9tAxTUeeQYo32WLRZ/cojkQLyqtSQG
oEla3bEccZKK/XxKWto/0wMXuF9sm34l2ckLbHotpEA+PGoTiwMZlTgvIef5WBqv
ciDD5hCEePL7+7r/nLC9AMv0VWNpkqyxu79C7jAOlULDApFNCfGDq8814uiLemYQ
d+viFAA8T3IlUEgwUewtBVmJv4F2vIE+xIdtrbbXvNv0epKyJVKyFfzCrWnwB5wO
WrePJUXcQmSdI1vL4QVWlcX1Lxundt6ptmvJ41vXODaPRXBPqLWp4eKe0cbcbzQz
HrWw6VsL1TseE7VON5hrl1AGtfd7gPmHlRlli4CDLpLCbxa3igHxDU7Y22ZCjwNe
Hp2l8L9/0lRvyiU5hEJrc0fZ5UfPnRwXXnHAVgNSXgasVuRy87oh24zxOWLk8opq
xFhRQt6K0rpQBaI+KcXmII9eOdcOANH7JTPCK10BgNBgkiJBN5evQfGZPC6ddVFT
pN3X0CJByp3T7QxHbWItMgqNH6Vx7W13mpvoNxct6Cq+g8ZkD84ORIeGBwTjBuxF
+ET1kXq2wHGSJhNTyxbPY65TJV0MeUlXlYwnvl1ETd3BjiiKMMMyW0ZZOtSg/m+k
9P5MYebo3xMwBTwkNwrnKiIbVjXPuE6fobYVKrzMwo0ib8O7iQC3NsrCmZluFmoF
hvs8+CSMQpcSvSoNecNdcFrx/45oO/lHIaZW86uGCqN1FZ4BmKHZg9cNUFie5Nm9
mFuvIeiOE3T1SS99ECIsOd+BKPg6kQTnZebMhnYLXtR+MvWgbcNuMA0eiCTROF59
nNVE4efs85oAPIBWz02Cfa2MWsve45fCzNCetM8hyS/lMyixCoixmhX4gOUllLgc
L5o4Fm2LiXLs0CxHFmmYGhX+JKt/8OhZ1IKxe3L0jWo/XAr6fMertA8yOn9FcQiJ
/+SWB/Mk0ZsqCZSO7PvXewTNNU1nqoRlQikNNVVF9JrnC530k492StCm7U45lZV3
X6LDfQtv/paTbih0qDd9rBHTewpVLni9TZSSVo5z71KK17Dhk0Qqeon0Oy/nHvqA
ThmX2jz2KUJwyDSlmKxkKXvsFqwqvs/I9iSfAwqVjbScrVnXOQ68IHWbg4vyDP8p
VgmeemNCMjAHlRCUC9/jyEbLn/4IFEkwQxaV5v+Zqunmju/im5QVPPmGVj4Ikvw+
hfx+tC83fvkNkXJjQlGq80nW33zAf1GmkODLKsmOViHTouoAi+/Qk6m6j+VH6ZgB
hxhYYAYKz/in9BJCFDzkH/6lBj9DOsTkAEW/FNlvnW7TCXYWV2bPJ3tECGBJD02O
E7J/JYPd6oUUWLbim5+7HOFNF8h9ydnxIL2G5uXOwiWOu7oae8wW7xHDL8nBMDmE
aNCpG4t/gQBes0BKlQbwrxkJgUZcs9VeZtGQlMfuiWjd8FRL3HqiN3nqYgvYKD/D
f0yrz+9ft7K03pLJHFYQNB3a45y+ZAhOmSNaXovAaz0AHvWU1f2QBnQdwmY7Nh4p
yHTuFY6qS59OneXvle8j0fxPHIDXkJy8thj/G55xHfMQKXi3PLf8XVwR4OtE8RoI
4DI0/l1S2ocWUeuv4dLGfvZGEkG72Ne2EDjukuRPW9T/O6vwaxlrD9mohqnlXuv9
qD1EUboO43CLyEAqZL6dl2HvJ6Y0dxK+Fp5hT5ccRYODnPq9QW3qTuBnmxrb/fW6
MjlrvP4VPoJhoBBFlWxUiT6CZSBmxn0BkY3QrWKeu+/TuXMTQxmKITG/rC+It0ip
gdbhGuGqW97WrHc9SfgyE7U36FCxYE6ZifjUB9ZVfRKxdGCuTcIx9gUbKLvt9Ys3
4zTQki7ZhkAlefIdAREp1pRBEnOHjvYEFNmO0aqc6RdoogFPtcn0fPro6I6Kmbs2
1SUDTD9UDXcbgaewAYMBkuBAV6rcloYeev+UW0j7QdgLNGE+SdQd5S8F3R4ngjN0
G0NByfIntxvYINTeKmSUbk47fGK0yJVIyu2X9mff7A8QDKv2T+O6CTGwkPKyjgD2
RD0iLGyNPmoG4KIuj9eCFpA7vOEZ3yOaSc1+cDCAvv/XWvuqQqkrdEYr1wieG2jb
XsEddTZo/PZj97Ef3P4kcoVciSRjPTXXQQFS9pL0C8i0QXAuc9cmIWvjfL7HobNq
o0cncaBI7d18AZ1PqLqftdTAdMj/zK7giphQW+qYx7SskCT17YDGqQDZOhG6jVT/
yFkkBeVQcJVHhIRiRXrv4ihzexMttcfajuuZMFR5JHNVuRB1b5UI9/ReZNOGjxLe
6shXPrDSoPLwg2PMuPhqtx6QPqqr/gHVU68SdnhZ3kceqF38fFVMuGo0NRH5WmtU
8SOTjnQy1tBI/VL0SY7bkWmAwdDnISOGR6rYS6VgC00Y2GHMbnZlvBCISz+l42FZ
u3FtEOjP49ubAURhOba16+ebVnpEGavv3SqHLMZj3iDMxIBVkf3Eo1Y0ysgC4IVc
++G2nEsSGdHSxkwtZcK3HW/Ar+AK+aThmYfMDaad8Q3pFRsv8ushBTPT+WnxdIEb
kWg7eS2+e/8pNeBK/bLqfq7uCigEWs9ZN6YYzyPxs0MoGM/vel3vfBH0KbIVvhO6
Ol/0cR2oneddbxk+ecPV5jH6o3TowFaTq+1BwjTByh+mTSVwea9b7n4EoSsTMP61
/3a+OGRfjWI4h7+4RzSMWGc2eeKzRw8+3sT/rzoUTwxgaaAg4pSBdP2EkgGUPQ1W
drJe88qwoETPnb9UQnzsbC8DqmzHZFrRjAbLYEuAhMAHT3V70BcL0jeKRQfwQyqG
TUyfjnmX8TzAbgL9h1CyCtYvq6p279RAxG3OP3Pi3h5Sr2omidXVNBWU1b03iIIj
CANb1/NaFnKfZRlDtcGru2LyllcjSOG9RNzdLTetxHDRuKlP5yCdnHbRNtzmhLA+
Hk84caX+6YNzirzz8SxfEYD1bu6oe+N4fSBmVmnn+oEecKFNHtqQB4/7k7qvG9pJ
u8ZWoYrGff6gjeYNPLZF7z7kRkGX9eICWI0yVMtSt2YUGl8rJBjkYcYy4X5hgQvD
Rhl82M6zUV7NJAKhVKmMOM2+hE+uuNnZRlybM7n1ocjZt6VNI5loS7oErP3iu4Dl
lqemAXtQjOS04n4Mb/BUgY7l4+xW1//tlomNc+fsBymomaJ2LZj6GZHGLa8s5xFO
fqkWSQFdWAadJyk33nSWyGRzHzBqOI+DE02+zNm22TlGwD32cUwjsr0s8htiBgVq
lq3X9mJmBEEnC7/gSFugUCblQidVDQIDQi/b4eMYzQzXEhHej2/3eCmtj3Sr5wdF
ARXwzW0bIHSJsNFGBph/59xNH+Z+W7xPNcD6AJFOUVwGTHjhVCrU1QMEAFrtfwTQ
Jl+QHId2fHchs6tF3uXNxXl3tX+L2QI9a2tCkH5idtdHkJoUaLH2cLWIh2yDiUGw
sA0+Agf0vTPAldGExmhe1qKBC3hh0Ju/f554NaoPf8V8jiK8+JdZ40p+Oyi+EK7m
2Kdq5lc7rshf2FzMEDTaFSrtaZAaw5e3UZBIa99fmn+od5IXz0rRO3/VKrfucgwa
PNvwcdif9eJ574xGk4mO2adtvgudQew7VSo9HI9GSZq65AA7Iu9scJ1iEP0+JWPF
HseDhXZAcPK+cmgdUc30UB58le1OpIuili9R7RcNuybg9CYaIhzpgug2wIsMezhj
9ayHhqbnE0FQBcrbijetqiEmwdwBqyPf57Fq7/tlZNgtvy2smzIPZnwkl00z4AN/
qgiG097fc9RjjNFBgrJeSJr8ZVgfvCT0QMMcY6kWC+9pxmPSFCuwim0wPGXAfQNb
BHavlo9bJ88wN4W6OG+czN21oxZ0GHqMH5IprWgEXcgNk1vF6Nz2HFz9QekT5L+3
thMV9LRttdsmfboha2073ZYphzvJ5aZGVS+dBKGpek+7y4L6R1t8c/0MSqJiLqAD
ecAidpwk9eGXD47Dpja/hM3O7llRsSVAuOANfieLtGkCrLt2t/3OImxwQXq8FrIH
I6z6ICeh5PDNMlXIiIW2Wl+FQh3kO36rbcakJYxuCziFC3GZLjgI0EnG3LFi/z9w
yZW9AvVafmhxE+sP2p9NWjm5tBGrEirAHT5fkXQ6d1Iyv30UwGzMTNpT41ITZJBf
ON/Z7HE/wIxkQcgVsMu4z3hQiadRheJMReveOhZHS5ii6mR5eZPIeWcnvn3trYL4
aXdSuPcNxZaoWfrl07pcqjtnafigv/wAEOwMaFw93mbEqQuyMysPavg0szqdWXfI
3WOAhXzwpTknGk++ciyKjtEd5bYR8CEvWDtVIPhPr26WyZzoV3GaTRyfEdSfypGj
Anm29BW7DfkWlGG4usFb3RSaCPaKIGUo3XIomNM66YGy8pWlPV5N0B74RNiWCsdh
f/QWS/OeJ0EUE7iZcS0CL5amP7VILPIZ3vW6m0Pac+LgDJtqgRYsoyqQh3bnVCJG
tsMbDPC1ERMHQQM7SX8HkdEWz0t8h8qvciiQOcIgI5puGXjrdyh2lc/XwZspdCGC
AJA4TRjfXg1was8oV59TNBAiFr3fukZoPSYGfLwWkWJNXbaVPoJVIzlYw0Age1Uk
FIyEpFAn8JsbqjijUSnWST8ODU/5XEBKrMQvF74mWuTJiRZQZshvkXEzOEUdutGA
uwW6qeO2OFfXdOee0pzjtzmhaD6L/jbi/114IeNblQpnj/50Wr6AsiI9rfwxoPxb
1zUNip1WE4Cwgg2sduIB99PVi2oe6IO5TtkIiBqONsQfYDvpS9bZBH8UT9dCYWX7
qQNLjDZwIO7sFg6NitqVC3zOPpwWdvgBE00Hf45lJ80PLamwtYhIJfgyqxZY9sjI
AedEMrve/NZHHpmhAhavP1cIP3usLOpy/lNUux5JG5TTcbbW36y0FSvWTO6HrFFC
6ZfcMMI839eNskp78TeWyBZLgVy7lCd2S7uN96cfP19tXwBmcH00FXS80bUsrR82
Wnnz2V1nAsGg9cBEXy8S5gXmZn/fVBKzWsZu/Jve2HOgV4sA7UikokHy1gxL6fdn
ML209miuf3IzD9v3nO+7STaWzNA4fbVUyF77XfGjufALQ6p/P+yebfbs9PDRzZrM
6Sz8YpdoLhyjXUkvwUAJqpKmMIK6pmyU5qARxMwxczyoA0mgfzjIH2O5Iks3h3Nf
1a4X0qQbViMHnhJ0iQNjMFTrK9KbhvfzEJ6lsWxWX1xL3/wRiP0kMwrBBymfQ93N
Ab30LcuFZHZd4l43bwP/Uy8ucZYfnsWz/ra+SVze0dWI+sPTBRU9nvFaKau6pEIU
Hl9r3YPHjaMlexBInUmiYB9WZKFrrYsak4gySKVACFASfJG7UKDqpINIE70RDSeh
KT3ao4Y4C9HaN+qdpaoJ3+9BtPoOL7G8d9CGTxaQLAl6Xja1Wi5/uIvvtz8pLw2q
LBNbwXaL4W9Qx8XC1xPv4sHyxMU3q20e4mLdCT77sWt4E1/etTN0mA1Lf1VFLA/Z
rx7DqacEU4oOfxvWw6so4FXDIPubssR9Ga35l0pDlHv78VBZN5wJV2Z5YC6XksYX
fXQvDb9JmhonlNC/Xd8lVxAMXyL9zdvzU/dOe/nQ9CTK0twNXHF87V8pU5GRCy7q
A0S78gegBuqaGQfd2BIaa6k/c3bNTtLBZN9Y1nySel8AeiN0Uc2jv2y+ctmTYCR8
8X4oc6zGeYRcDK25ceDuafd75gk+jvzM8YGSMbi9j6Efvqb6oAPPy3kLKjXTajzF
WJbhw3JfRsKJs35WSuuQ8G5lPVEuFta4yUNOO3tP9CV97aO/rb/ke2hIDlmEtmEX
Q8KiUZ5PXv5B5rLIVifq7T1T883i44JWoBAXjhy6PMspC5qz0cBR6WFKFUz44FeP
EJOA7paE6LoJbURZIDwYIHnASaQWrJ447a77wSmtIbkT6txqC5IOrO9hqe9ckC61
DI75CbjfEiSSaH5P64/MyhTJsfbR+qWxeBIoai1yequFhMSMSBv1Y0i2p3aunBH4
yPDOZJiKFmguEiKxvnFYnjmdcjuq4I7h605IVk4ojUlUO6xEeftwPlm0CmRdONdf
7e6ESEnOlBXO9hAQ0q0nDQ/X9Gioo68EUuHsWohcilTV3hE16qBThoS/HNXbNbZZ
YYskTct/S0IYkd1cps/6lH/Z7GDUDWbakJAFUh5/0yqWE8G4uwZ9tBjmvoCt39M9
RGn+TmL9zx31/uZUT7t57YjDJq7maa9gryyRPYuRKKl002NVsIvvhfW2RA+uKY+G
lO1Yid1GWRZJYqKgZZ3eCpV1HXh04RMOJi6ct4oYtN+YoBPW/bI8iYNyJGy0NGxW
qXwhZVFQfWvrl/sVAt+GKzvZ3QSv8OzShzhEbWdOesRvX+8YH6fZK74GzxrDKTTx
H7G3hKuyVJWikjIb1qlkS038YtzBi2bYlVUytOCaKOUfcLUr8XsT0xFIwAboOYe1
biTb8mvh8/8zwvXLSmSuUGLMH+ryJUJDYU7TGz/sGYhj9/FArzzzznT8nQe1AfUU
UVCNZciRYxoMT1bqNXNbS0jUoAQmV2W7Hh7e233n4ukea2p3WKJqAMXyQYT0vyIS
HlQXNWdqcZX9IBJpjdi1URSwUQoY4QHImXOZA7oiYZztzrb7evbHegzMxUs5JWEg
SviTNslVMC26KyJOnOgCIQK99ZNIztB8TPbJNDsQbfmvDouJCfc6SM+hfKGtxt37
I3uvmdtn5L66+9uDc09O0HJDcWegtybKkamfhKkkt2gWlAjMpt84Lflo1sjbRTjl
SvDffQUm/FKyVfFrhEB7ro2S9RI9V48ArLqKw2cZRgZDxJBTLblf2Op4BQcuel4b
CDVMP93rZFy4Ur78JsZ55JlhWTk1/vgT/zN5mLttn1SmPAdCwjxcFhlm1AoNCyWz
vY7WML7YaUReCsLS5NruL3cFKeUCUzp/iMz0VS7b/xEFnmVCsJbTHKene4KlyKlp
DBzCLp27ncIcPnIl9sRCeTAXG8PImNxJBGdbdHHDbL1yR49v2k+G1XJwvBmdlsup
bEpnwuxYA5cP3tR9o4088i69qvvx95PHQmwUKQrDy1r1OgqlunqHz/6bACpiN/7Z
aEC984a/txNEcS/kiXo8298550Fb7gdYszCtg3Xs51jUj0dgZzIfZHJzSjBNdhLx
JC34YS1ydpV90HL7ZIYOLJt8zy392VmlQbhj/fnd3FaEArzsOYA8ZzlvguTBC50C
cb+dKeUur7pa6ZsYZr2k4jEnV5Z1/Cuf7WJIN1FVyF0Ka6F+x0BCZT9B+RL58k18
rwJ53IYF7Vqx7CzfEExlL+VZAVLG9UB7zDDkcqMWTtsST+Qh9kCEo5WgknJElUwe
E6AdgWQuqWm2TIXPA4w0AC6wrjN885GpOl30RzP8n2iOqQzS9rXBgo6eeX9ia+LM
ZBluG+X4dnDNzr8RvN1jSXN/AldklP1rPNrQNhEdYPiTUmYxpEg9xFr4DwsYM4ic
RzzktVWdbBQqy0g0uxqAku3wOMnlCWdoBzAXAlsaOdTlwS+Ltp8olny1i34fbu2U
PgU0IHKjAQ8ecgSYLCk/uq4vzSRC5SaGxKkLa0vbKqnLiTVoTwU+eFjYR+gYJH5p
/DW1y/nsNn5Nc74rqrQv7GCwx1/qLVbkqgRHqvPIw09EKaHyYeXo8vKigIQbjBqu
iU/Gee50woPESG9MaJd5lXkVztLE2CBwnf5RLBC89B84msnSQ3g9Zzyn3o+gfqRH
lvRC3Vn6oNDfgFbX/GLNX1JGyZ3gVnrr6zGYI2IZ3ZZX88CEu5og6hmY5DE+P3Jk
AAJNsCph83mywuFG3j18ULCBewQ4jSZweaAH9Fo8Zul3alHDfua4EekrMNn/sHH3
5YVcnsA0hl+bj0bUNf/8HmnGfHyYeLRtX57eQ7N2JBH87thKefHzzcYiuEarrhJv
/zuxwVeUD7ngn4+0enwlaS8lu7Izu3skmpr74N8jxRRNwphTCtKUjM5ol7EP794C
yA+GPbKVinUveNdzpGzRqiKlFBjpGJ02RM9Exz5YyTkFkYxqUoFFrni03cl1eSii
bUJsbGnF0JKaG0XOgbf9vp8HKJsRpqbNabTMSvdv5UAfT9ghTqAN5Q5jqq5XtdtI
DjtUdYiJFF4aexmRNnsMfThWJIsuf4/VJFEOOj6DNqTimveAm8WQSOOFtyWFs2Yf
5DKJPaObVwFTIRqa4/6nhaWlelgSJ4Ahb9yUBFSWyZXWANDq43ujm7JSCksjOQze
zwpJMKNXEZFRLjceWPX9+uqfulI05pDrNfsHYik5XIgfPn+tT4Isnc+iOLQ1WA6B
oWkMEDUq/wiAy3rIMVWXphRf31zFGHDgOTsq74nSO+TfZq8BmL7nZL4BSk+UnyuX
EUUENnNWFo4k8WQdmthbMXr8FYo7qTn9pg0/8MJwHOlgnm3iXHfV7Iq4rlRL6X1V
ZVH1MqCytezP5+ZxMRiXilfSMTw+e5rRNTZEc7FhbqhW7JDn6KyWSQvhmnocGYvL
+OAwiLb+pwAPA3Yoijl6ZjAE58ir6eOqHjzRwesgU/IwQOqRJNjmlfcWbxDl1/jq
N8LETlW3jUFIJ3VrJ3wZ8muf9w8esurG3wyHgZUKyKpD6RRaV95WRw5+OO8GeKcu
x9pt/2hvW/hqdb+jTBfGZpEI+x0TFv4m4sTGIU/JAi+5QTP+dZgUU++AtafLtQr8
mV0hlCyH+I4AWjbyRqL1Wv9JN+aP1KE+LHlRXhgtXBXsMJzjHq39RnHpIMJFEBBf
HvrflCC4H8e90YxJ4mhkUb8OjfZ+0HqFMTofnlUpZd5j8nSYMp6DllsmvRKhxNXK
3HeTonJit7r0zgh6OBr+/2agj6i/QWB6aI/NVNYev8WRTe3uxHidcxWNGg6QiO9K
r8IQNd9KIPP79e38qTu5B+GvmWNBlewrBQbKZt0dsbqsCeXugiZVJv+W3RuE+unF
3fYTliDCc7W5w7MABFXjljkFN73FZleEM66K7P1Kes6LHII9vzc61n6yjIv5Pzqu
XWvAhWEo7VBIDNtkpCCGV55da6cpHEqN/3tIJIivYOcLp4IhDUUcV5LsEJZjpoX+
nvsJdVO7pKMKw7tpSFUQeLqVinpXmiGFALblaYOxG7L9OI8TuhGuNPKevHTG7VAE
2vy51WzwgaK9XNY63r+NApgA3BOX/S5g4NpFGHRUriE05/Yu8uOyfNHU0wodHVeW
39hwxJO5GW6uwSpCbK0Qr1chtt8vbxgXmrTLFmiswOE9qcaxQQuR10LFauPRxQ9I
4J9lEBg9VySsyTzCAjLUxiURDZdXysuKdACy4oqZkHE9rcHetaLh3rLkg6RTNMr4
YFVGAgRPCrXPletIIa3ervrEvnCTJ6uaoWqZ/+jFSFHZBzQ3Gg42uUgpNGjVvFMv
PeJpbWyjFFCNplZpjTUVeJeWGXvnp9siBa3jO2+t04IfLFIkfkCszNt00JKlR8s3
lIZzIc+BEuCzczltGzxRGHBZeD1z9ai4z3M+fQ3FAzuC5qCetHixS8jUEaqnNu7r
l42lI4zsSn0cOMNi+6dD6h/jIiDnzfrHulbMLbDceXsF12GOOAKJ9YjvbKXIEzbr
ybpJnp4LhXLDIKSvD1xKHZvSAZPjMSE+NycLr67ImSp623Ec51WzfI0VC3sYm24G
iF5Wvi/7hidkAAwtm7IOukWZUc+2m5nNENSfEY+l8WU9L1KX7t/friN5fcpPRbi0
hW7VhI/JFxNSUY3mH3B7lXKygq//S+DUYAww8JVLcJU3eOI+8jNAedJ1ZbAoJVew
1gc/aHBn+30WUqMlaltqAvv7ieUGjP8rXN/+zSpy3zTKTyZM1dcdX9RdmmaKqJHl
iuVU5940kQn/gvu/VvQWYetnl+GBZ3oCnzLOr7Ao1lAign3/C1n1ejwVoWrO2ki2
wdWy2jztp4ud6n+GwT4D6SuDrvq0OWjYrWJPdGUMvsnBjGNm17EbW2DAVhvHRQ9+
C2B+es/JQu4c/srRSohia5QtPWO0QvvmuFYZ5G52DgcZgNayrCz43JdElUxZ1C4l
CGEPU2XtsNrDiniGj9hvzICdSSlTH/BjRmireU7rYQUYgKzBXKF1e7v0Gu5KceJN
Jwel4c9XhJrYa/oEtWePXDV/yL97efwWGs6hwaIDvnPidVdBl63luwr/KMkI/x4I
Z7xrqfiWdlqYr/w0z8RXoVFGkJLw5ZExxlymqFCd/9IQnTrnaEncZTQyCpwxesA8
ZQPZNm99V+tGWmom7yM2gcGXtZgrZLB89I7+DnB+NtccWy9L3wOC5COZz7em5RPA
TYGaKqxe9i3KO+25ZNxkVn/nlTUTBNLfUixMYG6xmSRIfoJOD5LC+mdaEhF4x6A2
l1TcrHzKIlnFfWUBk9XqeLxPmp3i+HKA/0UChFJUodaIJOgb6vFAbphXI79cvTyh
AWpHqcYAM3p7jBwXnUWD60jWNpv0oedV30h/rOD8zPJVH73Nc3E8ik87xVUcC3fV
SMUAnleAlV++mAQepNq+bn6QjxeUeHZPH+vrkJkmQOBVk/a1Au5thcEk9tITa24j
JZgY9ELbgQyZnnz/6uvfdt5q9L+abrqxcyT1lrSIWMqDfDGW5MkScJ9T6P33DXAV
babSgCnqRiqlBbI8qQvULP1PQYwv2GXmVXqTHZK1Lucaf83oWuGIEbPAIxruPNzm
o4uY/FLDOCxrybs/Xo1+71mf2VepDf0kXxOvk51M4sJAwb2y/JVzB1Vv02IRCTuh
C5KPLFwtf7fz3aSO/TAcUnUeXYEBGtL0sWfMhphM7D4egZYwD0aWfFZXol0z2hnC
uscrU/+uAOCff7KUc5ougpoGYKCO2RVfHdkqREINDo5hVdo4KXyA7JWxmQCdXczx
DISmWlFmu6tV2dMmXPLNpC7y2a0gL5XWCm/Kyy9rDtZsZyugq5ci3SLOJvP12Nxk
BGmJDwHunRvHStY1Te3oW0gVwAAIZXbNw/QeJZIi2rxqg3jHoL3OcjXBfNp7M+JL
MGXkBIhGa09jgoX1nYA/k8cKhIBTAAwHrETTs3862hAdbqq+nooCTmRJNBheS3XR
hf/l3+HSGO62aA5WANY65BoHQgYZcA8G2yQXnyaY17uaPG9+bGnioUeHFNtSRMIy
EtxjyXcGoaEwMbIS0+63pYLwAkfKJwIVP7Ymu3FPYzO/M1UVkl5Nqs/aBdMn39IJ
u2+4HaUxNJockWEZrcpy7JuiVkI9PDTQpYD3D4ca6SFStY0DlvMUFa5FB/bkjP/H
W3KWV/8Hm5uZjbzsv9lPc6fXztKloOCjXpMX3rI4tpFPHLgLYKz9r/igR1sKgCKz
Q+Gj2Io2oCBXbrd6m5b2vRB4NWWTy4lKAp1BAbcNmOwxB81pNHeZNETwag3AVXDF
2PrIayFqroAi5e0hL3Fh6pQPEQB3f2CjFc2fcb+6wC2vnUoueryanmkfaDZhm+YN
oOw6YJ8l09G+SHrwsM4Re3kSmJKgJN8a7Wo1d/n70WGo1gz3/ljmKyrkXQjt7I1D
LerQhyCrEsugU39RV6fSLuxUqnrYMSPGwra/zI/l9B5psrj3ecVwMAEWoSt8Eal/
XOEFw0fYZNrYQLHE30T/8aXKcZXmk2hTLXoUUhIExEIERf8tEXeE4T7nOHtC1vYV
BWPUp8gFSMbH1TFUtXPkY9O1fZgYoGGCKgKM5lMIlEIfR8xO7bmWM9TnD+/cJLpQ
GQvc+LBeicKXKFkoURRLKPoW/RBlEVRUWOrvZC2IhJbrbQWgWoqFqiaopR1l4mcI
vT0JEJBUyx6VgH/ChNG+cJkbs6EtXbS4/a4Ty1NaHoeynID5JgWaL9HTfoYihbFC
b6lGTAvYbBQQifS8Fajq58SBrs/8rFkjxtshW6P9+bPjmN4JjPPV7qnWC5hfcyGv
AHeUGRtyRmr2CcoS1lAx93wd7OfeLlF1DoSUaPTn9U0Ywy8TSRKWIF/wJgBImw0y
b7/Hp8XNETvkAahabeIIQPHvtSzINST1NklbUGEi+Z6po0Cm0oDD7iOoy6VmY+B/
VuENt2CiRqLTctDazjmOIpB/Jyrgbvi5T+fCH79+O+8jYLPvStAdpRXr0zVASM29
5r/LDgefQ1pWtmSEn4T1pbkNuEBUMIeG1En35A7tv/ADoI6FEWkP4ZbNxOoQCeZA
uujBEW2eacH//t8zac94G1PdQrwBRN/yYiVnUmGhjCCuXIjNuT+F47jKLbp2ghtO
OUJFF5zDDxQ6ytKfCbtv4qIyznK6YSCUyBIZ1xUrEZR2MbOtNoFzBdqdrjXqR/cM
BO7puXiCfBsOYbw+GOKM0ECknmGTtvMs3CPZ6+jyCHpiiuLyUPcxKYhW2EsWhzjE
6gQ0I2EX+3KaHLIYWE2Fej4QVWOWeqs4YSC664gMBFHjm/ownTFFCNicdNKmnCZL
ygpbytQIVtkl7ILlEFVcIAU52eCEZa/M5gEzI/kPYmiBYyokChga2bjyVxfh7Pg3
SvQttgA/ucfJ0WrJ0K99q5R/titTmkTYrOxYyaAwCLRkPlkOCyxBiW6nc5K848zK
PLFTUsonPXq/ywLaTj5rRbzPaV3lVtHadW/rphuo5qxBLTsPqT365iztS+R82y/8
vUNnryeYVxTKdWMfrPhtyLiAAyCFb3yQS8c1/W4LukJwFLI+pFh8tR0qYUEgSM3/
VeFGJ9v8oZV+saKleZgwePgVxCljhZFY2CjJr6Qh7La6aGSR1EN/CztDXqe12dUt
bUcKXmdZlKG4z5fhdSCPD56Ekck2aR7CjCItX1vvhixogkoWcetpM6GtvPvfzNrh
O6fpLZnDQqW7z8WeBR775n7T3ZJYF2g/sATkKydBJwjKXCTfv/GDJYFSEXuTfHJa
/Wq24+qL4l0OVWajXEAeAl3mrpB8nq2MeRDRaJ5vcKj2UtbznqsqHnjT5qEg3yap
zmmENW/Ap+uFS8vomWZnnU5nrowJL5ouhKlzI+f5OUR4lX+p0CTQPto9CscHw7BC
pkd80nSfZbAiKsggwXTKM6/cAg1NimZFXKUEluo/UEeKDUEXyKAc62B3XSNT2I3K
kaD/GTrEvPGt1fXVyLiNJC/Emi+zxVc/nlK/yNxQMPT3MKADdDmTIGEiS9qvt0LL
Za1atO7Zbhe/V3kUQn+Py77JWlqcCKUoNAQ2UNxjpTwsne93IYTNmqhKBKRXOzgS
xy26uhqhHJJy1plisf3uiAp930tCHElXLUWPv0pnlti9ykcdx7k35RK6OeUpaNpX
B+YdFasfGTwT/PLPzTGr1fs8XaOFzOF5Wbuquv+ivePDKAQJE4Uzq/ZxZOO08Ojh
ggY5MuDBzRIfduopZV9gCBTjJHmtrfN8cDgCXCN3Da0oWoQr9fY1/adoBvOE4Mvp
L7Rj/20/BeNnnxG3jM6FPlVdNTwqFh8E278OyjmBO0rE+v5rd6x5F+bDZhC7GueF
yEHOZyQ6cmQ6XA83X4pJ+RTW51f4y2WuNytjEPgjH35zS7KJUg3t1q2LMY+Kb+8q
SyxZxPWUOnpyHbUs9dSht0ShvP02U4Kg9ArD7pSEWCR4gcn97LWoxYlH3gtkzQZ+
LMGZVggDnHyJdIwjARcZxOqNzJxP/tO0oG86kxibwlHKqjIJelvB4A4e9ZRoH1vC
RTQX4okdoHRwi+KYhAMJxxYOIp/iS8jHOgx/XpeZUEi+rLTQ72aQJC+pKvhC4pBf
pvbnfzl0AkcrOZwOBC7nWKDa0v+9/rnEC3p9tu33QbkgK4Ml+rnPUaaWlU6BGO91
fFIvHM+vCgLtkUOC69qn8tR5D7yMR0yjUgeFhqxFGxdwLn95YAXmEEasUYh2ldNz
Ker9VPq9BewPtx8egCQHpwUkCh8DPbWS4hQcmn+LCdFe1qWv8n/Q+wSTgAXudJ6N
/TdkYnHI5ILlA50gEqAC+zNiDnOaUMffYuIkntgXZJZVqU0wiQygzpbyNs0wG8+g
+p73VE6F481CT2DDneS9PDnecq4vpETh4HY0b4E//1HaGSP+QjAHkO1ixsX5FpRK
eZBLYUvU5ZtHBxaT7HAdw3s71peMK4C3mU5eh19xjBybWl9SjQj9BSIAYLAX/lRn
YXUS5uX4OzOK8jg3sKSgrJm1qQ6j4SOiIEvhSm/wl9uEu4zzzJsNb9/X6SotDb4N
bHBeAdA19lsy9sGMLNPbd0IBSg8iY04qkr5Jlj37kt/XR3NAjJNuisCNryjihJoP
MT4PjdAOSPO0XEFBxkjUXIejK1NeXneULENQzomTZT6Qk0giPzqeJaG3aLEQFctY
VmnlW4JsG0n8ShzUDzm45CfHMexq7ZSjF2smknp5oiII9stjARMf/d4ddzimK88H
DUzmE++DcN9HmFMuGEZ9VQR8jAUlwROisa61kOUzj5RE9Hr+SdyCLYYEjZb+A7xk
ys2pHkSRRFFvrEP47obGfS3DwdnSx577JTICqd+Bu+99vQQGz2Vqpfn3rkEyYBG+
xT1gTi8RWCE4Ps0x/1h9SXU4kFYiyBUZvPEbXgbMqVZZc7yCSRCpls56X9tyMzTE
ZFyJWAqiVuyFzUTtBNZgNclTHECppYvZ3mIBN0dg6dzAFCtgr54P/YebEI5AzXgE
0gm6MelzrjsnWn4eTcMGIMi300Bg6L2tUWQXrAkSdW6/r86Si7qdI+SpTqlx3AY+
6p1xDUj2fb9Vr5oQGymn5aGZtmtim7icPjhgSgx+wtBq3Bzae7eGZA5mH8DAAkLF
JknYNZYb4sCukvWqshDJsZYn0YtlsO9ygLeW2mVMsixzwCOD1qdPlFk/LwPkv/1J
dc6OGT9zNEqFLa1BGEXPNfvj76ZAfgBR1wjTrOJY2TNBUaqb05T4bs6YzhCOOF/y
zZpV620il2MbuaDzIpykU8uO7cSKnqkAbkgvbuGhR0yV1/TgFpW3rBElkeU55x7X
1kcvGnAy96+QrgpAPFEhs2wfHdtUcJUaHYceIVqAanmAZwfFPs6xG29h3/cm33le
EnLFkpILi2qYaUwX7IkgHY/ogFBToBeHhNjulrK1kmSjAS8Mg8qJ0W8nf6jvgVg6
gDqb/tynqNhBn4i5reaaN25akbOA4KpmHcNy/Ckt8vJ+W96BBJ22oUoEAuG3cgQa
iN2wfke0H0ziH1Sxxi/LsshlAs0U4wO3dTqAaxEnN/1b9R8SnVOrCAQpMwly3vnj
jePMC1QcyPnFYq17g+2nyBANofTD76FwdGgG6RKvykP3ahUHqiMkbvpdqjlxJ71I
tG8dcaQtzt1k6LLXdkZnUX/8YpZe6/8fqwuy/SJcWiM56oujPw0XaGsmVbM6kHFd
wA5BOOXvP3WV+83y2cF5wZs3H97I1LnHRKEf1ztdzGYxAcFRdnv5xsvuTQUe61Wb
iGjpIqV9uLLtwWGzrvGQC6n7nv8qKp6lLLLiAcj7qavIwtjzj+xVa/HoDxTLBbbp
/dJQC+bRCq/HxG9eLhPJwAoDzj3igKkfd1ihjPM8BVb/57kHdTjZGvCzXU18UY2s
VFCBN2Dnpc6K41zfozl9e8STjhGxD5BtfxDnP1o44y3vd+VEFRicaAlQ8JQwP6yZ
7WcJpJYn7YmbhJZye++1+j7X+fqsWJgb9XvYjTm69u1sPDe5Prsg3i4LBWosOdsy
IgarW8+A9wR3W+dg2Tso6bF3uuFq93z5EsGf6VrdpObatRLSOaq6EIgd8OHc5a9i
25Ll3qSj9vFDHG17ZgrgDcezI32pUvc8C0eJsVDD9x4O8TNnZTOL9OFR0PXSl8Gv
oOUjkXU6WaFW124/b5q9FC++sjAnjAs776CFeV1F2Dt4xDqEyIk82ANt5iHMcDqj
6c/1q7qXrl+lFP2KKztMMh97Q2tEtf2zXx3d7mRHKl9cPdh9GPDcqU3UWtjvZGfY
9DXKa5OXQsN9iuD3H2a+wL/qpc2vQSo0/SGnSMt7H2DIGSzbDqD5y44U/2bQtvxU
bibJuV0TCqtnPtgVTT7owLSMikZoRUmwJRoSfovbIPuFqdm+FaMXW1lM625vMYW0
2iJ4GpQP+ofvxYeYNrEuJoBCQcPjQA9YhP63vKK25flWtCFM2hXL0+1HDMjzCFRM
tVif1hcYNMVXDY7W/vy0XypLmwaFRBsxnfZi/pbBRvS3THWciF0JIvZKKc1zYeaO
5HRGZVqykFvCyBVUm9QpK+ORNiQ+2ryKTR7MRY/bWHIrVoR9ZuxXBeIa1pkDfOAz
zNLdC3sKJ9oVJzfNZ1brMDBBUVw1+XwKoSKHjCY7j7oZodGRUNuabrIvpUKCyxF6
9UgcBFz2Cnca3vl8von/DFBhi9s5sQ/l2rQwasG2UX673B4S3YTXvqXXMsnWakJu
INlgZ7Uyhy/de1NH5Oy3Ms9l0/cUkmR1ZQZ0D1lSjRVYMXZLVPw1cswhcKmDa3Na
3VlOe+UoZ6DU+Ap9xrQtASbkYKWIEWWRStZUFpYqsi8Jz5e2rRRISx2vK2+vwic7
6/Hnl4a8QqN2jmy/ghUEJW0RHXK0kfrCYheeRk4Xad7c8n2YTs8X12Vl5B/zs3xG
LnZwVN9hw7+DmpmU+umt/DkFkc9Z3oeS6mjorx8Scd8aoEPNhIW9wLCgSsBxnVBI
bkkIM32FwcMqqQWXTmvFodM+l35Bt0ZYwMU+3tt3dmscYIdjyNMjlqjgqP9zr7Cl
wcY1VAKSadJDWoXNL8F34FAc0TJdsrqS2FtBdZmIRC0tvUiQFfF1fBfHEbeamQNb
Em3iwnAvYZkPt8TZcUc/jrZLBiAmD9ijiPF9wPUhUOHN1q8Kei51L2AUpYIAep+/
ZoJHRoFwQTKIBg8+ctg1880KXVNQmgc240HQtDpBTBOVhyxZtzd5Devwn/GF6ZOc
gu29hXYk9H+TL9Sr2JXCDMDjN92gcWL87vyQUUri6gewXR5i7qE1oc5kevPJyG9c
SaUQZbBDcMe4E3h2jTLA6wyHtLvrrZNWrpnwaXHXwmkKPMOWrqMDtXARcSnIMwm+
QLVt1s7QZS3ucNkAj93Xs/KxxEAUoEORk1zOIrdOxI6Y8tcSSo/AlkVzbUBl5vjI
vodYR/ihaKcl+U92ehNlv582b21pH+Ftp4qvQzdYrye0fZva0bwUvE1nhiRUX+Xk
Ov1Ojxo8TAkvjSJ2Q4HK7x7VEixtpkTGtpkAM/2pTOojzTvbLbfyQYPwLzvk/JYF
cx0lEZXo0x/tfdVUZp2kkq3kJmsklWaD2tQP/Z9GxxS7tt/8z7RyoGgeemI4Xrw0
XUeJ26pPkjwFTsc02I/07yQMuqieGyObJCFkRwjVSUblNjZbhX/v0D/bKpbagtRR
QQyQjVuoQgRLGQVWfmNojXIJWUU9IRipfazQTf0m045suQDUZEqC8fZEqwX+zo5W
D60nbYpPFRkefc0D7PkSt9mYoG2aRyxxo4WOZWFY2HPB10F5pZaQCtEYHfLFjhPg
NYjXp0zoC9bnwdmCLMEfbNKzS0oqJfFUU1O2s51q8G9EAXN5izYh47gzXdVnlb1d
t/C531Jq+ZuJvChHelRdelZEfN27b1wTIKFq+JfPG1HRhdAlm3gefsq0ba532cJZ
0fKwcVQhu44DVGzMa7PsE1D4G9/XBACKWg1uMkxIsaDdrYjNsYcRNW6KiZvb5M1R
iDOWZjOl/UQjfpPmA89p/dTgIVTOyDZ+LJCxDKygiUrrf2gxgSQs4B9ueXXogo9+
/mKfGliXUCvVMZXWkscAo3bgSmtbeYSyyMxJTo8Pw+3aucLwqnjKFJnkHkmYghGw
IbLNt8DkDDwiZhPBGdgo42uKA31iSNlwW6Pym9Xpv9yDL/M6e/8z/COX0wVU71xe
PF3d26o7SWzz7FMW7gNEgZEnDbvbp023vxztRumrMWCubYZbMv/zDoSB4PNsudyu
wfOf33FbKg6+2wV2XpjyFwNJXdC/ZXamZEwiP7w++ZFuy2Z8cSSxD8dUtmI7bSVb
saOtjPPPC/o6PL8iibFjIRLEpa3WOdQ/LgBVPh8DGHYRf0XogKdYdxRkX+mdC7s8
Q74ruy1tZBbC1CQk9aMsNKsstSkQdcanW34BCxuPvb+GvL+R5g1ImiFI0M8eAsSv
HF6hAt2BmSwU1YMkJ2EntZbOO19MvvedRtMT+VDmByGlcR/RqkXAS4iFYSARocBa
03a7n2TkPLhetuYymlcqDKNVyWBc/AncQv1wRtZ5XS0ob8dt2knxf6b0O7HfIpK8
xHL/NLFQ97X1sfPWra/P4wAuAxosl1TxdCUbFp3bxZ5JGNplPLMLYjAYUboSYIcS
PrOvqdQRa2/vFPib7r90Aa2hFhnoiXe4I19sC3aOf4GrnduQiAKsJ8h8W/+Fg8Cm
UThxeuKgZc5CUGV2HyLFCrf3i+HdGryb2GTYmlYNpQXAY34Af1/ZJFJMJAKUzETj
+fP8E6m513FKfb6/Kl+ngRuaqDmM+nkZmsV9B5JN4asB1bNrdniD/4PyBCEGc3ki
uoooE6/uurUIBn5M5MNJd0hBcQiZ3elU1HCchy8ulZoCSQ18CWfosuYh3aaCg0Br
p1HetHlxarKcLianB1tNvb2/OFlUfsmX58X3BWOlWw496as1ZA//Qv7NJQkNSpiE
46WN826AiTUxerxFhK8Y4sYOj5qqwu5sFtSkBialstB4k7ElGVIrmypmv4EECK9/
6XNLDjCbLIvgkxcWYPggUDC7V6iSLomram3ZlkT37RSRg9z2fYAXe6AiWEwHHKmb
9nFFkG9P3Tn2JvBEWlzsHxVdQHlgAADIZvDIo5xYudEi4OuhnBEZd7CyVTf83qx0
XQ83jbFMRjw4GOrIgN7uTcnhdlvc7fBD1Bes+LRwKMgvyabh7xiOX+W+oRSmbtGv
1gattKHEcY9vsAFnCQjjEvPjCRxrVId3l1JCh3ipu99AeQ+RXMtIcL00/SbXKaxI
MRiHOl+BedA32URum9wtBz9I2YO5+bNpvVYGA3hZmgS+CuMa+quaWeHovS5Lrkz7
kmk44xu3Dv9v5mH9yOMo6ExjpeYHWULEZAM9lIw5IXk14ommL7318ijOhdAGE/lb
V5sPJyI+ndr5Phzx9bmfuYDkCPUDfoMt9QJRCpjjTs1CPQH/bxkeO/7BpF5SzQJQ
Lr9UF4eDSE+x647taO4RsVNKJ9uZqV+7TQTgxBAwmVSaN/ws9RYemfBANRzxAwvt
5wMye5/fPHhoabGDPMk88dplPbKWCdj9mPuOEBF5r3yu/i6ezzJA8cbbv3z8T3YW
YqTnBV8zM17vH1F115/vRahxOZXy9JRnF4VPTerSIX1Ryv5ZiGpv53mbGxvGYQ9N
xHO/fs/F7cyWFXTFewpYzY7L59UInjyfBOut+BwEtl+b25DIaql8Fp/0m2vIjqOj
3bW9obw+SFIoX/EbQHTBtfHyAvONXb7EwK5MB24VzbJ6FiRv5ViaF1K0Gr/SPTs8
gCOeFFf4o3AGAXTHfIUNzM4Tduw2JVrBV4RDqyKaKSGshyVaLBacqc4Sny4/Z6BG
SIUyGtoE+fLSnvg5O3hZo/SfEhmE3VNy3UjN8r2Qxi1WKOlzMwTsHF0mo9/a+GqG
Ismg9uRWA0/islZjpW+i1ip7f/yn8fGEiiJemYlJZPpokwfw5xSeE2DwSWOYTjvp
2RTtuwckvFWNR7hXSazY/n9V7UXZN+6JtCgeFCUNRJnvx1SmREN7Pfw6kgdn0Seu
mWzVr4tP4W6Xwpj+sLUj4OsrCO/wzuluPOQRSp+S41d2il0Tu0fUDdE9L/rOhl7+
4QwCf4EYcdLKzfAK+1LDWa80Yk182B14Wel9W+G09FPBtOt09N+Bcryp6RFw/Iqf
7KZkbedEetWmpgUjSRNZi3iibrxQBVvUwvR4NEEyvHJ7akMmDYN/c8wjkikgXWhW
SUAGO7fRLZsi+VxGIGaiB4Empc4KgIv/7IuEGHRJLzyXo0sPGIAySLiYQn0KBepB
211s2IvpMdNRG0OFOK5SMqJvyKL+3WKq4STQh5FZW4QSVyEMhcTT1LYkmDHsK85E
97hBBFrc6gC+POSRzZ3XU2BEGefS7vg9HKWQpW6mvwq62YKZY5GrfXJ0N8fOx643
lWcuWXE83EtR8OLz/UJIkFI9s+Dp7xeaXilyuEDP38Ttibm3T0PI+kI9QCCSCF8x
rhwTEozfso9purThJzXy4uaJYfh8d+V8TTmuZxKmw1WgPk5vQ1mMln5w8VCBK1XH
EA14WZw+rsU8x7x09afRizXdmBCY0MaDbKqp3mXiC1OE6JWAHNVVdeskorvoYPKe
0FB6/pQEdf16Fxo3FO08TNLaev2xlG+WYx9DxC+q0txB9tSu+cQvCJO8KaGS1Om/
iP1BafGa0maWHEg0YGSVok32ewFoAV0ExmZeW1jkGji04hIJLlXhU72Lq837Der4
J+uCr0NJiBo3jzBw455z5AcsMLPjHYDJYEdnhEuN2VKkrMb7GIjog3tWfDpa1zrT
RY8KNx8Vm2kOPpPLQgBppcDKDTlM7gxjf1kb3oe81jXUuXGrpDUIuIt8LPycBSBJ
O8H+a31dCYw1k4RwV/skAo/7pc8aZrBvLAhPENiKTbVKmEKaZJnPgIVu4OQPHOf0
TEGmIO6W27KRPMnbQ/BB2X6p/4v+gOWWuPxQ8hveOBZBU2Yqwt/Ys3a0qfACuSGr
nNCDePD1vY29/nwrrkBHOur2zGZgHAowlK8YoU3SGQraO+W/Q8klP4ntM652AayI
3D6krvm6oa6GVJwLpWycN/YaqMqb4WwBQw2NOvcHmX0FNT1oS6thO+iLPksL56JB
pvj2dvD1mPdqRmyMR/B24heNRsS9lG6UxS396ou2oq4q5nYS2nfJa85KARHDd89t
CqgOJhfNEeYQKJ1Viw0vAGcDbiZ8ATcj4ci+Dlu0dqKRje7Cfiir3IfRWBt702S5
/2KwNdy+/i45sXkRF74H2IKg59ONW0NXg+PdtCDV0iPR972qPZX6HjfuC9N2gloS
yzbrXkDxJLukkGfDI3RUuXEVGVIEdYtQNfrDf3kEBJ6f5T+8XbbLAeFKN71Jgipp
syz5J9IGvU450DXuoB++p+1LBuNIA7ubH8idEeefU2Lb71Npk37/pGxM4iW7WVV5
/nrShOolB4U+Da9UlTUXI/LGBtBrtUZnK1rNlYbxs609NrmPeDhjoE/BebgJuIRW
8Yj0GRGrXZayFF98ArUHlJkcCVTmCStN3yPmJH8AiD+LQi9zBhQ7/oWUghV5JJJu
fDCJeL+5AefFEyMv2wVeRSAo2j6cWWP2IKs9qSAVnOSvHAKDSZpw2L950T3rI36z
dz1peUn0nwheC0TtYfQ08YJYFyiP5RgB3KL1tkBoxCL4TXUzCwVJ/AKnUUmVolBh
McFGspEwIFcqCl4UkK30u3+Q3GeLj2hGoZ/iGU3Z69xEzDP30WH7421x0F/ia8QU
FgQFtDjBZ1Zc9z8KcbR/Bs9mIUBTwuTC+eEX/NqQdzXsS/09vkUiP7e5rZsKdMvQ
GVgtCDuA9rP0tOMYfl1EHQQvQotHhhtHF1Ea+3QAPMAiz93zT1h6CVZjnjEucE1I
4egbosgvCqPpBqTQDldeup6Cs9kfbRguIYnRbBAYyiYJwvnzzp7p3eu9PZThM5RZ
ZqbAJVvAj4ZQE21UJ+Jc5vpzVs8c97BGpLXSXMUCK2nql3rx+CXGteeLVubqSmEl
VN3jsMyF4Xp+Y/OtssoUvzNzvcHtU8AdEcg3FtXs574tSrlDDo6urKVFe03MMup/
1pyY7HDw3NBpCdaiq0W87wbuJs9rBJZIL8PqyZ70D4/sFWz5bIJ3rD1Lkv9DEbcX
8ESNH39n5Ku2Zz9PH/PJWR2KXy7CwJ0Z2+FxI5P49picdCk1MUfR3LG5UurSYwC3
K+qcLkMjViWwqboyfp2neocaaoiOGMfzZ2uL0uatiF2i/XsnhSfblcUf81UyCMra
yMmxQs4KBjo85dkNVySSG5eN5LGd4oIGNeNhN7x5WtiR/T6CuOE/YtWXoxYRzAGp
DFd7EkOMsGP/DLdtVEkJ8luP2NklqNmh5Z0f6IW9M9aIv6K5EeFYzqIwsgHmWWqE
8+9w7tEbQ6kqI1LZ0z0UX0eItLIBCEWiWchr6CQgcPchGjXGQdjcqG/n/P+PPLg9
lU60P+gEnkouYnsdWWAB16Qg6n+qbFyMo1ErvOqJI0D6RemPi4ZXDhd8yjGkkGCG
pU+uS9wq6d2jt+YeUOY+AhBbj2Vk9ajPXBvZq6GM+ASVwpytwVlSfMa4t0Ja0efN
iYdXHbiSuO8yNfXF81Ynq7hwEDIv+t2tFKgrnYnC+D8wswe+QFdl7gyDAy3O3+fW
rvoBnjHq8i7nEJyWjcH16EWkeMatod+cMDK2GqtccM7TKFub848ijOLErz4dh6SF
TTOBOz1lFTr3VvfkfuHEbtFfN2UaLNCgdQJKE3X5K2tG9s46KOMpGVjR4zzwOH/v
bZ1cHTmyiKk3PL1SFOcj3R9BCv1DfQrKefSp2gMbYGgHfejmeRe3odwLKf4U2TXu
4kuMdXDNCO41YoDD3D+v5vK8Nay5l7CcVn+QDDpqvWrx2S0uQxO5jbEC1vZz++Es
an+QjtG6i9q9Hahxr7OinNqkeWWGgl2HkDlvst8wESBdIfvTk1uqd3vFDwiq1357
Pm7iPH9P45KQeIc2OJmBFjvoggYkH1QsNp2zp+mho1FbBa6QGubmwLVyuRY8eHtu
7x52AH7V6drSH/C2TBtcwz7dBJfFQ2xDL69cPgtHzML1S9TAs+Ttfm0Qm1xwqfsq
faQ+SCQdukXotA9fpKAEd/7Zi+wL9syQlHdBEXjQxo10q5/SPAhQ7gaMzLPPWxRX
8w/ymaztAK43Nq45YdhHJfmrN3jjZuwNZ0Q34aIppZUKapLwB3OiWNzNyn1R5roS
0tc70U5D/0HWk19CxiI1bpGUBogVgL9xujcqMhwlizE1AdPGOEr7T6TsXCEcSoj8
lkXEX1UvTPY1vMZ7f8/pTjwtyWMrmhmy5eXgin9OBAOJSeeYRT71+72l1zqiAwQa
gSHZgUjuBjUsJoY8BobR1dAOV42aunbzgnyFxxBoLJ1YdLmaHHHlcRQocC1gAVPQ
n4zXx3xb2FHRMhDCc1F8uUuLgCyFjJvqBGNWr5sF2RsyWo3Lai8nG5MwbsbZ8vI7
To1GuNahUWghEXui7gBXTW7WJkFJVASVdZkxgte/vEUiPNYDxt8h+Ai6+05aqD1+
8AkMHXoOkHSeKytWtoZrmc/zg5pDq1sNKWcmODhz5KJ5sswfjkLFniVgW3/dZbub
Tr997eQbs8pVJg06joL5bUN1I3ZGaLbvai7cepqAUmW7dRF4e9lnLptcJnN9JcDH
c7N/mfe99kBsYwf4PE+5orQI6BO3IeHWTRFqNBv+jaz1Joyuw1bOLHR+xdgT+zri
t99uU50ICf/HW2ahv5Z6O49cO6hYYnfwTJK66+gHejY08q117Oooekf8m1DXN5iQ
LSLLL3GrTTEHn3EHSsNOlh5Xu9clUOms4gRLs/6O8OP3ZDOuDw9xH8y8tkzeCecS
k6z6RNeAs13qFx82ucoIk2WnjIhKpp37sBKFrkO7Um2OUJHM9VG9JXIvOl/dQPtb
eJsP3D3wlG8S7YubP3p/sCejQ/b/H1jubKiWF7fWXHBEjaNIhHHej3Gl7JpHnM/5
uWXZG3tzU6yjxOYWeMpGhwPOXdEDdGrNRjDi02qK1OskJCfqMFANBxPAUMuLec6j
CHWDiE/pIbwjmfPlIwGfgbuSrZL9O9DAyxptuexm14L3TiJs4jldc/ozJR+qOwks
odqi2J0FSBNgxKyFfsUtA/2S3tV8y54f5nV4xX5nIMqU7YklQ6x/lm1MAhlfP0bW
FTAd0biN5WkzqfqilViOgmhq73MsVwaYEyewdFNo/XP9bRyxFxUt9Nupn3PNluZj
Q/hhUXfcVdIXjAHaupIBAzUgaG+GbiC1jQZQRvwmVNvqcCSvQ1jkKyN0fSzkT2sY
dCejRn4ttdeb4gBQTf1j2Qwt0jJpIdKNJMQgA31KE0s67ODMQQ531hXWO3rxXJiG
L35KsM22jvXF2VbkqGCiVVf6SB0BA5DMZdK2W8lBORnCs7cONwHJhxPkBzYO3Byp
Hm0KtiNg/zSEHJEt5qn8M6YFCILT8K1xX0LQAR0PgAiEn39BhUvHLlRy9+UZ54Ye
A48af8XJ9HSInAsPugqTEzi2R/jF3drj5hgbjgXCsZvLYd62DgHS5kmhFtY64te8
mWPpEvwqp3cFeyIub22bR1Xz2teYxNpxe0VzLZrVLw7qz41Q91Qol9k4PHY5eTUt
SeooY6fWov7IE9WtZg7dczrKf73sEU33VsiHBkYxbWGMBohJkxE40sdjLBtO4GoU
BnQPqEX//5gSXvsQTQooiComwwajFtdrVjB/Ezjc/OyuDPPIwSidoSn1oe8UivNV
F/ZrffsMe7FHniV33WSokltcTVJqzObSgKTzHuGb9IfstXs18P9Wy9zBqgBqaQ9J
ZkchclCyKTV0VyUzBSKiMq6dlylHvDAqt7Tv9tkHiRTsqAMTBZmHnjJRTqDsZE0a
MgWnCByO/D+z/xdzbUT+7IZ96raTzv5taBxbvEVomzaR1D8YaEhIJPRGTjkWuM5U
ZIwuo0y6NO393VMMVyKzMb+nTUUY8nP3q32Gmt5ziMdwEbqokAx9s4PDnNgpiPPl
ukwhqFiU/fxdmITHQ5+BVYgngRvSlASPSKikhr6j+zeVvVQyyMLOqNyNbGP7f7y/
AMIQFXiRJ1z5wnQ0xJQB8762dwZ0eWLTcU9oqxfvtCwHk9j81RTYuu+PEzwfXPoQ
4+4ZwBcXXwMqsDJcM7znnz5htcymx7REbnq1Lj31SL/Tauf67bc64Lenn5VkBi8E
DB5U1b0I8iICSHQllkVGPlyTBkRh2lkhKz1igBhU5cLQifrkfvnKlVoTtWnMpHyv
qzbwHZ7PPLe6olcOqrQyP3gmU85SCiWR3JoYGhoRu8bp/OOQApk/LZrn/T7a6tAM
yF1oOT6lSU3VMfHBI1s/gvCt46GVeHUlUWS0ZVUPZpnK5ylhc31SnbBoNA9+vnNH
50j77I71jlwyxT78a8kDfF6nu/OvA1Ogb3zOrhhb0m7Z2oX4vm4z8FiRTnGeIQJ1
mZ+Tma6lDe3678FlN4dBdAy06KUAnGY6uUL7fSRxPk6iCs/obL3XN6roH70mwmOI
rweYZjSFEEZ74IbgyeUJYC3e3oBWDBKBvRz2GFHKIiCHT3AoKW5B8SGmFm+uXk0S
30Z+IX5z3Wn1+cxt7sbMSdaDZDc73KR+wAW8JA4yMCVFy5CQ09FZTJi3bXjZliKL
mDRxKCui5Klew62a/31YZw9k4FjwgqO3TczFqsratKZuLf66In4jX6+hrP1SlSgd
cmBTOErSvIzCszapGWExKCvdYsFpHngHJFrTynRhRUlbqdE778DJ2z/QMSk1qjxS
qsnMDD+gwtkQxGoontORuWOtpGE785Mi4Jt1G3da7NjFqyvKc7BJCF44vpQhZQqp
SPfDEjjHmdGe0Zpx3gSoQu7M/km6+i7DwiQUtwnE2xYUiAeixEBxnERn0PRDVDbl
l+WNVoKbB94RMa+9tl91XtInxzqSPfnw3JXzA9lFiHpg0923cUuO8JMHRTeHRyGD
2Css2gVIrldpvvo64gPNiZtUrT99voKaYiWEvkf9jujJhEbXPM4Fk7u6UZ1s736T
14m9LPezUrD3bM8u/u/TW3z9WNfG0Zk2H+b8WCvJx4v/xhqAX0IJ8IGPBuNJXNlu
Fsjkhepex71ELTIQqYrPLdzF22zKCKtGz7+ZnhxTMynumHefGlru1l8Hgpe9Ynv9
T3o6OaW1mxo8lu4TP7FOonXdMJJDVYIXs7nyaF2yBCZIbjfIZvOmzt1oh7r+SFGv
QVo83+p1sc7pyLc8c7MLzobY+qX8tyWI848kWUPBtyckCG+UdXldtOGOu8WT4Nat
7S9s0MuUwoNl2O38ERECXOOPde5M5wVz4wWKIJXlLwDSzO/cYpeApFTpFmo0dgql
S/3tq6jR6/DOvJYUv8hoS0rQA99DZIE/YdEC/Hs0hBtVTfphGlYWubQyhefNtzCq
0Fjy8492mkx9Mp4dQYxa7TO2R8JRz93MX1/Fee9OVpjk1uNB+NNEzj8jzWbDatxF
yXFNJpRE2MPPSPhCHlPKZ+WgYZGemw7dqwNiqvi4DHNx0Iwq9NhsCgU5jsZS9HzI
EPEaa3c9kF4/iwtIL2QKXBs50bd009GtpNyyA4yfgTkMzVdn25cy7k77/Os1vUpZ
7qO1IwDkCdzq9VsLkcTosh759MlQ2iretGIz1GcdFaCYT6VwzPBimlMLkongK+nP
qdSkto42KFT5AgzuSXu0lrgAQoemtIpUW5bVNlhWle6XRJ3WeW9DH8JFcdAlrkU/
1Qw6TQBRiuL0TqYMgK1SNP830wiL4W+KtbCLNM122Hya2Y+57ArrYxArFMo/C74L
gjrp9wr5DxWZSQ7mKvhW7vhiqpnkY/Z/AdwFwsxE4gFhrYOi3lOXK16BlTOCMC7i
Ce/46r455raOMBDF/XgRZUO2jUf+2Mh8K97siVx8ll3nc/22QD/wXG4pTOqSISfn
7pJBWk0yaXGTCO81ESqnW0TlQUWyzbwkrZZ+YiodT0cDfDV7WQRS6iVICLZGG5XT
MpMyikmUe44CZhKmhuHtsEme2Ze8/YRXPE6mgfDdF2WHyB/uFKuINWr0fayruQZR
9QN6LKRZ5F1JDb2lMMzvSG4/bA15AjZwMXTQlQ5fJEz8ZQU42eAfZYf/GQPTlR4x
JMmN3pbUT/x+xOr6GQmSHsJWS8Npic0TAXVqWxkctjD1hB6XT6q+sq2cqu0+vPb1
CfwV6575M2zpBOZa4PflNx2r4iq5jsw2OLAXBvo85x1Chx6VXuHwIFZWtEgWWDbP
1AcOwSbD69QCCyXhT1im77TZ8dHCzIm7A6CiSy7O3i64K22SqGOu9IbrLdootEBw
RNKzknppHgoGZYV/WA6ioTO/9oxtJyBbSQtHLmtWmTOCwjhbjzq3HUdkWc9TrNTF
/AIQOkbmuhlQeviEnMQDcAKxXlnc2Zg0Arwm27/z97CP5ZTSvcJG5F5NZDdPHQbw
yHnJj1LjypJgCMxO67LLM21h84JgUD4bGEoHgQXvhegnNCalDZXnK8lldvGZS59H
OQPENGCc/HhkhKR48b2tJxPx2USZhGp0nTXxL1ZfmgpzKsl1SqSauv4NGMt004wl
910l699foZHzrkizhBSvmc4dBh4PtbJs6cLTruGL4EvlMRCfVdTJ8Bn/uG26fwHL
utD3QqDC8UbMU0sXrUzs79ywMeo1LuEGXaxV7NtkPEiKJhAQe3CrNZoPMv05xyuD
CSsS8XZOuc+EtSJtscCZJkDyL1cdM8S6Qut6AfAoTDE3OLT073UOEk7lz/tNn+L0
Tn/va0qiGLmAmEhLqqE+jCGJxs0KQXKSS1/xDkbdlccpuN1gHmyiQryFS58XC125
rR0eT66gQh7yfZbZxSV1P2mfvzTGTXsKhpu5M4CNf/mtEvyu5heUutqveWkZTPED
Rn7ErNQ0gQKYrWeTOScdZEtKMDrOGrCfl+f16jsmFAmA1HofDxMPIPb2drOA2ax5
yAXQ5xdSJ6Pm3/6rdUqXZp194W52ycjdMI82NCMM6l1A8LNmwMTgdMDM/oE/tsc2
AF7h6fijHtTkFOzxJ1hD5mxsh/XScV4NpoKUCLgpGUg15VmGvMe47qksvBNRfXFq
HsgVX7+0I7BFFwunRwMoX9yWjWVyy+fMSwKfJmCkntBdsx3x8FL9D9QhwcMDNGC5
+jAfs4hDJzlpCfqyh6xH/k6gtssiHLZeL3HR3zpcV2rjNfeEI8aQB60MzCttdEzO
Fz3h/kQayS06HIirgzHNkiR/p9Hgh0hHzwWlvVixsPnZaQ2w1hlMvA7rFMqee6Ea
GVxe9W0fja2eoKX990TBmeHXfvlPcwIhynkLrRPKSrV3ucSdNEd2hPwS5DBnnhRm
i4KXPsvsCp9FKYR7Zz7M5GvNFshwNurTvowwzI+EBlNhLtJbEJCuzY14dQbAx6+6
rfmzA3ZnJLTqwxA+xECMXLGJRrJ0u4H8bBF6zP+dyhBo1hvZDafAvfInPd+o/gFt
pqhAffg7NqIzsXVr+jnj/6qzs5a7s/0Lk28QApQSfHsTkikZl5B+LmV9YkLvecfy
+HYlGA5FkLIb3eVtCnZRaNmYqVSEUBSvCKhX8AM91ufTX4Reizl2RmTrlHhxTKtE
nio4VZp4kejGynWLvWsAvBRCrXopgw5BseMOUFANbzrZZKJyd/CRKX92sSVHOe+H
RFoL7bmvN6IfYszvYoEl1jmiuOdAxWzT9wg+o8nuLFPx9I+1kydXEtQcj9Pzk3rH
Wmx0vhcWI0EkgZBfgyYVuiBbe2T+Ou0xJOw/c/WPpet9d1hf8UVY7NYREGsGoRHD
uYFQg0+GQ7CXCng+ikd6BpecfxleFP2yf4SEx8PQuFGfsHjXhD/oI76bb456d0w8
vw0mWAzSM7TwdrZj0+c2V22nB7b/OHs+dQETYxznRKLoBSOV+gMeaSFM67Wqzb/z
s83xiWPmPp9tdHAsX8QbCCVCkSdMeiALSfO4PLA3bAicQ5pkKIEGMiJOgGK0wM4F
OR40Crig9vtIM9xCydstoA77jnEG9s6Torm9q8LbmUY9n3HXSs68yxDoSA6fR1e3
Cm8IMhZG8CO9DqYhKwy6z3/qF8gzwsKXjsqMS3vp7X/1x90pGNuTuoALhJVkVy/a
F9vwrkCnk/O96C/vXDVzTHeqsi5jTrVEYCFOxbEnFD9of7NYiGUB+k9EFTddYNoY
BHNmGjhZ0smmi8VplVyx4/pwLk51jU5GG77ftzszIagfmmXW+fPtZ4s4n1VYQqM4
z80TWtpL1If+mSF6sZQAJujDpbRia/8T8h5ht7eyf+L8psTVRmOiKJbBSTpd1NDh
xq2fLmnBp8rsDPrNM6CBzSPzeC0SurqPdOrGqeZnJFKBUPmsuCMes/62jrsXz+dJ
B6sYo4Gg5MlcGxY7sIohRTD5x60dJt4pzRKwgyTPrdA6YnKYBsW9nmVz2654p3n4
uUNyeXUv5g2Ke3v1DrCJe8mLzwJhj/htIJouLoVFmptlV+FXtUAxAUIWHGGD/8q3
BnQh+343mg+ocR9FYD7FY1GnybMG31PX78ppAa/UjcrWurEUmDcC7YZMhRlwVgDK
8An7HfYX4ba8ylmhBfiWuuQ/r7G1r7H3sRMdp+AEJrAfWFCiNLSaAftxfg5kBS6U
XWp63OClH81TwA+DoE0Yuz6I7XjhPTI1eG4etstbJmPFcIb8M0GPoQ0RkIt+D9ic
o/UNLQIPv6Cfavociyqm0hocQEIplCrvMXW1tBoWlkyx8njwOhD50WI294cUr5AI
K6MJ59ubtjn8wyOKKWv4XTpp3Psts5qu7gUlxGayFm/iEjWJhTJ9WNzoTTx82sIE
x5BWFMMUJa6QRsPryQjzgKKHDsm8QgqZVU3JV8F9QA6ewbkBTH4m0jS3MJ5+06Ds
CgAsx+1T468jU+jYXD8PHSjC3dTxUg7FtlIeWM+lfn8M+ENcx51pMNP5TTW8Up8C
SNsnBcznEQo54Vr5Hmv0ozigIEwAs8DF/ChQLnoaFLW8+PqQ2WaN2n/eDt6n4Td2
GIbcb8U0L6ZyDPc/sGu7HheJQNxoG8spOPuJvjdN0RiSBe0dTc4g7qq2ZTbXsSPc
yeIM+Pd84QQ8jzUjsvrTrZzdUYzkx6oEAMr1x23GaXeKwYhb8PzbX1Kvf/gCgbee
YHXXBGMnvixFbU88qLWOtHJ3IR2hOwfs6lFWZwXJQZBNSBlZph2+mhhLSgDhHsQa
UPWZlHL/OlacCL12Bk14NqRPYiLKqWwCqyOaf/c68Q+p/PSLFhHuEF57IFNkltP3
216kOVsBsd7TWLj5oSzfD+HY9CqF7KrV523i7h8ufLlI3q/H7oKLNzwwBGPuhRk8
Zn8pMplUZ/GoW+MV1f/KspHeQQa4hKxMywf4V+UxkIHqq0GOjxrkTWs04JHE9Xlm
9VBPR63VJZollcpK/6XiRZA1VhjgpjlWNQjZlns/uNwQ2fw9GzvFgLCcjLBaBcBQ
V3Y/rRplOfuZouudZTCHfH8jZd4Dd4uGFu8ex68zoVeZAu/SFQ7ComihjT3oUjXj
c9hZDj5Lc5iHeeoqvevysfWNSL1i7Gj9dZURIJkogN23nW14aSdNU4Xi6sQleBnz
4ZksZQ0y+J5zv2aLqaigtcA3tfCkz+N1/e7aioheuPDJhnVOS58oM+d3iFbvRA3y
4YJnzey1hnVFuXUZqWS5BZwPFxtoGWQYZwzgRqCCjbDNefM5LPPdqTVJ6cViboxV
EeeHhYJi0RrLKZEhSn9THeAW6ctKMboMpQ3gOLcd62gSthhgpvI+iCp/rafZcFNB
ce6X1OX8KzMzSn74cG5GWG74QOZJ/mcaunuTMChpeG0aZ8kvDB9UhccLwJ0yCJ1o
N20on8LqRbV8oLSW8dk4P/UwQXDO/IyN49FFSLLe6nJuH1G9C6BqIdmSnYAaVqxY
mJlLvKh2AtsYY0bs6SXmw1l63eUGx6wGWeDJiOhGzuTz8peFYVbNz9LgpA5EaUbi
DakhlM0wZeJieys1QTMUu03ttkVh2u4pc2dE8u2jmK+D3qMm0rlxvQuZlC9UFo3V
hwQCpAncPCioclx7QwZZUygtqAsyGbF3YYLJntRqAYyofbdRqdhYDENPHvlQoaDr
Toy7rkNKf+URTOK2UeU2+McvMvEBZncf5rI7cNwB4RwVSOJWrdc/eGpPNm83O6Y2
wZTglZYgPU1/Wamab+K/yHcp669EfmB17PcFDlluNUd8JdxTE1Hm2lpRgrOAPA+Z
jQGBQ5HbjuXq32d4C8KbWi1nvBvXJMiTXyYV3XO3/GjTuX8FYoCwVrpZ6jiNF7ak
68PUi0TeL2na4Jq0e1Ym4qvJqdBAfU03H+CL31S6T7AutjnmSykKajlgZM2LtnFQ
NipPJ8c/fSYYpvjFm6l7s2KyM98o5c2P5yCt3eGgeOXzraUQrM10SiSu8TTp9LWc
TdHCwlFJsnnUqC9xkZqJloCUuenpv6eSgV9HbNGH0EsxDTDJaGQ/cYTqust1DI21
hQ2LqBir93LS/ba64Mw8xhmsA5S+VzLCqVAm4PAZ0xvJDaP/DoGt8aHAydYXT8rF
DDqvIgI/PRLLWkENvIXAhNOH8zct8K7LG4fwNy45Hvc8F9PNipdHpHDYmfhngxz1
De3TU0rbelrAxZPFRTIX59frK6WKgOadsG26DPZaw39m/ZDa3xWzKkM5462XsAgR
I0/EKplXu+W41Mn+QtBJdNnKs8lwzK2cKMZcySlFdn6m5ynmSBLrOMzxGiP7LwpA
SquMayz2bLZBXksQEoYsn6iax9zpmU/sMMMmW5Hkyz1Ndr3CpfFUSv7UawZ99X4V
RavuoWcYF0eMRFmcvdP3tzvgGtkmB5CfG0n818MfkVGpNvBT54krIAYjjb2t9gaL
KuMDm+MaO/I7iqYd7bE+e2l0R8LDtfZeFLEAB9bKwzha2yGeSMTxc+Q2EY1fAv8m
T1yJHsZPlDQgF27kNkft+0DdZv5OPgvDtrQjbi34hMYdY7cqttvaUDsyRPI1cE1o
KQ1B2xJzpSVdsGwrPlwO65jNy/fEbqNAaPKH13WvCjFM6uH+K+wU0uX/tWbDBkjy
Nu3J1W0rvl37dWLGuu7GzQoRZgdtH+uiSQkoc3/FKDCsj/gWsIZIJg/tyLJTuQ7u
SpgE952zt3io/mMW57ZJ8J/jBT4SwI26gHGTcywKh9BMiR0qLfW0/edtFBoRCuay
3LShwKIwVu9YVJTmDdR4983yngytV900I2tA8/0GN+N43NA7KSOw0qP5FQNajniQ
3wyBWgPIi4zl1dl+9LVVqprKhj6tHvEooxP/ylgNdIM+LWdnvzxw+kN5UlzOWFm+
JBj5Y1IQMIuGV2zyxhAaY9/h1XSDcMXQTkF8Z0cphWVbiyhSbphANLtzNv9dzpNq
CnOUV8hNCIP91OqtVpNDPBts9DKj1BTWy/EMg4RVRFySam9ZXst+b8trtEpCFNnK
uDQNMBdXxZyYSjTY5njgFoRTdUnIcHHr9cUjpj/xd6nebAnrdYK7+SuDfIzqLxPv
8pyLc3FvVKb1/88JuCD2RxjcqX3zgO5/uixrT3BDhZYEVLiEY2m4UsboKOwA/tZI
cLSDfa5rXl4gQB8kHHdUrjxHF04TKNKhO9XAWtaE5Fi0BfhoazKPrG7aJHZy+33+
lAVTAUcAgYMwInw86Wym7p7vkJA+VMFTiPwVRuJ3llurQ8MBzzGsFh+cGuAjXC9N
ytjyY2I7yHm3eD/1EZR4bXxKLqfGCkhf8VVgKpg5tRbcM58qsREomvDXuSIBMzol
ybuHH70gNtECRg41FSrKwnd4Gd1H9BIIjZJlTix4gNshjeVMWYn+L6nR1/5dhcUj
BXBCT/0RjFKQu0LB/TIDrcQBVyZKicFk7eJiURxyM5m+ejQxdRlqoQ0+YoXh3sT7
XR/hVOwE573kbEcOJM1MeMs7g0DBrhtUPh26pSsFRFB+wlqw1sEu2j1gmk1uCZUs
nh3um1RKgMnde9FFtGe9PgiRUGtPVQIUeDw0EpzWiVcxKHaYztOwkzj2ZMAt/49Y
CufXZBGucaVpkmOW25s+GCZw/RHIr4Uv6KMrJcUt0ehZCATJhe0PNulk3vOTwx76
tutSxeHn1jpoKLK5WT9knoPx5kBMIuzTrEOk+fu5OuO2uwTjebulD1nvXLObPehy
kEYNqUxasgvZRTMuwuucD1r9jvqP9J7uZT9eS4VHPJpbip4Sjx+btQpmDerr2VVh
jfdz0uvpEOpobAkahM3w/zIGzgwSp/rcmWOPotWDGnxWJ4ALYSf1jRnofmrMPhLC
uPBpB3q0MeeasANYiADyz0LWb9ucBzG0LkyavrpWHKubM+06hNKP7fPJk068uvvS
uQ8CUJ9mmXSAen3YlvjktWYLnAmVvkqrapqDsLSk51gtEIgCq5kZtlY3tTQocA5g
00cbklTdDakEky40xXyiXct2zdZFVgDE3iY0iRzKhsDgBo/g0MeGuKY0c8NpKHIL
g4HAMpYburtSHUQDtoTeGrfZPg4aVY10gZi8whkY2C9GCXXbTsjfQdOwkYOFY+LY
fA+BZqDHqghWIneaJvkWUPH411Gdzwc/1+rnjg2ddGvPNE83388eaqrHmYDTKijy
b1UP2u/c+Ypn2SfHjDi/Rh8gLXQYSkTjBu9+bc54+ULOxT89f1q0MUK7leUBZC9r
kX4QCodHwt2euNQjeOFb4nfoL6+7gMef2mZB+Z4w9T6V27nfqsdCvEdpdMlMgW6A
tn89OQbwIJvOeZvIpR4pER1/NCOnfiige9UkmtsGyU22fPS2ooIEqQKOETVPGkk+
lLLrgeTJqAmfzInpdxjz80M6Dm1tjwoTGypv7dgs5ViYjnHSMYY1o9WPffrXvqkk
kHCZwb1jKKgWDYm4eDdBCg2s77uzzRHMIUb6I3WBygEXT3a9++GrPbMIT56/+4vR
3HZ+zeqXJ58A6wgOpa5psYT6B7tDxXifCwDBfFaWUJpAYaXJTj6xDRHov4Uo+SIc
XsNPvfaIpwo5XqNEMjfUbbCi5fCWbt5b43sdqAgYpZ/ftE9L7gOkHj3GhBTPg+XR
fL1SO6Eq6evKm+nr63LeAy7P5c4fTAK8fc6rtHj6QjcVXNbnFR7aWaSZPOPSi70x
2BQwQZ0/ltM4Z3dZ3HiO8jCCA1pWMcUYeXz6yUrIZghSE8TKXd7E99k+Ebh+9g7t
kORcXjc1k6Y7DTLN8723BXfhUPHFITqPzki4xZZdN5wpN9sLThw45arqbstO+eWF
XS4Sabv17ay8edQfUHWYuCJ0woCz4EUNvmI8a0w3t8hMAbNdOilVa31G0cPy2AZa
7xHM7piYxjK81kOPiRgw+0Xv+DL9ky6nDCdEXTPStYey3zbk3ShJq4ZJiMhSIzXY
NRPnh5sHBTNag2uKOCgk4jHSp47xUx4bYxIpt8CcBKxxmDHnd1vK4mwjLjA0yL8E
h8U708JXB44tt5ASoV9kRtNHsMbJZuP+kr7nFW5yJJ/xt2lSJ7mhXkgXTNXPsVws
p9prQqHKXsApceJ+oWZGYXpge+JNp4tE9lmP2MJT0f9WNJzjM7gegS70KUfEs+P1
6FbeMNNpLs55cBB0U/3SIZE6n2OUHBDNnKx5rzeoV6IJ5eTW5bk0IgQwKyJsJTvf
VxKqNwIXY7a6TgfsZLZ5vvkK3tRkxsN0kQNcg4VZgLnjcmu7lHGao3Oqs0oWx+/J
6SPodY91e8MIka0DZ/9gqBdJ7oFCHvm+NBYch39XXzU+xNiiWn0jHuG72ljt8BZk
NoJlNy6myhJeT2LzQUSg+5nIPz3PqaLguFIVx0EywSJRjZdVzoBv5gDQSKg5FlJD
J4IdNdFkUil0/25UVuCfTTRfEp79Sz+wcL8uFcjk79uIvchGXOpyaDKZIfuK0dA4
rTFa0y3rmTKEEqLmwqxvuW5ixV5+svo+RABEO7qybNYykv0I2umNZEgUHocCwV6C
sJdXIyRkASglRjb1piDVhklsmezEkvaDm9hmVZM5ShEf1pMAoBrYSJQAnaY/gMVn
g+1WWFdwps8eAWAJFTTr9YI5U8NYKXIr9iepLPLXyAVK2H/vKoMzCFL5m+XmT1Sq
v1z5xR0/qoEZuqks2hSsOLUoQEpda++At6dO8kKmqOyY4ST6D73dkL7L8gDTpy5L
ebo0np3No/K/sSSb2KbGohSaOx4BNSdKEAshsFd54GkNE9HeyemepZPENCCmsClY
lIPK0sS9Hkhvxqlsbi3z0zh5GGkg/exfiEr239EmDh0JuVmG2EryiweMyaFaSKoH
FUhOCFC70vQd+GWx8aLsf0Ga4JJVcRBP+ifA0jnC+fkM9tMNNiYqti4+FtDxHjlW

`pragma protect end_protected
