��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_%�=��� ��}��v�����L P{u3��_�4�]�2(Z�kB�2�ׇ�T�fay�b�=n��p������1�w�L{+�+��b�8m�Xm�eذX����dF�a��ے)�����94�0��+{�̾rO��[
���/���@VrKFCܪ����<��"+%�on�d�+\�_���ګcޥi��>.�=+��p��E��K%&~p<b2��s��I����b�}��>Ҕ�-9O����\�(
g��B��)��P;� �Hi�|��6ΪȜ`���>pW�eGt}Ggf����.ד�[��JPa����U��9򔤁+'����X�s����y.�7?}`Ӱ����~	�+o�p���#�E�3l>*�?ϰ�������͚U�7Z�>p�~�R���P7�)]�эP�=�ii��]�"�3�F�N�t���B5+h�z8�)U����喣t�G��;�76�w\~+7�m����T��^��C��<�Rsg Ju�Y��b�׸CF�a�2�5M� �g�f��N=�����dZ>~����}@D) �)�������.��7>��Ҳ�^b�u0��"0�w'�X��y����Cr�Gn*W�J�P�)L~(���?F'Hp��u�h���z˵��.�!�߀o�]}��t
Ю����Ng�F��<���� G�O����O'�?�K��9qO��mu�@�0���j�]�'J�A���tƤW�c��.?4���~K;��*���Bj�ք��:���y�i��=k��}��E���'�7�u��;
�L;ӎ�d��ͯ��HQ�9��b7`k���13zh=�^�<�ٹ��-(��v�q�������8<U��^�ڡ�DDQ��ͺ��3h6�H$�^��T�)'T�cP�x�l�l�a��۶�^�Ni���;F����h`��Y�G���L���.Oe�ڏw��Rv�G�t��22��N4��y�������9��Y�ʪ?�jcn�:POJ&��VAF,T�6ws����=���5����B>XA���2���Ŷ_&�<�)hA ��)�~�4���1���T��JI����KZI�
g���)��`9[�*�
��ȅ�Ɨ�ᄩ�I�J�>pQ�8�K�;8鵣۲�#&kI� m�l���߆�j) �������Z���؝]��^���#b���|�e���]�:Z�� x�IuP:�*��
!K*������M̷��6�c����?Pz�.^3�5������V�e���� �E�͗d<O80y��e_���Ս�"��)�h-�xE�Mu/�CS�I��6�ܸ�IȰr��LĈ�R7��šP�i��^I��g�L��q~�@�c-㟛�T��x��ϥ�K����I��U�� @~�P~�/���L�Ȋ��~����Et���"���U29�Rν�N ]@l��Lp,��x�${�@� -Q%CO��
꿬�x�������p��٬ �(ug_�XH,��~��i�a��	2"����H2��i���1��o�!�NVEV�d�{���8�me�����JC�3CQd��w�.�+��6fV��[I�S����-@�bs�L�[HG�k�Q���WC�~�4(/	^j�j�����JE�]p��X�yѕ��J���NSkR�9�*�XRg�)|��7�K�
���:]DY��Z�L�����e�UT����؏<i�4�������V6�V,�h�c��b���v{H��Li��ަ��e:�(^��'O��&�����&Z��bKfP������ ף����/Xݶf�� +�7�O`s7���ՀRo]�Krx�>Ul�ҍ�B���<Cל��{�	8oi�*maJt�jK�F��{��9<�'�Y��y ��W|V\�mUJkƻ�G,���a�:�,h��9c8e�M9sV�3����*��21ho����E�"e/�~��NMħ����k�џ#���
=9bbƃ���3���V�Y�Sf��	���
��x+5�!���kq�T`o`�E�HkE�'�Q��G(Y�!�Z�0:��;_��@����������H���@AM�{����y��U�޵㏘��@�^���Z/>���X��-�z����N����m�=tH���&(o���y��o����Ȝ>��?T����|:�+���:i)��̚��q�{�d�ѻ���V*���n�V��7d�g�Ն¸}P�̹K�h���� fx�����iZ��c��"��J�b�|sT��#�Ĺ����w������}C���4���J_�j�D�or�21��o��_��d�*�Ű[&�<ꬕ)�h��R!��0�v�TlGT��e����߼�訦���tg��'�ǜ�&g��L���k���QS���T��ge�7𰤌���bW�|��I�wVN/��Rx��'�����6�.5,&ԓ��Ml%��v�`(7�c�m���5v{?�3�Z֗���V���-�g�O�6�,�Unn����~'����|Hp���P�R~5�9��(\4T��:��"d��h+��X|t�+�5�k]^;Ly-��˄Đ�0O5{g���<��e�n+B���q����f�`9Qu��C}��4���6�,� `匔i2��qÍ�S���w���+�M�0pAJ��|��{H�C{娬����l�#a�C.S�6j��V�|_����C�E7��S�����}�7^TPyk����p/�k�X� S{ʤ�P�����D�[e����M'����T�Nˍ���K�Bl�\�H2S�Ya(�Ȥx�45���&��X�RN����	,Wm��@\�@��`���fH;]3%
L�!C`�Hrk�������au Zq�P.D��׏�	�_�J�#(��2�����mе����S��/�?aЁ��C�]�ܝ_/o�_��|j��q}Y7�RK_���?:���o/���4�bF��q��p����?o�ּ�)ZU�Ѱ$���/�H}�ɳ�?Yd@Q��ϕ��,��a�z�O�JC>t�c$s��/T���<����O;c���*řM|j@��CXuG崲xP$�}'u�B������j�t�:��Z)=�/�joW�,r2���ܽup{�o�ճ^�(�ס���})t���h)����Na}z��L�Zx���b@{A$H"h��w��a��3:�NJ�5�L{\X�`lU"`��]���v�1ܮ��8���k��U4�Kν�઱zR�pt��.�D����L|�i��F+� �3�m�p���נ�¼סXM^v�D��т#,x�ī�μ��xq!��Z��Ȼ��*웜�׻��](�*ǫ��2��:�Ma�{d	m�E��P���ړ���n���0��0Ѱ���;�#���s���]����n��G'�`D|G�M:�`!�\z7�FK:9�p91^�* ʒ���/kD��­�7�$��%��M6Ƕ��J��n���lu��� 4�U ���}�R�<V�<T���:�uUnӷƿP˱��?9���s2.Z�e��Yz�`g��.fh��MTX��i>����lF���~�j1���f����������mQV���<g}�*t�+7 ��<[���Yt��q������K��<��]q��ۮ݅89_+�D]��E�OG�p���`��ẽpVC��H����l��8�q2��<���r����ֽ�������0D*m��+�%��z�"@8(�,P��7~$����[i��\��*(UT�<��i|:�����Z3��J{�e��H��ח��x�[.��179���S���SM7��Ü�y�c5E��Ia��!r7����*�¸� c3�S��ӿ�^(�l�W(���`�����Cu�!��"�/3ن�ғ�t��Gw�Bރi\�hy2��oj��5���P'Q{���۝>ݒｐ�uC�ip��!T~<�;�;�ae�օ��Db_�Yk8�B�UzR���9�D}t٘����#��:�W��k���mf@.t����㩹Up>Xzp��I�*_(rj�����4Ń�Y,�O�BU��݆����5����]���5Ce��2���#���/dEE�}ֽ���N��߄3�����䣤��}�Z:�{NY�7�;���vS tŮ'j�b�#ŭ�i�u�(�#$�
��\?�2	��S4��'O��|L[�� B�TmȒ��W��`6��O�]�� �����n�c�E:�b�D�2�8&$Cl��[ޗ���Ԣ#��̍�,�?i�C��Ij��U�U̝�Y�|<��O��[dqG�~j�4�pp�`k��$����r�}m����<�I��l��Q����h�!p�ּ�����-<�t)K�:[2%#���������z�}s2�Hl�����M�_��sCz#����B��P�
�6��wm�Z�xfDx�\!�S�ĝ#���m�,b���5��F=9��_|�x�$>����������(6���2G�� ��Q�Z:bU���ߪ��~��J���G�F,��D��Vy��|�- :��1K�������f�I̺��W��Gy[�x��Ps4++�	O��p+�?C�%��R%�nTˮA���u7��l���<$�w��UJ�#\�CX&��9���1F����ײ)MK��K�gs�tf|#�~I�Vm���5ߗ�N���t������S};�/*!v-���9�����W ��LѸ�x�-�V��B��O�q�8jM�l1�e�D��	�j�?*�t��O+&X���|��lS���g~�}�Zi3g\��!�WýN�ry
n���Uv:p��>�T_���H�԰��nZ�"Wq3Di>�`�K��U3hU|���U�����f���#� �S��b��+��8���ଷsdn53��uN��������� T��E�6W��@�1���ITO�c+���02���\m\@��"*����=Mo	�@�1��o��e��^���nұ:����"s��#���o~5� %S���4�I��<�M�8-Z=�e���6FM����w|��U9�P�*��[�����[F�����d�N���;j�Y\͕I���K�6*T��=� ��n8�v�Z0��$�_�]�O�D���!��5�N�lT�BH�����	t�]ȇ�9���t�-'bt�h�J��j�x��r�&�/�\��ƨ5���V�����k�9#z�bߍ.� e�!���9t�R��w�������� �$�Ęȉv���B\�.��Ndi��I�6,��`�ɘ˪iG4�%�~j�+I��D%*EB��$��M/	�c��~���M�;ni@E�M��-���U$�"ӄuc���1���|n2��du�%'��)�����&����	�Q���,��=����E�rM#�fj8�ev�X/����I݈�s^�G��f��r���PQ6f�W���U<'�l
?�}u�wh��b=?[���6~�tI���k����T1�+�����5�D��R���(X�d��ӭu�ՑŅڦ��(g�S�9щɯ�y�m���:n[��T�UV`���C]��.�R溵Z��*(��!:�����}e��/�]�v8�a �4>\���J��.�v�D	����ΜU��P�r ��+�*������>Y����X���l�B��tm`vsX�e�.l�I�MVG��<�ll.��MN-	;x���y�,M��L{�U�C���Ѝ�G� ������i����Ujب���+8#��$�X෻%Y����COL��&�tX-`c"�<���R�F���eOq�A�jˣ�1��t������.Uwiɖ�:�S_>���t��*��Tܻtl/�����%(�}�9���7_�;q���TY�s8z���N���n��v����oKh���������Y���ڻ���q[E?M�=�i�����y�w��
V�/�bjK���	�kX�V�z�ng��f5���V�[�zf�p�/�~�����ܲ~+
[��WgU�Ks�a��d�DfaQId�|H�+4���3�<Q�8_��.��rm6��Eֵg8�	����D&��!�R/X�ڳ��i�q*̙$�?Lt���D����|�*����(U�ZbSI��8]���ng����`�{y.~��ї;65�8>�7���^kE�M�[�:@������R�!�gm�f�mv�DM0�Dg�:��]�;}З�Vf��[��:�q����Y,2<�#�?��ȢO�5�9=g��g��r���jC9V\�ʠw�W�����r�}����1Lh��%K�2DM}�B]ѢD�>��ul�c����ӲU���m`�E/�{34�P���X�1Ǟb%|"��琵�ۙ�.���b������_�Mq�b5��'ѽkB�Z��|Ӈ�Q�8��n�a(�fô����X���P�TT�X�5+7%����~ >?tL�)�VrB$�,3�����ƓF�7MS<���4VVo��qk�S��$ D��DI�V�*BCM;��s80򍰋!SVn�j�51�|�����ʻ���C��*9�����I 0�8�N�0Ëϟw������7Y4!,���C�{�Cf����ă9a\�s�׃��S]o�4����K�s<h%�]6u)�gl��Ŏv)���3M+��i �{p�>77>�:Ï���wh����<k	��6v[q=	���_�&�X��D�7�'K�N,�P��J�~VHr�hB��`��E���I�x���¦>�w�&���_�D�B#�w#�f����7�䐞����� t�؇\��`�F�S։�%�(`XPGu�6��Ƒ��Ћ�>�Jl��5������0�-sD��\�3O{�fg1xQ���Q���A�`��FVٹ�q�<G�Y�-��4lIr�wK1��f]:��M*�����T�Hk s�cN]Mg�^?�c[� ����*1l0����v�/���o'�"}�Кu��b+,�+��/r�g�wH)�e�n���7�E�o\�yB�=�O�,8&E+W��傑A.Y/73�P��h�%i);^|����˪G�4u�'U
�t��H2#��4U!����~������z�������zCrt���Ksb����eK��(l����ۤ����6ţ�q�>�;�e�\�y}r-�O���y ��N?��^�JQiSͅ2L{�n�v�{c���ԗ��*<̝�?�kT���:��'c�4H�۪����;Y.���)�����ѴF���vc$��
� �0�l��+Q=��7��de)�~�h0��=BMs��}�h����g>�DQ=��Hbf��(�g���P*0���_i���"=��O�p����S=���B���MU���q{p���;����%�ʊ�X����S7TԞ4lJ�����/.zON����tf
j��`��s�Yt^�ސ��vk��R�v:qq�ng̕�]Hɝ?�W[aP�*T�]��%�{c��SuV�N�|�^ټ�_F0��J��*3����:���
�
J���
�b"9���dih(��90�W�/Z�*�I`������=B,soi;�&u|����x�^�O+�#� d2�<��F冪!��7V��h.�~^�BC ��@	r��ϒx|&��c��@��s��H�m����R<�X�������<�I��su�T���*�)��&�Dű��X2�g{nF�C徐�|�S��������������m�O@�轅i4h�Üc,s���?�L��m4n�z��ǠJyTy`�~@� ʚ��"��&�g�����o��F+���rǚ���_]jOقś;��%�+C�y�K��ꭵ�>��meoo�WF2��sJY���p=�e'�1��	�C̔�_�j���	�% lgm?���i\�>E���X�����a��a`2�/���D������\����	=D��4�#�)$���0�)C�a\�C�E�Eϟ�8��:��^9���=A�m�W�g��`~j�� �6�C��)\�F`P�PQġ���?
"Wýn���"�O�2��殾%���	�\,�X]�a�H�8qv�h����\,�:�|Ui���1/�E$��B��� �\��3\miʉ}����<�i��f�M9_���w�˪��i0��J"�t�uw�nt�����sOS������p��H�u���	'�?���I&mR�Wo��,�����m���uҥev��7��lZ��k��7r%�`�&���m�]~;���3��f?tڧ�1�ϖ����N�7ut�7�v�2��#!ʜ�6��E�ٞį�;� h��fv(�[#��ߜ��S��;�y���>����PƃV���Ϊz�§ߒ�k\U��3�gԠ��j��:���ڐ+D�6��_�2[��T���M\�,��8?���p��4u65A�rgc�%�v�Q`���](Q��oݨ�;�ߢ�bTc�����Q��2R�e�A50A�}_��ܔ�����}}�\�C@�������~��)\�-�6�E:�&��X�XA�GQ��-�&�<Yt���R�&$yc:� fL<x�)p�)L���b"�x��%P�(V�x� AN_<و�_G�f#k�����:x��f2�T[���.]�����I�)�o�B���.r7-VybHπ�U��&��S��#3��g.�q���=UsQ'o)8S��P�l�)�x�:��B�nC�hk�U���(���L*�E�u"��6����1n<��{c�2��bq�����o\%-h�O�1:�8� ��M;������0ho�$D�_�޼q�5�a�rstRq�v	zY"M8���i����k�!���`3�W�%���i�BP���WYEZY��vL��Mr��5�n�UWÑCm|8�~	��\��76��m�tBze>�� �4����-�� �?��{��,5�sdo����qo ��*�_���Me�W��~�d�d9kz��^\��Q9�(C�S5��\�1�h0tj� �y��Jq�a���#X~B?7za����O7���v$�?e��'�.�A���!�(�W�= ���D2-9ni��20F·�Aq[)�l�j�I���q�2���$��N�~�P���똌S�j��ɘ��*�9��{�W�M���1��+Z���]��>I��D��L!!��+���u,��K��9~"(���3>���1�s������Ԩ�B�`HL��+Q��i3&�3�X[�1�~P�;р,ύH-a��I߬�o~��ql�~��9�,��1`�N���يc�x�%@"�U���hGɥj2�<����8�--�z������3��=o<���Cfj
����@��L�! y�� ���!</5�~\.�>_h�M6Yr7�}8���Hj�3������V}������d�ͺ7�k���5�)�Cf���]�K*b�c<�g��� �|s7Rei�~ީĘ!�	����Qj��l�2����}h"a�Q`
)�*a R�X�D���qwq�%_%�pp���Ց�:���k���J~2�Ӳ�pzJg1\�}dp�r�S�A��ACv�J���V�Z�m �yAP$���)G�o0��*���Y��@�>,	�������=f��ԨR3L��%�:��D�f��2`n7��D�	�5�Z�Hv�%��a^6Z�[�Y�B���RA�[^��~ٲ�`>s���z� (��זhl�ю}dA|xT��Nc��ч�����ϯ�\z������=�3B�G���������ȸ�]��T
W����:,s��u�ሮ,O�W/,�_"k!�����"�:�+<�P-�,0q��~�`7�N�9����vk2��5��֑�t!��!Pt2�ҥ��������"��+�i��*~=K�)%yGS���Zx'��O��:�m�JƟ��\	1���a��$輭n�e
�:�+��'�oc?Ũ	����46
�Y�dq@�|~z/F��x�/<���4���fk��x���^g���C��	=��z,��ߛy��s-��V�ֈL�p�qս�Lg���yj �4J�Ûl��V�<��D�3�p�.��ABM�/^.���:u�}�T�N����b�$Z����ʖ��zW�D����V�t`�%2�����R�~�-ޱ/�#�=�f��Y0`��*���[��ct,�b,
�!~rg24����8�J�0	�F�0�c�S��tC1�g�����)/������Fu(�,t?�ծ��mM�I�bA��|Wl�e��(��[�IvBlS�6���_�d[�W})�r����6U��XQ��I�a�;�4,
�)�֠��<E�� ������䐀�t��ҷ��״I�cx88]���G�F�p�
T�A�!\��1�vQ��!�������� ���+[+��6K�{0� ���W*���,O�+@���4����pU�{6�4_�R�<�J�&���Ω�|���L�^.�����f$�<d�h�6<I�LS�d5~)�0"~��:1=	�c�.���N����G�P�}�s�,�,œ�h��@z��)�x7���@��іK�����;�)��}md0��
�\���,1Io�\��t̰�Q�������q���8kN��w	��SF��Cm���r��n���s=��v=���� �e�<&/�_�� ���k2x����u�.ȣ�͡N��� ���re�6�c�6�8CعH��Z��zen�q��o=����9>} /���f㐫2I[� p3�=N
�|���dz����]�DV[�V�p�h\Kv���s�sc�1'W�(G��J��TN=�J��Y�'���bi�е[n(��+���IH�N2D�/}L��F}+�X00��1����0�r�j��&��&W��9�D���Dm��-^_��oP1r_�2��X���zld��8���ފ��{��C@�S-�F_��*=5�)�"��ͅ2۶��ȣ�����Ѩѳ��@Ji�E�`=�`p�"��:� �E�臐΅��j�i�yi3[Fn�alɊ����p��0:���L��	kB%
BGuL4�7�%S,�fϾAb���־�X�0�;Ҹ����)����U�$���_���Ґ�����y�kic�5�TC�G�PvW����T<׫��)cō��9|�֙?  R��WH��B7iJ!��=�I_�eq�7��;��!0�����єԮ�oP^�7ИۻZ�	F��IES���m��'�*�)���Y���.����į���Ī|F̔z�u>4%|C-�|��d������z��8a#�f����[�� ��~���E�~#�kЈ�ڱK}��L[��Ix��q�Q��'��ΐf&�{<��� ���P� ۱-"��7���g����Ã�Z�^�,��9(���<���E�O��4��VKG��5���r��P�i�C�J��Z�j5�X���fc�y�A��H�	����Wv�Џ��D��P;�b�Uo�=N�L�֜�F����@��ɿ���@��+	L�-���F�2`�={���J���f�T��G���KS<��ݎ>IvD��}��Xpkn�KQ���26H[�+z�
0����f(W�u⽊�"hOGp9όǞ>�3����h�.Q�KF������ �$	i��^d�VD��L���jͭ�i�r��}�÷�VHʶ�Cc?xPb�V
^�r�_�䮫L�vNvgݟDM�k�?��3�Gq�O�Ғk��1H�4l��N'�*IPӨM�Lu{�~\	���������+�D��|�/"���!�ք�jZW��
�uV׭�A@�d}���&	a$'��I��_�` EӖI���.���u��(������T�+�1�u�X"1D�x���YI;�Nd�3�V5!��G"vM?��4Ę�j�5#��7���M�`�M��K�y�� VR#��Q -�k)H�|�4V��T�an����E�!�S۶r8��=������ܷ�|�5���7����e�;"[�K���X�&��1JCQ��X���݄�BXZYh�*���\�Զ؟�^�4^֠���J��mQ<⠾*��p���d���ͭ;̽���0.�I��'�Tu���Չ�8 ZL��trt$M��'�r�D�73;���7,
�}8�����6�Ё6� ��*�dn��
��չ�~J�W2�_�A(-�R�/P�Ĵ�I/0ӷq�) g�GhQכ��C��1؟笘O�&��'��~��[57�~lK��ک�As�8����x�o`�o\�ѿ�E"�b�u�t��i���NK�����f2��5��u���Ē�2Xޒ0ԥ��,O�r���4���t~S��J�y�<�T��j3�S{s�a���7�	�|�R	3�b)>_������-!tĎ����c�}'D9�(2b�lD�{��^r�~4��˻�|��f�������J�,�}_����o@��4塝)�A��BL���h��u���G�U��W�~�P��m���]�r�b	�̡�� J j��:\_�l�~��E����@4Å���������|���͠��`�F���!�nD&@C�_��<aԛ��_o!N7+��L�8_��?�1�Б�j.�i&��	נ�6�Sg^ن�7�~rtB&bS�l�TP�T�K��Vi�Y=��;�7����Pr=��a�S�3�����Rc-��� 8t�ƔM�,
�2�g<poc#�bp�vU����!�t�*&ƌ���y��C�^�Ċ�Z�_��:�,���Ґ� ����Y~���2��P�qBy^���6��=����dU���_���EMB�-W�ܫ���V~�z����IԼ4�ZU�K����gR7���q�ʕ;߁�W��)�\� !C�c>A��5YNZ�Bz�Q�M4;�+�c��#5����<$\M3�\(��鶷��ͻ�W!�D���ă��葹����Ƒ/�2oM��X��D'e����Ω�7�M��W��u���eG����D\iX]���b|� �w�$�5��0�[a[��w�G��:펽S� ��=$Q�
�۠Ȍ7¢��B]�Cr%;���W��`@�=��V������-k�x�D�����p�A�3���s;�����3��t�y����}/�8Q�t3�T�8�2�vM�&�%y!fj3K{��q] �p��?���"��!nRh+|��+�����ާ��������R(4���k���x��95˜&�7�/�F~_�Q������5Jє.[{��;X��2�8\j��_/ZX��!�b��������q�z��Ixi$(�wQZ#&ԠB{�RY>�\C�'��B|�b��șy�t��1�#���uP��q�럝�=�ZY�@�9�VtT�0P����b%�H��)��bn�#�SL���>Y�3���(C��r���:[s��J�x���[���)�I���	�@N�+��O�yx���w`d�2��YK.5+[*�Lw-�Q9ah`��.P;�M����k��d0�͈�?�&��9�θ��s{��W5��.Ul�ۚ����y_�HƇc�R����w�{gV�L��շa͇�����ve�#����yH������8pB�z��6�a�;�����T���Z��:�����������H��g+�F:��*5���~���7�Ad`~^�'�*�ty�N�+h� Ɂ,
7nO!/y7j?�.؉�^���������̜G7�b{��Ԩ�[��/����I��tYA��r�Q9Y�]w;��Ӓ|��e�e��}�KK�K��o���G��i�?��0��Y�p��]�¡"~���Q"�eQ~�ro����y�D��l��ȳ@8D���`�2Ít��SWhu�A��`�]"�wK�'R(�\��c"�)��0���O+O&��s�I2JibS3v���a)yx>B&�
��(`�iN��V���jQ֕})��C��V��O qCV��Nc���H�jF��=�c�>�놨�Z��Z(�{ڒ/,�}j����ޠ�'`��ƕz�g�C�+�����L�d`�%'Xg��p�+S+}���)�2��4�s�]ZR��A@����h�7{���b�6$2W�^�ݺ�ƯU'pt�8La# ��2�-�n��ҶI@�U|	�r�/�(gM�l�,!7 ��JdtZ�w&�VyZ�bꊔ���p�t@����tS{��W�s��0��*���A�Sa���H�yaJ� ��5rqP�H�
�:S��'�]��b]D�,��}�]��nk�^!�Ծ�:"����2�	��X�Y\B�s�C���O��"��v��U@��~��䏄7Z�8^� ��!�n�)���z������h}�zJ����u�(E�{�l��b�vW��;����Ox.��Fս/'ض|A��f	1$~���s�ӡ��(���k���_
Lq՝��ۅ��84���> �&O�ؗ�GUJIw�*��J��Z����<�Q�%e]�sJW�MR912��C���KD�م�Br�d?��]���k���R	]@�dot�I��/}��!�����آ	�܅�Sǹ��u ɄV �5�Ր�_�	@[�	wK�Q*�Tڊ�BO���8�s5J
*��vp�{Y�
}Q�0��ѹ��J�O=�+߳O�EEϑ��as~�pB�#H�ŧ@ ����k�Eb�G�- 9G����0T�o>y�o��	�_�߳s;�d�8e�Ci�㈓��'S�u��(SY�#��,��Av#<�`�e���]0.��ȸ&��"��[!�xh�G?×���0��^����h��4/��q���E��9��"В_c����4� ��oE�qR�-�/E�$LdxJ�7�v#��쨣�}Q�\�������vT��Ͼ2�6�"���Җ�QȄ�h�.{�Q�˚�d]_���~h��@.D��\��¦Jj���䘭࿱{d�}�� ����C%J#��$��������΂���=�B�S;�ʸXQY�S�X��ɳ�9��'d�e��";��
�4�,�:��Н{��l��Fѡ ��:��v&Y*���y7CLoJ����o�����?�"e"_�Fj��t�*�X��g���i�O]�������P��^�zW�)�R`x��� �����J,�`������n��'x�Y�I�IM���c�^G������=Hϧ U��n���Jk!�ݰ�#)�28/N�(��G$��Z�w�S����H�'a9���рC9�J�ľ���ِZ{'����/r��uk���\�೽�gin�^��Bu���-v�<�6�0pG���ƬX���j����H�y�H<�Z�byC���?H��A��������r���D�����@�ő����ׅ�=Y�cyE[�_�t2����C�Ms����z�zj��������Q_x��U�m��sP��:;^�A�
6.�3e�[��'J_q �0��&��#�!�%]SzJ�㼡��3zC=�U=��3G@F2N&
pX�|k��FYnq�~Lu��<�M��k^��\�Ak1ܟ���ֽ�0���Y��ut@�qd��g�i��1[�^��@0����%�vE��:XCØ�N���J�al/>vۼ�H����K�����k�I��~DҢ0�����k�����w:&���5�Q�=@8����6Z�'�aZ�R�^�W �ˇH��	��ɚ���f�v�#�54A3�^&���[��@��+���ܭ��܅�D+�ȧLF0�9C�Z�>>죋��u�ro�o�U���@pT�ޙ�=)�F��M<kc���Æ�7ʛByq���	� A���_�`{�D"��SS5m]���}u nCWO���o}2( ;��&e�n�vD�:!|=�E�O��M@0@�χ���z��<���-� ����-"�A-���'�?@Y@�ɂ�}�F��"��^�6c,��]r^��������C�2�ŋ�2�_[i8�ۂ݊�:���ߦ�M���m9�3�E�n���{,%3��p��^IP�T�j���-��E.HbtP�+9C ��������5U6��h���.��0����RB�Y�kf=����:>�u:s"+�ֱ�Fn��mT�����4�r�h#�E{C��;�8�ˋ\��Īq��%c��2%�VLrIJ�3P�$Y} �(����Cl���5�G�����l��܁��{�vD5}��s��+�|c��Y�*Ʋ�]-��"��ڻ�U�Z��{@<+E)��ꓫ��0�/pm7n��\��g�������ꙩ�܎��L4�I�BB�h��@o��"kx�@��\SB�����=�$ܯ}z`�h�!g�״����>f$���0M吥���y��Ͽw�7\Sz �$SY�҅�ʑF�K#��C��}����
�u���o-v��ݷÎ�{�͡BLHPdc�6d��Dx��/q`���9rj0uI�ax�$�7"".�kd��.��!�8��/�'���l��b�J%��� �b�n�r���P����L�[`��,��iA4Rȅdr��F��MP�~8G���ƎԙZ1V�����eE�OF��Km�%�	��+�Og�v�k�����G&����G�zӉ��C��Ӡ�D�s��hOT�8c�Ůng������ٕu50�00���xh��Q8�+���X����b�ɳ^U`%�j9��:ZZ`xRܰ역2� 'ú5*��b_svԀ��d����V�� �66���(CA�;YƱ@�I���X��Hn"�n� �G�Ly�j��� ޕ'rV�^���j�����<�(O�M.�fy�h�O����?��74�~�V��ិ\�%�%��˻��f7��e��ګ>\l��0��%~�_͏�~��;��5R�Fֆ���,���;��
cW|;�(����cU���`�(>�*y2i:0]P�9��NPtT�'^ ��J� Ap��q6���D��XkB4f�P�Z�M��&K
7>�ȵ��_� 2�uCM�՟n�� ٥�0�OL^:����8��H���>�;��]��ډ������r(䁛fM[�~W=`�YU�	j�9j��ߥ�W�/L�u��PcN.��,�Ib3�KL)�2�@bOL�?�$����	_6�քهz,9'�?Z��U�ɹ��$1��:��J�V8���t�U���\�^�0������B��lJ^�ܟ% 1]��ͫ4qP�-Q#�P�o%�2)�ռ�I�ǔ�&�/�;ac=aZ�����3 j�}�_zHl�4,���GW���8��i�hqH� ����㜑%� tV!��N��̷��w_jEd�C�����S������/KV�`S�˵>r &�=yF
=����v��+S䕭&���ɯ�z>v.Щ�𠃩)�����G� ��^!5�3�m�:�٫2�}�DUf���P1�鸚�K'.PHfѸL�=/�t���R��x;���j�µ]S8n[��̡���A&Y����l������#������[8�[��} �(l#��w��j=2��Ԟv�۬���3��QX��]*��2Ȱ������������@~r�p���1=0��I�V����2fSQ���?x��X�G�R4������w���dLT���$EȬ!���.Sޑ�)d���tEM+��#������9�r��iÔ&Y������&ъ�4�>����7M����F@jzǏ��+���Z�E�=0�϶�3x��.];*�����J����1�x��b�PA��������Yn�e��4i�:p����obQw�C^��ʹ_�Z�$��t39���
<E''����h����D���w���<�U�"���'�I��5���	@6�,�e����>vQ��9&�����Mb��O��<��3�B�ﺙ� OӅ�I���q0%���n{8��O�s�t��gH�䡞\Z�!sƶ&`eЯ�?���F<���e.X�:O�@+������vi��IT��W��5�����LْA���ò�6g,�V廩�����S9�Gf7�[����҂�\�*�$9��j�#����(��z!C��5�{Gdݴ�m_3A�$[�fu�]����'���t����ވ���a��f%>H�/��)I�]H�:�=3��у����Ì��v�!��FY{#��ü�E��-pP���ݪ�}CQ�7�����{N�*2�,5]���������2,�%��p ����K��遛�ޗϝ��]C��i�$(�c`��ߒC�웷)c$�$�e�G�6V!v���0�|�|�C��K��6���#�/����� ����y-&� �5���` $T�~�t?��n��#c�����L8�3\�-"I0(��m�VK�9�w	�c������`�4�W���E�/�'>���s�9l�����V�1���bRxJ�+͝p��
6�.)�[�N�k"��F�ΈIO���}:�Gj[��3��T�s;x���%.�R���>�_@���
`�F:9y/B�&R�;O�2Ҧ.�����W9�S�
�_]9�Dޏ5��������:=X�2a��m���K��
El�ʽ8篮Bu�KI�y�=��P?����`�Mc��l�d�W�ϑͼ��H�Jo�7��`��d�n��������hxRT��'�.�$`����L&��[-��/Wz����^}BJh�����st�i���|���T,��yf;SѼ�d���y
�3�6$͉�s��`�`KLV7����IP��D��b������
:c��}���$�;��LI�r@����'��*;~�v�������!	�o������"h]<���;y���m�搘0Օ�2�@׺���w�_}��}|�h�.;���>�q��2" ���=V~���,6�ēF3+=��V��a��0�&���b;�g�M��֭>��ٱH�88mq/�G1���`��~���%,�?��k4ƨdM`;}��'���ۡm�L.�	�i+`tO8Jv���ls� \�]N�`W�R�T�\�0*XL� i�D�_N��/F#�y�uP� �2���*0�:��Y���;��8X��)��d�G���)vPNyVWECN|t�$�d621v��E�XnQ���ݻ��z��J��6�(@@������g3�Cj���Cg8��W�Ҷb ��� �����f�5�9/�G���#S��p&������ZRvj�{��T1�_c��������
����)��x�����&�3z ݍ�x
��N#��V�Qh�u��� �B�D��~&H�Ϙ|3e����hHd>؅튍���mrf�k���}�{S�*z[]fGR%��y�5e#t��C\�HWI���E�W��x�"
�@)�7�5=�.A�#�Q_����!�AZ��'B}������I}��XxB�\U�z�hŚ���k��I�@�T��W����)�LoU�hy�9����F�|��=��|s�줽Q��)q��n�5�gB��.�)����~��T��K�`�f�⚔�w�g>r�a���K�_!�w�2)+IiΨ��9Z��VN���N�F�&�+��|��'�װ�M1Ն�ۓtJ&����G���n���C���	�]ٛ�-�`���|D1��v�:h�#�ӛM�A+Շo���̓��ߍv��.�Q��~FA����
y��YV'���փ���>�7�:@F1�b`��)P��:��ի�ބ"��4�뿝����Zg�&���y�P��t7�i��`@6���кB�����#A��ּ�S3p���[�bY���3���HIb�q?!�LC�w*�o�0�T�d�3˶��IX�"��N�לX���K�˺��A���4�F��8> �Z�A��B�p7rٚ�1/�����L14�Ff�h���^���M].V���r)��0�)�Ћ{������:���@��`s���P}�<V(*CȾ���`~P����0)�-�\�Bc`LxN��;���A���u�(\š���-����!=G�*��Ǘ�����®��Jr�OqV�[�J�V�"�.�]LA�J𜑜l���7�y\�t&˄���Dd�v��p���&K����L!��u����V
n҅��1���aTM2�V�X�n���A#��pa#�'l3��Rf"�1�9L��8	R����21�%���⠟`&�FX��)E6�yT�*K:U���1������;]� �n�v�v�a��5�^�~���j�̏G�5@�/W�����tFM�B�!5�6ҫXC�fA���V;�Qq4d��O�pQ!����W?zȭ���|)±*�Ov��8rq����։ג޾��#`Ey|*�8R�إ�f~2�l�(�?W�A В
]tM�M�M�ҁ�)G4P��w�AeϏ:�pp!�|Q��>8O����ρ9L�q{֣ד�����˂��iS���� *�=Ef r��~�a��ᓪ����n<�2�%e��-MY�5�Ƣ	
���j_�����ꪬЉ{$�3��5pa絨����)�7\�*�	����:���-߸���(-EJt%S�/�4H[*�'��`~���1]����+��OX�̥���V��#�d�4�d���f3saZ�3�a���V1K%�} Qg�g�I0I��_�!`KP�,�}n��i"�93�w�x9ºA���	Bj���,�������c'��NZ�u!�e��ľeo����#x8�hR.zˎ�Taɀf����&:���"6å*���������C�VIs��N�Y��'R�/"�ZM�Ͽɚ9s��Fݻ4�Q��Ȼ�S%�F"O��a�4���(<�����"E}m���o���&e��T5��ͅ�2�zm�G����l�L���K= �-=l��%[Vw��H6Zv��B�Jԭ���}װp��Q��
S�ZV��8m�H��z*���J~�"JP����)Qt[�d|��03��V'@�l3�~VB����Hm3���6���(�*CF�ˣsOL7��R �z.�v�'�<����Ԝ�_����_��v#�̇f��U�xE$)H]%�ɴ��`��"�v0aeٶ�?��Q=y��2��ҹb�(�t�:/���`��V&�/U����f�li@��O��%�Tr���ɫ +r�bP�/,��T��Z��y���O�2S�dc�eK`Z[T���17$�b��ݴ5��N��oMWG���.��==s�)"��0��U%`��O�.�@�9�]K�^D!!���b7�o/�%a^��5�����`*��}����4�8�r�[K���:����)	�=:�~Y���O,:���_�3ODl�'��Q>w����C[�Ot�yÁ�,���{�ǖ���?̬V5�yդ�.}Z��&����W��I���7�D���}��_�a��[I�j �t�*�8ě���3r!��H��ω@�i��_ ��<a�2y8ҡ?s���x�-���?3��[^9<�T3Yz���*����3�T^I}c�ۜ�!�3�Ԍk?,±;g��D��م�&ww���b���)��s��E0�桼�~��2oC7
�c0k�!� ��P��ڪϹ�	������{��r�f�H�&�s�L ��<v����R��75��es�H�H@6�?�x�"J�*D�)r��|��p�Y2����"!�+�)�-��^��"	T'Nc���.!��+|a?��lJF��&ڍ����s�ٷ�{���>^��W2JoQ	&�N_ne���"؍�y�T�G�͵��^��s*ۿ82�P���>��ej=N!ўp뛡����_�P[�D�]H��W����t�4�s+(�P��}/�v"�:�)j%�������^���/�]e����p�q�Bb|�O��3�
��<o~��\̆���TT��mi�,�k���N[�>f}�$��O���G��kƑ�?5?>���S����}N5��XݜRӈ"<� v�B�i�&�s��\��\��SqRg������J�i6�7�,�v��:W��$X���<��s>�M��Q��x�|�2�+;�>�Z���kj�n\�]�9�lcw%{�5�x<j�'�n�{!��z�Ś��� ޔ���Ȫ�z����~�Unw�pU���J{� ��������d���*8<�P��M�]������Kѻ4q�
r"���w,�+�-�E�Ʊ� J�Q�̐�f7N�hE�{s�ܮ��T�N��|��GH�[��J׉\�b����Ngo<4�+V���E%Z�R�E�&����؂���(4��:�F/��'�X���v�H36��`k!cx�n޻��A��:�"�T5�n�mMkϴ�Q���ѻ�l�2����dnc��0�1�)���?�?�K��ڳ.�嚡t��Z�|5�]I�w�D퀃���3�+�~܀&�{F{9�6Ź@iدt$'Ao&��kR��*'���W��dx�yNQ�-�uU�*����-�An@3���!�8;�8�����t�z�K=�ҤW��Tھ�=b<�_�ebS���؟·Z�B��r=��2�vW\�e1��i;x�:Xd��C#*�7�c�8��掎�%+��MmIb��R��ۀ܋"MK�`�M�����Xz,�s�R�aK�l�	�P��i�1MGVR&�A���E)N�����y�L���O���~t�F KOEat�QS�д��Q�帙d@
��Q#d���ӆ	[��XlÉ�A(~�a�zvM�u��a&�!D��v�87}�41L@��]J�4(:w��H�����	�> �U��\� ��x}iM?0�MV�OCM͓�/:L?�;�x�����VS�B��7\�-��f�EP���u��O~��׸E�������dL�²֬��'�fq�W�>I�a�D��qe�n���ђ��%�dM��؞��_<���#���s��h(�YL����O��3c; @Ys}Q�xj�PH�&��M�J�x���Ҥ��嗗[W��@xTw�a���>(�e.`eRm��zݘ
	+�q�l�7/����ذ��6#�/�e�'_W����3x�/�y�9�W�}�n���?\vO7�z�&�IT�=V�m�x{پ���I�u�R�����%�}У�r��>����������ː�����^�T��o�ъg��}����Ȉ�'n϶/�����?B����*����2}�l��e���=&�owv���'Hn�$L��;N�]PP��"��.jfĘ>��͌�,�[d��$
5s��g�gi�X�Z�(5�°4Mt�0}�[U5�lk�8 ]��AI��n��sD$M2��*5u*[�΅�It�R�re�Ta�TJ�����;����+��|�1D��-�JCF��I�l_]�V���cqea}C (΁�]���w�/M�-IO4���,>٦S���m������ ��_D��hˮ����h��zJ2�yp�ܨ�p$6C�=��Ab�#!yD�OҺ���;8�T<�[�7��m�-0}#�+�n�G�De�`xq���+����
�ne-qЂ�ͺ>���+"_��CRN��1��A8�fӊf`pc�<�`�x9[�̤E���m�!�r�����i���FD �ͻ��[��$�@�.UK�N1FsA��|�����{]���[��U�6,�D4���n/Z		�u���	DN�/�_4�TW�:Z��g^�֭���梙g���+ÖB/<e�o�7,��M��l�PY�Lԙ�g�;ѡ��P����{|3���:)Z��MMQ����g��z�O�ը1U��_KP�M5�cj__H5,?�=�F����^ՇM��z���!��><P���Pa:���PK��w�ڴCg�2kL�q�`�OV[�;���+[-.���Jp���2j6��k�s��Ce�pu	TqLHM��c3�3'��q��K�_�xFgs�� 6�A�:�HqOJ�� !�&�{�객r_��/�}�:i�vW���YS��m`C`_�w,DCǡ"�Ѕ�	
 ��[w&�����J0�\Fb[��H�]��J�\����Zw�,N�J ��;̎�Q(8dqC��C�,�Ԛo�=�"Nۡ��ɺ�O���܃F��Ɨ��O2|�	ʵ���kj`� :fO2d�'�6��JTQ�M���L�ş����36s3��
�BS�X�Ǩ��Ӷp{u��D$g��vj�~��;o��A�Z�0���:�a�&ý]��狞>�+MxJ^�,��Ek��@��>/v�*�a�����/��`|u0E�#���9*�V0��]����}.�zq�iK�N���UvGR�G��ä'��+7��Ľ3��+:���?�A'��F��U߉=�ɺ���z�u����&ቱ̂.N�u���A�)W�uV\3t̮5��Y6��{�k6j����<rja �#oW܄��v�1SSq�Q�4���W����P��D���?Hͫo�Ʃ�˙idW��- Lh��ӎ�*1��%��Ʈ�謵N�l����a">Jv��șֺ��Ih��a�#�2%/�4��O�.�@k��4s���#�ډDWp�-S�>hd�(�Q����Ɇ+}<�_.�uj�R�Y���t�?/nI;^ �#l�4eI*�[�B�<�t�¢<fͺ���D�� z�OZa�]�ۢu�I�؏u�����X r�����=�����ےf1��G��I�l�qb��������Ԃa^�(K�I�Z��_(zӸS��rFe�����Qdo�5]QRT��i>���6����n� mr�������c�4���E=9J��c�#5&)�b��	�X�H_�ć��Z��#��º���g�9^�Y����R�t� �Gڱ&�� lz����ʡ��M*��� b����l�O=�Ҭ_���N���c�TC) U��e�ou|�VV�L��@a�0��0V8}U���ۛpA��Υ桕B����9M�"�W�O8��fM'��H���X��U$rw�{}iWQ����|��ûD��Ʊ@.�Cѝ,��X���8�+�O`�u�	߆�.'�y�����n��zj[K�?�'b�����wξv/��ر�V�C&1��W1�����ڰ�\�p��s������{:G��s�Z�i��=���";�6�'9jGw)=��X$�!u+A􍮃�U+O�
"�m?j�񇍟�F�`�gȳ�a~EM��"(wu�Q�ر3_���x��Di��,T�R�X�Xc�!�V	�B��<ܴ6���ʊ�r��[i�{2�����'a����h7b�h%R������!1[��,���BA����a-�Ȳ"aVN��&c������r�^D7;y�_���,���܇������t����<���,�.���nI飄�l�_�K��R���f��Q���ׅ�,� �K�a4yF�'�V[�]S���Q����lv���G-�\�މ�����
�$O�5�E�+���Aޖ�ɳ���[F�6e�j����K�_V��Đ�;�1'rQ����ZnL���Dj�j��X;�����5�AL�?[������gb^�4��&.W ��>�[8沠�+۩�k���@���M�����A�M�Q{-u�C#}ƪKL���䵫�=�]�������Z��Y{_Q[G�y���0���^���������Q=Ϥ)����Z-r  �0��<��5
_��#����a4���m��%��i�@�M��1x�_W���ķ��0�H�k�$�W�P��X��6�s��dΘ Ƭ�ܾ�Bq�%��D����(ፘ~�����6FY������!Y?��R�X�Kc]Y���WA-��k�ia��`��cǥ$MEP�gFŘ���0�AX>�"}�H; ���X�.k3���B�2��x�yR���0Q�+��\��+s�Z^��I.���0� 0�6�f�ɐȜ�f�IGd&
q�&}�ad	^��=��52>aAɭs�8P��_�iN,���U��x�����tw�u���]���n���k�Z�
O�EBTF��踔��h�Behp�������"6��r�؎||��mN� S�X�JۂQ�|��N=�5��W�󗆁 �d;�8���l,m��+XBUᨏA�ڤ�Ŋ��x�i���r�!0��3	(4�`_��qhY\-�}����pi��C� �:�I�r?B�mjir��c�f�g"A�h�CTn0��P���?cr��ġ�"Z��AM��*߾���=���2�=������=zV_�p#<���nv��� i��L�a����E��n��B�&[{M�.4����gW���F��r�[�a�	�ҹ '�h���̒+a��$�h�SG�M�s�)����,RW��[���#�Ty^*�	��BB�U]q��J`Nl�91E�q��t)����>���pa�<����xY^h?0��9?�Q{�<���`���V5N�F���	V//O::}Zş"c�0�Ԭ��$��0�)-�	V�pE�H�E����-?���=�%7"�[�?NE�C�H�bY�?� O���:����۽�i ��<A��(�T��)X�ůy�d���g {z�Sm xs�!%=���v ߡ5���:`�����p?$���7�ɹ0�O��d��f�c�D�^���^:�6ܝ�͔���6ro�_����7�������ܹѹ��E�n�W�ƽ�\�\���O52�C=�a~���>�fp(����=�P��(�F޿���&��(��������2�uYdT�N�b��Y�7�����z�h`�)T�,v�fn6�RG�1Qc��_���@ٝ5l~Ky��P�����1w~�H�p��C#,>�p�9s�7n���]]i-z�;�z�z��Όc�X^�����>��L�q�϶#I��8�D/W(0m�l�l��J70��|�L�wR܆�9�����]�ϲ���S�e��X��q�N؈����A|I}!�>�$h���| ��3���>'X�̎�d�k�Ձe�B.��.z��-��W�D6wE$c����de-F��j��t5>�|�C���8����.ըej�����g_k;��ì�O�85T��L"\p�+
A]%@�B�vJ&�|N�^+|�w����)5x�;����,�_|�Uq��X,�]-Qh����	1�0����-B��vp	�Y#D��������m�yTubs�*�א��=$��bD����_��=V�{q4uC�$�N��|u��<�7���9}����R���H�Z�b��|�s�A9�?�֊���+�~p�M?�Y��=c�E�W��,�]�������{��*Y;!Y��	<�>a�q�+�׶���u�I��LM|1"@��A�w�	�:�p*%RtH�T-#�'�~�.�П	G�ܱ�rW	���3��h����
J-}�]b�I�1s�UG�&�=�\DC%�¨��0��>Xj���ڧoU�H��{��Bgjl���N��!ֶ��b���e�U!��`N3�r�ū!��,���C�f&t]��NV_���#~�^8a����J�7�.Hh����R���wT��e��*L�=���O�M]r��/�Ad48{m���u����Ma�wV�M���I��d���>�
�[պ?�J��{�]Dn��/����_�]����g'3�����xdHM�FU�����iz�/��N ��%���oS&3�%�!z4�(��e��?>gZ������Qy��xcD�c*n��� m�������h�u��]����-�n��`�]j0O�?r`���,���g�0�Ź���ӡ���XXZ�F/�@�N<;�����a+��y��R�<<r!R�4���P�D�K����4�:�U�Bl�a��`8B��@7ŕL#��6��W���aGA��M� ����=M>L��m��Tx!�z�2�����X	��H��{����	�PQ8��φ4M���&��O�n���ջ0r���rJ9�����O+����KbQ��rT�x`
�β�墻���)i�#_he�<�̍��C�Vwx�Bpn۔��	�	��qldU��%,�o����)��ƃ ��>7O�ɳE^˅�������:�t���,s�����ۊ{�!ؕ�3S{r�J��߸�3�$
΀�%��%���T��	CT��޶���D=������0�P�3=3��8z�N�ȰIgO8 �������$���0��#Jk�x�x�K]��j�F�wRs������DO}��J����?wC��,EEo��Z�#������<�;~��tv�I���G�\1�^{��z�ƴ+a�����eU՛��)2�	��FU����G+WV��ز	{]�#�0�pvk�v��g�oqX����J�mT�n��tX%+�O�KU� ��u$�@.,v;�<n����@Յ�&h�,}��6 �J���WA���!.����6� j�����a������}�B�U�1VGU�t��|�Qe471�jnB��9��
kJ#�븄ڇ�aS�k��.|�"�>.���Gy�r�
�L4�TQ���J���oc]�"5Z{��O���Ja�Fw5h�,wS8ǹ�!���uB�[���\�1��X�gQ�~d v��� 2��*�b@��Hb�1cOG���;ㄎR1�l����[Ƕ�K}� ��@�
���ٹJ!��؎Hj�DϜ����\S���C8�S������[�bLtݟX[	�7.g��K�,�������\c�<(ѵ3�R2������_�v ����jwa��_����>��X"_�����2�T��C���߹��}��M��&6o��քɶA~K4��W�l�SN��M �"��C0+�q�A��^�O���L���o�5-�A����C2)�y}_��cg�]��V��G%�@Ԩ2�sEb]Y����QJ���~2�k��N.���r]��ye]�"�;I��C:�;��{��L���hh�)ۅ���W�4�����%M�8m�p
N"�f�Ԡ	tΤ�ή���[^o��p�uH0z(�+T�m�f�b���p��lc�,j�AH��A:��[���t���ṛ��`V�����̖��G�Z�:W8N�:[yk��a^�������E���S��a�@��:�Tg�k6A�DG˭�܋'!�G!�}��b��i�o#*{�*�ߓ�8�&���Vg�SZ-���52��o��cV�`^q�����j��$��f���h$]5��*	^{����6Q�q C�a�<N]����ei��^1���I�~uU{�^����44��*�d�#@B��./}�L�i�qU��$���b��jĀ�ғξ3d�vk�5	B���Ac%����zm����� ;g�񿶳Q|:����	u$-ԞsO���E���S#�(�������`���	i�J��Ķ����Jϑ����c1���z��Ym���;g�_D,�	�����e4��1�z�!Zf̛
@fʗ���gکPx`1�ڨٮ���_#쀣��>l�]�!�#�U
lZ�k��~F��گ-M��5�h��w�3|����D��M��-��Tg��h��Ŀ���{����Z����HA�.��hc���ߤf��X�0��(0�ϟj�ڱ?VME~�iCY�4�P,T�rl��{�ن�<*i ץ7����'���Q�Hf�]$o4P�@�WV4�+�'�������ٽ�!�@�GW�k���k��NI8%�(*)yo��s�����.�\�̄xn�%�RYVm���:���Ͷь����6��pwi��Y��O�b�`+�j���W ������dco�=*V��:���N��+M����w���]@�웝D'}��Q[�[;����Ғ�7�n'P�b}Pi��D�z��t��epO�B߇�\�?[�o��/�b��/dz�t�T)+�R�A�h?7�xo;S�n[�W��=6�X��:f^Z�͌Q�}Y!B���Vʎ��O���р2�x	�Aʟ��T�{��(�W��k�)ދfվ�r�N�W�R�����-�o�����=�
K�:�	��@��y��3ɚ��<H�n\nQ�~X�Ԯ4�-$�����%������/���$�3ER����ZGF��xg[��c��mKKO�З��*�P�'�Q4�1�����N�zGZ��Ԛ<y���H�|�I�K�i����u��P#���rB�!�|��d�R�"R��&�9y~Ɓ�Ovp*��3�?��(�A���ZQ���0fM�z!���� ��G��j��3QZ54+�a����,�Q��;kұ�5���-���+��
g?Y�W@(	^L1�Th�����{��}��;X�b�D��e}��O�k_D�St{g�y���U�n�[��ZN�ź^�7�:�۝���Tr  ��w=9�q+��Ր�i�Q�mD��K��h��1�Gt��_����D;��6��C��s}�٘L��j'9yO;A�8��W��f���|!S`������;������b������cl7a��`��(���T2O� 0n�5$�O�����$ؖ��=0�F�$�;L�4�XS��>��%���0j@�g�q�k��B;~Z���^�\�?j+�]c`uI]���&z-%�S �Q��SE���3�͙�|g�JHV��v�AJ*12�'���^�@V/�����`Xr�f�߻F;�N��L辐�����+�\��YsAD�i �5����$˹������QUX���k��jf1�&��q�_����U�.�	��W�k���O�h�ʘ/|R��ɡ�Nl��{�9�VE��$�~��Z9��]��U2�f��~D։���Z?��O��^Vn���� eܑǥ�7�OO2�m�#��btu&�'[Zߊ*2b@P����9 �<k�-=�A}�MC%>��|ht�<P�&2�� 6� WB����.��RS����k��X��v�?9���Ez=B�� �HGɉ@R
�g=)�o�h�8�L��%��N�C˨��x)[׏B����� ��,���C�#
�J땬wD�K'�O��V���|����4��S�|3����Q�?�*�[�&���a��&�Ŧ���#���]?0�H3��D���o�$`o��C�3J�kh��+��&�e&ך�΢W�Ji��sޫX[�J�����B* '�#���i/{�gK[��]I�&	����a�R^W)�;h{�`�v�W���K>P"�������+�T���l���,?#k�!�yL)b`����	X���m�3���Gp�')?�u� XtSi ��˃Z� }����("-��Ky�'��ʲ�N�wDL ږCw��b��Q0P\-�{��W��6�tW*k��E�	R�Ud��M+{�Zd��X� �B�nH6���G7n�]�G���}N��$�T�)��}��=q�)5���FbP%���,����_�=I�ӎd{�H0<f[R�'=�\����Xڂ�XCђ:��^M=`��)u��I���G�"�,A,VCο������6�@�rx�Z�x��V �S��wM+��ő�.\���h�%0dF�\�tP���bX��PͶ��2D�-˘��{W��8�<Ʃ��ʦY@~���Z��=��૝�o6��DLa��G��4��Ҫu��0tR���MTq�\MlWU�!�+H��O��UP��qz���	���l�ʣ%��)s�;��z����F$aZm�rE{w���'rT(����!78P"L�o[��y�y�m�T�,�����ײ 3?)�su���W����k�$v�
J��`�C����a��:�{�q�7c�	�g����@&+�Z�7py�:H�"8l��������u#����?� )m%!^��fs�I����R�R"�Ա־о8L�=������!
���F�'�N}�@�E�;���ߓ���2���l��<�G�qz�G�C�i9n�D!*#�0��7��z]BQ�s����ޏ�$�
�o����M���%�w�t��HXoL��?r�t?O>A>y�]����'��G����	���kr�`��P)"8Π^Ÿ�1�&�`��]USl�����
!.�����-���a����B�q:�GS=�=v�3>���l!�A�����!����j"#i�n��pQ�B���!d*��I��M�6	�^	!�q<c0�x���m	���(����_���W�p$�@�����@�G�(r��k}��W�°�@�J�f	��zT�R�~2#r"�k
��
�k.������W�a^
}���i�.;��,�ʧ~塅��v�U;t�"��A/.�E�Ƌ��p?���t�
�.������w�ʃ�A�$AE�H.�I��c��G�j�����ɞ����d�as�����!��Љ�?��"���oq���c�ِ��yz]2e��{�<�>K�]Y���"�-RP�`�Y~���}��n�N{7,ۃ�,�{3p���1M0.��	��u�+!$54��7gH�Q�� ����K�~����!>{L�� - jK�xLx�$�d5i��O�G�=>����W\�����^$W��oG�����[�����N�D�(����������곥�����:O;��`���=1((F����{�v����̪3� "Q���@��s�_��!��Q�y%Ρ'���9��ܩ��xJ'P��?�R�Hn�ݘ:WK?������w��(+���S�i!Ѭ*��u��(@y�j�����FY�ja�n5]�G);�G����� ���Mtr��@4�Pu�K� ב6{�:+돲�s��4C��������w�I�Bž�C��3'�8���B��3N9-�5��<,����Z��������@ēp9G����[�F!l�M\��ʴ�vUe2#�Vۥ���W@d|*��x�l%�;P�t���㫛���Q����Kڅ���́��G�.�\1W��i�N-,N���Fo�o��(����7'ٷ*�NY�UR���ɧ]9���Q̋Q����(��`@�n�'�y|���mC������'�v�:<�I�|�s�UWh��g��_�æȋ��ݫK����