// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
rAA/bfs9xk9Wmk9+gg0v8Z9QND88SZeh1Ew+gu7HTBNkwENuW2dW7LXrKvlFYb8S
JJt8Ad037fMAj2S9j+1vEV3+Gh3H1cs5RzXLCObo838xLMrXDUK/h0y9WfcBgUeF
vgveu0SbKrln9iuYGbqZUToYwvOSL+76L/1LUiRgVQg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 25888 )
`pragma protect data_block
PpcJo3r4p8e0wJAzFAz8QcDSjaLBKNeQRs7bDpOqSLC/unEngcNr/RvRVVAg1JtP
sZQivkp71JNrIvbs1yFX00iXkMKsyE8HRe195Q04aXON2J6LAodB+zxPiFoLIGkN
+Hznfy7lXNUdW/kibPtT2YI+r1sJMZuSEFer38VMwFBFHjTrk+oUQg4ebYUYOJIU
WOe3+5J+cf0ERYnPgYBuOrCYwnDimnC+/mWCBYpQLIDIfdJMhbHHVJaCH2iSPNd2
+b8Eiggi5brMicxpubxlI4K6TMmY9LGkWd3K9E27QT6NnBA8Zq39at8RmU5RDKAz
BdRBq69VKPdUg8nW8jlwb0yonoDpilVVfkuft8YalImm4gsnqRdSWsmPLH2Ewmeb
r4WYkcI9Sx6izs+BMnuEHv0Wr19AVYZ0l4kA4CZxKLcsSr30Fcj/h3pOIrhYZn6F
k6pWKKeJJvalMqNlWPWRqrR9w0CIWpw5HKIQgbbxbyRyHJ73P71eb6t0lFCjOa7F
NmOf+XKn6AMSrV8bzt+C4/DtA+TWYUyvvL2zBmdEIimbbtJE09GA29fvLdlD+IpX
01EtcWBJ7ZhhhNJk7Cuq56ZOORpnFrTw2MnkRrjgEHNTmrfocgXGNk/VEO+UZ2CH
hsYVf+Bu+5nsroJCNJsMSxt9VIwgyX+y/7ncQYGUFb7ifks3R/rOj6O4Lky5fv+v
kfzYD/r1pSRKnZFz/aA0+Bp8D6H2g76HDn5pC0n8ORMTmGosrKcQn6UMlEYn/HOE
TM5Yp3mW9mB9KROqEIojskur8Whp66/cMtdc/i5HZau5p3J1Own+6IEKFWeYeQk2
lVzqBvtUywepm9otBW5rc1vd1wgczm08U21hyKkODYWhkqHxFN4dxQzk6fOl4Brq
wUAxckoENar6P2LeAmw4WUWxdd3gwtA4OnfV/SbrbhE36Zz2TtH4mTpO+38I81oh
4Lo8BKQNVTJbGFo9uuDPDzuRwtOYtUS2ukjPhaTezowRUQCtXctHAYI/lVdfXkCE
RUCHJbCCz59HhhR/RYAI7+VgIkd/xfDcWB6nY6k2H+WuI0a9wYqolUASq6JRLJoO
rV+GG3xD1tsWV2cZqGldSEikyO1Ao6LRkdYWdDcgmtRO7e55T6O6KuXJkdGV/sNH
1ncMI3sjYVN3XD+01n3sLZzhIdCbmEqP7VcQHDm6XbVR/S6S4hc/ifAhRu7dTkow
/SIQiWsz4adnXQmMvwRaOGFGytQ6yjoATrLEYlZp6Zouubo0K3KA3LMzHOiwaTPl
56RKzCfRLV5FcHGGYwXuRWNoQGf3TkdcQ1FPz8PP7TD+7RYD5on6rInHGb6Amd46
tFi70wxyE2fJKzpamwDTuOyFxkiK9WXafWknkCZob5zeN0qaN6zO8ZRrHThYBG/d
/Rk3ehXnehb+YX3P6oyRxhsFHdtEsnAZJULdggJFUsvRZ+Tkk2Ofz/e0HimmP2RU
JHNkRjxRKAWCuCgUG/OjYLDDxdjJHwfD7DlEwp68rOS7rdrjqpHOaB9RHc+W5mUe
XS2AKVrQRHV13Nefd8uQo6cuu/Kwtceutdg4gFRpbQ+94xOF6OOqumMWCjo997gl
YweOhpJiVoJ7xA2BRz1Jdar+SWWvmApi6BZnp644DbOnOOSS0/gT6wPy7pFcLHUT
fcukDDqIKY1+fCxFBM58CTgmuWU08br57PHNyhLRJy6PcHpDCO2fObSwCiDD14kW
6j+mse21Yjq1em3ro3SetvkQDng5ViY6LN/ZiLBIut9qghVHPj89Qj6Atout+bi4
aYwDWr+mtV6r4Hv9h4ksg34eAS1pG1RcCO0/DAKJCiKLWWZr7gze8I3TvDvLX6+v
8oMZYYkyHYldGtMqNV5IR/tqO3uZTyTaIYkscPKZSJu4sphgBkMrn7YhbAaqCdQ0
TnMPUqSeh3aKakAAH/PqA6z8EEBLXVVCANrlBstPRplK9pxxmTe/3xu7YEuYYXbx
2p8qNdt3fjKnDcNsuQvGBApqsTeZvzWoeEvOYXY10QFvRMW7vwj0j0rHfQGgOBO7
7WyVeEp8quTuESAOO4mARG11d4bKHfDI7eL1YP9Pi3ebuIYV7PepEuzRpOsFygiR
69NFamwtS/v58unCFC0KzUJyw8B9MaEDdw8AWBFWSkM6QNiSgxoedLECMOsa+m27
7+EVUhXeHgCcDrkQnV8TvXIGiy6WQ5ZYVI0yoK2oBJJkDKv9rNxD1ckOvSZVLtuD
7i5Y1P63PXwNCfZw6HFiJIfw7q79h0wG2sbjjYH0OngkOCEa3PoR2wMVhqLXpF56
AJ/0H94BYpAxgB5g5lVn7odZi8+/n9V57D3IcusTbNmxhOd/0eO7rh/tKUQKgGvh
MyGfcv802sJt7SbAAbZXepNcHBZbWSOnRH5wFONPi0NPsqvNotVvR3ZxdczhdYYT
4LrOcASeNnMHxGDEP1/60tkIm07bJpaX3JTXK3LilLc6CJKTD60rX2S0fhvcKwqC
OnbLUwzkPNUrofM4ilHClWsEOY2HoiJjO0kEJrwcG/AlP9Cz1lK1mRQbHZF0Y6ud
4AXohhY9sbPJ4FUG3yxO8WGhUioj3qDmb6NfRqOz0wW+8NFCDlRa78+bIyepHmeu
YmWvMEPTpoLrulEdyUmiz1aDBG1RpCB95OcfLwNVRPif5c/8om9nfAMwHmEy//Tg
bL4Dnhc7b5+NLLe3aWIbRNVnC0GZjbd78+R15+k7WOSyBrlH88Zc/uyluwivpEyj
dIORQpGwQZLJFZhsU7kMePcGcGzeZhU4gg7Iqxq2tsQzNdJ6gUBBqmQIuX3B5Bog
ivDWWcW7UGwLYpU8rRP3Xyp3uG5khlXC9ZKRgTssmoCC/xpXUCo622euUTL0udmE
0sHVT4pDI/TmQLueVyFsg3z3bNhwlosgJhMH/6df9lCgOGJfS/ycfPi/HuUph+hR
g/hm6aNvuCiJGMEEHNuwDkoPVONVu0U0fLZwbEHAeiGJGJIsCxTr1FjnbMOQOxWG
l5PtGykQXKIp92pj1pEe20rQz5vvxg/Wxh+xUojl9JcTI/6YVjn+aYDtgHm7BDjW
hVarIcJ3fKQqeAZOerhWLeVNkaJ9YBDrQjBtk+uZ0AJK5vphCUGL4SrmmsmwNUTX
FpMq++xVV0x9aPthh3TLRL5yptFY9H7e6DA0PCEQM00CMQkK+zyC4vcAab7pMpmP
pZ8ywJWktsucjb95OOozvRaBxruN6iWfDTFlBki944ErgJvhELXHI1SpoQ5yBrfU
wpxjGPQ9AaBbxVGuJbFSmDymNHmmsT2hwAneG+kEThiVQIaxjThW4t+y9mQcnJM7
/qvE30+tPuUIrdt6kfSbRXOuHxNYZAHLj9R2rGdCSVbDWvTOl1DIP1kz+HUjhkaZ
GomN9+e0jNQfqFgpGdgYy4h0yk0bPgLQvHV0a57DIK3TDIZFmC46iT5HgXYK6blC
4KSikBMUR24c1umO+AKYBaBd7vEj2SUwUiCjzt6aVP1iKCbz9aBxdViXeelrMeed
aFZybUWbGtb+mk8DgP3vD64sfcjtJitu5bydfGr2Cg2/04IaD/EZLUeeYfTITSZA
cXtbx544XUn2zsaEmm6KuRHeGUbmMYVOP6bsb8hrDcOO5edZV0fmuBoSWWuHBCsc
/ybFAbX4eJdVvs0jdyDChMpAjNnvQn2eTcjOoaRv8eoBuADiSPaf1aZA/jkBbxE7
jukSYEsByBaqwE10f763q/w2fQmuBfqQlX9sAPPKPJq1LbGmWGb+hThwrv/NCzdC
2w4N6onVsPO4mTAzuhoExM20QJsAHvLPjbqAueYpGHt5nJDzKMj++p49FJjoX5iT
DydUJIqUIfwCgyvPljsbEIU8fe13DTW8VQtPAc81LNGBS7kh6E6EHAEZ46Ks4pBM
jk6b7OTkmun4bmeosNhwvwuFbVkwiElSAujTLQnR1qEyOfkY2bdlU5KY3RWJycID
9PgQQ3zyWpKlCDiujVj6y7rJ/hTTQG0U10xYnV0pGt2h8a/HNwkh53/KhO99VaoQ
+cSqaqN0UBQsSaS/iUQg5D+rtvUipRY2Lb5QlrvJBKBNg8KdPmwGtJZPxNODc1Zr
xQDRDlHMFd+8TZccXv+Qw5RenfDIuSLCL0w+Cz6HAfYc87ETMaFQ0E6mie5zo+ek
1xL7sZPTCBFnrO8Q+bjywqV0E0AZz+HJ80hdydQnH080JXQ2zWpAfCzLVHXsPDug
OSXuVjtHQNrytHD1u5L55m3sTAdM9hwt2Im/hl51kbYhjBqB8WUJv6jcH1gNIoDJ
bGYaf/R+KrYo+SC8PFX3DN8ZC5R2snIfLCbyAHy3K5kXMk5f5YS7e/R4pFVHUvKb
ON78JbyqVuB75+BvOlwiN3aVtIJlJg7HF11CB/pkYYvLGbwMovWK5ASzXfVzIS9H
u3CQUxN1LT1BuPtnNWbmwQpNgTbJ3R+QgAnuruuI2maclOsKSReRGaCIbljsZwyN
mBtML7I+V6VJ3r0HUu8UkSh5XH52Yiw/k10hwRrY2rtVTULx1qEm37FwVU+PtP65
+myjkcL6KLUPUFdX7AQkcpEFtzrkVB6ayXmrKi9tzBGPVUjiCgKj4z1HTkM2FAXC
+oDGTBPxlDaEWkdwdpGp4SuEMk8CFiVQQwunzQI5/faqZ9NWIXjxPZcsU2+vLmq6
Z7MmaoGmU/utDP96QWzWHt8jvafjOsFs5TOZhY/95X7DKWujmhP8Kt4DTf0wYXr7
GY1plsbfIoiVTFRYwo0st5oAEouR9Eyyy9KUP0Mk9T5qXBNLdpW4bZGyTbuD09UJ
kio2OJ0/0zdmXldFUf+xYsZHe0LSk2+aDB3H3O6KSVqJF/gvl5pjLBAV0UyL1prx
7NUTRU+PUDJKXAUEFPyPs00WS7/ox4Ik3d0fErSXwspW3zeWUzzdIpFLw8eKCA5b
IpIraT3nxb74p23LQ78rj7CqjP4qGf2H0gqsjQbdBlvQwdERwyK0ArekWmhKj+jo
5u2jiWSn7KJxu4MSvx5bGCPWtV6c5mCUxsd3yadPellacFyeqUk5tltwxF0wHI+n
cGN148QfyyF20hUNrsoLjRnrKODhJfQcF9F0zpvw9BmQcTFU8hOwA2JvumNkjCOF
YrjikrmDFtueR0ULCo3aLDvUT0IZ5FTgMET3mSeHdtrvDmYR82wEbQty40yj0o14
xHH8cDc8z6Uq6NFZtAY0qKL0acbw6UrRkIv8cxy3vgMH/Mf3LBMXu6BH5+n0RbNI
9mHqC1LR7J2aVRXDVi/vU5EU6u35VODaOHm6zSTqxv/inU/Mw2qX0ksbUr/f6AnT
DpiFJXed6KU+NOTg58jHR5CUZ1Blse+GLboufYUZ6yIDu3djkD1ptmKC2FgBjtL4
DOKSAdeXpfUfbnKaO/FqWbJabYIZZGxTRaqVSxV9Ox1g3r4UTXb5vY/hoAL8cO1J
l5vM4EHbWhodtISTc37IED7xv81JMIEkYXT1UfEisGhWV9vCWT3lDd/Dmj5DEvsy
1KhqJopz9CWncI3O5E/Tm+3B6tI8Qu+rLkwvLOOUDdOIgiPMu4b+ihb3+6tmnpZM
UqaZ0pY0APOBSQt/PNAZ87+z3OcL8bzkwOZ+knh7s9XTLLqr+EHLVPVK7F0Tu9zv
qDj4DBAjytDGrgpdVeOpO3iKFOIXzMmi8Yf0FNh7mt5zsfP9xExla0OQ6/1wYkeE
iyAVZ9Tc1cSeCwGBt8WQNCpL3vOGJCCcQgs807Z6mk/7qCh8jPhiuJcjolVZzvX6
2LzBr9NSrdH/RWyV2/FyqQXmUdC7TztxKYdSOJeO8X1dpGf+oLYNulY6u0sVapvd
n/j8IZgDsWLaHMT8Y/bjPARKlxfpFNxramttKTldATyqv+P3XJK30jha2EIVh+UN
o2jUsfI4CwYznxlfzLvqAWVPB/ZHpGaIEN1xxocrm7YwxpjZ+4PD6o5bAZrReAyt
OXOaH6b1QGgwgThyuzy0SX6lZSD1Ht1SfgoEFwckXweL27AfdJLycfJGyoQO/4HL
/E1swSBx2DpACYE/kYe6p5lzjBqimVuQJs8KffHY8Ho6dpVChGLrm5iKpSdsXn04
yZtFBSMmrwtxPvRNH3z37xTU7z78cdjQeEEuKuGLXNyBEeh41RuLnfyMhPpdtFXZ
W9PXwUbsOerh32ulMAlWt3LIen7juBwS3TvhvsYf8i9SJCsXTJpN6YTuq8ccnJdY
W+N6tMr2//vMeiyyBlVMCnGWzPVgUWHz7GXtXuwcZud3dRUo0rlPPC5B0L0jiR0l
AtElBRPz6qosTJ3SlA68/1o1kTsfO1OsSX3YmzAUFzCPUSVYqo7ME5xMw8lNcSLy
OlmWovjBqdn36eLw6AMW5RfXB8fvexZjF7XA5CGgKqL8EXGjekDco2SQVJzKNhRY
1OA+KW0bE0RAdIhgGAKH8mmRFBuWG2rIkoR8/VPEBl2XgsSkaLGM6tI9C8oqk+eT
m6yO+p1Oz1hCAYHuzf4YKs1kyi4cA5Cjr+4mDO1WiSIugZBnX+/0tpPnydZCWSk9
Lz0dN+S7gU35w80y2I0E4ZEb64MRRat3SlnSuh90QKpnYNgJUwFzXl25Vx+JOcnm
VKnVYPK6TQkFAXMT7FgI+TAgRtNLUyRN3CkOFchYXFaMYWTOFWL5BOm2G3RqrgdG
mHniX3Ge0RwbnXrlXhc/+HMJUF3XFq+AQCliFRD+/n0fLcdFxFNWXDXD9VO5y1Vz
Jza3u/Z6tgWAm0/obP9t2JQkK3lsRl5SUjHV2ALwu3C9Qwh7zKu4FUATkgV8Zf2U
f59Pewy2jDj/hQ5+7mYGCtAa0m2+nHwTCl4GZ9mY6EK05DZ7OrEsMxnwRsLrCI8+
BKF/XLgCqU/G5+mVcy3ewjMeVUlQGyMtFuaFo1rQMS1agadundvxMC/cuD54aNLN
Tf118ZnCdmnnZyksyN2BfyONh/JRmTlPss8hLr3P60566cGu0hl8R2DVOyDttxL/
oXUGsWxLTZnEztpLX6rc04pt9bBfVEyJLTZcDypeFP60trOAmpzsHg3126BX1d64
uAUoN1z47f0ma5PyL8t1V92ncGd9y9IIZ9pz5b6OFORn5gM/EGh6WRQCmg+UguBQ
Py1yfM9pMp192pqZAnpQtLdZxD0HXeMabqLTApidF1nay/rm/aLIK+nA+IHr5+uG
rQV2M9zWiCupMdaNRc0npg8Sy/857UJm6zsqof1zB/9nargTi2CU3vCeVZrLS5Jx
o4MyicjN5/J5lgxC5ZxMZ+wdI4uBKodevyZAL5SbTHPDjilTnCpQ04N4OBXE4X2c
Cm53zvYhkFmhcXrlL3GyYGvu7R6LA2feM+OA8ikZoEP9j2XFZOmg3Y6aNZ/cEQZG
L3plpMDc9O6mwyesBP43YtVFJLYGpj+VGTOlhYX6M81RCYst9wLFg2/oF5odlLD1
4NbGBTTKiS8ZnRajWCF5jF9Aj0aApfInWzl92HfwjArb2KH+kIQ5dO+vq79Q0/hK
6U+VeBCq7DeM44TxcBq9NH8i3If+UEoHfZ0n1/5NmOwgoJphqNiwJCMCqd/6MVV0
oEzc/XBux7d8w24J0SueuNmhlUnMRbOMmr4TK2NqZWE8io7h54ZNkHYwRGM4Y2lH
pVDUL7JSxSuzT+TBpvUxeQGSKeOlb0NN20Y0SBwpfhAZylZ8IAsqKIpIDBT+u+Kz
tCiwEjUZM0Nv4PZLdOwFYt2w9Z636+R/AgTzA2mij9yRc5QEneyrVKHVMhUD/MRq
Nz/g1/wPIlouff08Nnno3SR/SeT0ommq8hHG2s0r2LCbMY5g3R3yX22mFFpJmVFv
eJJs3I1UskXfABZ6EQqTDVJltTvvLpz3pnh4I/JH7LxAMc0Hbl4Nekcebfyu/CDF
kzbLlJWyOWRxUxwDQ7MghQ7PwAcfL/V9+srzre7q6ayN52h7lEDl5o35C/6dr+mJ
ekOYo+8BFOZIlRB4QOQ3wgao7CBvb/5EQCQG4j2TOCNFt+ltTNGES7kdRn5yChJt
9JZrDHMkLXwvK+F2OCURqpqtSDC2wP2dNhpwNnQGwPpzP8uYtPJnCrOO0sbY2qvb
I9OjrDYBKz4eCZU/dsixxKgk/yexM1V+rZXjuPW7uoS9FvjGASrC0mHgqbib9sQ3
vJrU5/qvDp+pcrrhBB9mKTULCNfXkySt2WoZrFSzKt68fHQR24/nWfPqHAN/akrD
HJRS3hy+dQdfEcWkW/2pWDJ6vIrWPlCcsnHuMCSvJlEFG+w+p2vPLUzeC/hZpMUu
9CxTYYyh6gFo4KyD1g6P4fX7woxoJZ/PCOw9aKbw6X5i0HPRpV04BR8Ayz+xEFZh
rHO+jbU+J9JV/87yHyq8CTgiKk/JevJldq6zqPMulKIG3mc1PN3FoGgoIScL4FhB
wl4FsEFajZiYjmBzyfxhANikY67iyKUnO8CkCp4xU47GZBAiXdmxcXb4Kmhreipo
BU2vJX7rLZL9HXkX2i5CCY/RJVtwZLeH5cHPbdXuhXWVqChYUHztZ/mgNPU32vEj
S2LqQZQyi7ARp4JOMI5JWtr0IG9EJringa4BDH+Pkai9ax8iJX9Ve/0QFM8AlLlZ
QsZESgenslECVdIdQwYfcvuu4Ux9q0d0RFrjNJFuwVaTVsRcv/+P6Ph1a0IuhFd1
DRng7XpCJaL7Q7KOtGgqG1ZBYbOHCdirYWxIPsLDuYU4EJpT/n9j880F6nEFfD9J
QNm7/VNYyoqGoPR2zA2LWlKX1myWVwwQ7cswPn/EgUDhI5ncb1REnbBL5te+9r+T
pwY/EZWUBm1VLQHYe2hY/vMSLzf4EcZZ3Ep22/HlojvX2y4cNQSIsYa/0EVEjnII
oUisBiiDsjUCbNm1ajsBCl59TEm0CwycS6HmIWlzEFIi0klzQYEyfzOikNm6qPFl
Zqf+RT8KHaMEhWvdd7ykU59eOaTxBBAZxSenWH3yHvkVZOLeePEHQXAKxmZd7/Pf
gi+KGCyGkjnZ7yq95ElgpqfI1rZMgBUS2ga+6J6QCPaT+qiYJOAwVmNDMLLu0EyJ
OdYxUID5ovQvokxCpPNd7+18wjLPr7g21vOtYXE7boB1GIgV7y8mjfYpmWQykRh8
VrPJ7rgtgmx8VpVo3FMXnJoxdjnu62eJci2LAOdFH9DWKln5yl1ZTvKafIMCtA88
SUSqmsu8TgEQ26UYtRUJSYWgY1BJm9XQZiDi1nKmIu/GIhaGpn3+HxOzfQlWCv1X
GHVH75gAnb5iToSYHotNvx1zXKc40QhWvFNZhKB1+9qFKt7659I1Vm4PpzVJVhcA
JxfyEpsl8+YAhyOinOHAn9jVl4XjOmd2HBz9dit/04ZFeN74fFpeGC1w3RP1rz9N
H6Jtn8fellMJ2uaG3zdiVvSVAQI62WXwVqDRb1WAyHufnDFy8VvKyHuUBEK3O+1M
v3BrOYDhxYKrRJ/XfLmO+tWMdWYOKvE+65/XVTd66JDqGlK6M5/dNUMBAOuGTYyZ
nXpr0SRdE4jK1IlebZ/CQVZZNKlWDjEUuNVzQ6ELyJ72qkDZEvz4Abfyumod57Aq
99k8QAU9pYtjxET3enc2AGJ8OHxQWWSYsFCUT+X+oWnp7Fmb+kBzXCfvO62EyI5S
apYdlwRMH6WGGlzyp2vgo8BGMNdXyW958W39nvCNMEN5jkumj4RlCBrfNgYFTYYe
XGd+NBv4ZrMWcC4c9ncD2rRwZQ0ZfF54v/Xvmy/sh/TEFcKQNmxh8kCPWW53UKv+
uWTtgrOMeaYupaDOtghw/50lJxIICGg59fuQMItw7fsWT6WsU/9c1lPjGz3o4FNH
mS2HAl5OzPtZJqrM8o937zbUsYY/JMEfiNeREB++Fg09Ah4Sm2B3EJAKWcoVs1jr
l2+DwnphBgbf3jY/UmltSjw1pTnwMOaCRErmJ8hdoZApNiPmC2UDG9+87/u8oIOn
ROXfTMWF+bdWJqbDD5V4DVkRRNyYCwOLYd6eZEmAYz8V7jJiunTUd+wk1FFLlWnT
vRzd+9LcFRGxP6HTFPx0jfXiT3yxcaryOhyHQOs7zsCOkE74wunGnr6xVsZruJwb
LSsgjvcfoQ72lTcPEOKtPDT63HONQQ+4PCer7UndyD0enSyvP+i0ICFuRKWlSd+G
46gyXci4Tv9WOY2xF7TLeRGqKJYpp4oW9z8h9PkRxej5XQFkonQcHe1dr5sYi7Zj
1kKeLxT+0jsP6XR9RxG6+umt5K3WEQe5fUeGrC1C/CtsIR8r9xIxklzwzlvQDMGU
g0iSBM4/gbEYuWBGdq/+OZyfub4Y4v1idNOYs/Fq6K2HDpzBmEjGp/jPDCDZdb99
HCdGVuwH+m7t2xTK0nlesY2PFn+c48B0Hf3ABJhqAqtlM+b5CcyvasiRxP3ysADS
qxR9rc/J06S9gR1Rl2W/YpmvwCX203VI0Pz5q6WGJIpd0GsdewAY/O5O6UbuqQpy
COYMaDzw/MswrRCROwvWjxAuYGExHQhv9L7KjNiUBUS8Rb7t7eQt6To6SJL7XzkO
C4XDjn84IlFMs2JWiJeBH7+8GW64q+UVkHcCjxycUNdmfNanNhhkk17i3EXHmfVZ
JbBNqnsUdNNY7rZwJmAVoT7x5vcsxGK/SZjKQ6JsQ5Ium1LMtrVbQZDDqPRps2fK
ABbeqVUZlbgC8Cqxu3BKlcQhAu19hDOBOkw0lWXbPJ91wt74Q1fEAeehE6EaK//r
Kp8WM6qJtL5TZR3/FXClQJu/qkNHSUmuueyi2cCBJQgcKs4VglHi6kgmnwojXjJf
IeW71FqHIvXgvwx94yPgxDox389RSDv+YBakcpVucB8Yzre86dkEDUaytwF8rWI5
eLgI3pI+i0RcoNGVypV4DHGjZio8TdLF22pMkQaMn8gkRkQpcYdUbmnsXL+HI2N0
8ticfPaHaO2vkGlrMVR34CaPKXXZ22pupfOp2LyZX7FQye+2mPi+zUphPXsm5F6E
jfCsfHQJuX5SPk82f1n91PEhQGy/KntJqTsbYjMdoFJYoPw6iO9//13oWdMKKjHc
oT8ZaGL34hqwiwE7ghE0xJXRzFcZBnk0TKJqfh2FnjM9czkqmGAzuSng9GClkdc1
YWDm5w+VQxJ2Pr44v8ulTXhIAiAnxjvIVpHV3In0mQr4hMaPvB05U2OHJSNjCQYZ
8rxx9gho12H+VmSWPN23kdU7qXQ5VbvAfIeIeLzAj+B28guCrphPTg6KRUrDYonN
VV7lDCQNrQUl0dFSYZE9bqpj2pQfoADgZY0yOomjhTESH9X9BWQl2K8tKXzFLGzX
N+Ijw7ezWtgdByWDIPx6id7JrvcEhDHvjwHjc9SbwMX/ve4C67qKsrOPBK3LlmbK
h9sNFXKIjFG/TSlI0pIxKLbiVRUmpsba46exzPii/wMrytqsf8Y0qNb0vH4H8Bfi
gGeu1qk8bNqJ4tlTblR1Q2smEW7Gc4Des76nveEHQp+mwjLYVB5ycwlGqnZHtHNi
n5R5mVh55ScnUfEiPQO1SxWnjXRZu/HjK1u2kCSpWXEYNQc+KKcGr6L8HNeYFzZe
qhkK/S6F9MQyrLq65YyRr6Pl5DbpPWx/Pe20EbRm0htMUr9Fwa3+5/G2lRhBjxH9
T8DIBmO7ijy7qixwNO5pFQakn5sZmOA9zQLg+PcmJinZBe/XQErajQYTxXWRQAbB
ga+88e5E1dIO1EDbrK/GcWhT+A7LXjridLIR+hYMWl31tmzKaG91+jTWUJ8XTTNF
pPNOzpKdco6hdCbPa15C0c7DpFGVBN/Pa5Gv8FXBmtWU42t6Fgc2bV2D4y5d2Bba
v50EgSEm095B0pZx5hqdjvRO5qzq5/3tGE9zPZha5tqb7A3KyggGjR8qyYU27F7P
JOrcZZlJroL9bpxVWdVh7YvMLkEg/mvydkzm0H9Ip0ruTt4/5M/y4pL3LZz4t8Cd
vFFrv2ytQ2Kz5EdVu4VrEyAeDKiZ9S/l10jqlbHiTDMbLUREM/+UrlphPKfiCnuv
cOSJEfEQXDItwz8ELSNbEW/7HlahD9TbtpsxQ0SsEWpp/lgHhBgxPqOys6mYvCp7
+u6ClgXGjm/EBPhAfp/FccRyOUr5uhYlhXYyr42k6HywPKmMieNLOensEKOl53HD
NrGsB6jXTHGBEOvEp1d5gE6oLyJiQrAgF/p9gRB6vB4LP3apizeIT5X4z+nxa/Vc
l3wvO1D6I+q04UD4KwNOSJYHlpunlcziETA5WS2i3K35TZdrZJ0aku/jSrD8Phev
eBEEicChkxym7mJUndEm4+ujCtBHVs/Rv5fMkveUyQiAMBf5MeUyVu7+UC9BSSne
p6no6t3/t8B8t7ZQmGbdaRuJ4ozp2jpW/ddJOsu4ysnM93PRyusdWzbrcHOdWvFA
Kd/EeVoeE43kpq2f4+s4tACTcKysKjUVdTPDFXO14EYBbEeTpPSgIhZJMjoCkiBb
lZryraKYNdul7/2XMKmzfQ+xgrJWjATz4nGqXpTacawODYaMvq5JbZgrZ7UyhHvM
tNOKxenTse7C/4QqezkHg1z7duPQc+vPoBuJDToZMJPELp2dBD/oReW8Me+TfYl7
DjSqvIO1CP6T1CzFyPtYfrcSE9w6cpGWfFwjRdEq4D4VMQqc5TUn4Hr52FtsABiW
o0Gkkg4wrD/0gE8JifsT4lKOvDaqgnpQEuCy79fnGV5covEpQMrioKK23vcGllz8
9S/Gifu6PESU29t2Ighqo55yKSw87hNQOHzFWRdKx0yNapYSrDFCx71E8oM13LWh
pL/3/agFo0HANSt1EZMYLtaMuwiaktgeNykk1tVqDlKD7iHkKQQ5LoTXrsQClb+4
lzJmTNWy/u4b/r21XmO3jETjpkr87i975OBV0tW4PiHIKu5y0YYND2F9EpaoP9+J
kQh5Oj3KKdiMUzpa3QsG83TpFg9a6xKm4RgXEJkHtPXma7PZIAJ1EOo2RQp9Mlsp
8kY7Vy18hA67OKaMTHnWUIdMYwClERkwN8U6Jk9+Z1UE8xRT8E4Zwb56664uFh5S
T189hJlInfI510FgHDD1KwhnoOHyhMCN8A44EfBvRiC5ckt3C/PZNh/Yj1U2a890
M4vW1U9vrMgzfLQ/E2NeCIQ4jTC4XMdhDmeI4fo4P+ARTOFlamGbQw1diqsG0Zp1
kv7A0a2vaRt476rEITa6IrjV825EPeV/Ql084mszcMVsxCIzG3Doa3yQJAPBJFGj
nsCPIX7sij87WbaB4Bp3XxCi9fuVZofBs2Xco1F5sIkFpTPQFzGEWCC2bIZeStfc
joCkpPbcGZoMrsGEE8M5gMcowlV6613j4d3c46K6o/633cPck6mGvqCSnKQutkDH
P2abp6vZObNodVJDrMiGmWRSvdlKcImAfnWeZHaJzOuKI2QghvCYjl3J4n/AQoNa
NOrOLlxn4IwWNQ3AJsgwPseTG9ibPotK/0hg/3rO8rlAFgwxp1vyuTFnogLcE7WX
B02wya9w+vwQnl+UbPF8CicwnFK2wY8nVmii/iaMsWdpV2sXv377I7lC1mjD6+bt
ZTPupevovZx4GQjx3WzIySBYJO6WEapOcExvHYe/jGAEXlq4gtlIXy8GQ4nJSr2B
bV2++wWxNLXyEhThB8lfP3FFuhWjza7KJwR2x0IlRSMTDyMgqYLCk7WIThLEhDb0
lQlyl8x6kRPyaUFf3y1K38GeVS4RDfhhvjeUcaoeUkNgF2BP2THJ/fLlPoEwal3k
wUdSSR/pNvu2cYR9LsAOodv0uxTQRWpxxRG0fpHHLHoDBnKQUX/l7jhkbry77jdz
Kk5pN1CJgLCJvvLr0xbBI1XOJLV2lVR/7VQfyz67CkZpUGA8OVu32wJLEF/4lCr5
7a22MPy/tBiiz96njrHXLjb73bQfbArcV0h2Bpnswl/T7mom0HHLKKyDBgqWC5ur
giyHPJNhng9JGlUVuNp1pv4/2f1RHhUQhNdMxjSjbFRHn66ycnjGKZPIMwY0yPWv
DdhWICb1k6CzKxi9O6U057P57IwhCrIF9HeK4ZYECydAXR4/+bIXKZGhCgEu7u+7
vbRWS2m0aFCQjLx3uOZXyqdKCiYjV9GFEvkUs+f8/d6RZvwfzuYxhWhe6EUHDpYN
h4CogwVYWDwg0otBx4lm1GLr5+sJHMOr/r5VLJ6b3hv1N9CNT0ZhgY9s7hxD9w6m
gx37xfs7w3gT7EhG+M3b0L8I1aGrakg7x34Nac2JOYvHD268u7AWWT3FnvJqfkrb
wE0uurnzMY6xrCVl+/c0f/9gE3Knboa5o4eO7zHeyPKG1H2sNSY0IT7XTwHOp5bm
Un+q2LmHc1PdqmoFPbTxyVII4MTUTJq1JQY4mGzSeFViBgnxZdS6ffZnvB7QVcnB
gE6k9C7ujJEnyxSLzVA6olA+AiUkRKypPaIDOYafVkgbNPC52JM5KYV+BdS82p/A
gKXvr8nzx6z3/n+r+1veM4yGVQyotQxGtx73frHh6sA5KLpo21wkFyS1O3syMhJO
1jj+JibAH7VJlDXvDFXTi83HG6lQUWA+5Rg+2FZkLNQxT378AHnJVWUwAH/aDWgh
QuBZeb164IS1Mo3fzK0fO2Km1RhFHG7UTYFQRcvBuT7dGeIoG31ZuQcNrlaPIwWE
OkyTRHAn+vaOSxaWVex46xnf3qX0ehlJNkZgEhA0PEJnx7g9YUUdu1XrRdY93pmE
uAUP194vsCtvuEX/BbdoClVWqpiEWReAU+G1/leJ31cOw0dwCjQ4sFwQnZTPsfiP
Qf55m1+2qaW3/CffxL1MPSWFkDNIXwKm6rUwU3FaaYbzmggTs4hyVBZDaddhGPvK
0ptJHMOC6qCdL62BtD7qU4nWhgdk97eaFggvZdq7ZjdB+F6Wm5u9gatwVrBzudW9
LNpIm1qKgJis+oP57jeJSz0cq7NDZbiGZTwoUm6WfyAW8F9gWDoj+MKGekyMJAv9
M6SITUjCBMaXYTipywxBmbncoC0KJnXKPPyk30C/paYgbwLUidot0Ji70BH/CVlY
Ge1YUEw6D0kgXBlm/Leocb32LII8cAKNlYHDwThX5jeDtYm0WOyFmmFRjdFuuNu3
3DdkJbFvlsudgn/FfpqgPJDBSGXplKtwOsMgRtaGPQjFkZjHHaisbZrszDIkGwiZ
eIp+CTNY70ctAHS+VF9GSnV0StHkQMOIb5OwiTXG3UB822TcdcyNBdrSrp8Mbe/x
LgJbJuCbsiBBKzZjSLbUXqLAiOKLcyj8iDPy9BkW1xrBNIx+jH1QWRGFDJJQSrUF
KdJVbbPFZuhoQhRfbaMLZxaCsUojg6+WSbSv8WSa1uuZBwUyo2S+QldoL53aSbSl
/JuQcLh1YfeWWyPdPPfHibLYmIwWwkm6ZKVrCDQ1kk6w9eT8xaHbZMY7mUUmU/qD
UvpXrgKg+IwU07Ata8C/TGW95Q+lF6J+uM2ERaTf1kT4vaeY1Z22QgWekg2M3GP7
mCnGxzTsGZLLn05NBbklDUiCMpZMNYoyWcO00gI5qOQdAS7Z/0tBMHj3Ou8rJw1W
W4ToEQduEItGFG461pck+N1ovDJnhbxMCcKNH89ide2IDmM9LnJS5pCV1mlVOsCn
WHyZDAfe05x7YUP1Lsv8atSG3IfvWIu6IfVwBK3yYKt80UcVhY69XzGDWKMl5xn/
OU/sRQlXx9gEFAI/yA06I6RH39Ga3cUHnmGRsRsEWr7U5cM9FXTpEEqPYR6y1WbH
jaz5pX+i3xVJVt9ZItVE+S32OEIHiQOWcQlfTpKQA4C4Qleh542bL/FBGvBZOU1N
dkWdRqQDyo8kYYS6d6eRkLKM0uVmbcuMjWFUVo2E9sCcAPU29XrqJrgmwhkVLQ+u
sFYD/BpZj4haIC2ndfd0yUIkWYJ3yPSQX9H0FcKLvkuhIfmKlj9aqtjWueg6MAYz
UjqRNAHl3n/NeW6+zguhf52XmRRRGW7B2Q2w64xCSvzHslUhbZeM3H6Y/Nq9ihW6
WF9tbl8QiCBI5utlS9+pMAE9bEn3HKvs8/pjH5Eemc9Q+dnGs9zyQAK8e5FcO98c
ESXhcr+tHPby319b2z6refcWmpWF4F2sjScQLcpbw81h4vaJHVJMMSpiYYGfgQaT
ACWRIax9Pmd8lFl381RvT4UUgpUQ+6xEDagCuBsv8bg2a2sBKmfAIB3P7nhKuRCb
2dNpBJh1rLDa+GL3FiRPfe0yl4PiMyTGhyCkCxkQO8x5D6ZB2i1hdkSwPx38E1Kb
DNlOTQZPYR0ji+t1TBnVScVgF9lDCjYEBJMlIiBSLAnK1+5I4n6p8LUhQcKFPvdM
8Gg0tgndIgtARrnHAAAqqQNYh1XeyYtItAjo2fls0HS5Q/kmkALlCDGPWCL3qJfF
R+bJHibRhvFoHL6CMbRTkooy+pNTTdzEQhMIzWTIBO/H0QrrN37DgySPfb2e8PD2
JxoMv56lxQgnkOX7HjTAqd2A2iEOdwUQ2eH+pHU1BFMWgKmA+LlcBEbjft9iqVcP
GH6JLTo5HdDMNnjdjrVqMwi7rv0O6lKsIPq69Lu5Um4mdKkwbg7yJEw1ySskYXew
AaryIN0dr7rgTZbJVrtU7+6eWg/aQx/O6Ag1lT9Uzv6nTmYianw1jxZsqX1s2prw
IZn2rxzawTNM9vmcVe4SSx7p++Yv3ja4w2haoCqUuHMY2NpcatPVML/Bc6DfephS
yRCKT7Daflo3/4j/dEm0y/3vFEM+mlVNftUBiwqedlIYvRUnaHPqg20sPylL23BM
ZOeGChTmcZ6PJgF2ETIuyztnwhlOXfSjJJfU/36h6lktikUGuPYLQsuI2Td1qs+I
TPafSWI7LlIZ5X/A32tpLkcwO7bXaPTE32wtpO3bJuQpT/d0PlyemVQfC/WTArHB
ZNpbOKWgDrApfRlxyU8EEzSykfwJWeVZYgjgsmjHYMYZIYgUzdHd6Ocqhuf0vtHm
jvjK6i/073QwnR5fqrz0iHu8t81YNKG7rKUoc+BSlyzuYAtuzARbT6vYrnsdPSsW
f28SR31SF1IN6ph4dg8Btp9WcVVAaLqLnADYkY8AghAE+d9eIC+XNIoAqnQt5T7m
3aCiglhql7XXnH0vDt2yFBqvnsd1eJ/BohXrqwckSHOoFEsBHY1MRfSAXhjBKGmX
kaxrB9vtfOm7s1wZEDg4k5rztFx/6HJDPAh3tftyRHtcMVBYm67lgsHTWi9Eyqjo
eyKymQ68SQ6v3nCkZa/PtujmkSZrpgg9uKKP+mGyD+695CSQHwAB3bQrDVT2LfM5
xQP/N/IyGZUp76x2zaSTeb8mWMWW0ZmpJGn6qU9C08Mq/GrOYpwvBjn9rvS9783A
Q8oRnbp6jn5NlbLQaX2IjT8CNBxiNYbbzpX83SN1mQ/AUtOm76aN7vQQzAoJQF2Q
jLAx9q7QDMw5UIVnjXmVv9FqnB65p/9JiKHSQurWGlyj6IyglEIP3AJ177Jtw5BO
EIMRU1V1mNW3n/09ccNYY4UJupfKAboVsSDoUoRw7JA8x/ARMWClChQh5Zw+HvQz
EDg4UhKIqFfg9sK5N9YO6xhEXfIFUkfpKeBCqcPfj1oQydjIkoXu413WFzRmQCzg
6WyEzYX75l4wmIqq6crCwy+1OFaBEehA9A3Nahzs78nkX7TUTKd+EzRCXkIEmum7
9yDbAqtxxh+K925hbMjD12mhqsntGyxYRLnhHhf9R+hULQWFmq8RvcO8IkR+X4/u
/BHTpS9xAsA8gvjPOXVPQgaZRWvs5nzm6vbYISU6HuuDYMgidw+RbyOdngzPOXNn
o5FQOCRGuuY2DQm+IsmAGiSehH7UTtPULR6qBQXxI8n07U6nFXOSCp2LTEb1AMAJ
O9O+LthjISB2MwygE2vZCPr7mJJsrd0x+ytjg7qsbmF+sA2EMsnS6eKQ0EY5+aOE
4/dKVLeU2ubMub+Z82im/n6AdVXjM8GDsm4/n+gyFnH2iZQvvSf4cHk4m96UoRpy
v+28JbB8n390zwgyuX3XhIgFVuLp4wXvtNwZNuNr7aTrBN9Dkvb9h71tpeOzr32F
VjoRiRVqAcTn8PAUjcBS0srC+l9ysE/bSlZBjoUh/2v/AWWbe2ig8w1q70q3pibG
8vXEjmQ0ZcMxY9ONNP1opkJ/P2ys0oicTWoU/0M/wQLJ4FEZyWm095tjFUcJ7idb
GXVL16bTvMZQS99Kd5GJbYz2Qp4eOlKd8wACO5mAys7rXhBjemL03qDv+P1w47ts
aDtQ7BpGMNL0iodoqzUjjPsxisAGsMwYnvHY7aP9D+OGNRzTKnwtbxHXujd8tDj9
SNC3RsuzoaOdbrJahVO/esFP5ktd6P+iblcoQvKTd2xOvjw85ib4Yt5Q2OhmRTK6
5EvcVALRQACqxkcU7yCr71fkAnWgUCFdCivgyeSEnTeR4yVk9tvNWhFCF6S9+iCS
HS3uNi1ON7fp/MXX0/E+/VmZLOGG0NK0XIKhjxegulq3O8xEnXfkuf1j3CmScE5v
lXZZgmRxewKnjIT4xzrfgU8JEwOJrwXxJeo68t7S1qncQYd0AFN/BSHxHyNkERee
WBGotb3r1he+P5pMrlCIWApulbAus2M/wpyoUspS6Xf5l+oOf3sMIXmF8Oo6iZY/
quVw1OEvpEUAzsgMbiiuQClHAUdLqVNh0XShQtPBjPLq+XLIchNiILvUJ2LBehb7
9FFJXBM4bRmtSu+3j+iI4zxBcji9uE7kzTdNaf7U1dXPpJ0zB7ZXjwfl5H2nFVE+
lXUKzI0gRupw+ku3ImPfHSF1T4u9AU+X18EMoCUptg2zP1awSQLUps5xu8S05fJR
f8m6NlMrkflWGaEhbmNqMJ45NSxOKb14M3UVBG+mUL/pU0BXsphN046tQlufMn2u
CxpGSHaDpsLjqJQJ6DrpE5WtkoJ7LYrsjUNiWDVojD7qk2dgvwb4J/4lEpxQPbzg
wsTT7RNqWbOqjWAODNUJUajgB/phZXMpFRqKka3h2yVNOst6lyRgIYDT+cvLi0l1
+L6PAZw+VRDuX9EvgEcgY6wiHBv597vefE01javKegkXIrZZWjRHQExWyvYLBuLZ
6LGhJi7MJI+/+Frezdn2x3ym3OCyHxkeei6wAGjcXXlufII29t9E/PsEZXN7SfUN
FNVzCQ6DZqFBVg8txI1rdMs01iJGF9qI23Yh17WFvXJzAViu6cNMwl4pN6nFxF5+
kNlEDuilBOYNXreU+duc2E29vYzGQDlZ2FGIu0JqMFJP1S8ivt/sqtuGtSiDltAu
el4Nvjr0iyzspid6SC7gjEBTA+LmfdKgBEsk6mRcDaD0xMabYq11tggRp8fTSfaD
JvDNN80jgpDNmKN4zN4zX+hg6+IuJND/9xlAtBF7SswWopW0RLyDTmvhqMf5/FM/
WS5VeaifPYJMx2sz87DKI42/Z3FW3Xhs3Qx8bM1Ymgm9yXlULYbHUl01XRRJtUfY
5eLjns4Np3oa/MRyR8icSb20OBhoGA1I8lWbfoQ5sjKZNTMoJN8AAWiTvzpm9sDu
zlsjKYI+CY1ejLvM99nJHxNMBK19+KLi9AhP2QeOLLvjDkzWAA0psWz9CjtUHuY/
MH6/PMROBP+wfejGkEHNCV7CM6a5i5liv3HFogFEeadCmwx5fQcxI2nIwTgfkxot
cNM+SWwrXN1bWi85xwJarfLzc6FnLBBggAOZnm69MbkX/QeqZff/f6StSKJzgZ5v
flGsaVid+XfryT3ikcC9Q/rNR0B1MRz15bFeCmS1ZRWMq6rXtD1A7jLENnaZmQ+A
ier3DBYvGDqFpxnqjrGGpq1RbOQX6lCZE3bSeZspLrOFWYnh9ofghEj2jfWVjBD2
vpgsF91O4IbKfA5ScQBklBJaaWmnsgnU9gwonYbSEx9B1vAYmwHdzi+/zFPvcC6O
fg9Aw8dSB5P988k27SebhWVzl2DhH9hVR4hJx0p0M+4JVPOwrj4yCmvXtuzD/OWc
HCQJnayzrEbr2YHT5hvrTd2WHCpNNE9u6wjVo9+A7afMjFYatHzeAMo9PSFUHCQl
pOn48u6XYix9xNS9WoA/WyrLsuGIhJNPO+u0z+f5huk715TSanq4UO/MvHbGDwSI
6MCK9DKi5fXST4H4ZawB7Mr7sxr8b/lTSv+L+GOPoCQa9DLf6yMnfScbX/bxvRz5
6mMmcATvlju3+TfCFNrDSPcOIdDOwWThxAL7ZlhwxR61B/Y5/jvxPIBkvL+595Ue
xO13eongqi0PxoSkf9+lWNIWrYYrlmY2GYmoZI0HT+uFfQlah1XbP2ldIiIR3fhF
qcyGAUJXfOf4n2HEHEHGjrXQDfA/V7GvUVCTWt3HRfo2L2vPKAiyn9KXHmhCf2ja
Zdu9K3QGGVnuYg/2pwWWpu0NTKK3ewmoNyJVzLdtS/z6qR6nYV50rxLY8Culc40k
4CY8qI2idFHr66V2PbKPu636rFOoJKMneEcC5Dy2xCKAPLp61ijiTGz4cmTm4Az9
rWCvDAKMvd56Z3B3T3x66cv7bYKg/6x5xobbuEkHdLQ6jWV9dkOXq6tua5i0a3Oz
NzdYzu4SFkfG44onvjjUu+Jsqz5BLSACyf3hZZz0Dmv99JnStQfzc1BMkGs92rq0
xd27hUufwoBn9JEjYRdLBLoP+IU70h3z16z/dYtFQ0apXMfXvcy+o+z6lguOuoCv
rZy6Z1oTux8gIR2ypA6bVBzkF8nmvBM9HAGUZPdnL+jKpyNwDrv5adA4Iv6Aj6x0
914ERnkcLReGFG/uwqJHBmRbX91EWOYvOErXGNyORHMiOGeo73s0qOSaH0YKgZYK
BcHhg9QfLiVBfe9Ws42B9/DGJeyvqlpac7fR2RPB8qY3MICUuSs2C/5gVf5Nr3RT
lzN1ntC8u+J7UDZO+PzBSrIgi82DvFNy/Xvp0ZiO5zairIaREz+PX+st/8HDyzFV
LhWLO/y1giWugrWxmVEWpdC4qkIwZeXWQvzyX8Yius1Lv7qPEu97ymdDwVjMPhoN
lc4p4YoSms4mEb2ThQeWNYST0sAeY1d8eNYUlfqi22H6YdOQTEaAjbvBrhyDK0Nt
ZYrcRw0TUEetbWRmCCXA/+ocn4zoWNT/HAdNiUXBIMOucrW9BdqnPgouHG0PNnkp
xVV4ioR+rY6ZDKH6beCUGNNGiNadGrV7pBp8u5kDLGavCpva1KiFC/ddqqxspvD1
hocmkj8aWYf4CBC+VLSrfs46g6xbj499jcNXebsi0gBe5w33pAeqJ+1kfhNM2d7L
QH2xgRdAV96M5RKNeQa6zm2noiAPmG0ZfnROtmKXIZ61192dF3nvLO5pJtFGdDhl
my/jCMWyeSyeFQ1BZYAJw/cQ58c2EJozs/zR2qVvg+BOj801C2u3rQi3eX40O8HY
PBLF8E/U0HO6JDXVIMXAV0ObuHJlVC2fMT6+PgYz3GMJhqqV5vEexbAUnRLCpOy8
v/BySAb4bisEoEeXe3f8WqTbeK/22+PfaTCzEXktlYTYYzMNqiuUA8vxWkuHH57G
WmJPfCpMXXPI7MGWjqLLSFHT3f6iNAdGQULBVoPPC3VHJwq18b2rpd0cF2GeatOx
/2X+0Hm060iq6gOnychW/4KRiDwkWh0n0sW+Xd99pPNWSix21Y7z1JrkLBo8gJAp
dBHS9WADjhTf73QPKnRRKQUDzXQ5+GZ6gkI1mbLk0mdO/n8ADQH2dfAbagdm4HNw
+kIz3lmPBAIN7rasv349HZXilRTRoL7qVfS0rsm/LZOgqNVYVtTYedWflmJcME46
i5b+ZYHnUihtwHcjhIQltnZ/X7fq8DE723eWupY0fsqezno17IxsSUc8psOVMH3i
93yUl+AfXa6Ca9g4qkwkuIoJmRhYkFQbUteTL1pest49MyZP4umOkBaP4liUjwgh
24GbJg5PJgkBYm24VuTgkrcvLC5znyGYHzMG2HgN9fh34WSDdd9gNYorQtylq7Ri
VGwfuvdy0Vd0Br4V6UAFTAYUK/DjfmnLf1FJmsjVaXVwpuLPNS542Cy4xcM/nhd+
9DAXbpLgh86WKqgdug5412P843EL8Y6viMWmbVT+48GTGJTt+hPR7lnf1QPfLlGe
MLr+A0fnFN7EebrdEwU2ObBMyEPC0AKdkRtLjUpfRMDUMCRU5QUcLqTz+5GzkO0A
F7MTH0YyYOMndw8CjZWQGK6cQRsVwjOeS+cCxB3OoAOIZPRfliS4QXYSlrmZHdvp
ytJUmFuqx4Uog+jndzOl4WukRLOGVLglxuoDQ8+7nOUS1ABLseNokKxMt22btUT/
6BYARP7A4yBwWgEzeWUWArI044SBhXNJkEx/D9Sea1sFO3fnFX6V0mNGFalY7JLb
AixdiUFGoFfAdynUbaYLshosyOAON+Jl8RZAR25Oeku35YIP3Po83rtOnQlvDrVT
sbK0I9eu/1E3Y5tcMvZy28tqb6K8U2dzBuFWSW3wiN/5c8Uei1ZqQGpJnqriLe0j
hg7Z2uqJcP6yO7I1Wz1opIuxAXLwqZhrs3voI27/H21u2gtCbhP88KCXiAoUaT4I
XUlvslTaMp+BiQhdBLo3ws9VC5cOaYkCve4Lns7q5TXBbqQw+8nappIs0fZDRW+9
+nQDa4cnTB7N/SegY5WlAKT6yG/c/Tt9FZkDRf+naxdJIIzRdpCPeXvsmFgDAzIo
xLfWUe1VdiZJPeCtAlJA9c+E6RBNDIJFA4wuEaGvxmI+7WF3XZoruzDPCCIrH/NC
HLW4qpM0/Sf4NABG2N1IAFY9gdjONGYv3IWv3eBIPsVx/wsKo8o6z4GCZOwA+oQ/
/5DveBvm6d67cPBKoY6ngNyjVGjDxaf1hMqSe4MtnQSylAp5h0pW8vJaQicH8Lq0
J7EsAUAdEASYACMtrx7sn/zgpdDRn0gO2vkcEQpqrx/iTMVGc5BrrpoyUTotUx1C
ApXyDH2g6H6dIQ8NVs1EN4QdTBL/giDJ9kdnur+9GUszxxD1LtwO3yKJZ/fxIuNk
1wYLb5kQfTEyDT5hNR1XQKXsGD9S+253L5GBVQh0jvpfBLhxAUgmTzSBDy18XKQl
dShAR2eSnTGE4J+Xhz83nR4Wy09McR5GPnhEMnv1kSzEMVK4embnkti3M5DpkmPG
KujjwBerXpYjBdxrk5+jkGOK4YmX1xeD9/nhDXEDSvTQipOI2duQEO7zeCHVQJpH
swgxk8ZkFsqPRZfifrPHS9gup0DcfhMOrHGcHhE+A60GJTKxIgctJ0DHLHNmgVsG
QZ58vhMZLngsGdAObOOdXsoRIO+8JXTIeU/rG5Q8BG5NiwHXMduBhjVt4N2hu9p5
2FZp+BXya+DaCwbkgnXxaLGeCzAoBEbDvy8TY2HtC3kLvMkRVvuTDJNcDV+Q57Og
cHluDyt86RiEzrdr50DKi6G84+nr/Q170JfxM2roGXiZwl3Noy5ln7TsdrqRHac1
ZA9xGYYdJWbOJSCtQOy85eNuHIHUCnKMMcemA5i0dCvghVb73+DHSqqOWJDkkytQ
V0y65RofPrWsT/bnXTtnKNWLu9+hOnZ4UNi1asSfuQmFxK6wuGVZ98T7SwfqF2Z6
mIAvoeYmqO/7Cd0wlJnmjVBbP1MACGMnTkwz7CNK9eQ/ZFxAbACHJZagCl3xfa/I
zVZfE+49brc5l3NAPIbAb82B11snjDbzluvSMrsPZoYtnrKa2NB0Q42wUg0z5Vf6
thNUs3EVsvr1xtKzwTZrRzuJrEFg0QLRcEQh85rtYS5M22qsePUL9G38UJ40YoG8
o/iyKV2tQZ2UhJITUS6e0XcWblZDrYhW+Yh+gI8olgpGOyKFQxTP41hNHLD0NU0z
4PX+A7JMfQfH0+Hv8EwUle0ZdFqu+MnWFcv13uTirPbEL11Hgj3hqQmnBGUlJYHX
FnIE/9iyTuthJ5eEmgVsWAyyS2tXt18VN4tq0P1Xtd11VFg52pSKpcuPLdyz6wo3
TafrYE/mNspQMvGPzSKjKHBrgMDWb2hQkGVjzcmX8JLKpfFYQNyH9w3rvawxH53Q
7/DElT+DlE4EKGHql0FhZL5v5dK6loEvTKrLTIo3AdVnuTe6VAxG3id3JH6Qnlbm
juaJSK8sjiB5mX6zPcWLhms62HkxB2mX+LPTKDXgKgj6emvkampNiUExU4CteLLk
wkLiCITpcvQ6UT6iUC1lvSxBLUCBlvY+Z3uSS4ul1pSQvoo4CNIyKdWLD4gX7kB4
mlENbBUhXFydeoV8pUxzFXwLsq8Twk26fY4aFfT0zQIB9iDbw+2m/Y0omPGt/Ydb
Oz8n6z7cFFij7/7LIaIh1Szi180wn1jv+m4j2HTfpL+UE62EK/apeUV0QjMtJX0F
HYiUvQt37LhsF+Hua5/OURnVcgFIF2CMdPkMYHGh4paTOBrR4+anptx2J0SMHNgs
1ljSDDAi/GD/1IyM6f8QdwiEcdHQhYxurdJZiVz+tX1zGzgitOv7qbZ6d/13WW9+
VUY2ot6zqLh41DGUI8btrRLG6Us/gbsxdbzqz/ircxq+BgGLQNx4k3Upj8nJVLUw
FHFgZxz/Zr4NnvZDwvgvERtNvdFVkj3WmxpfCWq5p6swTZeCk3IhqhXErT87HLrP
lo9OOh3LGY3DBoDSN4P3NEWOGtithy1mT6UQqkt49nuqhu9LjlgiTvPYjQjrwan5
smsFBaIRH7HU8hHEgZO2r80h8vt5XBirPc1TKBp1LWaE7uEgg6u0NLKaNnFZaart
DS6zjnPmKJ+cIB8km0HmqfIYxkjfFme7QO3A4ITpCjIEdahcwBJUIxV4/Chrn62Y
nkKqFeTQn9w/1FeJl3jraP1pYSoDGebhk009uk1A/FA1ssi1/DRNZDytUvaIEYa9
mGR9WVOrjK0yXn+seG4wREzKyUezAn4RONd8S1i3hLoFb0PONn4qtXy87sJVRHM5
J/XtZ9T/bk4NArygbUQDJR5PcM/P6QrtUhwOsrwOyYCKeIQKkbQFDHHkXQ/2qbvg
O4bJgDdiBmw/1zwmhn0b1EOdBU0/+at9Xw8Kv8r5AnYrsVycLPDqOK4v48BCguk3
Xh/F0zloq5VKzQnutRw5KuoLAtNacVvKcZbymWDhlTejkmg/K5IG/1NdVvq+/u+L
QKTGvIhWRjT8nmJ0cLLAiyjTzPScRUkWdj8VsKoCT+0a29kWqk9ihnbmf2t7iEOI
uh6oTb4ooLseciZhkCX7fHsvX7PccYg7qak+ecrbiJTzp5ATvyL8GqZeZ6aax7YY
RAMq3/wCPvN8Gq7e7JSFi0dHl3Dv/dtjqAjvChMiEFQchkbWKZe2PZ19izzU7nLx
ty13TZ1CNBXfsJCz1AYOWQi7wQsJGEc/76Yq4aWHCfkf968LCJgl+PdgU2YRQXf+
NK2doxb7yv4WnN3pGcv6+4qEB8a2vVh8mvXATxEkpeWRai1dCQa+h0Avkz8lF5fX
kRCmVoslid6ZcaflRsxT8XcOpoyWfhA+XFqjsP3ASEEwxsq7EoJLAv3uG4ctc0At
uHO7P+mODIgYp3AQQtgndtL20Cn4qlO/5660J4UOtf2k+5Iw0o8TvoaiupGgbSLb
sQySzGijZjKqkCY1dF4BsPKEgHzseo+m6ZmwQpA02n/ufRtQChzPxx6KFZ9nql0h
g3AFwPFCZst7CfWOTRTkvnZEhxNeE9wcB0uaM+pi8V4X4tn8lWq2X0n72uruAPaH
8tduGAmgoWfSQMxtB/hw+14LxCyHS7JwdhIhXU4Hqrt1ThXboPJ10M6xoawJQW+j
VmxobAry/uV2ff9UsGjAO5Hj3m4AqAouBBGc2sQbI9vke5g+/9kT1Ke1MV6zzYk0
DIHSbgSCRBXnHK2OJpD5GGTIfss897R+/UtBekaSG8AmQG1PlhJ7Qz3T7Hb6n6a5
lSO0/7/qbF035olpn6JOYpmc+uk5+qwAVvjNoTH3vXj7HwfetRfH/A/DfFCMT3Fa
YB1LC98BuDtFCupv/BJgxb5QS/OX+Tw19Ehsitod8dPYOdm6sovHfD3elXbg2FT0
6Vz5DC7ZiRCn1ZWPw9dM7RdNlpCrbFh3VfTWIDM1a86kT9Qp5t+8TSnJSGnN8V0e
qIEz6G/aqob4TSNSfBv9H6BPqlqJhAUuuy6UP4o/1+Jrk+2FXK+ElrWK3C5ky7TQ
PVTUuNvrAXzjIMFWsvAwy0ZkwTT0gQARCai8esl7yxGlZqfTkDeN8LPnXTjZbCjl
RPaZkPkz1mCDcY5NHBch/uuRtGb31wHzV30/BF3OAZSguJNpqwr6N8f151DexjDG
GhXppdO/eAWG8i4JWN8k2TtgzEHnr10oYQ5cdCDfGBAr62+ufIebd4wiTjGys5Na
G4PzjbSuDeKDHEDWH+d8+Sad4YFyAVWgTheUXFjLXRxNzN4WQga2+gt4kaBTyYrJ
P/GojV9L9BefQcSSfRgedFDpZcCQPvBfiaF1g84lRSy0+HzFxJenMCv083M+iOmD
Zlq14UeE/13Fy/Uepu5h+5c55JbycZYfqyU7OxS85FvCdpepyvUDd7PpHaT59xd+
7eK9VzivtXOiu5x5eYc++xYOFc0KHWExJionDqMD9yBlJvR+ynTA9obIy6TguHye
FRi0qdFpfEZE4DjfB3U7RzsfKXkdGC6m2nvjk3tugcHvNbbzagGMW/+Csrjktj78
NA3zTwEcCJVgL2K2kwCGNaUfp7A8aBThFedr79FA/BpyI+fG2r7n+qhTtEDNztWG
p9IdjOsPF4JjxVuuDyfKlCw0KH/rN7fjIikIiV0ii6Fh3UyVmdmbJ4YY2o+OoG2+
o2CCkhseJGHcBi6fhtFGCSsYOlL3Q3ZwvgLJzh1CtAdOp81E/hMzQmell8oY02wC
LH/pSGylD/f+KFweLceHaPuD94wFKRvUD+C1+xTOD0fwNM7BwhAiVToRvTC87b/z
FNYDOcjLunuFc04YPammKWeUkTUVMzuvGywMAaJ+8w2CUqLXDSld8VT2Ue/TP14e
s0GabX134fxt6euutql85YtVJy9L+iTafZ9YJkormfh1trVFxclc8hkqJ5cz32om
t2T2n/+UH2Ai/BDFv9vJnhyaBVZYfRRQy19P0EQClkn5iz2vGDScTOWGI5HPL7HZ
ENh0dqOHC8+59/rJQcBMplFiiAmNkGO4JtLxdSFhfayI7H3BnZ/SBHFUTJgtTjf+
bmC8I3mEfCbjoYBokFvI1VJwcRe9bC+uihypTzUK1qKZbat5bX7B4n5c8et1Pkua
fsjuQviqv2ircY/lB4c+sDwajmGc8lgQLbjkX9ReU9d1Eu4s9kTll+ILekdPSzSJ
5z1YqcaKerXu9Opb2aPlzvFbKgfb6HAYdfDSWBDgd2+BTaw0Uym1CJyuFELktPld
wFcK6x7KKjB7jkEQjCAa61mTCjQdLNoOrRervo+OKcuEWynJWLAcxKdhZ6bF+pir
a/a/x0DhwKHQlYuJxIumSxY0JonVwdca1Wr8iM+wf2604vRPlDf5fO/0LyHLLBSi
cs5z7bjzDjwtX2IegrAfJ19TVeTHkddnoHFgQ7JNgTrprYkn2HMBXK2sQ2m2D7vF
j9+Jbhg1wM+Olaw60NpkMD6Iu24AIIJ3lvr+HOTuxCqhAhMwFR/nlr9H83Wx/nOE
t26z5H2zmcg+wMLVU+twl/TtW8A4dLxMmwiWXsWq+c0sz7UlPGIIh49fMQWEa2xi
0e2wPNSGya379oiC5rO2AOuxuk9DHCfyMwHQK1YDy+uBmK+HUAKDBL0Byfb8guJA
UaKyhfIY2kzdVolNrTEmYweAFcupUM/GaDKKM6v4pygHOB0gif7oiNqaiDKBiskw
1dskrrs9r8ykAq7X30kh7587wMsBOarKG4cDcxPCLaiFb+L9TKjYixhIF+4ykGyl
VRsDDt6OKsIoZNFdp1nSgfNY1hMdiWxcUemYfXiCCHANbjwBBwVofRexdXAq9U3/
Phfa2g5ZC5XSDAhmXoA6WtHF2xTNHP25C4H4l0a3ymeZO20euTEq10ikFJHWQflF
jOHbDOqG0XxkTuDgy1n9lwXHTxr6iU8qe288tv/4zs6Z+M35h9ppyuXwZZW7RASG
Oixch6OcGeyRoNWWorfb9Zvg91ftvk+vbKKeuiC2MUcklV6e2U/5Ym53J2VgljVM
5Ivm0qlktxw7XkcUqqBjT01XXZS9fYM0kPVnFOBZSapL2AtgRn7QwZ8YeYHzDM7d
iNaL+wti7if/yhGE9TmfrtHFRxY1I6IozHL0NaolKggoL/1rJKrJwb1zWKnqaNmn
E2Bv8olt6336MUWYjbRqR8EYRC312ueyzOoErH1MkcJZERx6dwhQd5sTTLt4VMLl
0+acic6QEEpdy2x+KhMRRGkIeRSFL78fhDNyxzDcemrmaXmSnI0hz477yLc0HmFM
jDyMvBH2Q6kKhugM//6kbRgA5GjT8FUN54cjZKiNQnC443PiA+TAu475jeNnc3cM
y0mf0/xQ0KQEBPX+v1pt+VWyksijgXjUqn8hex2Vrw/WIXF/r6qHu+Lndxxfe0Ek
vYnr8G7F+NPJdLT2OMDdC5/Qymi6dYCQcD5Dr+UGAbMHoHSV+lBgwxIuK221KI1o
Op3zykyJxtChHAynHwWMt0Ob/FL3o1kCf2TDwPiCnRnRl92Yc+qF8uFDw4H3HnLv
fm6fNGTXGaVxoOC6h994sJOJXm3nMkU+LoMxHrF23/7huJy1OkBADtX3QjfWVXNF
futQS+ZF/qEMnvpwfOWTb5iUbnDAGpSE/5+JsalqFKpKkySNs/aA177a+57s47XL
XU0fPQXL49SADRvIWxI07Xra7C1YGceps8dYdkPJ6xMQITjKDS4KC3JRPuerVDtT
CuexZS5ll6NhxmIgJe1hbixhAFOevisYrsI/Cqx/SGOiEm/uAnw1GOWpCIZjlCoj
IAWcLO0aVO0PjAMw+ouSWEoK9vaskw0Xy+RCdAANaAAHLnSiHbS8avcWzhOA+pEe
gxC+fbspgiMak2qTijwvYjTSYsgTq0GQPnG7/9aEXHNhscY/AVMruYRxTGBdbn2K
UFKrdAXE9PuQVUR3apQvrkBbygD/bM4zHax/ncZHJWMgEjo44HUynldchgJajpbG
AUkWfb4KT+esAZkTx1K+fHZOtnhg4GqREowUP4bD+oo4SqI8dV+vgdYcd/1dBrJJ
Ps9CLhclc5YbDinBQXr8x0WmXC+6BWMScX5rGqLUrd/a1Q/3B2hM0YNdQvLYC8Ye
Zp4BgYVyy7v8rmioTvtWaWBk66t89Lcf44dr/MX7k/eyvWHkWqJdJND2ZeP6AAK6
nvTXpFRDVPhw7h8ctLwQKjFwV4mFEtYhvRqOd6m0NPkqPV0m592+2rfA+Lb8oMT7
+KnLniP4htbcrz610X3MxFtWbY7e9QXG1oV/3XVmNh0o4+6gd5lwGDP3VDIH+6Po
6zh7b/DhUcw6TrRxNZn/kHD2dUnDNA5NZNN/wmxRVP338i4tUy4mrbQLOkYAj00f
FH65ue5MCx2A2WvGEURr4TB79DjpsM45KpufErJQPYcFgiY5pclGt0FoGFYPwihg
hVyLla7LH0mdaKwF9LodKul+vjZQZVISGXyaamWc3oUFf0R3iedTOs7MhkJuBWv5
obzSiiDTo4iT2JmX2gZbKOTX6V1eL62p9uVpL3I9iEU5Kwbq7YbErrCRTUiSiA9i
h588IGVXeQJmrmRQRO5neamH3XbotDeFdjplFCSy56Bkp21WnQXUQb9vdQz0urlb
8taiRKed0onwJ/qNFQR2dXamO6Lo5ZktdOIsWD2JB44dFmNW50cbvW8sq3nLHKhL
qTyJoz7aMSzeuCuImLa2Cee3DfYu0AKICxGODU9dP0r5epd9qdlnRDuwVM+/6k79
X5snv83OCurRJqLcioMRxJwq+dyFiS+sq2252mCRd5CvtW63KQ07sl/DhNMsvDrx
0Vbs5lKbdrZ/R4ZTWW3wdpZ4snH0SFEORWoQhik/DM2na41mg3GLFCwfBUj+u145
5tG5qgJYbhGsIQHhDVP/I3eXCTVG/P/SRgoo6EM+tCbUuSiadlgHHPA5Y11kDRCT
++2lf6JCvDnAQ/8vYuyzQFYK6WJ4JgSsIHHwfrfaQSTgdkGGqLaukBlb2Tf8yARu
QFKMXKxD07RUbAGTpzlrVtsGLUT/6HWBLO7JtbJi/AZY4bBU4HseHI+OjUMFlwxO
/GhUMd6grI1V5pw507yDRcL1S7mK98fI7q/tBxnG1BiBwV9Tas7rLo3zikmenWbc
el6vlvGBVQHSRkENpEqDBSqid7zTDdgo8WDJVMmZtcy3lyj2DzogGPynPWEp5GIZ
aeWqCOVIbGONdrjk52Kow3q96yPgpbTNvMOPsCx4tn5S65zO9GsA8zMyXCjhHrvh
MkLXD2QPhBRR58QvGMs+n5yMvmisnsYheM6ymCg4KKrt4KrYRRhVR1JEVhITZ6fr
6TsaZlIHhstHACxl0/1XOvFtccEXWzmAYQQNgssvICyi99DmDuga/qy4I+KbB1JA
uO2CwYGx3styO+uUz9LJQve84Mj5uf7F8qqNXIjvnaJUPBThml3YeXst+BD8rqCP
idw+KuGuVxM47iffGTGI8+rusK1RQzPVnugjHLBJR7J1NcHGuTaKLx9ul34o0QuI
oAcz0ktcyPNnYFmwCCfpNcfKo86zm8+Z/c40s9lpkNLM/+1Hp+p6j8CYeI1/csgW
zqyZRkDTN4qIRM09lkhNc8JkelrHB2BMtIvqRaFmc6EU2tn6RUi07iyiH6V5pAoF
moUQNwXnyi2EepZEvMeGm9C77mL2Al7yh38J8heFYRzgfQEvBabQvjXEYHFvhdXW
j5UGiAT3W2P4jrqwq3MsoKW90ut6ozgbEcAhPmyvBgM38bmcLZ7QShtML5CDccAc
Xtd7/cuSZQQZWF/84WLRafH/LFbZsW8wXD5fGNO+kNXvv9d4bE9akJ5UEefjstYV
5D73M92ajBf95c3GqHDP1CiG/KbIHSMoI3LPfj6cx98Zwp7LO1Re9BkvTffR+8M9
mBoZ8kezKT+iiG3Efzfvekc7vPfKtTJp9Z8ip853bqTQeJ9D3I4np0mQP6DFFXA/
UNwoHbV1s8U+ojNUTJtuuSW5UfrwEjphMbnEu+rbCvRQygB2kZZz6R3hgKcD2OEc
nYHQ1kK95WlaSJVjYY9iaTZ8DMjB/+Tdjj60nGc5u25axvz7zw83NRH6UUDuKRyn
vcUtojV3I0pAdkx0dTPUbg3xd2QbOkuvRPMQTnRgFDdC8jlA4PgXrw77JTOAuq7q
YDeMfxgJJQtfYr9hr86IMv8QuLwyreINdjZ8rOrlr6vwbI8Z7Bf4QajsvUqAv6/m
lbBtI2i7MzUhDudpE98ug1h4rPclym+6YBVbFshSjMi5RF/CGBbeqVI3/hsJl0Ty
fuD9k0OXdsqxiv4BlsTXu6pT3YKyIm3afeAszaog3pG/8M9tmqtLkKqld+mLIIxw
Kf6wQZXRpOSmbECW/IWVExnHOlFp65+22UO6o26Rl7gvabzFvu4hKG6QWoq2zD5Z
DZUgJMnFuQ69VED44tMn7oEPA/sDXoxDlTJFDAYYe07gR5Ar8In578OhcDWSgKB3
cbh8m36APgpILRyjQZ4FSrCbkldw/1ruXIm6IisP0OkdxuZtLOW/Y/vk4U+Ms0b0
kBXR2m9kZivnxgP3s0e+Q7RFRe5SImYZGv590LYtkHNowKoVAaRZ9xmJJvI3XGEt
05esTqrklksTEBzz3XfGkDImTnKDX1fCPXQi/kDSq5JZmWIjzIX4R9sMd23KLdIb
7Gb3RqSp4ubDEwlz6Xwkjp+MgU+67mrHqy1Jt5g5127Pj2KOByCfIkTvlCmsTKEy
d2ZW2gTUvEL2m4csmeVDTAbk2e3JFlTNucuHICuEmjrqwI0HsxSYT/L2YbFf53Ex
9TsBEvq2EAB/Tk6rhvhQi/legD1m2CgoVF9Rb40KJbwoaDjvmfj+FzNspeAFsXvz
UXM3ULWdJrksh6L/J4So6O65IYiU4fVBcqJ3B2hzsc1KYDlTLSMGWSBB+6rz32Bn
go5R2i7X89qYawppTgLJ9HM3s05EAUUOof7xlMwotdSfT1/k6JG+dci9V1DES4cJ
yjE8jd8IJjeCVedhoPj1bqyLFEi9NxNeqCDmFv3o3xhqDqn6sUTmflSLZ4n2s1LQ
upYmUDweF+Gk9NIyJV+cWRvZtWZ21oZVks23xH7I2vysQ7t/5NF74FaPl7EW1Mnv
oPz06hAcKxoG9gcZvTmjntFPV5Ewz7oKNXdh19kPi5r3HLLaf+mpVOocLZJNJYzA
YDAfFlkN+zOTK0vVk5xIm9CSTvjokxnh+JWnWh9inr1qhcznMO/9AsocVNa1HVwW
p/rmc2wGAUDYsbNfTPdWh5nCqyX7iv2mBwK2kdzZ9PrdAan4m3rO+vtYUw9NyCj5
ZKYqf0O+cLsYAQnLWouCdtJ7rcUiIWRsvDx5eBov09XToU8yWC3ZBoPT/LVbLBe6
qlc2MbtsWg/p3Gi7w6Z+FMm3SOnKQ4ZB96P+d/z4HNnTsILDYhxYWNQZPKMmhHK4
BQE5asmia3Q6aZjD4TP0hcpUOB7R/T4av3kz8iTp5095QryGqbePtCFprUzqTYtP
el5Sw5qZc4h8aJZV54znGgu0BX+RssRLuBUov/mQ/DO7w2rSVbBuGn5Une9zkMnN
lotIsrAQKWyungs+7IkObmgUREECrMezY2l2a/JuSw3EM/NsL+VpOI3C6sLPd6Ti
NgKmQ4hlabR6X4cKXRtPLLq++/zNIt/bEJk9CNasB+sN1+OiOmvYs+IenFFetuvt
ef67vcYDAtgpPmCV4cY0Yi7E+QmnlY2JIb06NZ9WrFv41QbYYFWeA1y7YdewSUie
Hy9WWYt67ZLEFxW33h+2EvbSe/4tj6tVF2KxgBhGhLibiSYZ0oa5JjAPWLRDoOgh
JCDZrBZIgNekdmSg3sHgcl7ZJjJtJocfL3ZGPL0iCIucPnPvYceSQin9BEBhtR+4
0TmTAwKkpd8MmmE2WDaZdR6CLsjESC16RUmi6vkV3fm8EI13NI+LJV96rOQlOCQZ
pC+mxRkwWKGlsOHPL8w9hzrobrtDlbi9/+9bwC7qrPDdWAT4lZkehdpfc4m7w4qQ
UfVN0OauA4suzGGlpND71KUpK1h6Ge5uvJ52ALfOm06sdBAlN14LS4jpm0FWm4gW
Q1nwuJeZwNeNjpH6dO6rDk3jeQpJUYTAEi22fS52fubhb0K3lzVmGAh/iSCkxu76
FEimuIoxfA4dfU/hVF5GgpvXy0uXTEz5u5oxhzmkCjoiL4vbNbKPtJ56JhPzd0ei
UYCva7l9ZspqE5iG3wJsYDAkjAfMjmGPL49Wm5WginJQsWl56PKRyRZt550bURF3
mxpYGK+Bi6gwaY4eZNntwAODV4MeQpBlSfj+Nss9Lxom2689gwDySY8jyr29zvXI
C6wZsnFvTcLZi9d7KYub8Is20hUKxxbVhOwaOw3TO09Lq6GxD0a9ikBh8KhSjm54
cDiSs1oseiXbNHmzU4fWpzh4pcL2Nyo9RSLlHpKcyioTakerXhwNG73l554ovoOS
anoMoXesO4MBxeDXTApMFhliCkM+qNUZyO1HvWTppRJYEF6hKpvKa1UOH3lQCLOq
PWU5R7Y+ZIO537f9VyjzAxapro/gdCuthXgQps8VZYXxYky1CFXeyMFq5oepae9U
1DOf41pdedpATzUXUhlu7eE0LizJ5Jh/4uNUYY45zt5RabjyUF3q+fppbENf7zVK
Ek0DOUDFtCLgBoziWoUSe5EBM+udHHu6mt9rq2450mYVbG+O/GpSM7rIy+NpoxIJ
iugFHVgQIdreihjKZwiklJUj4xChYpOhqH+aD+ZMeu7ZkZJ0od2QxPLLbxx9U8KP
tf37qF1SnbBtP3WwGJFkKO3k2q6ywyI+1GApDOz5Yb1TeJqVgCXW0TIpyNpoaw2Z
MNI9w0AAaD8rNGXuViICFFqHm15/+BE8MfNwn7paSJEGRktzUmN+7+zLKEvs3zEo
pGVF462iSx2tjUYTZR0wifT8qLWXnoEKrtgnBe3d+zG62F7cEoEDxi8EjPk5CQ1r
aAKN8+Ca/O/fZPL58vp4vnP+ZmGRaz3VmXUzLdPtvNdgZpFr8rjwx+IO7t4sOHUl
XejjgBL7LadBlUrs2XLV1O4OvV98vtyfEyUJzThNL5S+GlKLgWfNhWjr23skuXtf
lNB14UfK3cS1o0xIkfifvQ/emwWsM/+V0IugIYypTN2bw1QhFqdpcYRldF7NtXRg
7E0JFSWs60IUSsWSuxYTfI61UBhTyejGQveE1dd27YTQB68pwt9s+mQq8xrYn1Gh
9S8L8jDe7ILCPmwIimXkix5I7rrh5Yr3X+Rnmsbev/TD6spBj02uXsERiuTiFEud
JGadzC51ErD9T5exuD7aMTRWbja3JeQecpvnxUi8buwdiKV4I0Ll5JyTf+YZ/geX
XIpTlZYTJsxea0aSqzmJUB+71FU61vMlb239glOSjKcvVLHVLSkFXUuYm7DoLmFj
loZHjOBLeNkU1d7i1FjRTKmb6s8KLw++yh9UNs4yjJDo70fTCvYnmJ5un1+0QPg0
XYowBZx1O+3c0lniYh+f5w==

`pragma protect end_protected
