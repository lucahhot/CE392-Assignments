`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LYdlCvRCM2eIw/AMrP+p/GRBMxhKytahhKslQFD0Sv7Y5ftBXbG4HfDsdOxHhiqY
jzvVawchvaRU8m7Q9I1SiSPhOYEPAJMxWwfDn6gmHFyQnfjsVS/lp3bjNM7KffjX
9KoGcvt2AXbCCyYqE9d2HrFCPuOGvkgoHOwVLzriy8E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3120)
p/QTilQ2gAYOBQBPz3mFsPuQ1UFe0hi9zMMR5QiI7C4pyeD9p34ofDcnRrf6MedX
lnb1K/MqnPJPfwJucsLRNtGn03NFKRJerS+A0GSWgSG2dL7oVVN1GE3hlTHifAgS
jr/v3Qd8c/+SvUnyPMVwfpKMyAk5CgRu+NMXivMdyTH5nhqypHA7avlndmoRQa1d
KJtN/JsCOmf/zj8kb5taPa10AkqQaD8tdRhQI9SLKxIM9xvN6r0C6lIIY8ZwYYy7
sHhWWWxjbPIduPBDOq3MTwMZgRKY9ALylqvx0TfJdAZJvQYkg4LLPK8m+wHeu4pR
PszzhM/GlyEzNJ/g0VWcjHjeYVOFkzG9i6eawptYlp9BxDuNvx+4RLE7vtbFzU+h
emomGsHgv3Sb4prB19cWZAuynL/hGeQp+WTaeC8KhOnwCBgRGkRk1aK5E9pxrKzr
l65PX85Q99ae8lWHJfjeCO7Cjf01GM7pGlR2HttpiuGse8OikYIhBLca0SUf0kdu
8G5tS4Rqy6WTmrnO6powUOcTGNsH2C2wBQicO/ucbpjm5EwJMIRHyE0njPd3R/WN
ONGi1HMZaAOJbo+1I7OUY4+2ZBkWLT3QA2wyL+5vpv7cCEJKilAvfjtmEsAF3ljh
V1IVgYKQsHQxL/AaA0OF5Ag5nQ6x1kOppY/1pxGoAQNIhb9xCs5vHD49DaxNw/8I
JreknfBjSxpWVAbjDfP6YbhHMxpxywdg5BCxS9+Obx3GfXPO4Hv1j0lSuB/+0ym7
03PPaDvQWYO7P+IBDZZf4VTdgPrdnG0G8wZzNmTcDCw13Kj4sgCfhKATw1dYQZ7o
yxiwAO86/K3AAB4hKNTxJVx5TfKQ1RlhY9+DJnw4nFBfFKo04YdMfcTrByHaDkUR
PHlIWYeuFBboXkXdnVXFDBfJ84gPtNtQgbp8qd9woqDD/TQaelv5yxElTt/Vargm
GHUrr8+miU1nXXlhBwHNkahOnyAHsJ1lpsJfY4efiQxdpq6aeXDYxOhly40HivjZ
IKgAMTbZ1PxqcKcLn5NsiwHjA13ySOZiLBHhCmW86NN2nYyxc08f35jFzTdsfbft
F12KVTPD8A159XziuI4QzCS7n3Oqpyyb77rLqttE67M3F8tawJiPhkQ9GO4V0J9A
Sg00P4NAhF9DfgUFZxIjuhX/BI0TAyhYr/iEoCCKrIxVA1JH2Ntt9hzgPCfkZfWt
bwcu+gXJ7dbR/OrfpsVA6u0KFxa/KLIZz+G8fyxPF60fQtLFnjGsw0coYRXkWG5z
EUdRLrGIAHN/wnfF/gBif6odUywnCS7R3r2zHqVImLnHbsiob/n84gBvZblW3shq
mZ25l4Aub6x715i/nkkD+sJK89U0+J0mdSMJTJIIn3Y74/cPUmxiugB5q9pfn3VN
9WPEfE4+AxX1YvwPI+leArR7aXAf6Xyhpd2ivToyO9Ci/QJAklWKE7i2+d2zvsKT
4rDiFKu95cHUcwkV5egCcgZLiCX+epbYD4OoVAuH6mcSQ8ie31ndjXhAyfoIbn3Q
kxRTrGqdSrpY0sO+MZPOXiD5F6XFacjrwNOVw/uZP17lu5g6nqQCjW1Ny5qsepBk
6cYINFJvYRj7c/WWOUcHt8vA9lfOAY75w6SRO33GgD+OU/4LMZzMzuOlqdFrbl+9
N7zOnmL2sM4BEdzggD7JUM95a1QZx7EHiMqSc0psgRY7SQFbipJLoNccVZovNBe4
Yd2eYfCrvpD7jcYWttQzyseTdps9q1SXjwbfbBeyr4PN4X3nZzs/4ijGO147mXQ6
MXqs+dCurpK7C2h3I8j3pMC1AHgQBIwT2/sDjMlO0DHTaokEasOEKYgQCdGnEIct
hXkkiaYEXtmUxra9ZcRoUhIEABPBKKLem3KaFEKc41AYmdvVQxonm7LowwAzOEDa
umFP64Ckq9cNiveJn1ba3jwTJEWYGtIHIPYhPP7GjFBFv73gdGjf6hm5LC2EjPT9
34Rs7PiS78jEmqxscXpsT9GvEVKnCNH61B6z0u/SARm3BzHxRUbSBnJINeTVoi9E
wclGmc94/XxL+tbASHKg8Kh75MDp+ql+cSRPpycbyqn3jt575KVjYs6w0XuE6JLt
MZFC94GZsTWAM9XyQLin+rM45igsBYGH2jQRwEc8Gb3DHlpeeGWp4xlaGUp+cCCn
vCMDmBsfSDa0Nig/ssftm6yd/viZfHkPT+MN2FssuLMipydsybftfp1MDqCzsX5L
a+TeIKxFnab/mCBTDRrBFqh+BFWbewAnb25DYqaHMeXgIjeE7VlxgfcjDTxpHpat
x5ae6tzM3S2gMxh4U/6//L24rc0bnMzBxLhkFInTnTjuMBVcd9WcFnpolHrKlBly
3/OVRJYegZTDpSvlT4n37XomZP/P0e4Pav1zl1oMhvK4+wYpvaj+V2etPT4VqYor
9o37m1i8uiKAcKWk8H47TZ0k4Sws9O7l2wWGqppVnVKBVxosRn+qY5/HwtCdLrAN
QGBbIDF5xLJ2l4NClu6/UnHl/kALZQXItLbFIT1TmEkWpnHm7fXXAuRKstCdTe82
rB6MKdRaSwDQ0jCy2iVp30cEdKgV/H4/7Vc20l/mK9T8L8Y60qjBdFG2MSG/Ekfz
F1jQ6CI05Jb2th4hAFhdkIZ8IEktxRfKdwmnekOBwc4fSlby6oLyZ2xJA8rYg0e3
lvJQm0fMsaW/LVGD70/065mueuGrtwWpotgO8t4hggUsmTNbrlohVILoEGVltnfq
zZSwt/oTA5bY9i8R2Rxhyclp5sxl1NY/ogATaj2lpq+zDxyMMv0m53SOJ3KWpxkg
RAncReQjYqzHRMgV7IRTEG2HQdbi0d+zoRyhb+IyvUQ2TE+C42yQhNn2gIdNQkgZ
vwOrVNm4HDUppGaZJdY237Z5WPMlQD4hCwwOiPYlwQUrKpuL+IZjSZ3TYm8rAQ+W
vIUldL8ytMByxY8Nt0rQ2BJ6a4ErOUy2eaW3Bhm3hJ8jIP7+4NEfFqP7lqwUDeWr
H8S8tZmVnHh9tGwN97QMj/aoDw6T2ivKE0ytmAJktdvEfsaEZ7qqwYWIcwJ0kXNA
k8EQuBhrVRVITsoq7L//WTSkemjTWQRwnFTyD5g035NoiiGtS1abyzVQ3+r+k251
ZBMdkhw/G7dj1M5IKg8GkYdgm7mEPYHVBkhqoEYtPzJLVQtOI18aiphfPPbaOjOv
ISz/GZLcgvVmabi5ElvJTB0wSbtNSuX6A2tgME586gotjYV3pFCnmeMEeY3+0xNP
ZmcwwiEwZD1vj6NKut23DGChaHAl33lkcEN6wKenA2SpFl0kETMMz+wuBB6aYb8w
RNco3afMXgL8i9Q2qMkhkBr/dgwgnt8+8NNwf/SxxlRGomIMAjNMEunC1LCm7xqi
EdG4UCVIbDso6QlxPTroA+WNdkYkYg5RKKH6VY7mfuj1oUTlEf8BBLd4L25xU6Ci
B2bMpxi0PVs4+XxB4Jf1dD6YvPjXVVI+YH0vnkrI3sJZSnhfuInTof3Hu8qXcKd+
Vu11yFtFxIaQ22VY0gpAEXpseIBZ8QUBUa/wQeD41k5h2H/8ewM54VfD/Vtv+6U8
K+EZyXEJO2EosDAVww1+NufQTZR/DQEeQOEJyTGHFVL8H8xeN4X80hN4NIZGIRZn
/qZQLlYWtNhMVnS6LGtvzmg/3L18u+1zGgK57H9YBF2GL3gEXrznayjhpp08Ibdr
viABpdZUW0vBhfmXtB3wSiwrA+eilqJ76bmzxfJHZB/4CA2jl8z1tadd2dGRptwE
i3CBuG4xQ99U5139QmJXoLm3BwkTKiI8qlNogIxoaqOBc2O/mteLTe1irj+2CvVq
vKH6D5ZqCq0sS8PHkKUYWe2xeRIjrHWY2JIvuh0Q/hUEVRJR36dp/PE3sw2vC0Dv
10UwbK9H7m3xZcf/mojdZjSn0TGqn4LHxWlSitVqRGfjubWtx1rpYYFbFqvxcZIe
2Dn7OdodhWpNbgBZa2UA2yC7SBVondHb6yUHG2nLcK4v/WEPCYDztmAi9Zhtrbj5
ortCkMf1dDEFRlexVji2UbBVaQ0E6u4APFshpwoi0UFpK/wZtYHootVqLfuz9S0C
Ly60kVCL+PtSI+DOqt1wgoWH06jjOmIWirHvIGh3ARXEkb+urElwnPfLWtM/4HzM
`pragma protect end_protected
