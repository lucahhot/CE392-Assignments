// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
BAs+G3UkvqTkJ3WLTWrsvNjHJOZsWovHVx7W2Df7ACQYMEMYlifJ1VFyaOgyVfvV
z9FrNiaRKsikCTaLYYCQDhby12XxVyZPJ2BqUBI/vzmuShGYfdGanPDMnDglffD9
2t+vpFNJzM/wEcdJgQS2I0ZR3p6COTXeDiZAe66bLSE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 78976 )
`pragma protect data_block
TO+TuW1EqBQwgLly/0U0PECD85JTZ9hbqgTEdQd5byKXPYPZJQePohlH+AffvuvM
/RilpJUG5/q7OvcEIpUrA8O7OCqVuq92YpWTt7S16OVfcVMEj/5kdwPYEgEmZ+do
XPPGa5iZH5c/P1RD6maXVoJnPzFon1lpfHQpJPZhEO6mJT8E5Gk9BYI3PMp6MR/N
My0HbEB4fjZjbxhDYxB7Y44i5JKs7M4MHsmESwZ3yjl2wi1BDUnb+AMZzWvgvHXP
fr96LXBcazLXi9cz91BPx/B80Pi01KfZgT5T3StMrz0GxjZ4s62ZWrQP6ZOPr8M0
YOr8V2HvXDx98cJoW+pMWCg0TBnHChKpgK+vpYqv/hYoXvidnJ2LUdEB01ZRtJAx
BOyK6/uQ+Ul11vGW8eCFzMtVgixWiJ0uV6a6OCRjwgO68DppNy+rj4FyL+/n6IEd
8aLWhLEg23oPaqdB+5SZpm0W3deqf+BBJyK97cnWugu7Y8JcTz6mAnoQ7l6Y8c3b
MFC/Czl3m/1VLceKgQdGNbgyou7Hbj9vahMJvPT4kRFS3k5SCAJ6JQXX6PP0iWbL
e3yqvrPfyghblrzC6OcylG09q0Ty6ZHLykn+cnOjp3V5dkjY+vUEwj492euzcQDJ
a16J+Rc91o7S0BINAMjggzFAkJ3FNTCXb19/lap5av4yvZRDcRFTe6KqMMv9Wiuz
726FNJAGflGtteqclyoA1/7X2iEM36hxABecz1fpvIXlT01PDG1MknzTlWT0m5Wc
6t/++ZpdODO/B6QKo6ttHVwxeiZ9fpOQLte+GPJuSCYaWXqdjwvhSc+Uhly1u6nd
z/Oxpco+krB276+uoG3VqyEgF28efXleUDUnOQJMwcaT8jBe+6039LAXxpHumEq6
1tmutgX+wiy49igWcB9Cj38lnKyOsXeRl01RbdKnzGnhWZkOo0Za6dZ8UaB6QN9e
E5huzWBUFbZKc5iYlSiadanPovdp/5plfe/xB7rJhsr6zeAoWeH0XNv23pn7XLtH
7GEjKs6nQdHWPW7z/WIDW3Z+H6gUGXlLZPt0ZVOSY2td2Mnc2w4bAZEfWMMHszP4
8WJO8R9J87Ake3YEJ7wt+6epTx3muU0+UHF6JcWCitX/LB4qlAbJ84wi4vHpsPCR
0Yun1qixdJku4cw+e7KLTmWNqgKLPxpkq4NZuc2HVLukRYUPQ+i5BVgVmW7FlzjP
AHLWeXff5YuTtTht2OBcJ4Zrptd3yyMkKcrJng18+xcpgM3YqtliH9eRGkNSgmSR
2VbZzoFo39LQCvnfKa41sJ+Oqb+LlCHcT5qjzhBLfGO+TFFAuWK9ds3R0ZCmQkMX
OJ4j+cCRAlx/WI0GRKhJfbcfgB6CvYhSGa3AaSuEDrf+QcqnafoQRfUeg/YUauSA
boH1ZCJbYme069FkQeNHpDBxwviPBNJxyWfy0cdTWv7gHsgy1pPqkvaB4o9v/v1+
1l4jKuujjg2gUqGTWLLpHp2PoP6zMVfqZZw/50JO+KJtyWdeTP+GF5/IDJAdmsgV
CxWJbVRimgn6wS+zJdr+2AOyotMmGOnW7yPEg97Q4ak81E8rd68wYteU5M5JDI8/
4V+FimBKVYXSE80ygdTOyhWxNi81PLv2ivNaPRpbJiQ6XmTvKe2l5KA4vN+w8EUs
dkaapLHJqfimXuaKp5ml9DGi+yd7TCfzu/wV0+dwOvtS6O1fBWcUS0vL3jj9O4cP
KdLlEdrFcCEuQEJrHZP2dGZoR/auF9CYexc0H44VcRiQGtZNbLJLYvkxNz4jUvFH
WtmzOpqRryAmYwskBV/PRM3A2tWeYE/UYHidE59n3JDaDOWLvRDCmZNUdFv2prwl
y9WUDVrEQQZb7GJX4G/IjqZWglaEOLnrFfe45AY/ph8vry0wPjyi0sBladm/Jw/j
+7D6Cti5TiNIb20srEWWC8KZTjjYj21JSwEn21E+b9F9/jJ2TMtq/AALZXYo4FGQ
cG4c8QLQP8DkKKFLqBSoNCzVqx270Y01XLy+ES3nG4lmmXpfJ3EOEVbhkNIO2VT1
o9ZD8tbJUIVpapfkrDUV+NfsbylwuCFhbISQuncK3hwf++A7lIXJuHxhsdUiBEQp
/YM7Hr4w+zlWRtwVrqQk2MBuAksGfGnfyed5mdhngLA/qlP/65wzc7F+PPTDxNMi
xKA/uvkXZKgImGXs2JY5JdtIdrXElzuUWA/Xiszx9BFOkW15c5+MtLE9VhrZuAIV
IoFr1LAGx4hfxGsHaTnCQdqLZLkzNDdJ1WBK6iqofLVcO4WWQAww2fQ9uFHWTjiF
nfYqHq4bNhlOII9ksatLqon/ISpsxZjzdzgwuGSITctmCN6t+3a2eC1/VtFeqrmo
RVn0BT/CA/5AXtmZCrzDMyJ8OqK4MQRz9EQw4uJHd6Z5YkvN7lRIjDDbmbKB/Rzu
Ys4HgNFTaxQt4DHa30XyI2Q1WBIuRrnybkpUjrJxyUmh9GnSpeXOIhyC+c/mZz8G
FIy4PNwulr0hQN6Kggj1JBOV8KKq8d4R7KAq9jmnsPZBbg6744WhAJR8842IRzXc
mNTneLsD6Mfj5cL3LKf2FW6nCuatyNAofwakvmvlAhqHklG5+pkEbFHd+k77Mb7k
q91187LXleF3jZwic/JijpwBeFp+OnOzTjO8ojv6Ztg9BsZZy1shBNDgAGMqeXCP
j0tCozk6V5e/lT04M1GaPlFTHeT9kdKZRESOOHWL+0POtZLvadWaSnUzghZ/I9hs
TZPC6cYxiXsnCDxWxXbSWlJ2X8vppA07FACi4eX9cLgQWYfo0RM0QZAfGyI2LAXv
XG5NoGZboR76/omS0IDD7zkexaRlQkr9olkpdVre0sSwQCsr2lOVbFrHW0ZvbpT3
MhKaKQckW9slNzWEfqbFCAumOVW+eOgeGS+Eb79Xr8Dl4CtjBk7dMIg/kU6VEvby
1ZxDAlIdqiIX7qkDiZxfEuCA48Qk9y5c75sklLN6rAJn8eDcQqcgx1DP40VmtKRw
kzmdD7g+jfO+lHFHrKdMy/1QZtliAl+Ty+fH91JhCf7c9LcCCZq4ON9TGE6w7DUK
khBlTDtHKip69m3uXn9CB047NeMTTEh5ofZs9tkzkUSC8P7HgwN4W72IuEaqI4X9
1uv81wYfS9HYegwDDF3RCv7uW9Puzh8WKnbbuXU1ZTDnloAs7nCsAjCidiXxmQUg
9R5AVtuL7vas7XRacJZtmr5cAvAcTAoPwznlpgoDiYv9RNUupN3LGknQyszETPNI
5peRaytlqYKfRoHj4Odl4SaXlYS+9uQ6s8Nb3FfithoHBnOXAPvxrXo9wJsc1ABT
br1EgoXPVe/RADWmmozwRNIGT50fgoPJ1MtSa8SzS5fYekZffhkxl2MgSVl49+/A
3Cn19+51U+Djwr6Py26w379YWnM7DJ8EK5HM9yEY8/6JFpJ012S1u6GP2n2mPXhE
MflX4CQLL3j/RL6Hl+c5rcY2R6UByhv+dW0rkajHnmfeZ0ytKRK2utu8QTnBFBp0
5ZOKGTG9JVXUeY2DfEK6nlZ3DHJXuvCkrkw4Q1Xgt65Mo3/vt9bhbog4eFOyCU0i
BAhKjkveWUA+mXNKYFOLXNFwpaYjUQE9qymDT5V80DelJCYhh5nN74TIeI7sT6Mp
7AVC/cE3KCnJFc8d3pi5XpBVKJ38KO2rF0Plc9m2xbTM7PlZT2tJF7nYMnrCLiUV
I4te5yiN7Ktg2OJS6JRk9uhpsnKNq+2n+i4XcqOHocWk5ATTIkGKcj5r7Pv8zi59
639sVBvp5M19twMeLbroL/b2kPnaEOuq0lDlfkuHd9/nm4t2D4d1XhVuOLjPZNhX
DA52Duasb/fjLAXwPjmJG9aM+V3bVsN9Lyk16F6D0FQXA/SV/QzoCqAkRRoI/7xF
Vly8z84BZxxuZEr3Zxg6rlePSGsG9Lb6xq0mLrq3gmyqurBonvSFXjOBCBzuqleP
920gKCDo7J3dmWxRDnAYeHR2usLY0xxiqruaTjkO6sT7vwkhZsKUsVsBlPnoJwWg
egK9eHIRFpq9Xj06fculEBOPP+CBQ+FTmqHht1snG5aem+W++fealZVNN03pCShB
syOTekCEmzJrkYRB0Gr0pfRD5nRILIJD2ArQKHBGxE+wz2UBwmpIRXIGDo/zfu8v
34ZRdG+b9bLYLrq4A194LOYIK7ZZV68iXCD0bxCHNJmVGdXReBvXCspSYrLm2scl
HcL2QN6gXxanE2ArPykxPlL1a9TGyuP2gfTE2/nY/ydPoYRO78PxGWG5i7EQSXFi
UQkIcWK4ylPmPgyXmqxQKgVB2ZFFa0FYnACQpTpjPp0ep4PGROG9batjdvbiNK9o
iHSP3JSwCYUy+eFCv5y56mGp7Tti5/2kPpE907Xom5F8m6xBQKz8sjqjJZJRiAP4
Y8VBoa2tlW+k6RJ2FlsMdRXrd1I3mZRu2ewnaudppWr8CsZQZ1L2aZ3kE8hfxbaR
oXB7Vs2sN6WhN6rdpdYRgQsnblsoWRCQnvShZkLybsChVZmjqPlRUonf8MjChnT+
ZbaNiaNAbTJvpu7Ia3kxkBSa9d5jzngObvocizsYA0SJA5xERR4bXaPkKCchVOkN
vfBHzkdqEyJhpTffW7zHlGzWiKXl13Mw8hODwsYnlaEguDDEpWQo5i7LwdOeuk/t
G53fI10R4wc4E0Wx/H2iaYAjoloqtx3heCwLtL8w22N92SZP9d8RMB2qQuItn2wk
kpiqU4fWRDFiNvSVUPKj6hcRqv6MZ5Sz9FFlJYmmeT6y/AX5SNfbw2FQHkhNdoY3
4J+/0OD5VYPNlwBT6MSB5RnFEo3ec4tCfrs/FYu5QbMOXMKsT6odvOGmiFexzO20
yNfKrsKc9sqzwS79uDCqRj9ZwFnaRzLreLUWi/LpGOc9gr0e8oMLjD2xCgBMtq69
IQgk8HeXYnHjnHhxxR6qdMPPke2S4d3LKSjsNSAMwpZqHoN/VjUHGs2stmZde3x8
U0tjLpToaWMC3Pj7GoFOyKQKxFkbJKkb0IxF/BrdzVHq4pnyLeuAzYrlqH/mi5/Q
q8LqeJ5nPB8tsOIeoUmL1i8E4GPw6s4KhuKCXvAM+XBBn1B1kAY/5qfppFhlT5Tw
D8AYqTogsAuBg5F0aTmIol9UK46BOIC+RDURUoBcrbUhvMoLTsVzBe08OZ9dW3I9
DvsIbrysJJ2cCFTE7nl0q1xZBhn95IIIRVMEAaYGXSBtKX68ODQLMG9EW6Dwl5mD
1yUbaYrhJWRPkMv9ZWJ/tZN1lzaRJpu+DA0IyDlWRqg3c6QPJ9y6OybQpZ8KvNZC
yiklIa/kMunMfQotveqbgmNqo8Ppvp1SZ3TkUPBGG4MrUX7go0Q5QGGzN+hEoCQw
O/God85FFEQ70ZiIdaUN6aR/wzk7irnh5knhYy5i/VjTsWf2mIMQkwPwgv5DKJIK
lpEoP/feWEAvXilTR5Fm+F39oauLvac68s0uPeok58RDhnac/uI2XgEueuHu+f2Z
RiGnQIrYalPFD0jQQsCILo1d7GfQGmD9ujJ13Wx0XdyaJinG0SuIqse7ZW9p1TIS
ic3Wl6QWfhyYJfl71SD30k09lZRJIe9VxwmxUKe2qS9PtI5mt4WLN7vCdnyCL7vi
PkmxLU2t5pAoNjkPA4vPWQGfw7GSmmywlBSbdEgWV/Ij7i0dXOEWr6nSJWIQ/RS9
T89KQg4V27p5OSTjJktmFaP09qBz7iW/a5GrC0IpexN0ih+/fHAZet2xk44sd8fi
GKaECV2COj5njqi5+i2IOtAyNl4oLZQHZkRQ84RG8ABzJCCySFFbj0NbuFqWtDUx
9YUjcSKfvSQykGobHf+4fQ66xK+YMetFUHtylykjnB1h70E4S0U5aOzrdb0IxlJb
f0RYVGufonUM0NMBW8YDGartNGhjM5Sm60wn/P8gKO8BgucsL9muIPGYxAqibWSY
1SSVgj3uTq2pVvSGE4XO4EbYqZzMFw5ghh86Zmj7KQsLBnXP4qI9pgTgc0TE9ant
b8pRJQdDl4Xk1SISELuSRNx9oCIeaVDaEmcLBftL5pclBRdhT/q1lE54O7e+Lv5d
5fKoYDSARZZDQF5GhkF4KrpvXk9ZSGbVgiK2x9wJdmF7GFhz3pg9pIYcxeNbO0yn
9caSuJbOsJdePz0AsDIH2G0vnM+u/lDnmHb1U2izhBBbw+Dnjb0WTTElS8tnb/eP
q90Lm3crGmsb5WjvK+vWre7qg9cxtg1dQ3q8Fj3BgUxtNDBqFGS2fYU1M0BmGVE0
KQxVZt/9jwsKN+g+Su0mJsxc2PnY6v+FmqqMEqxWWkU3WBsV5vYqvGvn05nXlXO9
0Q905eFVBE9fqe6r7jTMktVeX5rGGO7m0DvbidDpHXFhZKmaelE0eeRJ4s0emoon
L/PjZrHrLc3W0o8DzXbGBkLiVjySv8atydoKTq0WZSWoP9jEWy24N07Dg2QSk0rn
YnLMsigMKl+HWZm6udLym+2UzxXposGZBVZEf7mDj8IOnzivjhh2PW5mzkOWop+8
6dqezmjgm51HxqmfpaxfxM6+3pRekP9BkXh9NVTDzS1jVc3zmY5ew0Rd9FZKsDS/
uuk4qFpDz3JuRN7NDRW7ijqcvX1Kiq3EHEr4hjf67U5KzXOv2aXunr1Y7Lsbo7eq
Y0AEyfZuJ+AkRca/Br1BIZSWsjJoxTkX/8NgOF3na026ZsX7SSX6uOu+exlNADw6
/VcJSOEZTJSNt+wCQJftYOP9AYb35hS7iKYseUnM8AEyoBy0CUf+th728fouO0Es
HarNIMtzOt8NUBVCALq3+a97xneNYZGUgPyatwVC2cFc1DyIa1GjOG8y3itnDiaF
oXNtKWPQooNwGaooedHhObmmphlekxp9+6zD1MdASgfyoAN9whqXJGES7bn8o+3v
p7Gzbwdsu8K5tQ7EvdCZmyxGJaGaYG7RUkmAqsL/wSfcJIqcLL3nOIP4bVyTLupY
TrkKMRLPSU4ISruF4VTy+fCmb1IZPZ3WxmAX3677ugPtb2fvZxa9rEfUpAEASocN
n60jHsmUJcqYo7xJzfn8iqPkJShk+bHc25OWbD+rrSIQszmC0s8SAG8cwzPCNF86
TQEvGpyoeyhrokUMHZFOJXd32gWp9Uh0jgJT0X+Lm6B0PahMlzNlMjOxdK9DTdMB
2DwnWkVI534WTtPFc5dMAG06pcXtwc5t9I7ir+YY4EQ4MfVL7rZHv8nkk2JHVRCU
aZAAgKGJ0vna19bWUh09edEs2s6W/RMiJIfADWP9RI5MwHNaNqDtWwexNSsSPhmU
5CERnj6KMD1AfIQZegCVlNrPuSY6kRmr3u0hA+hozpgfarw2p6PjtBsXdyvBx6Cj
LAIES6pULKo2GI2LhhRRm2fA6ZOz/UA1LHHFmK+2T7FzGZb6vXJoF+qwo2W6v57T
fgCGuIzkiNoheNCafEyHZJuOK83CyVMtYY2f1qrGB6F1U/nzGrpLentYHhE/fo5Q
sArpM7Qlo8r10QDJ9z+I7NLDaiOhA/gHE8R4wL1BF91izMcyaHTDPVhS7zh902JX
e+5QIooLbGwGlTp1Mxf/zRIss8h5AGFRwJMneoayi5CKwjKl+u67crF9yKZ8FSoI
T25M/oWeMZ3d+XBcN2aJFjp02BxaW5xBNL9QHQ9KlbS/oeS0atclCfmm1c8GO0BD
qR28E1TL2YPgPkBOkL5L9/ni32e3UmTvWIjYNE1S8dfgEnZGXLnO8pOJMPijSgKe
HjotaSVrwOEP1d3jTdJmQCKk97WG+gOT1WcmeLmRdZbJUtLVKt+nuyE1xQdaJZ0h
Z7ac7IfhgK20nR4rKm5VXuIcbqw7C0vOw0+tJWzCFs0y54KVzCA6e+hNdnbNPKFl
BN3OSJJklmbe5Q6Z+Zrf4JnFmq0JEvLdIW8S8eQWcAJ8rjrCE6WAgECxuzBoESlC
88DipRATwjq03iiBlKiBiA5/77jEmdiScsI4N7PnNHi/18Q92nzpUTit5j4E1Z9F
r32H+GQiNMzy0Td7tDjnTNzHlw1V5ly2wX8yf8guDR0/NuEoCVafqXGiwGwpnJdb
lNPBZtPquQ9Ngq3FJTDc+6wshATl7c+Jzz+K1sJJeIZY60fCh4eGIoY0E13B8BQH
O2u0J7pdEdBtZl2EbMZ/Ei039ymBl6k3DD2xy0rWCrikNbhVgTNtn7sPpfvYoykx
GaUrTy5eF0RCKpwXOlXsdOfgDVtSuiFOCYxSgmBIR418wLlfGjJGV64FvrLRPvfy
MutNhqevBVIZLaR+pKkIofH9i1UcDJjFbvdPgUT+F3Ob2jpu7zreQJPjGb/fe+G4
x523y2sYXtEFnRw9qjMDAeB/4qvBtdaUgq+YhSWOeGScDkylwlA/PVQ2vEm3Ooau
s7Fq+8qTyyMkq9RhCM06cQlWdFzzn16OXNILvjZvf8RfOBWPJHmh7Ps62Z+fHzCw
CC6edhCYqp5DJrIAtv9oZRftlCVLOutXH/kyzHRofiPVv7OnoHGO7rKEUriWtjZh
GJaLEQ7P54vCqK4Pyo2g+vMsLCO7WaijnnBJ1iBMcJx/JClLW4Li63C3bwsXhZE+
tJF2mPSslvQR8hzWaPjn7KZbOZ8yjL1n+I/bJRKP0anZDf+fBgDieXoNX56bX/Rb
XGFISMFEHpQnoWUnIRlkW8rmOts+7UYbX+yyo1/kXXnpiazsjlWHHpW1ysn+2PWJ
jL0qnr83Ae07ra1hQttMoexV7YvkAy777Wf3JOwX/dF4ZjUnP+8OmY7mi+mEtb3j
aItxJ7g7jLqyHN1flyCRlzGqcc8AA7N9M5ClDYlxxUvwShWTABuwXPpIYqj68Rpu
DikyRiOT54/n1DVtWObhWVVx6RZKHsXrh3buKLU55avgAU1YxUCVphmq7qWIRv4E
/u0uJO4hRyNDD8P4yi4qnQnnhIn/4h697PQJ5jdWAiH+5T464V5f+w3cRV/i3MgV
yIl5NWcenJFnCpING2IMgJ7cjpu9hQ38EECEk6RTauWNFZnk7Z5Urc4T57is/B/h
ivNOGEl3VlQ7WL6X8I//mAWTmkC/Hn/hi8YI9Vrwxo82rQzMREffcLMTfhRidlDf
TiQP7UjWA8hI+fHLGRP2g+s6hpcnfsWNtHrcICkkde6GuuV5OYj0jzQvv1ZLiXbv
qj7BJYpDpemvXtioqGpy/PpyA0vUmAdtXwtTeTEN5XD9MwVyhkT4x3JIrxoIj3sb
f2gSQzDsBUWHE5J1XUTRbeN5MJDOn1nfr1F7+sIoOfwgscqcSnSa5+LdIj2LY9Yc
BUrxg4vMU4nE/9GBfYf7N5ljiXWxyhssKFRggmXiA7E/kItU0qSpIqU4dGy7pwq+
SqN0Z9oMUm7EAl4M7G0kLG0JaUhQ7SNvwkOCT6oa9Ipix9+JAMitUaFQcfFPz2vz
kWVCnYQZ1npdMu0GIo6x7aMK2WBZBKBN8OFHAP08pzY9KTA8MLMOh/zqUOVZLlNc
/j2z+Xoxwf0v22xuDji0iUCzZCrLtbSIzsRv64g3gCYqfwqx6pSejGcn7rkJDWIv
7WAC1DOonMcWVzB4dL/kQcyXFfN8bWj1Y1ReDSrcZVtMVAfOv/OtriXX5sLTNNGF
52OQNx0eYfmWeIXyy2+U7BchxWRTAv0+0Vr4Bzs/nBr6HGpWb8GJGPe1tYerPIAm
BYeDnAtn1Q2HyWtiW5E2gpFroknu8FUWux+5JwweELUheczIAHH4JF9AWohparei
qmdErQJafbfwDI9GWVpoIKxEG++OfWjNk+xMONpAZOpigXfna7OV14VrWgyAx5jM
bqOJEv+NW0inzUlDMd+n9hJlWS/akbPsihb5CTtk51xWC4SaBTZQ5QMiBjOc3hw9
x9lMS6W/jljpwfLX8KP65HTQjfHd6K7Xw0gXoR7mWlukAsFKV9TCy5d9U/+Jx4CS
0hx1b44qJL1hAIFOZvqHT81IUf7sWn+9E4ZkRDhmfOzmEgF1VjE5PkpU0xRdzcOr
WajTUiE2/JakgBkNSjLhZ+5CpzREtZMclwEJtmdEmWlzwo0xVKH67EEjsDk5z7+O
yhwZCJhN0se5iLmSHLhSwOITdsXU2kbsPS3ISyCpd8vPTR5nv3VdwMGoYjCVj4bZ
k4VTaRmOtLw3YKTcRjfDpPBjZ2wQfYOo+7OwJqcliUJKfDiDXncv8woC99Y1G9oP
cObq3Xo93oamnkF7rdwU6Cl1GpN9M2iQBgzbgqSX3VwuBtKwWSnH3Cti9gdRNtU7
pN1PdDHgtnnGZdXzv5QQnvuKScVZHTenYE1+KmKofSXPbPjL2f+Y2IH2ww4mtPOk
FTQrm54WfexvOC1Fx3+FbObLj7/iE6obiWDKx2GQJkWnR6wfXBgzwgWwDQVVC+iT
XgzCxZQJGBUvAf9m9DZpeJJRMG98n7jfwKvCDlrs7dMDWAZaNntDWqYS1tolRCWW
+BetVLicvHfPXYv3CzIueGjHIvs+Xz5eFxsKDgQCs+lc6Mw3Gkh0ESoxL+XA+kJW
JNmXCP1HsywjaiUt9esIZITUMNqkmw0YIoFUiVb8+CgN6emlUuRqZnzzvcf+sCmT
5cHDcniF7OXMAUTLWaAiclE0XCn9+W4awmO/564s+CZSi/tO2Ns4197xKdUxUSaZ
3U4O5RYRtz97gYHnUjYlMmsHX07VntAsNeTAe6xLthrcfqSYDoP0MKa/+oi7Wgwl
AsW33c0xIKMYdYadfmKM/S2ex8I11wJ7c9FQIgRRnbe4ArcCIZj8NU+Kcu49WSQ9
WlG5eWeSoLItrF/xdjET9k6xArbCJGBQya8tSEwcFR73FIdpZfSvef8WZ3+Bif3T
Y05vVS4DnDYwNRiJtXsO2C7vcuDqrL1d1yVizBlRIkIL9wc//W0c3gUQJm9zu31p
MtjRYH2tT+goR69J/y1r/8fX6HBv6M86db3/ynyDc71ZhBgKdFVrU+uBiwfJe2mq
pPFnL8wS1K7TM2LnF4Bfg3gAqwvgx0ukMMhog5aPy9xa8cg4efjuJSetGwT8uuNY
ZxtPmnWGKtnPK6oFTCvC+d2mkKOfpDtWjyYM3KpNs523rjm/6m8d8jOsFx1gYhel
zjpdLXVOA43J/kPqH5Kck8KpY99DlixGlaI922ZOnv1JidnCiOrqzWboiefcfm2W
SsB1vlUAGts4r58ldIFUfqKM8eU0tBQxKZXzENcEJX07u2ZhHeKXi0LFva8Doxp+
oVtsbrPWQr7Js+MRJPfv6I0sEbJrZjOsYC66Ga64Q38nY9d4863uBaJrngmd2TFa
seZUJs9sFMii4I3rhaLTdT5V3MlLSSzFE+E70/yN6Vf0+53L8OIkf0hvjZbK5jEz
UeITAk05/VjmOwz1EMxxO5e/BZCtrnho1peY9XmHIDUQ7sxenNTirgoPRDP497mH
RM2R/rD3F4v/xo9RlQFrKTRf+xvCzyZZN5p1g21imH/8Ocvg8Q3No8RF+xZ2p4Lu
Xl8H4909oyM07BScsVw9rAEJEXV2eIljTj0MDp3xzuVYnb3zlCBDI7e34E9JO2+R
XvJH4Sb74tTsi+tApjKkRX4/YbZjc28Q4uyFxMNBgCaKLYeDjVHeCqbcjlpxcnd6
r8/CMRaqzLyckMjbDydkWXd5qnQpqdYLEA08MCP8c9lCgULC5UlafV7pPveXo+Ww
WeFe7v40Xjp9LHOtOLSTVCWwZA6z6qvCqBCLyhSMFsbOGwLaLw5f2gHqN4r0l/a8
HHasQZrbidyP7mpYvwcR7D4IbYq/0FJEGVqMRnZZvVVf6lc6SIGJ0BOKXKP2Zj0l
tHkhA5VfgKsJBQLHEl3Lsdg4OC0jtqP6/AJGZAOmGUwfTKah3hItr0vv08azBHP2
ldvXAMRxlUxl1sfo499jtN24jsnTIz4yFo886hGmflqjByJt1dz9bjlHWlTyciGz
ePCDLTe9EF2AUFsqszFx5/p99XS7tBfm4tOJCHh/YEhJ1KdCxV/ZMdMb/ruQoFhC
44NNYeogRXscmCOZThA2fBPoM+iPzZrJrLDBE6ix9Df2dweuZ2pXiKC3Pv1qQV/T
F1z6gojptfpr/f4IueJxzYZVBz4nmonWVYKZ6+go1cofbZv1bGal7gWwsn4SSIJH
VE5xMSHpjRT9Y+PEy+tBvqUt1ow5ljsAjdbX1QdHOcdgGHPXxXC885cfUzOy1sw+
RT2IrcedgMvLgi8S1g4rTXB7nwx6Fk8OmJsnZCWVgNMni7jVdsuixu5/69yunL7A
HY6ID4dcktGxUqaHL1YUzZCjHPF7tb2du85u2G2pNbT2+rFDutq65/YvjvwsACdd
X6hNz5Gsj5xCJUqYb938CFGxPb4VUB5syIVfC/nfMQbanBS3OMFr98HxvyfRHXh4
boEkhWypglE33KC0xVFmM3ySTGYSMzWhJnNEvjWVVchGoXxph1X3cEg+KDY3ZIg+
Fj0+vgHEsIcYbQFET2kBg4DH0K9lnRg+82UUg1Z8SrR/NI2osK9cBpCtS7+Xpe/F
xKDwk2CgBxuf5aDGIpCWvm2KWkYViqjh88NNUAApf1Icx1e+G8q0A58BL56tpxGY
+WqN/OxRGB6E2I1sQ19X1P8/H4qmpNVAxE72WwuzAqOTWi9SlyODEH4uh3JMeTQ9
3+L3AGMLVVVTQoDyQ+UIBp7vhHb0acUs3we1NthOyw0f987lIacUMoQaKhIEBFHY
reAGAw1iEJzK4pmKrFVyUjXG02/hVcwHMnaBrY+TjNMjRbPotbe8iqqSAgHc2oKu
/hjyBFBdmjrVbUFXZDs9BtIS/EExG0AqKM2NfwQTWUWZofQ6FvTXenCGUoCqfrR6
d6eA2vRtcLTOXWi06dR9ZorzNDjGpZywUMIKAZX9FZJu1L7557d6WBgArEY9AzU9
irIJISU8WRC/gGnb2iS+r6sLkADnts1eYafFN5wjcD9tOoVr1uEY1KczT9Op/9/j
hmjT/mCLTnPbEhLzqJIZ0xbB9pMU7nKYJFRVd1iRWV5V8eBZltZIH+uoaNV5qsWU
o5Q4xcYFKSdf6nfUqu3U2Rpa/rfuXJSlIplLoUmV9RqGhw5MFzoVzgsogEZmkyK3
WnJ2X1yfznGluY6jauDP3uKGFQ0hH1hXQu+BwREkXazEaxDaQ+ke9QVwkiulGHR3
llO+0tzpueLng92pykZ8pYonpNS6T4evpw31bLI4l0nhehu2gVbythSeh3n+paOz
kD5DBtY0uchGZ2SAYGuRdNvrM82hswgE9G6r7bPYEnkvBdTIZXlr+u82A7/x8jPe
igWXvXJr+jHERuf0ooIVJuFjFCtt5MSkv+83uYSw5jrFCLLZs3Q2kFKXMISY+/qD
etffp9MGDMN2H0vncy73DkjrUu+pJQnmIOj+0AdsLxN4/oF9T3vThN6ZROrei0E7
i9Vy0BETA1IdhB+5MyDcuo6cwkUownFALUPL48uhi2d5IZvtBDdkQNArV0CnsO8r
R/s0NdfGKdpi1DXTPP+cuFbJC/cNY114JoqqmdrMkJPTgeefdEsHHev4btuEEzR0
UxXqpPLUOK2yu6746w+B8r/5KokNWn6t1zG8mfkM+uLdKdKdrXo2jQ35OAiI+Y6N
gXbr54zfLKQhNV9+K3pM3Ck+AJ7fWYJrCymwDT8Er6pSylMifcRfxIE3xVzkuVOR
p1QvIXjwWkGvRAfKiBDHZZtmICrzn95yH1Ip00eUbKIeXCxHsejU5KPnlR2uBcbo
6Oz2nXJu4Iix9MSKpkY2iBTHBifJbRF1GST10XHBpj61tKyIAhyCBpUAYT/RJByG
YL/vbWqNM86y6dc06UkZhKn17XL0uYvXaCWuxYquRi0g3pVCLjy0GQS5OSsDFBOx
5+/Zu0tMPYrLy5iKjUC4yrSgIdDDLkPBHol4Bd7VSCA4FhSp89+mz+KkEMbL9OJw
8XtrcRI9OrKOg9AyV2+z5iYOVxRv9DzLWpUqS/ggYqw5N5DtNVfRaOzqjhPoICPE
wubp3hq5tmse6vQBthtCUM+VFjtMNNgZ6Nn54cvVI5pB/KCwjo0DPXtCS7nBC7YL
nUS9qneEcPViHoKm2E51NH8WTYVIuuXWndkBoktU3jMMK9Vr00WsRlHZhqvUHyEz
QMlRKhvBPeCI6R+4fJ6GLX/dkdG2voPb23fUWUznxqBgui9n3oyS0ZvSsQL0tCkZ
pEDvKtfkDZw4g9089EWecqSVvZZmuo6EngdiC5XqjA63iqbh0wuZpy0S55PeF9ye
5B9Vu+xn22Yq4+MB3pk0Yr71vZ/Pe8cToAXISIa4CQFVP6wWQr8LNqexPS9G9+qE
wfJujGmC67bx0KDZfQmds2hoM9/uZ9JngH4baL+aaXgCApDRe60/m8gLeFYVBVqL
cL8S6O3dRU77xKF6zIyypFdE7h30nYGcyuW54qgBSJ1YHxapw2dj94jChHsLOtQZ
0eTjzJtTDjusMub4ZnLco6HclkHoIWIKHQ0iqzq1puTRJnCCx59pnKF8ibF79ueh
PQuCkQVDRPCZZdo7hezfzoqz+Uwu/TcG2y+5zNcIVZaC7SIvqp/7FQZ6KATsdXMA
sH3ioh89DjM2HFGX/FskSW9YDD2iA844lWVE4/PcbY3pWlX+sGgV/6N8zgaVrnFJ
BJVHFSph6GOkmOaeJ4WduO4QRO2vsKM15THaQi6oebncFLJuE+nsNcOxeNFJOEcm
pXaBvJqQLtyY40d/gbjdvW9hBDI1BskZfAVM89QAv+CP5W4+c2NLEOa2073BM/bq
zAzTJI7eOjPpI7fifaHpL9JCUQKdKBBONXM/Ll8jqVcURypsLFJ1BMcD7AvMb/wl
7kj+0bQjC7vgd9EuPdvLjrfTOhJ5PQ1FUfqpddP6HngQnYkrCH6QU0NqcCCw52qT
evJ1vWo02KbNTt9rwqfC3p/DlLZZMiIYdhf9nYXk+QsP2XyolR2x8v9chspX+p1I
usaOhwtnFAQN5Mec+piyrzuIPd0kTAG3LceaXCcJFIirRr07M/wO5QeuH0wOQLlh
ojAbgEX12sqndetnne0SpVhb8geJibdaf6XVakSQdKD3UF6pg2UNVfJWtzYGf96m
0h2+czklXTSj245P7DxXd8I9n7QuP+wZCJFPDB8jLx9sJN9J5iUFBlMBjVwGP4Vb
COmxnFMXU5/o6d85B8gLN5uSzJT85Xmhp4KWA//B1Briq4XHLFs/lYnZopl4aR7L
vqDv0xcZZBe3DlkH+9IA2oDjBVze69B/Cz93iLGMqekWkhNPTpXrexrTx8ykptdg
M7P7ok2r9dLvjsR10It6H2Ml++z3CVX4EAJwtpVZbvHS9ZNtcNkFStoV6m0HBCQN
tKJ6E3tG1JcvCdIgFmxIEgyjs9eI5uSvKqqqpTqfjqpLH3We6cs3vQR/UirKLEHU
gTJoAJXWr49mmmi9Pv1Zt7DP7Rhsf8EBFxLgSz6zBSFPno+pYTQMJ/1x+MKhlU3t
9hnOkErognKpk1k33ud+9VCpMpw1ppktyF+KksHk8zNkzA+gfU1asDtrR0JrE8Vw
Y0hP7RYho/gAor++1AEd5fpl7Wl7O+37YEvXrgpzyVF4YZ5Au7UTq477daGkGusw
APGzl1yaar8gNNh4lw26XMoxBBm66xuRDFGv5opZlH4UcRESya9d+dWEPcUt9XRq
/OEpygoHqW/44jBBL2/mLdDFe+Z4/YOJbb3GLVcLyMPQa/paFP4Z6m0ABa9NBmoZ
1TNr56ujghXyMOPCwkAcYgjq7X7moc9nNjqhosqcoLLi6wcJ9knCM8puyyrWt1PE
0bfniZxFIBdsrdyhvWENByXr1nqG+fMB0ca/1G1ssYOpKC9Au9+RlU9iy/9zsIkA
5GP25fm2ntpNYocFXVPUzQbILDfg+lCbwv1TA0QQWqPSAsjLjLdSL4PK0zcrqgLH
baysR1iAIFewkxWiQbRQqQkOPA/F9WJSPrl9LrhNE2VN4yh9SmTA8legM9TynXYI
mGdSA/Jel9gXNGO5qBqlc/P4VvnYEUHaw6CyqqWQPpCO5O5NguucI5Kr4OPSLOWl
/ruLNRAqn8qczXDmDo9wrfewiyZZWA0hZUNtFrA1i9gGu2lJ2xeDVrs95jR1DW5A
XPPR7RXrjl7M0jZPkEsEEcqqIrjNdVsXfpShlTRFlfpI+s/PjVRtntTzv0rCLRpm
MGqk1n81flMGK96nM7wwjDmWy3Uk4ixbDZihPVRnylzlS3/1ZPAKa3pvW7i4ZoUi
lK6rQbUT4rH44TumJI9n+rGbZ86bcF5+wFeXtqkRmiWkrOwDtbt9WaGyOI4s84ky
LtB4zYoL+94VYqW6edBrBxr3UT02vRZuBGeqBwx+QiN0HVTkKrAAdA/Vl7pWL+tD
DJsAi5fQO3DVLS4JBzN6Ti06TrLRIsFijX6Uki+B+li7Jfgf6+IxFB8PaiwVNdMl
gVOMG47v5cIBf7EzKh1SA/iQhRHjgTZGB6bb+cwgCJQX0pPGzZpxMzhUgwFqah7D
oSLWgeaUIhk1Zoxk5xXqlCwTmZi4MXGRC3JGAyyAeyAvEoVTA8F4qfDgdNBd5tbH
zNq8SxhnmEVO+jyWv+PFWpwPTkPC7WkaKzciUK+jCHEwccYPCnaaKi8L8dZbaHkr
bAcJRUSXHf+QD1H4peGZzt+RXbAqf7q9OAmfub5LOaYxWkitq1Oy2Sog2zq0aU5x
CT5DwNg6RnZM14JnPFDIoZw56eSSWpcWaDqpVoRkSq6ls8cKSDAl/yK5GJ77+i1a
7+4Zv3XO8MSUiy/bHcm3eSvZf/4GxM2oHA9O53k7p5Ve8BVl6nuO6RroKRNpt98S
XdH+4f2v1sWeVXoq4YywxDePWmEMi38VFWEhH0pGMJYvFEiDU+m+FAdBtuzFBAS4
zycvCnyLNehdzmuUmB61LiXxd8rZrQSFenNkqBkVCCDJdyfTZZV2R3LSMM67h3X+
tUTGfn9KqvwvW9RVhWFEfACBlDgBEBcElueA3uJVbEPH04m/2kwzmFH5odEzW5xL
pCw1risNapHl5xkTFA3EeSypgTOt/1sfJ/6yQ7uValK8DCstzkK0EBc08XRSkiwE
1sqwlzsCQZ4PqK/S8cax+7MnPab28dOcXmQ6fkKzxkJ37m+f70sgaBZZAOdmqAKv
bhU67TqavUeL7KYUtWnLsht9q9b4dJHV0fNC+LC5PpYGhf8x5S6EDaMXCCqs0/G7
4tKuUevE8fMsj4GVpuhAioN8rlyn5CuPqehIzQoKWuSRXfAkat/6HfUR4EtPXiHu
flrXtMJ2hLe00rxg+q77bvaYVltPCA2GuBEtYPusG+ULzLu67VHsVbZRyfO40feC
xxBDLzDbsLaiEHJtKDVf5poNszJJDh3Ls09Y0w66bcozLaGr7E08BzPI9mJxfMGq
QJr3L+llFz5IMK2MCHnk2N+LHWQt5k+UJAUkQYQ+WWjZbwqLkM4yck2g56uBEr76
vUgWv5RTLmfczguKNNlawuH0zie1gcqF6J2dHB5cJEc99EGiLJVg1/hNvbeQhX4/
VFgIMyMZmxD+BBOhIHpQIlUxZXGS34MCXgxlldhrypL7LlUaBSztuJj7oPnC/70i
1/6QkH8mnmBtjc4XkJ5snBfKnODL2uQZbon4Fo93uX/iSnwJ1Q+OBfhANPG04xjs
1EQKjCV/OybtGTHjLIEnJHhDSjx7nYGtWdojx733/cmsex7wYZBqMFz1hyfJOWaH
FzeY3PeKdTFx9pVthh8PjBQcn45zZPZIqVr+W7fDlDjwPhFE2ytiuhkRvSnF8OEE
flmNmMDDv0ltPX5NVzmbTUBcDzNea6hYzZVsygLNrNc99DUHfE5J5vVu3pcXwpci
LPD8V402nNtfYl4tog2DSMj2dorHZqYhqJ37b7Oz483AT6y8zqPOWHbIyJmyMTLG
VQcMvdJAEDP19RQb64LKjChE95Aa4aBFMBK5JDPPf3E7FApelrxsJ5mj/T2YQRWH
VLjVir0CQrJYy9OGBVXB0nlEITRP2qcuKCU9md9k+XKDByBM1E3NFEYlmLH3dryH
Dpv/Kyk9PRMekuEu26CKfH+fLbMOKfsictmDNDXJ62yMADCEW+t5YDqpbmBhGfZO
CR2YFSs4WToHMTRI5USNCnJu8hQ0VhU+wwkQgkkjGv2bEC1J+Onen51oscUXB940
hoxJNGPLuTVyQswWukO6EEgFR0ae4o6/jhvLu9NdfgS7QNy0WMZBCFXIzS9lx8iq
m27ur1gIzJyHjQrk4VUMNnT8MJQv5hALmhEwZ1raEHPVE5A5zLvAkELhhD7piUTl
6p/7zKyTfPTAEQz5gte1G71hJD7a/s67oD5IgkV32K2lktrZlnTKXYKJjsczaHNJ
c6y5dqI4cddtEfUXWtVc7zurkPDewCQL/+7PCkSztntouysn40k0/ArSNUyaxD+H
aOxt3/SiATUjZfxPlHXWHafsCLcojqDInCuXWEc+D22kYR4koSVihPhXIjd1pKqP
+2t2A7p4kQPiyi/DrPVW29D+xCBvp5AfZm+2zTi6l9PfsdCTnykVNjj0ydZ8yvrP
DGI/nXRODNSpazcUXVreGaC9OY2cTAUlb7Qz9o32Ge/IRKt9VzQVM8G7l5MQ3EJU
CWVlelP+uQqNi9vG8cNvP22+b7VNZB266V9R9biX1q5QkBYRYdL1ymyJUcjzuOPX
mv2RaP8q2jrIhvZTMO/om/UmDQGkSKtfp32WvBLU51s7gRjeqfzBM/FstqEDl/jI
HB48W3MTMD0rvZ/lh39dUl8kq//WYWUQs/0GWdiL1svhtSECEXQKtXKc+Yx880Zf
QbuPrgZwvz7cpuOzCA2o3qw17w4JukCBOlW+x0oVg7lhYsuxFEtEHQc5W9Df/TGy
wfGE3NiTGIAa9ToB1gpk9B5k3lDZ8xEPAspkQWtmD0kqktACNRsvRq0HXgKx4t/w
VObk8+PmyvBNG/WK/2B1VcbaW2UZ/YJwidizz+wISgj8Bel3k+y9qM1edJ/xlUa9
HcqYoNcKP7RLhZvjHG+oklzedyhGBct28CCXL0aDn+qjL5Qkdn11utDaSouZK3Rd
AZTc34iQAU0FSlKk+J5reOXrjggadMoQ6iM/AyApdCon/MfL0+HBy3BMbWL+BfUT
rrby45EDf+w4mPBoJejaGRMh7sa5ySQddeNo8Tibz5DxT8w3FufQwrLEvM7MWUMq
9YylxiWw9DY6RUXVZtrp3J0dXzWCQ+eYVq2Q4JPEi0nwdSnzjftHWkzHQR3LL9Mz
yrxJIZJlx0Z+xR5nuDtluol62r8Oj0tbHXslyzQvMyqOby6yfFeqUjopnp85VS+O
YJDviq+FxK8MfxqI3u1UiKsu/bM5K5kHzDpcsYCOT3wn70xnIHxUkvuRCn/zAlv1
uq4JvZXNXkHwFzXA9sWGKgaZM0siFugUA3XAgVA/ZTkqG/LB9awps8CUWDlJC0FX
Wpr7GE/m4nTQhcgQ4WAkWUqCfwsVOByGmqYsGn9OVkwIcBAKmV93HZ0k/XPS7dy+
RiQ6otFBEpd0YwvktByipB29tU7ugTvxOPy9BgYP0hE3ImQjYOcJsCLRW7/9HHIE
ieYGMVIrwW/uHergNkxbieM3oSJVv7+zfjUj7ldAYcphL6H6wipdgVjXbqV8gVFw
95clqOXhX4M/OTHqy62hIspFXpskEvlRlMY+5cwGrICjje+jWaYzJW4JMu59v4g1
BdUThjX4u5YYPBzIFgR0oGohjyYeSzbllHT2McKbYpBE+ugzm40Qj83f3WVkuNWR
XVoKQhaxwDoHqSBLcQLiOZ7QNvdeRh2SwNo5XXyyLtF/YmSjzzZ1lJDYlwDXAxAj
xlJi9Y7kcP+GWmcIA3uzsJGR56asNGbH2lsI0/ST8cEHMV6wShQS7NghUYyu74HW
o5hSnkpNcF0r4TAfHWsjUZ2AdJVTIqwpPFdcuL+N32RBxRC5vJAdeGqiW0+RGl++
Q4mkWW4+3lnpiU57dSe6YakAhK0lBC2j5VQ/31iaKzmdejAcr+IrL8Wny4aibw4p
tHTCaY+nxrdG3X7D9N2svlPunCCKzCOKVxMwqDJc1+YFafO/zqnfEEa38ajXvIMQ
I1GkIOu9/XZIO9MYxa2bmYPFRZvxGcylabsDa+aN218620w1jnihphbRv96IGYXP
6LZ0TIX5RNnBdJS+cpWSvQsdDRgKR4E0EAHxwE9ypjy7T4zug6Yx12t9MZbC/4o9
JO3a2lQu+GilPgKPY09oPvXHnZZnXDNe0iqOWdeXkEzzYGeVEi2p+Ow+GTAX3MTZ
a0Rq6Zb3FSVdyPIaeBS95GZmhCvBXjJxzHrxRczLLs93AFsYLaek7Eo+AAA1EEzW
HqtviL2jDGoD/y5UQ3mnctIIX4IaRkU+VNnFmoWsUgYoDI5dyQMKPKRZNildNQ6q
Qx7CLcUguQtQZ9DtSjluHOZYEiJavzwTrto87L1LYfVHUDD7dq6bDChrXV6ZgPFg
cNfoPikPLMfcGj20aJCdJMCtInvHtiQVTXHBlCaSbys30JnHpyyyjyuASml1+AYn
TPOgatUKVRafp0ikKNdyyQ01J8hkfcov7bEtHVgIAB8zhUsD4Mac3YBA4tl5u9Ku
lJA/Ieaf4XnvlWEompccOGUgSNGCUQ+XZJkYGZYdpyNTe8zeidNvvWYKWRrTkCRV
eF1FGPaub4qNmUpF6dQqS2SLU+SWQOo/ZDcC5FeC3JzkpAOVAqniKXefavPqQvws
1Q9W6eC+Epm5bOC8VKp2TmlDaZJpSwU1NX1SiMqQJXxVzyKolNtb7jVH9fESyZ3x
lMM7emTH68jPy34Lg2QP5XkG1hZFXp1j+hXzwNGwBgyZBHAdyGatpcJgc+tYa46o
hNzuHPP4w9RyX7KFa8H84DNH/WHXc6+YE+QukVOTRkBhKF/QcIyOJnyibY1FRFjK
PgLt0pXxFOpKqsKR2gun7exYQosNXPzth4rBKrs8p9q9Z8TQyhNalnr6DFhtuis+
Kj1To5W2UcIvezMz8Et56zvbjKfIsj+LGb5bVtPJz7baflQrcxt4DkvRCVWpDdBS
Yg3IctG3Jwq84uLaMFaUYEhmQnPh/uz4qTN1ZZOGDhVOwa7flQ+1emzk8SdQUAyA
ZvYg1NRbnWyFOcFcsZouNepInQbDljxQ3bElyCddcdBk9JOidMu/WlkyXX9wbs5e
VcYZ/kFCUK/JdEyUsr39JQX2PYr+sp/wKtIQGIomtElILZz2nXPzr0K2LIDts4Ku
NBC7qnVv2W9wh+SvUsRhs09NNBAHMDpRwk6SbSe8G1nUVOhfZjUNkVApjDzrL+Ft
XE12NV3NukAxhJu9CZ8i82KxZjL9TDiVMsWwZFgm6V7Ax/fcUCNUY8+E7pUyE8hO
7n4z3/6lxOul6M64uKIWeOtf3rXGVcyZ7kyziTm3CfPe7SqgsFcmCqlv53UcyQ2S
mKssz/jBIcy+n/2tavF0J15PhAtnRTT4uGKLnW0HX8ZtwML9n+O4LjnaValVEPcE
10Xs1uavK6YvTiljyvscKABqXiwVhiy5Ei7IMw/+e5Np9N9e+JaDRaVD0lIgChtE
c+WRLs8li6RQcEVpTgaKJWKw7MdIy0z8ryIkaSlSDCPgOn8nzPRjEw1Vsx3yy7Ra
L05sQqvW0atfBTWLTtkzXFQwN+1TS7zgc8rLdSxPx+lfP0jbaRbylQQtSdu6Zoah
0tPQs53eeQii9a9d/7qUgSrl3AHiTbadLfTYQGeJwGCCpkfRTQoWMWoGX+6fg3uM
cInIHGdKahnOU3S1ogjBMH2xr9rnOGAqlN5+L+j/Ay43D/SO5TDFzsnENkwmjjtq
OW+eG7DBgsR+927G00IrHbD2cmX3ddljVH+633CePOyb1PrsoHFV9GGRhLAhrpJF
5riIg7+fCBPh63Jt6vv5mkzeopDzMjtUDAcL1WLxE5usmdCqz28tpO6oiA/Fg6GC
StKWz8BZ1C//rILsDTzRfF4NflPH1QkQP+r4pm+M2j5FdzGZ0E7q+AleIthKoHuj
YVI0nROUE/iawE8SMgUFSQG6SLRaBwfHjtlr2dkr9o84281QveqrB0AWmlnNQl/z
eX86wJtzsMPjYZtiWb7vQC+fQcdHZGjt8Dy6dZcblbL0ZC8KVOrn+ZeuPUc9N85P
qvqXdcr+ToMN+/RrdYj1aZm0rF+LJd5Ag8DohqtL9H1hAHPtb6dVTAhLxQwRxJwx
P5GxY6UZ+/mhoKO88XKeHCVOGkQfg+xLtR8Iz4pE4/p0yKfeKH3f7W6nWQm4a1su
CnmQZjVU4aMD0cPDFL6FH8KgGZVIgS5ZE1mhHqAhdu1No6h7nBJwKsesSLUH2it0
KCy1ACWQFtDFmqzMHWy8rRKv6RfiHJHlBpbU5iCdB2oMU70rOsPrvVf060WDB3Ro
kdPWNmcPCWLjyUtSr0m9u/n8P/+RLvtxHuUjV57bTofp8aKxXmW8ggiIE1rbWYqJ
+U5jZMJRs0mVqlE/lK8GasqX35PVvy6Jgra/FzO/P6VtOflgTuHpUpThZ7ZUqFmO
6qFKOMLeKxGWgd7JBqP/5tG7ZYlmzOm2VtDgKOwSbzW3P2W5LnjYWeEWC9JvuxAc
PeSshRQYnvyvamlfNEboZZSso23WetxAlrd3xLWi/fY+N0YJ/+vHmleJZT5t64GE
H6G9L76yaIw9HJ3MPmJJRF2YTESJPOK3oDhj/vy7JMnaFAxXeN3QGWufeP59aCCA
pq0kO/33XY0snoYz8LYIZHAdWsyq6ZQyL70zjPqR8atVA/WtuJww7XFhLHVjGtWk
7BLtlb+VDU+iPrMuWD2ddg7oy6PVmFM53d/wAw3mh1DSX8D395iEQLiJmC5QdPDy
JAQURi6fTc6OlYRag/gO5sswOzrMMInavjvMjM3HKZ5M+M1hBMrHauQLfgYUl3fY
Vu6IsGUEdSiQc61u9aKscBoZ752jpZhZCp+AFqQSiraBXJVpjPG0wXhZyiR7/mOa
rSbku8qODI7+F+332Vo1Mj4s7Uh4h5VhOrM17yB2U5wrqMlqF0jSO3zhx5OjdA/U
Ve8PG7UHai2CurKXtI+yhHIPTDI+I7wqeK6d0lo4ARwiQLxLgpG9m78rKY142qiY
nQQSaQaTYwL4tmGfiQ/gjWQUHpL0bdOsKQHAO79iIqGJPj3Kyp7HQ/XhOyiaCepA
7l2czTun3J5XD5RQfEwg/Wh6/Upg9h6TC3Ig6cBK4i60l29aVnGxsbRh/wWNk3R8
qAQu9L6X4VP/kptgbvS3nqftTykq7txXvzMFr5VScwYNIr87R7wzmBm7A974q/1j
DNWveeozUCzPS+fteqtuOBDmJCZSFdNKi+1mpcfEYm9DZwMhaMLdkPzZw4UyQs2K
E+vtrTO+el3lQ9emFCHeXOmwrQ8tVAxPDpTol5+h/WyvUT5q9OIuS4hh0YjwO6qD
uCSsZtt/cR5ZEQXZ/3goWoTenWf2+jyZezUp9EaZzbJRK6kCC8RRL9VC5AMTGA/W
vfvXrpg09PrQy4SQlw2c3dRio4LRaWQivrlxdds5NVIfjwR8wmXrA5Cpf8/z+Lon
DvyyAp8sC/a+awBS0kLTOPluWElHaniqwLCL0xfnnghqp/eI23ioWYoMDv8m/viy
6WeggY8SzyHiTp5wWGeVOuPo5zNut8SlwefcLqs5iqBvEUHPjkwcy6JrtGmb8nsO
IYZ3sC6/vNvjJxlXx9vyXbKfyFFDUfmISLBGcri0kYNoXeSEleGlW++5SLApgcN9
Qqe1UP8eqpbxyDxx0SqyOcXEfH/dYrC0/9cCYIQaPhHZ9RjU3xjXRffXD/yco6sS
i4dZFff3vYowPY5PmgsyjRcaFWiaKMW5xJqjXGuFDIfK0GrA/90yZ/+t5J9aYhC4
ru6L/MprI0XpD2shEwFooRU5GH0bViqD+84LAtsrGdzrHI9J/YcceI+Eor1D3Vn+
gdgWYNTBDM+DxSoQCT8FT3nvh2JJAZQx4G/7v5jiW1BLInYbvlXQbWZpYrQbK3qG
wD3tYLPldkSAl9mECsjbSHlj/1p1AnOq+MpoOE4YZG0ndYjunsPdJw2sqvCvgXMZ
0G8AqMONZ/jbKG7yVYxOG/EZM80iAEiwF40pgwaoWN5Eb03pDmAg0LYwWl4xxEs0
fD2MBbhk3KlJ6gyETQKzLH6X+Y88g/UNhNiTHH6vpYdXVfrzdw93JLrCdZaWeOjm
GaQ4sjEoulltr6NCgoNeqX2KbMSqZUsOhbpCpE28w1r5Ewr4qBFisAOkuRekOK9y
PrGW2mrct9Rl2Uk80Y2kwG3Hdl+jilsFOtBZlRSVRywZmPjVlsJRVaJb2u1NyAJo
H6pUGWgv7kwY1pgB7xY1b39BBLzmzMZHYm3Ew3Xvh+E8LP/I6EdepaKtwfZmKiAG
gK+pkk7BJB4wbnUWDntLtuPAjYt9jsoPotqpA8ngZTNq/k1dUT651MryrpQg4Lk6
BWZDQTxXB4FtAnGHj99kTtzQXfxWu1uMBgfMTw+XL0RK9B35R3W+Y4q1XQjJXYZL
w32t7IWEodtGZHQss7eCqZ0REwaouodpn4A0fKjsNcRy/ZR4/YFlyFZ8iCivy/Il
UNXiOq1z5AjmleY7L9iJyXPnlaetYOiv48UuF+xccCAL9hV8ZSqB2AJ1SFM5b3WQ
X1mxBnQZMSJW9HvYC/s7JFMs7zGGOf6SDIig599cgqH7LYhgrilH5GmLolUsKOcm
+37YxIDECMyPacgmdwXywzrLUzklH3bUnNeoGXPBsvgg3IqzxdGE6i0nFEYcSen6
zfSUXsPubpfMC8Z3EClZqyhOpP4R05LqxiVUAq45KkFd9rumo0gPuJEREnw9wZ84
moKeKsBIA+2YrIlDX4kSKNc/R57ogttByG1iCgCptvapSoN2ozH9FcGZJa6jft7C
UpAQqRpDK1sjHYsH6jR8VehTEKvfQZQ044JvKN82wOFgMt843tKKetmU4Ov8fAF/
KfSGDonLuDVh3jpyzBlYMC4wzgVQk+OAai7+9LApgz/2917N6lb1NFcnONWPk8xM
aquN3I/DIkkI0UunLo+iF9EOKk7QxTY/Zxx/0fEa9CoSWFll8p1a4bPLKsbjbEtA
hAELU3VpkA337OuUZyICh+t1rH09Ez9S6BPUcSDWhaFHOWv2A1XNMHxusa7zFYm3
oPxeZoF0EZ7E4682sM6khzfyS4CEBSqiv8lcD8l85+8I0S/PKvkwy1Adn/IV4P49
2XBIW3KQAs7AmU1SuKwXmlzxpmmglufhYPyP+3PcWcstubM3ypVFgSGC4G/Uq4wS
6DXMH9726Lmm9U+sppZSKWlfd0saufh6gtGKlzOQFnWBoOiH+S2aLcBvd2VRzxQl
y3okoxUtgSxNP0waQfPjC8cne24vNYHEp7fsB4EKLpf21tyWKNP67M5jgvoCx9XP
iihjJdTF9bHrbITEBLHxOFDlRTRyjObmmKNaiavLleQLKGEYzXF5fnbNFALXrIti
YqGB8/pOiZC1wPfeFsrYztKH1aoZDR6DIeUN4/XhCVftNTeNgtz2VR3Tk81mFp5G
9U88VCsy06yxozEPF6OU3WmRmjbziC7KkJh2aL9HxJa/wPvHB4eVgmXWXz7XNoS2
Et24iS+giSqvS75GK5hrK+eJIaWbdcfMsYybDlhdkE8jRsC80dWKc7EZpxd+A98W
Xut0mX9Ryn3X8ZMjxxSgAq3UucUJed8W110lbo65XOaKMftz/tDKtWHa1Ae6A+Wq
qBViO+CiTDNJM+pTRoqy3hTKryIAFdwkwh/uRvGqFY6hIcydsSQjne6ijia9MH37
IBGEzvvUx4uSqM27Wm1LdHxaI/1kEicj135ArMH0Rodn5F01va4cxTIY1Ya00YkP
R6Em8qfGV3ReApEgLbSA1jGfy9NomT6bJhWmcMFUdR1cG8l89vWZEgzEHhz3ITwc
KYkvH5LN+BHv3EM2tSNgR4I0OmljSLGhfSdZruD5NAigxHKSIOg7Li/pTwmW73WF
cn1U04Vz8iG+hatZC1wN6V5aTtcNg/XjwFrtTdc7AQTfwz4rt9yY/TsHtae65Iqz
tUgoJ8v3+5MHDMiddasBhz+8G5+8r3SPJcUHGZuDX1nFsFfSE8s7ftUgFUPuwfw7
1qs8CImPuv7NBWeDxh99aEf/nc6T9h+KAk2rRJdjDtygHrGxOOer5NxQv/cC3NJo
MjhCEycm927eWm+iaCkaY7UkY+FI7zJI1S9S3Rvu5+CAeCwP9nhqGvE7XiYmlc8U
uHiEKcfnSOfXdqBwgbrkwltt7EHisJoZe0i7MZ0D0MuNk62J1TUMOBzhML7ot+OZ
iwIhFRwbEaJTR8FLcuXUaWiOd5ttsGYWRMDzwvpgL+lXPDY93OfP6lefadWK/JAa
i12qsNYfTrmkmPte8FMBWR492uAqnP9DC2HRY52D5zrQBR5JNtzq/7ZpOlgMJWq+
N9fJ4aCUfSHaXWE7xERzzbr8/VH1STJQlgxGor1jCEhE7GzVHu6Xd3VT+3/mzYFe
Wz8uht+JOO7GwqHbZG/F0IgMs/lkHSBZTkGWMlzE9vo2rrw+Srg6LhkJaet8/CEL
Y5mP/Rif3a80IdVTLTuQhZ0RPa90GkFxs66ev1dlJhpqpa2GNFnd8XP1vvyQrVQO
xVFnq3HzCedItIeA83atDjtDgAtwza32F4rrkz+YEH2LdTWBaNUY2BRK2mT0wGI+
VJO0OIEUv8i5CqhP3YSBgYL7b7gy0aldxnfkmjZq38hhcFoWR/afjDas+1ayyIcy
xWrNddnbk+a/NiqFQR8idBME2bz4IzV462F5Sm0CUI+xtPfzHufG5oweYrMCG2pF
sM7RlSSnZVfiCZ4cIX2KIuttcU/Et/ab0pa0PHxAfszZmKDkV443D9JEN1HxXaCh
puLqI57wdh/ceXlW/wqn/63CKYGeEFPXwFT2h1pD4IFkhcg0njpS9j0wjBOAG6h8
9QoK5tO34u6UOxJO8uJsRKXrUFdqVxVjR2Jii97wr4D0dVLsnwEKtQ2N+FrMinwH
jap5LLffIJDJHxpXCMVLtMHdyHKaklB+at6Vxsqo0v2LxrsYkk7/g16U2/+YSRds
nebdOCJs419bZ9LX5OjuhdJbotT92aj6/PUnvIrYRM4zHB6K7H4p9C34vKGb3c1v
6lJUjRKLElZj70jbtRtzM6Wh7vhujDw069a4LApbaWh27bQ0zskSGlD972EuRC+f
8X3bg0Ihp7mvz8GrkICy3WdSz5geoNyT15x7kUyb3zLqqtzLyZXqo+5EOkQfD4Re
DUBKgS6N50ZUEDji5jscl1MCvpCD9MgktiXJNsQzYuW/CN0vx+FMqa7xegUUVuar
Nx81eSq0qdgJ7nyt+Ghv2qYhYCEDwvjxt21GFuQeR3h0SI3TR/EH0BxS63JjVvNR
sQXuOYJQ44r1AozOSGCOq2d2plrW/ftsKgdKlR1X0s4yfDs/l30/LR0ojlYbBPwJ
aNXXmVXUialRYH1QImvVngGU3wPYgXArsfGaEXqlhtAHanWbcfK68ZZcTi2xPjdB
+xo6r4gCJwmmsXCkV5nVsOw2qrIFF2RXkdYoD9Zwp8tjRbF3eYYO0m+mf1gkTZDS
tWsVI/w0+KoTx0EnhxY3vNCiucD0DLsNiCsEhRU7asm5/OIYtjQ62RFLNyedu0s2
mAoWUQpenwu+bHJsrUIs0Rv42qVNyQ3K0Bd9iKOLgLzhXlbC/oEnVQoVaPjArOK5
wR7yeWMhzGwO2KyJ9M51c9eTIaZNouoofopmjZD5B7SCl60RE/s5odOOIKsgkpfn
k/g4F/2D4xyzmAoT2AYKf3v/R/8SVihMZGVREEa7ag/bZlOXougB//3hbAbrXVgz
n638Kaw9tPTGgEs1WYWh+98lYGXDi7eNOD/zOEpZ+OPDfeNUp/GJo3xLPUBNZd2I
4s94+Og21gULcKb+c9xGTRtFzCDNV+wxmZaloA2F9ebG67UyHYcXqziYeJDCHAQs
WSYbTMxtsVGpfrlsojiWyQZQfQ9LFs4etkG0txidkpfya1AxiPSe5+owG/6qWQT+
sYmtbd/4RLnbi0/RxcW2OLBrqpNm5VxNYinwqQMM7lw/JPnQhgRA/YM7rA8M4u1Z
vg9pBBBca7KAIrbqGUaze+afiGmT+BKqzQrX/rsrpTTzImEhZ6MJP/dHc8BuIRLU
VxbVYb9I/QCv5f1tin3OR1RYRQ43O446iDWK0jh4w6NESVuQXBHWnjNzB+xb4gnK
tW3oTkKEq9ytora1jIHMTHt9B0Vs0g+6x2BSZ2nWqoB2n9PPrIY9iKowBxlRqJff
Zu/+Hei+D/AQbf6FE8fFqYHWd+zTmm8uNl7Q+S6wLcqCFSZ4NpBs3T2DOJMbH5al
KYZ9jdF6v2LIRhZmEwugrRKqucPF0hJXfsxqUXrdddmG9wiviMz227F7bsfEGIF4
lik5YmTvD4U7QfYUdmB4/7YoPVojRaHg3iyhtnxByWLaQi0mMQaGGiP5w3OYPE4f
2Qz/tzypRQ+MbXN0QwvljpQpbvSXNqUDoqnxkSnMq7JA6XL3l2OAhBGMcVg3GUYC
Ok6pSUvGUGUPoORi5IpyhP9dELlDHlj+IP0rBPco4tz6gcp14AOojMA4vMJAr2Cj
1A/Bjo5UYbHae7BOks1QIWfiicgjSsrB1wR0mX3Z/QDnYfrw6k8pdezCi6TJiWSM
Tcwq5fgWBcd7WXcKWn53xisozEIqHdcnVw412wl4GmsTEeJdpi56wp3FbsnJG7bI
nTPiSA6c543Kl0r2XURo6gdrqSFzQXNWghnDt74aUU/bcJLFMpR9lvynShP9+6Xc
18vmblRYO+4GsJTpdmOQ145Dy2Kjbzo+c/6ABuohki4QvgD+7mNRcMHSpUGsw8VJ
koYez9t/OByMGDo2OOi+B06WJcyK5xc64aZ5MeccfCIqeb5T+dtYJs9pTqv7c71O
NoIyED0iZcNF5LmffkrA4gjv8d8heA3HcPoAvt5sYHsKNcLkDb3IbQJoznsU2fIc
B3kSO42HxBeH8Leo2B00fVvRtVgE/OhlbMMAEZFCR0Tcqis4vImrL3BX820bERs7
LYAz9h8snY34dlhMPF3T8gyBE4Pm+P7qP+rFSKrR2981PmvceCAdLAUxRGD6/S0D
0+FFg+eX4djGETZ9IBN33yqbcQBcYhhQpar29IloWKSv6YgUNcYnZNsZrk2HL3q2
57i3geCuIK3pCPB5dXT6LdDfmpsEz8FyBgTC/jil2uNwpVrokluVJ53EpTEmfDI6
8oLYO9Vxyz9l7KnE57ZaBESa4rR+qs/gXIf3YICU+3bUvZ6INrNMAm8VbYU584nY
EsbWJrYRSmiqknf7Pq6fkDViOWtxHPg33GGp6DHMEAqdd/C+o1juYiPyPQks5NGc
IrgW4/2xvMchdoA6IJ9/gevVmGwcC2sRGtdU2m0QfAyoHycB1R3BrCoLP0aGlM2Q
3LwLKVznkIs++UWNfrZVzPoG6hDTglkMnt25NikILhpLw5uTn+GyYyKSF/OahtUe
44rF80j3QeyejK/yuJBU8w0Ulqzpp0yts7EJILdzzZDeWGS4KuMkRP+8ALRVA0EM
hxMtWNPKzmiKIFlkdFHWkMZrLfukaUVmaCSqyLClaRKbonMihOx491n0fQuMi/9X
rpAqFwsqpFbGMmZKGvxMYybxJ0HsPnbDFaMIUdd1Ep3wnih2UKIzrAkCPfgC7qu4
nxqvIud8HUJq8VlGWejBFdf8aiRGLIgZDRC4qLrafP6MnRj/ftToz3b4csWl9DLa
Q8ZVI+9zAAQTQIJfrp3cNHGYeJdZk4C55FJ3ZSFmRStHnZzOQUeho9CXSUJDSY+u
CCosJ9DtwN1DZLnP87HSryqqSONpzEGBki3lGnsL/pdt7G6jZl7ysag8FTPybBbG
yjb5rcgM55Qh4t6U85R2QZ9NWzRtlLtY/shJmaOLpwJJniMfzsJxUJCZRZIA5Rxa
U5u/vFcnFmoLGL7e14vjmJZv9dhOXidf2zUI6r32KqnqV4+fsxUIQ3X2mUJMT/f+
95k/3+3scdm9bAcnD4BS1nd2R5JY7pw1eZkBKcr64zfYoPW9PL7aFCdnbiDXxbZC
UedzgzO/ooe07fvme4ITBTFmMFNKOknaEJVwyPUR0phbLg98G0tf9cjGt/uEyhNk
V+n5h/Yz22Ppn7wOnv4w+G++tedUFkWuja6cB0bXgglvyOwWzLLeLvmIJEfY7MqZ
EUFl8SCYrsfAHos4ac1KPjG0lv7z67xme//qYN7qni1d8Bxmjyt7w7+Dpez1fIKI
Pu/b2YFdfyVuKSjvQDvCsJceTOrk3ZNSCnGWFiXs63srmESUah3O/PF/M57hBZZn
9DBVsOEMr1+BNP5g/u8y3CF3ATsXiTKxST+/f8MKt/pfqBMizoFyhkp77bp0muvu
jtUrRpj12wiKh5ej/sTrqoPMadjPGkCVaqcLY6Fns2Q081g6PWCPP2J3AsuZU8zZ
aI03tbVsBQDjckgg+RjGOYxZuZNAo8Utz1X8NSgsYD3SXoD89TOZhfkDicA6RPvV
c9Cguu7/MSylSnN21g8p4X7zLVXg3/3zDbnfeZVbKsuGDDy10hxlFR3TGH1nJ5xM
4NWlu84PApCFZGiKXmzcn//iQLirbMWDCN881PeVI6a8MEuMS8dMqPzAueZ9wIBJ
5lQQaJl75Is+8CB9c7EG+UxNxTu6eElQBIUkn2FzvloygLe5+otMy2VcP+j7xEaT
Pk/1M0P9oDjYjjF+ARKlBXfm4wZbqghm4Z+sRqOzp+zzhRTLRUiemUa/0ZUW00gc
OGi8HNKeXDIdKnTN1sUYq71cxz9hhqNN4M0Uz0hgQMtnuFMROz4IdtpoV60s5LxN
EA7cb39kkoQ6Ua8LLykDNmeuP5nWgdpFMvqfOXW4CEu6Cly87xJLgbHzGoL1ny8k
FI7w63Hl0O5cKQZH3c+gCEK7hT74hVX0m98ao2oU1ric7kj6S6dVoHBVMqvIx28X
egxM9VRCW80OHBC2u5hNtU6hX1jdcPT1SsaUgbW0VnvRP09BxpQL1Sn1DZWSeQEB
O+tqZB9TIvtIlpHPmKox8CsRp75Mp+9GxzTgSUFtlylL4QUmemOnx/e5rTzYuDiw
FyoEsnnkpq/cDaQRoZRUNyyoALgX6UxtdgVWliYNDNgg8f6hygPG0+xogojtOnRX
h+uBumrLGQfmkQiGsmdbnGTh6D4+BTsVnfbZx+UqF7BvdJgUVz0WcBIoclQvodJo
wvtF7dENuzmziu8vNKNrhKIDuKKEPCP8ktE6YzCRBDb28CsRqNpPW3sYyDy1Fzx0
I9aP8IlObvPBA76m4DDN1uTS8f66I125gMgr6y5BJEr/zpif7oxoSsSutvNrozAU
QVEcid/K5KVBMiaB5HwnbyCged+/56afZWxJQyam7HPV+EWZbX8heQ4LHPFmah8N
m/3wVSpnknA+s7auZ1KEDvxbiFB4iKLmQXAHI6dyQCaDGCqXhU8QmYX7ylFny94I
NanD7YU7C/LaeEakG4NjRNtMzXL1iG1BTB87WB3DlVFNjqwsPP7u80h20GfDjQKW
DlLnArPjCpH4xx5Y4v7c0gPXYWRrXT1zEmtVpktVvgNrxAlV0A/CI1YBh0QDJV5t
fTshrKww0+PReDHFQFOJ/AU2JLrH6kUJKJKi8zCs9hj8tf2zeYpL4BwxDHXHrTG3
9cNBU8uVr9z4WZDxPrTYJCMTezghGMEjcTq+6d/UB9LVv+qNFLhe+litPO+QWdPO
DA3LIjb4usLO5xw+nfNqXZ1/jNoTOtexTJIb4Y25XwZiVxJmhzuzT+dEZEKJtMBw
dgoGpcYdlv8Eou2TJqwXqdPYGH+rfOCUE8vUlWhk+PFaYuRNlKbkyGgnJfB4n3SY
0H19ejXzjyQdu6CWVm3gpGCSxDn3xzleBesJfXuxcOCGVlqHNIxeX+X1QtENSgy1
txJUv0i/T3qyw3nV15R47h8+n4Vb1AQWewtp5jLamLi2XKdbHB6lQIjrnFwpJpE2
JmHL5vhxJIz/nmKyAy6YxQ0Q3pTqRJ1T7RA/M7CBQPVL50mD6AhtZ2oSMmdC7vBO
VcaJeSIdVxumxxTV80yUloXLXmLfs5L3Q287rBqUKShCQrhimXyDZd6Y96K7ygxg
UfjWVJzIcrg7IALogdK116JuFxf4hJQ7JjU41v4RFiWtbRvyoTy9HO447RUAlZni
6F7KzCVWn0vQgB9BxjT2eNn7lb1Wt4Lh8uJp3RxrgUi7vIvjMXbMlNFc8PyGyRIu
9CAzUvPeghnTG/t7HofQ0uzN6NF+5L39lQKwPeZZ4c4W3sdI5HPBuLnDFQiPSE45
LCF6r1MAWpyJV+fczW1Lylyt8MKd3kxHxdFAzm4I6Fk+v/HY3/wR3q1n/J2CKnI6
Un1H70gdLfcsmE7ED6hj8j//28K1rHVQe9Cqd65q84u2ryKHHBrRRVrQQ15ps/nB
cGmTmMCrSL/QSEMS6ltEyN7EcP0HqfMhJ2QOJKN2TgQylnqFSgj/FYCcu1Ut/DrD
5d3HtLJZOIDnP/ZOHUNELWkH03M1CoGE+imJIAGGIVzjSRfhd1WJKczW2QFVOsBB
c8x3TTTTfMmoelhuk40qH0iWKCiW6TREtHxunUYddnD2cOxqwDfyDnEzh0oAIjHU
K5nJ6+KQEz6BnUsXmoxPTEwclFZgLsqlh9G75aHHaETzyKjP2g0mC+4+qgN27xJg
y863DcslMY1DO1gWu9LTeKZ3B+dw+Pu9tlgsmxguQnOGQ9axY+S7tKs/GoNZqyBR
4wkgOmMRpqEFWQFcauLJstSaknTTkXyqCmynNtGy2eRfZfwrvrnoOT9Iu6Xu8/Sg
FbNfkVihVfdyjHXXY26nirLjoN3FFLHCY21jLi7a1IinVoybd9f1CzeFWjOoiGbo
f+xOUiLuuXKKW7F7nBHVYmW4y7QpOKoVH8005R4Eu/OcE/gYQDhs90D8zqawNYoU
NFFQ2p6jOBbbgVf0oBT1iLKCeJAWSyJ9JL+qI98YTcCMCHQvDIk5XM+N157jeVPX
+KaxhOAghVPDCeZ7CB63oZnU0t/jt2dBJnsKgggJ6jXfzaECP5tLpf0k0S+iGXAD
sBAx6lNZNHVS80Zv2vEUMfc8XkQPZSs+DztSPtAY/VFSpv0CVzmznpWrq2Zfv6S+
zMk6ugo+PTACu8ElqOamEmysRFVvgUIDcionKBLAFaAfKSm0a8fjZIMQENOgMSlE
7ZYTzUukzYv6NxVPO6imR8Ky5ILXlhzyqn+0efySmFY2pYhmtyO4USt7Y39ciXw5
BYojTGz8rwyLucswphCY4mW41d+U6r+51OFu+A3zSRRDbdrig5MTGYW28Ydd4POj
+Ll3L7iqul0KcHKF0otYNvZN6aB7je1/egZWU7MUYOlaSO4UFllrYmAdmbYNyb7s
8gAmkVb0y+xd0h/njRYWzRBrecsamcN186Af2ZGtXn9wahzSSj+txRd7pyaRGLWC
HBH7dkn064O9aUBhs1LRw79/IgjIQhNNXpzsla4HoTMr269m/48sOg5glw3zev5s
kEWO19nMhTNHPoQcTCuFgU7y5ofMz0L8fIEZ50V/GtRLJfYgLcnrf3vBQ3Ivb0At
CQBreVtel/ukUcDldBr39a7kf8ba05Z7f2jaLd5PX+pPCZ41LwFFjod5kU6LOuL/
vJamOuJY4yDaAuvT7ENelKwUbXkhSk60JvwGQKLNpmag4emP/KXUGvJDhNb6ep9d
XEAq+Kgd4IsfRRp7rgL6TafUs/8yw0gSiNjax0KPlEU8rXiz9Jq6Crpzdz0k3sY2
5bYKHJMR6Q2KDd1guHu/dxY+MCNI1aE6QupY32lWtfKG1XvsnVQJf3pbra/ocf45
xa07NHu77SzqNBfsHAelOv1ROg2uXBkrRVR4XAWgdGOzE5jsxi7akICI9iM2xRw+
qQfTUd+GYmI2Mekn0F7Vm/ZmkcLbpdUQQIe1/D+ELZ/c5BRHyMPMSgBFHUkeYbmz
YbhcTo34JYR7sl4GNnPxwAdmvqrfSKpNueNA/0uO0Mk6S4Vz9HX9pF3Wu8wFr4+B
dQaMtZgacZdCI+knQmj0kcg0xC4+Z3/JQZsSPUM7t4Ge0Wlghf4jwH9EAOAEOIKz
6COAQuGNClyQGpdYQ+lD8iy7TAwS7RwhJYOCrvesX+eY5eKG6CrJ2ts41PjPZBIV
YhacwG9uqXoNVOZaXk7JSeXU1tsD9fTgNcEv+X2CUh6EFyJ8lRDMixs5p6Y48ChY
tg/4KU55VrPYXVJh14FnX41nPIML0Exke+s1fWAWHiv0cOQ8Z5tcKyeRnCmDGkGZ
8Z5OFZyAbkq2GW0XXRzo9q/RKCUYTpks2A81DiRMAGxcUlwfmEDFYHwHNEG8h8zD
oWefFA6NEZMoyJvl+snDBLovWMom2hwuK1iI8nBJc56ppSVln8hrtHNjUbb55qDf
vunF5LmlWlVfs18qUElr9OwYQwhjOwob8xr95Y1LNT3G4IQOR7F75TaOc50ZdxHH
OSQ7FS7xjycXnvJUKAIM/jxP7NMQKDJLKkT0pITvS12J4Jj/+w+AYhwGEdNyMYca
lIjb5DT4e8zxtmGPxp86dt9h1TXWy/cbRx41H1qocGgJETTEZJmHNmY/mrRN2gEJ
lpdZPCJ4/oi49mTWVrYxt/gcdUE/q8a0SVjI/CJuBEltHN8KjF1OS/AYM5l/BGov
RtHIby0pANGbLJTl92sUTpAyhLuhFiE0ul2uP+t3hdg/TB1i+7w7CnX89Bf1ak2Q
wZ8kqDb6OAIu4TlOzJlV5CVF3NKVBFS4aXN28PfIGA7PTys4AL4qWLRJj4RlciSk
25qZXwekAiLyo5Xunh6KrKt03Zjnz1YybZAtv1lNJ3b0CV987JjjWRKuE5XKU2Ef
2lpzteZCGKoLcyWCqcc0htjXNIPLA85i5ohn8QUlKu2QV9oQ306qoQ6dsEAEnGie
ot7uVxbtNRoNlzqLleXwrsri8D3/D9RL22H1xG/PfIpckaYNc1v28ZiL/zZGo3Xm
1TX+ZlPSJ26A7BsRYPHu/bp3RtP0d1UMxH74sG7IqC3P2BN1XccNyrdbnJY7WnDN
rDpdQoHEFnPQNGi+MyDA760A8WINhBohqBqBDeH11EXmFF65XV+jgvfrw1FwQ+Iw
Ptn6BAdOuW+tIldCTvZT8ZYjaNaNvhvMnhHZKtFTcCOv/ln3X8Mt07MOMRO5dmt5
RBa0YBHKA9cPrXgqIYnCoZTNIOEXe7S7PXArrUcWTVk7GSbAMEzWhp0GOX1F+LSe
ZhVNM2UukrMFHKfb+MuXNBuDD88fjSCaL/dmAiC0FjxGVnYKs+rBJkINPju0L2Yu
iPpXV9nLAh/vrbQ31+K4CVN9ititVNTt0wHLBSwjsJnlJUgg+731bytWfP9OsfGe
nkQLqsAQOq51DHEwao3qU06N8zVNMxBfA97HxfZb6UZP3lLf8eGUIdqrxzRqvOaI
+eoVJBROxXRT90/IJiWXjNNaf09QE6NpYeFo9pewar7fy519zcZPuAL2NNZZ8MTy
LgEziSZmHTnI1YEtCXXoslqC6gbeHPwgDiYuGdMQY5JhxggiG5WEg9SMIt7KUKEq
H+FeBM5VQKrOjoeQMFmGdEDbroUpUdbIF8tTgM747kbYvnUWRqBqGpJ4wzJ5x6jh
IqC5F0cxdo/mNUcmn12mQ5UK3siHh5t+WJVHjWyfzRhMZxE7qBcGf/Q5WzMEf6eh
yEBORe3sZMXNTdAGHvCs3M29RjGMgmG7Jbf1qX2nYoMPFvAs+V3Yh3nV8NhvpgsY
e/NlTO5K9WbNpKtQ7B3Lws87iQa7U+PvF/4mhIVvLuZmgVa+tnG3JWdBTIFnuwNv
gG0htiAXVtWBpOksLvIg4RNSJePjanSNY9mysVyi/hETV21eIbhS8yEtWLGXPs7Z
UL/xwgmDaEPqkIuIoE2yx4XQjMgpVjiy49yAUbSVmzlyeBpNzCMh6NAgaA4VCA8g
isgMT7buU+sqtZEWDth94A3veiagfgJ7d+iZAUJ8lCtJvusB7eluK1UnQksKhLSJ
ImjmDfgbntktxWL9OUirYaJAFGuAGAF7clriGpeAmdYIHhPTu+BOJc3EotB/fM78
XVE6D7me61FnrJ82PCt82OvcYeDwwFkjzS4Zg9C1wpbF3HM1CrvrU/+tzA2WPYKj
d7VLEqiGXY8USCso7iDmQhg0pmhqW9mqqRlivCJlppzTNB6odk2vbvt8wmMpb2vq
+7VwoGkgQY4IcJfHmGrOqZyKrs6HyhRGtawm0vjhl2UJfTzOLi58Oc+O7pGoyylR
vFcdQ0SRvtxMkCLBc2dpafYtDlEaqU+KT21wznWsBF7LCaOA5P3QTLrbA664FfJE
BWGcJdqFA4WpfDZmMNNB+klYert4SKcA+IyzVhzDhbApIOqoKAB2w7gbBV8R2SPl
k7G2G37LNvouTaMVfKu65HOqyllKd5I4hxIEbkjXPd1FQMqNzlVqEa2PAGII0AoE
z67XSOdU/rE8/c4IDnoQCKUctW87MiD/iK1cNSjpbH87imXDtMn+pbVpZQntEfMg
UjKVz6CSQhaELHMuIflKB2RakvowjSyf1pX5M8LiGgkbHOoMTIwNQxLmWH3BE0N9
pH7grB43oWcREhNDN+dDfzq856gJPi5DgL1QZ/xAKm0iheXUgGsQOZYOsElLeXcR
KKaZ8VwneImYqmKW88fLkjh8MxcA3EqUR5TNiI4YmoXDI6uUGwY1/4zKvqcoLIGi
/xGV2CfIZ9BryxzJc0db2s3Zr4VLW/aGCvjrp6qNh14qyUBOOmgaluCP5IVl+Fna
L4GSds1I4NITDAzp6LfchUjGDKqyuxjUC3hlvnF41Cg/Za+fpVqsrAOR8o9pmpvb
gJQJLt31CdMyycVBZ5ND7qMjlWwp3NcyuxUHhJHDg3jJ2mlD3fTJVxOemHPaen4N
OH2CZtCxttOvhFxs17TNbvP6FW8BLUyVKvl0Ev81KKgjTKQ/IQ/0Qa15ko+UiBMM
ZehupCsCp+7LAyTeHFZDLrkS9ON8+PS5uB3ixu3KmAZ1AMmkeXmJczNhPj4jWbiX
W71WrlzJknqyprQYA9D8R5E8MQJV90DsfGsmH8od/cENvI8s/BsfxG/C0goRRwNG
PYh9iXT2k4LnTkpRlMjYrYpW8h5UR6hwcXngFYPwSDfr5jPh0wbzCJH+Es1Rr0jl
slRj1ZSMfyScb86X7WvQy87w2RmHXl1BpAkybVqjgOQVSbgsZpu/sV5XO3U0JxNT
OrHTy99VWo/bo7C9Bcm14Ag4dFF9tQj4E7KQINwVJTNg9wrh2xxVQHmPUgJ6YJ8b
gr1qPycQRPH1v5MIqpQq3IfqzDg1wdTvu7JgANrNOtvccuXhS3YbTA4u8Ql7pSof
WbsNvpQj3FKQGZHksjoeeleUTFa3YPdSk5k3qqDNh3+mtAAOfe3tcwg9A0j5xA4a
dMeEDiFE7taVoXUj/jVG4naz51FhhP4iEiLHNrFkb2a7U+h1r/NwmWYJuSTU/qQM
5CuB1p42YdL6aV2+QJCddJ5LoThyJI10JZOHptg0RutU9LpLjRFjfhIJ3RcDSH2q
Yd6dGFMQUpAaGor1QsE3hVswdKm/HsCljUj8gfCSWE9Lgz7maxkx8kfxoHs13Rnf
CVyKwUFi6qlxxs2ta44gFn/0ZRO9SQpdnAdqvVUtNpskTkzwmFw9vB3dISEl8yyf
gbFktsQR61jrim0WpQ+p7EKk0hLF6q8WQmzp3rNcB/JKOiCeB1MUeqhUF6/0fYsZ
B6XeLJ4mknOFctfiC4SQ9x2IKvSLYCedEZ78ike8sesWj3YnUwuLUeqKiN2BiFgA
tXIhwp7LigorKgtCijBRV8ubG7cscnlesZhCjddtx8oBlvmfZ/OzsjqUZVaKGbYB
Ij5YetGAW7PMPw++33RDGjV4eK+9Evh9C3NNEs8rQSrTiEOe0LeYa5K1un11zEHD
hri2n3M5004ZlOI1BHvlpd5AHisrRHv4N3CmOluTfvFQ9MsxoKtCut70rpUr9b3q
uDWg67IczkEW59ymydshr7iQDl/BhKpW+j+2qrEmWs9xRaDnwlqnrMvF3V099Wx8
uuSPRSyhxd25LCbHP77RMlQwaBWbkeorvOqTdrTQgSzp/FDM7rxwoLcnLQAsA+GW
LSqBFKOGQh9ByfxkbEQG3Xer6Bxd7FLDRfrzCD/HLsc4Sx6YzVqDwVKcjnsvPhkU
c8dsXutKc84DTsCyOkjIp3HzgKLlVO6lP1vBtCG0xBuTZoEXcKCBOWOv4oFTmCJa
GizKqxcv0qVKVilsCTnEy0KviG/FHY8/dPPyXKNlDOjpUz4WlNjC6UxHhnZ+GEvN
BxO1JRkvPUhVKpMf60Ec4vyZYSavrydHAuNxMQ2FRkl01RWB0mKjQA8ny6NBS1AF
ieU0uqNwdFbIPjxkrI1BjKQ+507Psh87qrt0146U5qIsYR8zPNvsnD0gTLqPBNWK
M3vLkZyrtRxGdNbBoXtHRMRSTjqHFjwEmT6CaMqqlhOpIqQ54IGKvOAcu5FoIjLD
BiQwBeqynQ25w9di0hxcFN30PbAgcZ9MkgoS0isMPon7iinGdiKfJc5JjuDtjQY6
PugQbeUQ4ab8dwKUoF6bkFi7ZvyB93Wbt4P9DEx3hGKQj668N3/ywN9vuPv7r9+X
+zrd4XJfKXXi38z42SsXdtuucQjmXbLjFMdOttBjqJjBVPQp+9zrXjK3eFdVYJl2
lV6DmH+I4vWfO0q4rPv5tW2/jJyhM8E378+i44fd5yxuLKl2f6VlBZxFlsji03OP
jptYBsHNcfDcdoPU6Lf/dRX6ho9klbyRBMnk2OJtldesM26vLrY2u6ZFpH3aPyEa
JWWUyW2vzNOQ+k16HDL+gOA+eUIqDg80k/qs9ecVuChEdCCR8mFw4KdfUhOUKmlX
mScASO0hcqaAyt87pT5nJwrfWMRD2K1x6QCyqz78cBE0vF0liBFE6T5nF0H+paUa
vERQjigHBr4BoOwH8Lc+t6sWyLHGm35GEbYnuK/5JlRuIxIyvS9UL/F6Wrbff+HN
ho54AdBh28wX2QvWNRgUz/84zQ3ZaKKuzCAYIunVM3lBg2hEEUL85Ira1LOnNcRg
uk1+qIHD1Xe4eIzcHY3HfFH0fboAroEjdnlF1q7MgOKo3zJ/r8J8pu+8OldOgUnV
WLrSqMnWzNh7Twe8tlF9lbqwAqzuDKLHCH3FrewjBl2RZYZgMPiq1vWzqWqS8GTU
ikCnRb1PTfmImjwrJGts/Mkte60RObGa6wpNjhgUkahkm1HSHqtHiLc29YIIP2Ih
/MFGblMMffotTK883ll0HEJgipu/lpoNeUs1yS6zIMWk+wxAuDGBM4BedPf/yW1d
bWe5RyW0eIECsV8oAJWM8DyxBj2WB6t02Mk5TW21G3bcmWKYuGYfXr7WeAFZqCBW
eJxxKXEVziSHvKkhEqYCX92AU3ZrBziwlx1T38tL2TegLFlDCuQPh1udBCUH9GQF
GDsjgPMbBcFvU1DTHqb7I+0GU6zg1tmCMw7/RZEpsy61h7WsdUXHodHRDl1g87GT
hnEkMQs/FlUD1z90Aed8BRXSvynYDMCrXBW+fnjEUXgJY4sRbNNAVFrzu/Ubn2/t
nLuJzTTQnVPy/BWHkdACHAR+pePbM4J5HzsG4MUnhS6aGa7xYB4RpqGNZ9Ze3Kke
qRCVv9MZnUgKavR4WfQ1cCYvVBB+ZV3m4Lc/WMntuZiRofsWthtNKfEDDcgEmZIC
9qh/APlt4WBwtKG4a9bB9pn3z6LP51XFYZXnhMISIOTKC0nMKauO3Df74kLBsChV
kmwy2lRnmFwPrLb3c5QenDML9p0rmekmiAN/SUzxa0dinYdU1H2nAfsvSohupaf3
GZG9ekfQJBoFwi7CzDYmvFEGVJ8dg9MaUyWsBX/bsnxemvoEbnMBvBdl5lVCBCsg
8JqQ8c1VVs/R95N45jXLn91DMvPDzM/etuSt+79fv3UYB+UaoLyXw7HlmoyfV9m8
cNmOdbkOcqUmUjF6H9gFpSlLNvn09JJLXKs81GIEPMCLsArjMIc33ZYlp5RJNMIP
lM9SFyxtVPcXA+i+JD0DXxR9m/ugxusf0U23cRVpooNJMonjvdZDtJ7J2rTytaUE
JqqtzBZUhB1rhqyiIYqFxsbKpIFZ6U4t93huujTqUupJikgGKs6muTADs1KJtVi4
Ru9VWTl9dNrizndS+mfQHaYVO/gx6jlg/uM0kiiW86oZ0lCWn48Y4g7qnbNEEd0I
JNWV6wUeJRgogvQX9Li5Q9uyVjtkS5P9qVgkCQTDpYjfolXO1Tt1ubreLPItHQ7u
tVHNwb8fXKrTLPOpfX1QnTfytZXJ9ahfrDTx3Lolua7YwXCwt4HkbVDs4H+mf3sb
YyHOrCM3fvgCM9WEW262jVljHceLzBYBI8UixgwviUaLOqia2tZE/idUjPyGJtTZ
yPty6FpoHzOpgMCD81MQ5rsNOzMGkEAA+O3noK5f/J4Qh5C5fh8kBJeawwmdEVux
tjxWUofSq2QcgM0IbrQINb2Sf1/Ls48M+zgAGUJg3USOZcVbUkdejo+SfAhMYXuX
FpCMoD6b5YPrvczUcI5FCHK3wbxIro0gRct/AWhs+/Pwng5j5uEvnuzAU3x7DCW/
TlcziOITGK9Gg1ILZBrHz8XT5fiM6ETmvwcXZ5qF13YumFv6Z5V9mWKLFUwZgFtR
i/yuY2k85qyeoqxjKTeco74PkXx76XzLyNDg1b8UnRRdwgQqozDmx+ODcvndtkqB
Vo5JTDOoFrM8ii813J34hOYziiFbaaJyFhT9oAvzEyaCAw9hYbJQ5w5echI1eGnq
JzFhRPAghlAMlg3o3hibaxaJueG9ZPK+h8RGpalPH1pvfQFN/ddYEXLmzxJKb+fT
K0HTefy66UgJFA09aiTgyzacHhq8taACBlFjmet1oHHZJBWr+5EMyPoa3cC2eI68
jUKUNVt+wLE/Uj4R65pwf9FTQbG0H2v198Y58TYUUyySoCOG9WpUPIfHvT8OxTtN
ii88w/nlCGBuNvfUtzE+2D9VKbf0LxS15fHbTWdvjGzE15aStoAWLBpviDqrV4ej
6dIjHBPcosDpM5rvVJwz/osy9gt7WO6zUhjtpmsBU9hxfXotUwEoWbzO0THdrojK
m5ELxRnRce3aR3iVy4Veu2NHmi5ZacpgtxohuZigTdj3lhZIIkVprr2MwW0vQVJX
A4vJ3r3BbXKAoos7ac/Koc7Dom6A4MqFi1iIfcVttmK+KTMkjtemWy617f+GBGtm
3JX13pwD1FkP+3NbhVLCk0IeoiIed1MejnKxvzWo/aX31wkGUy6z2hjkqZJABZMH
gL0pBMk6AImg9j9hLxZcG7XyeTneWQfyXf5Z6/iocdaHZOW4c/l6zdvxozSc0lV9
oZCh2TTKW1wQ46DyG+sYpI/AiwXUeWrOHDiqVTkuIBsRV9sOlpwehqTO5Y9gNBV+
vrowCKA+WrmsNxEs2mQBUieThEZK+VN5DrPhLY6EZ3GVUtv7LNpivtxJjvXnXX2L
L8gNa3OdgUL8zO+0VASZiQP6ha8VFQooRaFIotxPvnjaflltWzulCErfCZ2h5E0J
eVakvtS22xjwfFFRaQqMNXmA2TqK6GOMMUeGF7IxRr06rlW1CBKAw5cTkrPffwmc
APWKIlQvQDGugOMtfRjbLKH/9GHPGk1Hrj0MDbLlSWiQnQipcJO5mEpV9QDgTdn4
NQIEx2A4BuPuRV6Dli3l+jWTYXUCje4pD54ILEdg39rTozsBnGGemmt7z+1djs3E
aYCAqHDDJ3tpg7hgEu8s6WKpDmoccm95TC5obr/WCcowT0YNJQR7oYnn4mFO7+Rp
fRWRbgTOTfWLugia0lRH+C1SHld1YiEWMhCgX+rwhwFp6JapHDVmgrzPRhNfPhdE
/nXkeHSVkESyN2uCvjUzS81I2leldgZPYh+ONTHaouqR8OTZys1GPOfqyobGWBhq
ZlIbvFqX6zSX+be4MGK/y8FxEhhVaSvXlox2XoyMixHLmqjZwGW6Wqnn+qzt33NG
ws9mWwz75zEg81xn/KBnTNYTi3NKkVpDAsqYHi45nc+U/bcm4VRd7AHz7Gtf+LtR
AfA41cZbsQTyUCHXSyxGUYssphh+Ef3Xv7nsVEBczyrsgTjzxaRhn5Yo0ZMi2ptl
hDLfpX1aXo291Ff1RSdeBe+jElYbl1snyhVwH731unBfYnPFqNpyd1u9+idZqXdd
Gnv4/Zpjdf5EKIbIYHvhPlIirPcVMy2VAFZBG9JxmKYWj11GA96Am6hrkuTAugvN
eDXsPYw3mukUvXAsmtweRflddCAoFRVedjfiFnzkThfxPXEgUoD0i83vKzuPUaNc
wuibjo37DjJvOTBwtihLj/oh9tIE3JWpebZVuVqD5bgkep1P+6Sacy234iVdU4pm
pPTVdaKdDJX5NiAmldfcVfMO+OH3GU8iejcdTZK+YXhR70nv2m+6ACO+jKS4VRp0
k2C9ZkwmTl5ePJjUg/4DwquPDmXtSkyDZNdcwtwqILXnYWgqsJkpVPwcsXVHn/Ji
52H5MocsEoCBEO85fQgInNn4pzg/pHE3HRAITcvX8+yZn4CL+Y+jBLVaEwyu7XBd
zYe2jQBAjXcsBrnaJLRNwMis+iclWffiJ3253R11HcfqgUYqz6owXyJUGncji8x9
NOxxdfcAHdBLaOuX7Z7Grokq1Xj8W0GXvyXH44u8CI0qYslBo3S6dEQj7wK1iyFS
DHb1u4wbRoYwMmWk75P7olyADg89yoOGdKd67I9YvcOFYOsjLQc47FlsD8zDpJeY
0b+PqXxW7CS9hiRFqDvY6fwf43PKmb3RD1oayDQ83uQTBLmJolakzUTLmBvOZSyN
hrQqq4B/U4CfVCc/4VVQXY7z67IO/PJoZmBCr54gVYOT3lrLR2qQonRFrRDwJ6Ir
gPo5as7mllTd/kJzIlHa5PmLqGBo9KTx3MWIuIu29s9Z2WMjuqqNMuGxbnRsPIcT
4P9X68GgLkl5D1HjlbHAShmzTrAnK+EMmDzSvD8vkvIevaWcQWgfuyC9IS+DhDz9
dlN4A3sR6ZoQ2yvk7rDsoR1xV746yaRsBqDKg3+Jmrc7Xhb0LSJJTCf8FXTNOZVl
6ts0TojIvdPBVl7LAQYNXjzWXuaZbauyKyrNQqlS3g59dM89oQcBjGNe54vEcP/2
xwaWPj8G2QvX30ZuvO1JYaG3okFMtS8T7H4TFIEjlyW1AQX2t93ddovcIcmO2BRn
fN6yRqwNHGwma70pTR4crGE1IeS2vOD6JvAGmPaSxzMSaG5pWcSRCTCmEJhLyv2G
khm5Qxy9ON0gdRGshoQCMZZ0023ht5/AJKwvwAJGGVy6JxDdunE2OJIZwhuNbc0k
BD4mXWtNnyfHxHUQVDt5idGIhc4Y+1sdUgUIXKvtsigjeUYEtaoprywJlazksO/P
QhaMtUXJ52W6qFNtpKQtmGuv8iyYK2pHhfj+vR4dLfGaxEM0onS/uBW7W2aUP6Ud
3m13TyyIuJ9edJe1SiTtSXgn8ZCprMCK2bbuXIgRVImOvNWMSJAfYv5MkvPYZEAh
o/6PArHozLWxRpJ48wFC3845u3AIm7XhqD/EkF0HnmDQF5MtUrqjD6/wbn1wavIJ
QtSdYo9yYngcuwD+aq1NZ7y3bFRRDD0mVaXxX951IRBf5kDb/fdCoHftgLt6NUhh
AcnogMe6s+wsy5GU+rMGLUt5mVNSgeUs+swtkvXf3dpt6LoffgNNOyjx88S/Tphe
FvJQFoP0Gv8R5MoxR68LgIcmgWNTBxB6nryeUN9v7Se0N169tnB9NJpsGHW/+t2d
RfIcqkh7OAxSITu28PDuZkDktmaLuOFZ7sqDE9qMkNBrSmi+F4czaIo/F/5Fe+ce
dRPk48xDK/U98XY287xIfiad79XzbDrwIDq3awn5vGFftEBOz8Av7gL8YZr3lf7V
o5LeYP9xyQx1v0VsANtm3cGK5Fr+SJIVXdqHGSMUU6wwHjxyTU34A2bQnFulycsc
MQliWldH4pfr95k82JPJT2wrgaX/4ks5CthOzJrsFB4pueXgENS9KE7IZvlyEepI
0cdINn9vrzMQCrPYdaROQvm0d3lgApgGSbQ9E77NwRVmkh/CZxyrOy/ftVww1QI2
JMbscTLup362EvzSEws2M+xxDThH0GDGuIVjsHRTvTqXsEOrWHFYN6yuSKaEf5Lk
wXLpoFNpTMSN+zXIXXUKWl6rYBkL/9PSoyHR1YesA47mYGXjj0cQ29HrTEk9rZ55
cOvvbCqACeVy20XTsFoSHus6VZcqqPq9nwd8zk08+0WFbzWu88E9DbASMk1aVfgu
elt1cJaC6gN9FH0h+MxRXJdlOhQUfdimonbZ6y6cdOkLs59yrUBQJy0bREZeD57a
S2oN61x+IJzggw6wu4AiNZMtOm5//T2zbAOezvqevY5RHDayVHNml2WUTd1q/05K
O/S9jrtDnyqWCgKexk+z/eCGJ3kY79ToYIY8X9cjQERR5RUfEnfZxtayXW2MJXie
MIiIDLXzq13j+5QDdmH7NsdGnayZdO9O2+qlnpGzuc6wnDjmLdaWoGFIOmx1HDoF
LQJbUL6rIvMKc5sGA01B24LRmojfn9yWZBurfpuFb+Kyiayk0XNCXsfJzwTMKpvt
lkyUpZWdVe3uti0PvRI9MhRzsQrKzfA6xrP6WeKxjSQlIHOM7W25qiCGSTGdhWKH
kLtk8CF3x4IPP8dPEFCXQx/BXSEm/7pVQTZ7JOI3bnhtQfhhYN1cQHG6qtbwuuPZ
nxf0CMEm4PRtYtAlQQAxnSTZ+mkgVrGvFVhq2XWWNDGH+sc2iHxDfuZTkcIkqKzI
WmbofMWx2FmID7Jwuu+qMx5XCxZK3F9v7K9gaoU+1QiB7K0aCEnHBJvGpJsm4k56
J8cfxMTnNfFhsAZEBUh7sHwWC8A1DPVgYY0/c3OwkdHggcCXMk4lsfXYJKMtoHoO
Q1FrK/eJ0Gu9vK7/ApLCdakbkuEc7osfP9RGuMBDTU1mzrPfxhE30EoWMcZxHGTo
guMVWmZqnr0nKLSSYFND89xIjOZk3K9qJwbGFe68NbLUAAWtS1b1ypihM+O+qM0r
702K+JkuiycTB9HWuG0/I9oqCFONvX03Udz9WIvqHvDsqxG6Ze+7B7YaKgqahl84
pUnOB8Ork7RsRcXEDQrqIGHduOY0RAHrnQcnKSd/nBb1GecZnVyvZhwGi+ZWTrLA
60qWpGgiJaxEOLGksd1IwYRMlrhQ3awxjqKi4s49bSCYujXh3cY3vQxWGSrF2+ST
NcKbnHP0aNBTlelIm9FEvf3u7M7yFgnEl2+Cyg2ERnpQ95CXBjyHjmT3jYbVlLBc
KJrAunByFtXvFgqZPJGoXsTTvT+31wEPOp56xGpxHgMH0xNdMScp7Z2NeiQ6oXOT
k4jnixMGTxii0Rdta05tohM7Vw1RqXlkpelAMq1x1W5DDxe6XLRlgGRGkLnZbsiK
IQauhXk5oAbHcsP0+Gxu5jKo8zvPSanXY6LqB/c7FmSfYIr23pNjSr8koyNa/e2P
3emtyoy4fCdHqfIMByy3D9z8Z9l5v382Dx/6nR+b8W4Kf8IDH+UUjXrbIdywQ1Ei
LdWbSPHBCJMHvznlu3kUW36zeKCgcxNIWQzMMmDD6ivaKTsjjMzlsvjBtNCq+1Fy
wpSIXWFXlWVcjTEGkU+YGRlI73kEWXU5LRHcZK9fMTaCwgagpOnW+BmkFmUQLE5Q
DEOd67xth/iOoOQrNCuECu3VOELyA2lXCb+dVMqdCLF/3rtzEsamIzaoB35zJtGY
gihPplQUzVSR9vGthd2C8BS0gITE17ZwdsGC9dQMFFg1ppdc9PAesmrEcAmQJ1ss
iQfvAVz5AaofshbzRzogfFFBMQdIGGoVnKeD8atXSBW49lFW4YaHHt8aa62Azkjt
ZqsIa2AVji1IMuk2oQyRmTckMZbPzgBv4Ck4Kdy9uNvxU+/ld8ANwnSXpoThlFSR
YG3BbavL+z9SXp4b9V/ppuVqWryzunJcNjuNh3wKHdC7BB92tspLzbpXNqKDZ1tN
16JwXUQmv8+bT0u71z0gY8VXDELekxYzA+zNXevZkOEI/RdTU+syAjTU2uyFzGt3
govxM0w/dG407ymPlo/sa3iNUdpTPS/GJD3yq/QjFozX+O/wOAvFvgcc4T6Elhtn
EM+SuZ4IRju9ZWQT5Yqd49xCEHkssNfaMCM+yR+/YHhwZuyvHlBHmTaeDGUNtKay
UYjn5WT7nCekZu1iGARK4kjqgWtf6EPGKPcbYkNiPbKIw6hdyQJduwuxvzYHuW/5
BO1naFJMx0Oj+4m5CnKwHszWgu7UYDlUVzr7SNOI3rF7hVj/AEtSkYXxaUNqi1kO
IQPn0DDWshXVCVwCIHJIX80aafiWPtUqfSd1acRKMu9H/Rpn9D4KSRZs+jbmvmnl
xeanuQPGts5g8PUaLk8ZyVBeRas2ONijatnyXk7o66xpD3yT6ddZOx/bWnVdn94i
7pwPlv15Fj4n8FoTkEUwdUVImXNDQHvgXf1VbkZB7hWjC6wir74TMVCrtLtrn6La
j4himne9m7p5sQbjV4IvHPblKgajuquki/Hf5xkUWAfpLQa9vFWWUx5KxtKC9Yhr
HTlLCNj0zhCHbXkNNLf3YPHnxA84mG6dRxMfDJaU0V+m3SwTVw/fHV1imE9hVznv
+CCy6206hGQ6+a7wbk+a/Usz9LXQYL/9S3E5g1RL4QN6yHn8DGCXo5sVTnqbnN7B
vc/QNhDvSIdjNoPRxcdPBVG80Mvp9rEEvyXaEAMyL4Qo60E9nvML2tGaiIwQR4Ub
+1z0ViN9CYOVU1o5OtVb0sBF/Gm75UnzZV7MoSnJWP7CWwGPNnll0Fkg8RuZhk1Z
cOIiJTMt7jFBefCKREuMJzrqnZCXlwO+9j8m7qYivoSZvxEl6h5dweOooYDNMBWv
Qlyo+kPpUkmMZcWSgt5TwpCkwkaGXcG1qTvU7A/NC8yMCyzMHUL3BWDeGGvUK24x
72WXDzu4WkvIKHbzh0EJh1iLd5tkXKh62syji5NMFWYliaSyP0nAMlrmPtuulHpj
2n6GEfS/rPLs5f6MZcHnIXzu+OH1i06tlrU3aqGlpX2zyAA83Gtp/DGOI84PH7Fs
RSVS63KxOwzBkKy1uXDjmHVnQ/6jyCA26Wb014IdkAlNPhYSByaBvjk7tOHt+pyC
X9adhFLBAqkFs+hS+3XWC3l9BX8SPWD+GCVK14tnzgHw+Hn+H86SaApMMiyCPwpV
FDAaN9ZLKEAQtHAaSmsC8QSh9UidjrmnWboYy6xeTlGbCbEPuaauEfXx+cTR06zk
GfbnFx2irG9wLYE864OH8ZjzJ6FQtF68AOGtmTjdLQ9YmTDBj2XuwNUyq09JnT/e
AwckApds5oKcpM+6oPXq/ke1kzob7kFa/EgIBTdOJgBy4VeW1SJA3uh0xnBE+CGX
AKq3LRdH3ufVzuSvUuG+y3yxk9f1rZCXp70wJda4RAS47QrI4YGPHCPODpm6Z3LN
w8lIVUw2PEn1Y4pLoh6pYd5U0XLycbAs6PdbcZJSrVqeRN1AMFcqK5QnGPoGeQlu
VFwQRVB3I1th6LvcgMzPUB7hU9TPgPkIB4nDvq6SPMIHiWua+haiM0SNGYoLxLg5
jAM/eeYhB4zej6Mmn77WabcQMVUCFz0C9kzqt6BoyK4GPDh7JorwbRZHWrlLZTg8
eGqsnRMK4qnfnhbHCepYYPbDmvg9kTu8W37W6XBq1aDEeu3G8Z2aT2aMfBGHmX5H
hQYnXPCDOmZYano6Z20Q9eT22wfs062rbcQ5rSefHpIZbwPa0HM8IwsvIIk3kwOU
bkGC9ZdRRrEEkztGLPPot+TtnZkskBc2QqIEjXb6gB8rS8m/ATISgFmuY3tj6hQx
OeC1cNqKomqOZ1KYrwKBr4dVdY1rpTnWCgBcSDz0pZRUG28FQPqDbh5Vx1iJ18Zj
jI5q/9YJgzgFiVuRcYToOGKwHaA2GPOHd1NjYOvV5CydGeCm8fZte/ZCYse3R19q
ind5oRu+qL1Ia1gxmTMPRWPHTosvPbLEN4k9snJSyINO8nhc3OXOBRMOeMyvoPeX
pK91ND2ZYKEWFhd5aDig1+cO161Sn0obeeXcmKo/mjOBLGNYT0/uAsv4nWvwFP5z
ljWxFDm/vNliYLXT/Ae7VrhSGqd50bl4qkRa6uC731XuUywa/AbgdJa6wG8Z1PDa
CXPtD49l/OQxkTTW3JjOZd1V2HmN+M/xi1DPLdfTfbhXFVlkASWjvOr1HjNlYo0N
PdFHHd153NKjKJRJaApNVL6YbJXioUCvDs5zXqyBcYz+y05e0VI3Pln58ck/Bcr+
DzLzdN+b4cLUtl2lO5r70OwljoNWpt7dOnWUHYMnIbFEnksUXDu6Z3YmPCCn68ED
TsMHbPou7IXgz3Z5FitKFGJg7PjPm/St0pHcuReVVdN6DAEGPefSXTuhCqS8Mu2T
d8TOgd/B1erbFl8f6p8xdFlxeuTvPxg1mCDmrjilALyXfwTrgQm69Va/iBTHS/Xf
I9n4U+0F2O+JbUAEacghiLkeYKM8vOur/vKBQTR3CeKzT08CuOG67ZeD9LsJ3Pc+
3TRqzZHInDmfUXlkqmL6EM2CdU2yNpfd9UBLKUNkCLSdp4oBOVOkT7bYWuZUzRQp
ZuQRGWxeH07gnteCLR2HDzHZCLWJfLG0aMceONLq5l5RYDNxp4x7GT7iAjBAJLDb
vdgUIT5ic+azSD1jiOd3ajyOMGPXQYN0vYkbQHHN5i/VEft2WzRB2abeFIMyUqVR
uWqUI+vSChgdlOo1pXSm+qYCinU0lmFc8DikFLJdQnrh8eE8DOVgkBaQauhhhKU5
qXc4z+3K1VDdZNGmIBq+K5Ts36C5WiUcOn4FHPncIzNoINxGBP+YGawtvQQEM+ep
Vg5c9REdyePylXiyDKVSI1Q/KVBvpu4H57kxcEWhmbbiJ8CVZkfls9Wf6jLK2VVE
xZyo2ZxvETvDOzhUqiSIQA0TASSzTzeb+kIIs1/LrQTJ7SllZDR9kUJIVf0Qu9dp
0G+iKLPbG2XKrsP653AU8ibgrs5nViQnYgMwPGUAgfSG3g1MpuTUqdPmmDvTX5D5
iA5XUwooFRT/aUcv4A9ga9HhwPUTBAGw9VHbI7NXkZ0vggqNmAw8vgS7o54V4m+R
njQvYu/oZOfmzsGx0kYd+3/xC23SMD3Mq5q8iHsHDq5XbcjyZ+dhDSTfl4jVxF4e
VQexxexPCEDpBy57mQNHQWKqZHRTcWKMQH8Gxfbf30GVWpO1OziWb7LisVU0lv7F
ubdSjQZmJpTa7ahGUizDf2wawl8F5LKXeB384ZoW6SyddXgwdxRQzm1iNKtEj5jq
Nq2PHeRb5h4vfRBlwDpbSta4yowLVSmhKKKLgkHjwnm0pW4eJ4ukxNGD/G5IVhgK
fvIaxmA9V8Ap7B7fwriqwbRehV719TPbCwi7tiLC/OxiSEt6AIJzCQ2ps0rYFRkE
H2iu/58TVVxquFFY323RXuu7g/23wQcGOnw0kUAzdcqzG5Q0xtVTc4s+BNt+Lq8Z
uLg7WUKYYWAFq+P6Ui5nrUmI5hMT/kqcLatXPDebya5VJbxoQGcta30LZ95XHBT/
LG2Ypp+jbCEG7D9UuQIm/gNOTxFAExtjpQKHWZU+I9nJSLHegCYkXdm3GD3fJfsk
gqhIHw9LVvRl8y1Ni6mW1aoES+pxdhnmH5thYUf9pq5/rFTHjcd6UyJ6ZIOqzZOP
xkxWSpblIqQ4NEeeKb7PpV/qCgakYu3NUBHFECJtB3/oLnSchIAC4tbmX8UX7w75
VoJUyGbbqSwPA99T/fUmBDWGGZL9z9rt2zqvxxkI7g/jp6uzDv8La/nKEI7m+LZm
W63tSItQ4nx8CqKejN1e5+tfzRPr8+/BQKm8kE1PuEKU9RDlAFbNdMOBz66UOoqp
I5VkY+BqVJblP384lZ9f+jIARigE7vWp8XGLSM/q3tlQRRhgoGuxewhff4fNyzxH
64sG1zQVfED87r4k7v1d9rASIkerleebMVUz7q+gdMk4t42OIDFdBw7aopKJ6aSa
B9XApxYS47uZ6XKYQZ5cABg5nKY0mYDZvPPsnIXm3ucCfD5jlFubtqwdBz0esoI/
Q4EEkj5wkA4o1w28mKnCkP0RWs1VMr/fbmmoM/IO+AaCnTUUF/r+g3SwcpLLLJaq
ZMpTeXSBRHO/qm8qrUK/7xt76QCdaoRwaelykdhwsBqdJ0pVJM/rWZ4C6lRDVvwF
61b8u+dmQNaJ9/WB05ldE3GlfwxLeabI9V/iBo7zjy3ZIeuOuKty/aoiQZED4WZS
C+oECGaCJ3A5iESO4VVbQnAdBvOWDqkeK3IHvugAes2f6+P5wXSOUMY/cIE0cqrT
tIXbJYdUdN2XMefBiLVmxvDOM+96kDFbRwMb8rVW/kJTSEBShr621Y58djI4s6ts
o1Pzi/9geLT5am4tXc3GY4mEKTjY35+OAvubA6tPWyd17yI4f1K8MFKOYEO4aVRD
0tWe5r+JLoImxZip+xf9ylAlS0oOVVoQ0Sv0S4jmvkJWYIIyrqzGLI0fq6wAzPPq
FmKT1Vz6p6TbANEUDbU7PAY83pNH4PFK0bN3bYO0ZyV+58uLbkZmXtzs70Vmn0G6
yykmmBsImBhs6jwP4Jm5KLrluT/3g7BcOP/H/fatw7F28NGXISbe15dRYvU8hp/v
8gvmwTnK18iMMHiwSlfMr8iii7AuF1TP1EMfCkAH0PkW4Ay3/hRPA3NsaygRREuz
KIpBVhiiQg3whCQC6/DE8ZxFg/T4ZA6Ktb0342sx9i2LjFIDe6t3mvh6cq1C0HmA
G2tdTCZj19+24pHGKfTi8CuhP83TfGmEexPwCctDVqWB2tYLeRB2h36xq2mZurdS
47pLWqJyJ/NTJT1gPa72mU9hluS845oqR99JKRYwkeBYkn+8wpBPearG5AB3kVJN
FKPbZ/NO9tJbNl7gBl44e74rMfz+l2UJbnUZbXz27kNtOWOzDWzQ+vuykCroINlz
sF7j0IDG3BTvLKMUIAhi9qL8wvCtVjHdIy2U29SHiDvES/QvoHwovCuWfXdIhO7m
5JT/qq1JzRiS9ToI1FKXaQL41ORb4yind6FYhLmwL5tT7bSmzVA059QasPSFYvMA
81z74Ww2kjll2nGsm0leyvrArJvMkN7UyLJFctyMiEDweqQMg6IJczKPEDQJlSXX
IELyA11g3vIMS5JDjsAjCZ7aktOtpf0H1I6fdr7f/bnqxwsWEhOjhtNHUvVwxfO3
R3tob99BVB1Oy6Q88DL4BDbQ1cWfaFXPUI8nTyMlemrQRg1SalUO7qy9ileTncsp
VCYWWkKz2Wk4Fyf49IInBUEUV+KtS/2Lcyncu5Q7tj4TnuFK7mqjsKXFgtP0INgg
E4ZkXl5sZB2xolC+ukRCIu9aZQjI4nGmkM2asFnPH3voI5Sqslu6kx+HPIYHezx4
w8EIVX0LxRQthq0UmShfRLFCyhdsfZv0FsWm9eXmNn8d3TL+hwCUdmXk1Dl/c+ll
TCrUnln1FMCE1EINjbecNdKe9cxnUvRUIPCy7VP/kFBYpxLrej+TJe20eTglnQIr
a/D43H8hj/41x7LlPNI66dMgWOc8wmas9/F9vZDqKY8HplvGz3F52J+rbe913nEd
7UeijWkEmepZWs1l+33pB1P/g3EizNV1+aGnBnq9eDDn64stZMywWjPUkYXchRPS
2fcyJguZp/3zr4/BXwAcEaSX3VQjoJ29wx0quxQuiwZVVgNlJpUJl7ecS6pnO8MZ
6qIVGfjlECwA7ov9MXU+fJvg5FgYClqiP0uwL82G6qPP7ypVprwa30HGsc1pvvpC
MHhFqBxcL4lufiTacTm7Sf4RU3JXHImXF5By/5yxAcXGMVhQrWd1JBkF98Lsk2CB
mcMucUOm/0x9SbpxKfaMR9b2uJfWBDonmyuJt3XsHJdxi5Jl3/3RIVzm3AQVIcJH
EemHepiyyqWpjdnGnD2N9thgT41r7SEKecBGVkBhR0C7c885tM4hSdf6qkX3F4yD
Wx+49Og3Rad+zVxXcx8j7Be1o1k2IpTEfq0xNj3wRZISJmz0J+z78Hc7jMH5W9wp
kKZkJwmkmjgUozqII0Lq6affuoPxq1W86UEOgd0++UKhMBwRfMjXAduSdccs0Kyd
xq6crKsQIy8/tvsYS6BYhFYk+ZC2Fc1gU6mY5ChLDDvj0eM85l+cnNAu+gwqiq1M
YGgcNH1QQjBEHn/IKECgMNA5kBJYC68vw8FoajDhzzaBePNPOomrHX5Zl0m1KKdS
S4YEsYyWa0Ugb8w/YExU19xxYRbmPONkwmJXkqeU+n4IriDU+cRRqBRD53uva4vQ
Xm4dNvMj5o+fuhwnF8tSJv7RqsTF4sbto3YPhxtCW7mT3lfrgAqg7UqkkF+2I1Dp
8rPUzSu/tVS89O8wlS/L4LRy9o1srLLjE0I3gO+d5XEcUxmOI6Ite1Gwf0nar4ER
i9DH8qcLw1dzEberxKs/9ddmqwfbIZHUSlV4LzA9uGXb7qH4JV6QzaCXIQNdk7Vx
cEvMIDBYwZFhlIU97KmrPTza7BQq/zbW6Ia/HF04mFVIXrMO7uvVjTqu4pdDos8X
MKn89uX/ZFOLGdCGF4OPPZwJYEEphvDY+4hL3ltl12708IboiAQr00mb8wWMI5BV
rfDzXKb6VtVEWJOEQv7Ni5QPUiAjkJIcwgbRoKxmKRuQJEcmV5U3zGztvtTREHvC
veyilULRZ++1tT1q0FjnsmT04FQYu38Ol+BnNcSuTT3lLEbOlS3LV0bJrQnHL/Ub
3PlkfPG1nl2OBTWICcpGsv+rInDxFIWidaOT3ph/Rs/NqktVi0T107frT3ReAaJm
tDwx/A3fc8UOuv96wy/LsxLMwJdurOuc86Zt4Iyn3JFhaX4OmKORm9rm28lScPEo
iUDbmJHhX2SorGqhTXvZ2ER9WElCykLM4ny5JRx4K7Ge3gVfUvNqIMgAuIjuEeuh
NRmKnWnW6i1Wk1TQQxxPR3O4go0/LSXJKtmV9lw+hUczp2h/wMDyf+u/iJBL+peV
JtRYgM684YHwqcsICDuKq4JE28lBMrf+mcvWR49gKkqghqv/UXTRAaRAZsFsjww+
9lMeTY8Z/byNK88mx9vp05yt2o9tOTWZmo4sPL6XXIXWnUDI3tKc4OA3EbbcwjZn
eJy46y3iFpQ+tfch+LNT/W+WeYv4L6BgZCBgXha+MhHbMONj/+PhZwNjy2lt9jF1
XWrIKCFDgLITh7NXYWOcRtBeZCbTnaHz8PS23qaA1YdpN5mC0ALfMOFPTBBU3Ezv
kXWRh4hBfXCtQp5B/GoeyGwpdRFcS1/dybXaQzgZuRRP/yKQA7GcYeTvpiyPIFh4
S71IF8WhyI5bce3IB3TAYixdc/DzwimigS1HwJ50eghVtS/FJSxSK9qnGoSxT0s5
ic2UnV4TE5XI+0Hu0EbPXhEBx/wIluXJErulUuHk9xvLtGnTRVzygG1F4zrSCcw8
1D48fqGZylPB3WSqfjR6iQsQxS94iLHjlOI3uwuI1WGs/8jhFuJTreBN+QYK0ohn
jNM4QxRlj+80w8o0hgYrniWvfzoMDhd+LdJa67GPtfmeeiu7errXWSOEIk99+LJz
PmaIacgGReCMQv09wXWsYKprNNglJ2gHMle103B2ECHloJD5t+v5AYKpcG+FFuvz
7vSTeWWOUTxMleUFw9sJiKX/JxTnM1ChrWO676dbeHCvzLtGn1qTllp7L1zIcZ+8
ahY7jCZkRdFbQ0X6yQRSftIk18ysYuZ1SPeUzXEORdLizhSCXVZ/6WLrCuJWbhjX
mdZGFXiM45mY4FMt+fSMV4DKmEonEhDGf2AnkDZn90f5fsr+4G8ByMhrxiEw0Vb5
TEobEdNgMk7UYtwrpgWt7/fnGwwax2PxpmaT3sI76FrfFYE3m0IeTflfDo7D8o3A
Q78xdhd87yKh+JOIIouAbOccAmZNdL3+UhDAyLln0CADXb87hEgx5wjuGJTqgqbM
VItNHsryEbDwy9Tk60Qfq+mnqZFFsl+inOsun+dHI/6EFrA/PNqNuI420s+VkqQI
EEhR3zrP3/JZ8ORQJKzjE63u7E65zUm9mcx6J0x8FBEtxnDHhJDCSrN6d+Zr1sAi
EZfnIZUou/9MLxrNnfoknigbtFTz0rxfsND390btZbfaqSim/lQOJp/Vu1NAc7yk
YaSLWSPDT922tpFOw64sRgVg4zb8nQYVPAnLNWM6p94P/MLMIDgm4nxrt0+oqrcG
pqQC6ptI+9TFCN9QemK3SBwMrZFk/kwekoOVRofZItXRUuZwjFnnIUj6F9cv9WWi
cJcIXN+i5bq1jOg1OIlmPpb91OgRkJNA1VB0bisXZBfqdja+gUpmUxmhl7KFCEIH
w5Va4LfzfKwL2ZNzksTIupvftVsJ6xDf2ZATiwn9IxBvrb3WlChw8LuTB7813gRu
fACbEMhsNXI1BsWenEo5J3AXQ73h30blc6pKSOQDReCMxF0aBTpFgjhb99nMvTuF
OUk6hJw0YBGRaLXvLBWjFs827KSL7uYex3N+o0JMYJgx1iH/De3ahZ47I7hao1VW
4IUI4QJY2nHECE+oouzGfnbVRKWtLbmdPbbBuz4GPm2K1bpmdoDVLagA+/vgxwiX
XpgRzmE67/j5+ILa3BcI6SxdJd2LVDNjfpXyuX9b1ca4FJ2oDIhz9FlHNbSs/wGc
XonIjrXaCvdb9X37VFtPLWMh3J0AdvHqy8ia9wytjWsIeLrMA+ojhKuS3nIYmiaB
C+5lNF511f7WReOobKLqbalb2lvA4e60BUD+HxsEggI5UJQKDi3ia5mTHx3kT/et
QxNgHe5rENk6H43eUxnuNovEWnh7Dmx0VMEBzYIlZmcTOsbTO+tv5q2MZVuUH1vA
qLk5/CbHvtk1D2we+/l7KHsClFJKPzaN8Q14ZpyHEi6qkfW6fkwkV3IAOGMupaxI
sEIM69r/JimHz41ozHmCszLjcTNOo9pUY7vBXhyMubwzEhFgyMXhqW4ayhJVs+QK
mynNhWEEVzTtoO0Q6fGNfLkcRsQHGny8hRMFdoR0exp2cBFZBZMPrDE45iozLFsJ
eV20zcOD7iZ4c1zIWj1fCOkcPaqCTCmvouN01DL6GItV3qt0wb32ylQ5cM1AgY/E
pDWz/S5ufwNTRrIW0cBlbda/WFEJNqk1U176tCwte2O8jKVG02QJoNwInnUogZiA
3XV7zq04llWDNZJwAuNC0AQ9crvpVeqPDmrH6UER3ikPOLGj7gd1zW9GVx0RLHVQ
+MtADpne+L0Tb6CsKZ4VgGZebecx+V1aHeTZUtjwDJzFrIqKjuez2k3C/y8YR+aA
Qn4sLXMj/khhd59BAOMcgIVGtjtsYoBOJr5wKX2Heo4BOutY6AEyf5WeHwzgP80I
IvDJYvsfyBXnV23634Sbm81SHad4Fdc1NUXRNMhJHlrdtz9Cp2QtOPyMqWxumkrA
gFN8asoeuJLagcYyHmtnB3PvMo0mf/oEE4/186rT/8/Sq5HW4bpNx2njFiZEFhIU
GJt6R/bfrxqGF26gcqMuHpSMpFCtxYLCoozyrvDRYYeTIC4vbkcAdV3NEeoyYAQp
tzU4KQQW5ilFEZAKCLa2Kdllxk2Hrh6Zprr6fZ4Mgv3Lqb1YpOYxaRaQnMXuuh3o
LO3qeFABzt7Nu8rLDANzIBaK3Ujb90GHYKeNmlHTZ4O3iZr8uKxVth3OeVN1juYs
7Z4YsyToicLZsLM0MsROKeKW9VvpYTECvCTMwQLC5rThkOGvC1yH4wo8BVcapd++
b6zPVSIMeQrOmVZtDyviCUqPINgkYbOY9/yyX4wysLVEELO9iB7ys6udnfJbR1zL
9mhGiFu2XcurOP5rMzow2jNyZwRShUkqE7cLmYdgb4DN/eQpCWjeyhseje7iZQvs
c1j+TinQotVQeRJ1wx00U2C3CRN70BhxEo+ab7SHZM2WleFvKFrbSxCB0umnoKk4
Bx2MX6Qt3LUQt8x1XyIaVLGc5BA7atFG7WhwyOLrHtMq5juxJdN7/0K8Bq+jug6p
yJ9azTajDWr1t0fZxov2pglGORXCvlDUKKy3odP7nL0EhMHhE06Q4V7F19hqn2Vb
W9KUe73Qv5Y86YISX8oXrPBcTQHEK/s+XgjacOIOtSxRHeLOhYzMjtXglEmsV5uI
cFvSCkdc7Qerq8RtWpGsJjNPT60lZLE/6fHDEokcgTTfyptVhrWD9iXqET5qdVh8
cgoIyCkT8v7QZNgysasmN7PI3kkZrBIElLA3fI/wCLgiEuiVj4Mnjik01Xf5y/xs
GQIHYQ54oHdcNZemFT3JK8U1F3dJ9KAJmnmG/YbiAdF6WdOS6oDDuxkZKRpVfAEA
Y4RIPdobMW+KWabMTsHDHQicNwfXb7qUjSncNhlOKvuIk4RATuWBhqWxaORVOmBw
dpS3Ud0hVhuz+sf3Oemgr/Ts0wur/2r+ajQAjab4/8zgZ3fTBMplvtOY4WjvHvzQ
6DkR/NT8Dkvxq9x/4wf27EUL7TbXdgQRLKIpvFOb5L6Gg7danKTwniZPEJDLe0t7
/riNW7ClRjDgJM5M7p16jQmF9or9bsSDtAtOZtXK9dgCVziu5pou21Xm5Ryfduj2
uTNEOUiX5gWrc5ojRbt/Q3U2+otieMJiuCAE3+CbpI87kp5rpeQjvFZ7snsScreD
L0AusI8qlNvyRqtTQCiAAQASfGxVuh6mwTISN4bnv0TxAWjhLJO/PjParDNGyq+8
Z+umKH+zHyMYoK5Q7lyiDYA3LxQDtDebfMOzi4A/bvgeZA/7HL9mSjnHqjDXvoJO
De0hUN5obxTaCitOe+bK30ktrJmUqh144V7/ve+2+zdjzlKP/1aQE+/Oi5/aeuYZ
aeSaFO8Z6SVf4qBhi0Pwg0GY+79ynXBDgV8WLGWBaqZxOsVO3DoCd+NvIvcHl1LR
kewF0sjAazlilb3jRrr1r4dGt8AQbMByGZFvVvl8xgmJjXLC9PLwLlN9TDaIQQV+
QKB3CJ8kF6qHfhpspd9bYPB2Ky+hCOdxIoDHdsEXeqllSSoq2OG/ZqkEJJOa98xX
VLb5ponlDl22Sm0w0bbREQH77SKxxuUK+Ln1aZ7IbkPLf+NKCt9QaDck3V47SjvK
zVTHqQSOQ17+Psd5LxV7TAhenzKdWAZrFzLh4AuR0dHCue/q80nNmEk3uvoIt759
O0qTBp6dq7/eL80rYexGM7+BPxeEXtx0Zfi/S7j1Vm63dGV5fzmc8CuPRKO5Kmwz
PF+2tZk+YgDpdbUzuUmXsG20CvJhIlCk0b2c3VWvDW4ilmdVV5XWdlhZAHswcXFO
CZnGZyXyyFgDd3oN+nu02KgB0Y3oeZIafLFyH9gm5zd7lmvjPgO/7M3QV34Z9mis
f3BY2lGrtWz/A69KdTscX1IMEy5r/3IBt+YB/eisQ0l/BCsB17/NDFlsjf510+DV
BI0mkVFLNbCJABOPTkADPFqSRbgCuIQ6HXdxyjQKTqo+GRJWSEoclGRPmxf2nlZD
bU0kL4vlt4C/cHM3qwflF45iiUSit83JGxFlsrVbzdh/yioKLHTx9dgZ3um3g8Rp
OtBAX7ImdLb8N0f4jxXePhuRrOlanXF2FV69sVrln5hBJVNco805U0FAdL3RfvaZ
UnC/XM60RbHWtinTl2S6o1bbyc7F/IGQ8dXG7HaWTc5t2SkDtFQ5picUZNm7GDNI
gKPlUjFcki6xdCYQTmwou/ELVmP58yPcR7UUt9LDR8f9QgzfdcM192xRFqvpndiD
TuJH0E+4WrA+oZd9ngtyi7kvlLZiQh1MOCOr56SNairaYm+bCT0Q9q1xbIlyD0oa
TVvdVXPf9M3CvVcqGJqAhm3vptODib5TVpRlDr2RjAIshekfgYDSWapJkq845Tf+
GA9GrWbQPm8lDdmGYLxIargIz0J4uApaN/WQdhL+uCk3zeMEX+DVz7sYxq6w2kqA
JBXxpZaJqsb9g+ctLcbGdLMc4nKmJ6Bip1lnHKPvvCGvAO5/XIjMiBkFRQfWKjR2
3tL5gBQdwMUgvjs3q1Jf6yvZDnjqfXMP/Hfw1c589IEw1++R65FSvTRMwN3ZjG4H
Yf1TOTkumFkjIH3OlnrI+uTsIN0bfDtmmxc9TEPABX1G13XK+tBZvrbOyhQD9qjK
U+PWJCrYsVZw1uG6fB/HoXTuheEHazG6Idf2EljJKJQMJDTE3gFUdj7mIUiFCPap
qHKFdum4dYFtjkxcKlJXcpd09JFwgWzyDOZBL37RP4FXZ+SsQNHHwFg640ho5jpL
nWq2xf9EwpVajEZ/6AQPwjmpoRo3r06k+xcbhu5QLfeWOBpODSwjGr9H/2TVjk1x
22cuoJZmc1cTcqXzsLZTapkUzJDkHbxJlEOFhtbFWTj7JGb9tadCzFsRg/Jk5gt6
8koYTw7HKp4Eg+JXCoaGMVxeEMI8JvJl69VOzfKBUt6ZvRDVaYhrTTX59Lvzsvn8
DqE6yxsS58K7tfh+LBMZUF4e44Z/k1rtV/F0Of2dMj4/PNFUZjppDBeFtSqF9j1+
CHQGW5KQWY2xHoulC8Zon53UAsh/M2ERtpyubqSFGy6zTNIB+W4MJvB+8yBZFmTH
gemuEy3u3eseAwuqhRW9zQXqTEMac6GGdzKwGE7OeVC8SbKLPjX6/UWYbSnuZpmI
JoW8i7jkWSjX5zGHibswzcCY3IJlO6wO5W+4MYvgsUfVB0Avc5ItMLzzH6Ib3+Zp
6c5k+HLdXm3J7NfsSdnlN/+6tTCzdoeqgndNuV+HAXeJYu//vNA4pBjyfpa6n00z
U3qUL5jTLaGAl7zpDhs66gUTdPGBa30utDaDnZES7+ykMAm1Lk/HuU0YygX/SF71
99lm1gCH58ClV2ILoqFiFuyAk5Nsb62cAtQvg9GG/IHCMlyr51QFBHLHtRuEce/j
mPECYfmHWBUn2Re3QFIoHArL5Mbpo5BTWKSiZcM3L6saFsoazxSysgb86/2hMeAt
NQ6yuP6gPiROndXgyYwlQwcpDl3L0yfOmczqV9agyA1p1LuQj4zitt06yu0F53FD
MKnK/gsDABbiHrqQK77jGDbkHmKok5Nx6g5KzBNqdAEviu2hE61AJQZ3XNJeHS1P
YfjbKdzw4heJYfQPzeGQ/BhKaykZ634+XGzZxv1t63EX6z+UohB0kJLQN3p55FDa
a9nM4H5B6OZoSkiX0apqn4q91vc3b2btyr8/iewePNKaWM4Ddz4UkXOzfAMLta1U
QSveCORj1/OYiN/X4pdjfdEZI4pwmvSZMU6OioTBJcANhNIl/KengsGjT6g1b+kJ
p7piifsytvMr5gXQrlEPk4SioD41E/OF1wIFH8Iy7uz/e0JDvkzpVWkbWND04Qnd
qJcMBQF5l2c3DdVu7T1xt7ppjNNvljiDBmqf6RRgr/FKKB+9p27DjbZ66SU0su3R
wybOBGPi5ny0qqarlOnpyfNOIESRHdQU6K/tv/M65Hc7T7tipCZ+7wljORtD81Lf
RPXEtbdNskEtro67rK7szMAEc1RyX9vI+3cWcXkare9P2WyoL2rwJ8SWAtuUuxdF
AMwZq7kHUgZ0eVVvERjSb5MD8LiWlRj7hxQZb8cI0GeMpcXTjKf54XhJIcjmf43c
2MUpec9IyYydHimalr4lWxYl/NfHhd0h5QRzU9jrSga4ESFlmK5C6Qvhpemt9LHa
N6jcXpXbvab9uHbyBr4x66QVofUCupWX0gTMf9mickT/32x4adH/6tEUcoPPmw7y
wxZ6x6dW/sO5jOj+ChRRVfXUYj98Xvc3ruD2LEvYMBk7ivDUOuVI1A8890Kc6b82
viW39JZZLYVqaLqSH8spQyleq6Sdr1HCoWR7c72LkmoTWMewIMO8MvMyww11wLEB
rbQdp5G4YHc2gHCXocMDdDlcs8mr9qalZeAvVNY9gpHy6ULc51WusASg6cxL5yh3
eyFYSWMCRAmaTLD4/IT+z8cDqs++tNRYjaP8yxMKLOw9cFn3cr6h10vtTH7NuXHw
jSuA4TKmIbcvM3SmmQnkWJWgPuPmrj/nlWe2Rt8rTh8vt1ODl3lKU2ObPnpG9Uuj
WNqQU2GlJf0asgKDZtXhonoKE5faOE8JzrW6JnTMOonWqBs2dwLmvS7I4+2Ki3P2
lH0DPc/NzgSi1ElOFfLvnLnNZ8bMclcpxAc+gcmzme4yaOiTBLdujUrqJ1eRGSMU
vZS0YjHao/+Jh2l5jnmCCaKmqTk1fo/Qk9087jYKFRzZmvzpybCQb7pvWCymOoLF
eJwgsfEvMlItfYQ89y7hbC7XP/IQhHjz5ms+Dw9jEq/CAFfU7MWA5NE1w8wsRST6
sqsI7rdBV8ib0s/91MP4zqqOYXOwoqafqpInQmBPtUeTommkoYKckJ2q65J7WGzR
3XdMRfwKCf9b92Ze+mdVtzjrgJL11KDpHvLbST7T9/bgBTVdswpJxy7ltxgPdwQU
+3IR7+SZk7bmqGig9FmadCu4HdF2SQ/AKbaQ7/YwURT1XFmPbcu+RrJocOIHdBWb
h3ldrxzUL31gsZ4F0QTKLQRGFTj6sdZ1uFHf0sb+QBrDjhKtRpepLhyeOauR6sgx
CW7SgMofB7Glcw/FE3mckhvWeQTJ7LPZ3H4clFLgujdadirejl9FE4etav4mDaqF
5VsG2dwbygu0neuAzgd5jatkac6Q37A6aw7DB1UT0FqAdZzJYAnUGxco+rsWOcN9
cPN/cnF1bxHH9LphC7P0q5+fonn96vI0DnulK8YSIkjTXZk0hvO4i47YLasfDFv5
E4Wfr4DzzCGvSErDp1sz4IcX1qwWZCxWQ1g0Pxhza8U9XBdw8WZ6byzewvD7YOMI
6nCvYqD8VEEwjQP6k6n02YvKTub5NjseQNqs4GXR0qf3UA/bBUmpVD8F8ENU7PY7
e3iqhildS8w9UmvtJRUYrp9SwndbdHuLxzxo9rJfi5Xo4Nw162ZHDqOjIa0Cbf5Q
J774sm9IkhdWvytKu5MIaovazsCkbQ81A8hNf54ZEmn+mT8DRGvx38D7+asr4AkI
o9NEtI1s+jJEp7dFrxgS93ciYogzd9bGSZgJRMtdGiGFWdmYxKr8jdKV1dtqYOmL
DFmu6mNXCyLzNpAi4ypbij0oHNJcEalPUlfYR1kUU5ZmUD9o46fAVre4KIl5zNd6
C/laPgI4brLLQ1xQoXHqJatoq3qk8eMLU+mg50zx7ZUkF5Tz51aRAdE1hg7V893V
m1W19cAhKqTNjpUh9SUgpQ7zAeBNduW+IzqYtFb08gNdVQgTf1y1nHvhLk4mH6Al
i0vt7gO7bLyUp6NKS5Qv2fesFX5+nl2XKVEwSv5qc2n0ghUmHSHYlOX+ydye0G7n
un/72clKPET82jkYKiBldXUNmBLmXd2fVHLbE1yCXRWDQnlrOuegYq/dJs3NqPVi
jD+g0Ro3Q89n5+saH6GN+HfIt3/VAxThys4GXJ5Bw/w6u8ld65lQh+MsJT1dcfRz
VFlzuW0RHLejJ5z3TMMTgXHsRqme7Pff0dFdmA6BRo+DHvvKd13R9gofJEZ4RB/7
nZpdnlt967kA2Wua4KNE0+rh272sFvRUA6WWK16ScFqxTAJ64NuWqi/AKMJg32O0
0IU+56jHIi/1oUmAXyvJiTHocmRQar0AAFwY03xCwPPPP5cnhatmCPU1PLzxdbgm
5yUxsy/PW6f+zUDi6SgWy1pNYhEHmZrVek0q9rpBalxLKKMhxoJ8ysukZRjbanRP
wpf2Agg6uQ3EXWfcgDrn3ZfIQxey1scr37yqOnwGPZs5wSpshNRU6rbQFS3gFbKS
hcA5Q9OPAMXf09UoWfmJ7OZjG0+olCZvSuQhGkhSW85A7SYeLO/EYJUDkK5rQR7b
TamR/717F7OH1/0tIw3U+BfpmYL+jNgb8PUcBRCZWbo6KUcUz/0ivBTYxRs78Kxx
HuFL2ff9NzyrY4zfB/LqPxzK+60ywG+ohsg/QFW0AX4fIIbWV8jjkhtN2V35whUT
DOKPOhDdepH++6p762FTRpV5/0DqWpXOrIHxlXkzaeH/L3b9vkG3wgGWZXncIaIS
JksVdzysc95OnVTOmjQ89JpnBWGHJXYMDcf+2QqILJCu2GwnNN4YSnQvxOjZGe9v
VRdJy/sH8BSa/XpQJ3J4oNz8tPZ16uothzYMfdiTehd1jFaie7oiiRyynC9oLlfA
G0kI/QktRkBEdS3AVZ8aZfXsrExbtlo1Bz9dv8PrO8Rj211hA3J5HWN5HOZHc0FY
+RUDZV9QyzFY/GJg9Z/0SIYOllVSoI/EhjBoFEfLYkmUNRGv8o1zrbHjbNvau6Xe
K15JNo/riHrjWpQboTV1Vzk7QgspryE5a1whrTeciTpW09nnRNUk77efOagV3rU1
hh5sly+rar/hAlyPnR2owNN2oIrW+zzqElJqGsIipO7xXwtavmdPGWTYCxUluarB
y+iN0WW8XOTkfLXt3zAE8b1OMDXcQwzq0rvZPaTd12wDSegWtXytMaXgMQQ+5f/T
oM0iKX2sjzE6sJdQZkyzX4sZAYnddd2tkadxqSxfdgRntNv9feHi/8OWPHro6xMR
P/fSlNsgB4wFoNj/Lm4QKyy41dvuL4wwSIvfVJ2ikpA1vU3KassM0RNxRXNcZ5zO
OzYP5Vjq0z6kGSmWU1YxIl3/HYyDWbLR1UwcI6c/fv4fAEzIl5jSz66Skrl6roee
xlH1ojChcpB6hIs56oiQ5m5YWJmJlYru4b37OemVdF/HgsWM6cu+b0UHDNsicR/C
mH4Fl0LR/7mOxhbcg4eLU0OKmsQeHuP4rpM4jZUlW3DOJwWiKJOEkLKrm4hUD2x9
a4jzLzNIi9FPmAtP+OmgNSZyT04tXDHo/h5KdA/9cDPDEvAOlDGOD2QvTyahBki0
ReChNk5omJfjz6RLU1R6W3GwicbcqmIh2t3ZCQt8DEky+hJpC1RuPMliJGufVPFf
aGyzyfqIER/+RUZsEYe0HBuKKWzk8B1Aq2vs0vtLiSgfYn4vJ78VHkL1QZ+sUXEi
FERsDCBEi4dFNa8R2RXzVkha8pjJazPKgSuXUPkFPOOWqaV8nBIX7NrGVwXBdaLP
Fs7YFBC8cLQIt2XAaqlFBxjbAN0aR9ISXwTUSqvCl9mSoxGgGiFXvH1d7EA3ykWB
rVfQk1IiLFXfVLDh8aVwoEW98AsVw+naKhO2dok/QkNC56QyPO/GfdHc9hZ4gEPH
VdWhSdWCwutQxEQvSzrAZxD1RbLM4fZAZJ/GBC5JfDmW0HmUq1LYRMqRqArkJARP
X9aLni6xgOqP9EHXsxgfwuY9fx6sxssdZCXaPjq9djwbBVTI3JjfSxZvmqzsO4dh
PoN+FmMw07olbI16G7/HeGbCABsjCMbXyJ12EMVxyYUaTBboopBFhTQFLAGpioYN
1PAqiWOwdw2WE/IBr+7QJf0pF2pwpMosGcm1EXT+tWYsMG0v04vcjhyYT5Bs0Pio
cihqkeNI6jFbjYFVilv6LQaRaz4x903tyYYwAaPSddW+DiGDhtUD9rCqUoXjabIi
VhiMzIAtLjrpreqs8uc1DPbzKUKQqV9lZub7fOpWYKWVx+ws2NZV3b7CgJ+AnSHC
HFzlGTDpJLXRrWPW2rYaDvqnUjlYF8Xr9gX53FL2S8Jdol51SE1RSPHxF8+xCsWM
ViUeJ21pcz3mNjEaSiFiV0vKnYGM/do0UxEfMkSFf+UMCxjijsX/t6gb3juYcIoR
uzclAxdmiLD7kGUywH54QVofuZNbF+S2HOx6u/DMTxREcerlUbJdJOHWUQCk/h3p
GWd2z1MD96NGjtZ2yQ3TozMO5hLP5h/Fksb7I+3kWwISmyhh9a73VoQhDhybQ7Vk
Pf483BnTSfyDsSGixfeVUzGRuCcyWC2R+2zv/kW1yBn99jCZ8fdo3bH7+yOemeiF
nsUho/tHJ5dyMRg0CsKUi4F3fepYBkwTLwsnphNTA54pvItikHnIIfOEUSnFMe9V
0TiWUtH8oshnqy8IhFEikTaKPTxH8vmSfTLd1Mb+vytuR5h48mfqBYUCEDJrdsih
YU9qIDYKYfIw2dNXj5DNf9Ph0JuTjs1Izq+cg/Qa6v8LUSuklCzKcfPP77rSyeyy
a5pHAoHr/98KriBOM/YBwcR5sbXcUjbRUdvgaDcnbP/OQ7OAw3Fpbe1WVOYIhM0Q
HPPBt8U0OovBYd4muEIbofBQOHPdTtsXBkhqQ7alYl+RzleEz34NUbSU5y2di7ZO
k0o91nNUsmIkIcHdcNWX70EvJMzYzJk5VZHpV0227lSKMZXJwiNdF/fOEJ0rzDth
7X1Zzf0191JJQ/YMEy0zhwo5OXYVTOp9g9UgpV7+FK5zDD6Grdkf05JjcuVoGBWW
iK0thl50+GONDPocrhVCeiS5TaI38egI2Hw5jxEPa4ZiFTmG0DptfqHiWTFzKQNM
bqZYoVJwis710flif8gaaZ4CtdtPOjL4Pdj1k/rleABk2v+jLea21UpISLIUJwlY
fTNsEElbC0TizjgAdIGdljTE9AZ3NjdQiWRt4kfJC3x/OHJpmoMMzjFXYLrR+Ua1
5YeDcRRGz9BsE/acnStig5UqTehTbZ6Q6ob3+VdzxTwd7KDlR5kqlhfMQTW2pg4l
RwhTHFoKXd1aj9W6H5/ujCc5nbSYjLJky1LRWgcqg7Ws+ZHCuPDjlbaGZliwhhGf
5SbdfnphaqY9bkK55U3T/GrWWXzr7ETPU/Z8Gjr54Th9MC0uAwDnwHvr+FGEQQLg
73EAVC6cVUkmD7jUx2ELdJGdMwmQ5fJn24r7D+V+hK/bsa2z2CTUlAk8Mi8iNdZ0
XbAQjR340dVdZWTrNU7Ab9ibvdNqw9W9g+uyGhwj4T8RiiFF7qvsU/9IZE+hzbpe
LdBxXt9kosNi/KeWe7QF33ThabU9cF425dX1x0Wh0mUFZBr3+SpukAALX/ioq8HJ
YW4ALgknm3PouQcf3KkDNQvRc9x8GCzQt+tuzjXFkMPTfePm0ObpknVZCz1NALn6
0Eg/UhxYaAH8+OSDMZ7+KUMPaT063dyKljyAyW5m9xeCV9VNtDIDjY8mWpC52IfV
xbf3LJG3cnUuUW+xZeU9jLixtM3UVhuZc8ZN6uGDrh7uiSHITAQQQQ9Kx6Eqs/1j
XbvWmSY7pRqT3tJNjW5Jg5mS3L68Y8buZYwi96gPVcq51wVeCwbSmLOMy+yuV/vv
gvvPRQ3HasXtLcOHGWJiQzos/IaEPUNZWYqyrwRckjhH03agJqQgpJJQVUM95Xeo
0ocJxVleexboI62ovPPIYapw9ilBK4wBOSmSqPFfnHZbBQWNQVkv8GWhpZwO8Ytz
vH+2stJ3ikmClArdbN6fPHzmq/mpaoeYpb/LtwkfcgG/E7A/ljBzNzA+pjqb+r3L
lWdbsU/1K3ETz1KCl/ETZhjKI6C+vjI33vc0P7S/I2kZltpm6Hz2Vr5mWRa+t3qS
2ZlqPPu8A+GqHyIpb0cCrv1jfRd3IinK5FKJfStIakofVfKRwHT6Qltt40IPzJTs
kLIY9OFbWbgzUAyiV0i22LKeG+MOvtTQABV4ycA5fDJc6Ucus+lkbfD4gUWcfWJl
Gw8Vp/NgytOJEZb1HryZVAP0K7jXyUn64Qakan94azzFkvFr2/f0MmIDY4gZ+HSc
Aj+qdF//OSZt+cAwsvpzzstddAqE5cFHMKWvgCHEmb2rqeOx+oZoeLXijTIUlXSe
7MzthXaBR7GZp1gDOVFnRQtK6JMg0NAAyIaYmBLjKCo6DiihStpMCJFc6nJEIMDM
Lrh1k53OLo+KsVaXgxt26PRVpv3/KawoffFy9TxAKLJeVBNw7xShDuzTq2kEzPUr
P4bLrwJNox5fWJYjSqVCwziGVG2lBMvF0jLMVGFGw/fQ8X5rvUFum7QkLq2YIn4q
qmuB+FbEJN2XKfMAXKVLh8MTgzA1+xdJ+hPhucXcgvLLYgN4P66DzdLRVwcQ3Wyr
2nl0X3Mg0Dmb8VP7zKI4fu0m87xpdoSbweJXCFN1W9m9ujSijsDUkVsPIq5q7EHs
LXWHTk8P0ni3CytrYMQ4cCehAARNgXhv3S0wFKHrpuHa8G3qhAtTuyWdfqLH4aEh
vsbcRC8CKA9c0cnN5HhVp1HCF7u2UHy892+oXBUyiDSC8Qie4LCFYhxrm+nxySYV
/BvVZ9Uv1lphI/LWNgQ5bosiXW/TITIroux9gE7/R9Lfv/kexCm/tGhlv/zT77XJ
Kpplw50m0Q/94vF3txmA6VQJDCQSGnngtzsvFsxA/Y4cetJa9mW9qdxHOpNKMR76
U4PNk8G3Oyt/8OGm6P/NMZob2pyk27vpxbtgxKh7A2ZMzuLZfl47sBJ3u5evOknI
zJNGiiD4I0MM2Uk0eSCCV9sLiv/nWO5sxXEwmSd9BP4engYC3o7MEqgo2chmyNUz
UOYLQ1APlxVlC70887a3Bm82qFoV+HEqaqDIr8ml7bttpFppvvyCqAv2qofSKZEE
mNoppTOughB6HSGmFhptMhFrUg28Xl1eAhxrFe/zO6cUqn5xv2u8IWGJGFwOoBki
UVIX0bE7DscPeWHepwzjMBPJe7eIZCxXrpktsm0a9ZrlQtcHanUovzoIhXLEbal4
iyngXZAFom+FVgCFhbSOq44mWbAc77sXwl7PbrMkAfb5LNqwjBtt/GjOnKEUzz0q
W7pa1vk9mGTOcm950LdvijKJANq/V2gJxLWnvni7Ed7OZF2gZvu0QN/9hOI6iXZr
Wz5udqFjXnvyWYbT4UWZX511cVCuCLSf+nFtD1fiUYDw+8hTha/xWPstf/p36VfE
wKdj/ZOXUAdAjKyAXoedPFXIOSNqESd3d0xb9z38yesjsCR054CklteLkpxcadla
YL0+CdkLrxhIGttr8rF0NitCS+ZmUxuyNlJAayTXdDBoMJBYANJOa7R6duJhShOa
qIOZjCCcrGleMjaOIffFtSkGPWz1RGE7iCPlQA5XkWMf21C97cMg+Da0crsFE84G
PiiaDgcdA4lsmfYDLGWPSDaLk7vjZ9je3zofvVVvwC4MC6DMr2u1em6XSaqXPvcn
UkcPwddwJ341Vhj0xf52JS2s3iZI0V3jJ2Pzl0s0MPUN/qKHFAlnJLhZnVMl7omb
bSW1JZNF3SQCQPQBvG/jzgGKUcTgTkPkcQ45wkJCrgzPpRLosNFpwSAGI8jYGcDl
i7e+2FkScxEgOrALzptZQRlB/eHkJ4kkZVdoaGn22esZNmJ/GYoIRc6r5PYae68S
YiEV5pmPQJgIR0ca067P3iuW3ubxgNJX8Jrwi2CvcqBRlevnezShTbyjkrk6oBEE
9or1wU3YhipZ8yYraehqXFyQ0wDqDMFQvD5DETRwOPfhzU0H9zL9Ml0RBseaYvaw
TjU/YQGpP4hlAt35GsK2kHqrsZOmiizA6NVl/qD4F7r7bTUbp28JlpXblTvyG5rW
QRqZPTe9FALJ9PaqGVxO/phcRciaV+nNP1ihdPwVOsFv5+a6jfCgw9CWgUxHxgja
xt/Ec1+mTONffbJAFbVex0C2jnPFCh4nYcZekHo45Q931hy+HIgk6nvaSZ2DGdsD
FtS/sF9sqxdXGoZiWPObNWk0+z3HupUJzAZLDlI5s3nCngwc+mh4wM+rrdBNJQgt
b68lRVqU4YLaGZuDd7SnK5C0TWnyNLfIkHaQZnWjFzznOQf1ohsngpKWOGH3p3sh
lptgYQEze8eRljcI/YB5LaATEXE0VHCKeugfokohkobK6i5wZk+h2VJOUTQc2Tq+
HsxVEbRSWNDUp6AFho3xJzfHFIXu1muG9vBo01xZy5TEfRUbQqekdChVGyyk8j8y
lhEj+4xhgA/O2e0CF4tTdOUAyVPrQruc2ievXRHN6x3PRWy3QAvbLnoFcRo6EJ0E
DXVwH0OCn86HZXTg/5LdiVVasq446xPWTBE9mHaWkixPn9Ut11gNJ6hLxrTu8vxg
E7tA0znRCoNyUvpgUVcZyNhj7mWGnP5MIqVJcy9MjSgCLqwm2Jklpa09fEALHEjT
s35WZIfjTQQrZaAm7/4exd2052QV79qNIYZ1dywPUB3JoMilx6yZCTksd3661G2P
hd9+HCufCf0/mqwPH6E0IKVHSElst3Y4+OOh/6CgBUDGzBdyOxnNKqhganvW+7/M
aKXOUgtMQgXIaC7bykOMnw1UuvVo95dm3TOITZUFetQbyfimy5/r2ld6vwy7yXJ4
QAKiSeZ9bGDM/cxmBgJ55q7NCjfz5YNOmOB5OYRWwXOyI2Pxyl13q+oSR+1pjUe1
Q5iOW/H3UZ28DdW2XDQ+qxfx9KUHnLzsef2GnAXhSfTRfphtZXP5JoTCDnuS+MNK
jaYJS6h5NBGAaB6bWz2DN2SR13NLV2WavarbgzdNWbCJWYqVM1r58JuvKtBNyP9K
5UY3aD2SBt3lTBHLzBwWKrtBs95Y/Hov0+aA+At9LidXUCV5ec79Rvm1KnKRESmW
Iq6lSOwiaPRM/+AHQhZylidVaKJzTGjsR99llhBAE/3qCyWFN5I9+1MNj7+GPKzq
VPSC3zq/UvZldVSHym0/s7gc9TzU4hqCPhiO4ur6Ylsk54GemZbrqy8+93QJ3F8l
1PeDzjy0uuzyKofPdYOPTPIE3zxVbD9OqfI/H5aroiN6ePc55tcsglrXcfAO+bjb
ylaM1G8D2aZzhkDn7I/fnRbQxSD6UUqlublbUB6gEPzyYVrAMUKYG1PsDla/zA9b
dRu33IPfa4T17BHflX8kIYo4E5K9LgU2NT9+qZXog35odpvC9DKe034qHRj6szka
pBwYTIo1QGUsg6/Dgjc7ofBt8P1uXGN40AfUvCA4dVLPXqJ0YlS+4QZPwHwBlKiD
z42AztE/e8QUVfzA8OOgkk2Meqi5MggQmGBZNVdsu5B1uAJDRi5xFDGSkEMDWzWp
mQ579cxh7hrVFgk6SnbpSd4zajG0M4YIJ1w7NNJ+JK0vxo+VqF6rkPNJxdgun3QR
qDiT4su9aBh380E2S55kI7eulBd6VYGYHJC7daIOQZUnvFdPfc0rblZfPNmnFsjM
IJ9f2+ZAuZX8n+jMV1UvJKZBgnfeqTKqkGvQm8xNPwJzgEWN7E2RbPJaO387Harl
Ly3YQYSxGZfhri2FDhP92EyYvZOrr1QkC/IHv3AxKy0W6l8+wtRpgV5ZfLN6CV93
KU16xuNxcv4sp3eSSdwMhTHmZRXScTzk2jJGw84H+s8TgrkNrSUM5tjDkg6z5jQQ
OQvV+2vDqahkuGq7ijsWiLOFEBVa7ai00ipDRzkeVkyXGRMBq8JtyInfmOgzWE2T
hpDWdrxb/vM3zLmdA1hfBpE4Q1rIeRNx8+5CkYjrXHqKyzBLCiF1tsscIN6cS6zc
wWGYj4dibO/qDIKuwPyHMOk886QAWbIvWuW2osryOt0TMh4Jz8cQE58mIB9OrHpd
T9Zj2RW8SU/Nbr/5AYmcHtU7PK+EH96V6mJ1gUwMgOp/3E2F2ptgDJh/QwKLdvP7
+6ZowRITcF0yJtrHAXn116IouSqGur+D54qLemzeJU/01O+phvZlOlYASUoVdVnn
Ey2J2jOjEfBGs0X8Iuec25oT0WYX+rGRpok5WQserq1cOInehpZCL3vYBi1nHGAP
Kz/YF/rbRoIXPwlj8ThplKiRAG1meHXxaxr+Gg2wwVVT5+15ySas6lX9jLFpGkEd
8X02bxpkQaFDHB7kJQV62QPpUWNqxEzIVbJIAMWepU44Cp8qahlCuVNNz8clgdP+
PFBcLdHchH+KKHIrJECod76uo16nm5jm8vTz+e9yDYPt8KeRCZILDGulArBOBJyP
bGR31/HDezzwHlCCfs5VH2K4b6JI8/YPA77uprlaeoN4QdIPgfgLPV8zFGYz9l8F
IIysTyCn0ONBqUmPi8rTYW0gboQgFJ9G4qzKTX/h5pRiVmeBg4WxUPKgBacqowDG
ggyBPVF25slHrRA0WXYAJdwbxvjQXNk6D3Ims0OEzIu7L+ufirfw2LlwoJlCigFB
stGyepGqiaZyO8WoJAZ913/Z21aMmtaT2M3GkT4XVQxt3Y+4N/5fDWqhLPAwYbq3
pYjNZnfk80r42JTIWZWk/pEPswk6bvr7uDoWgkCmYACQEGj0p+EZH8WGK4O/D/d+
8xmc58xZtN5/TxbPfaFumlEFqXdWzlglIKg/jRwqbos1ITKhTLabyWOyIf3f+UC6
yONUaqjkXBVZq+Aav8KJOS8/Wz9i1SkL71zDwUnyDcUsQVhLgOWMOZFjjUVU02se
y1TgL79J3s7fVHCtj2gElHAkiIcsmEgRHsryR1xoJTq8YbTM3dden1kyUCigP2gL
5npQBUBlkBcSZiI/aMwi2RgFQelisMImym89QGCU92jtGNaajJ0KvZEqNAcEgK3W
mcmPEsrekzFENtj5nuXLpJi1zAHlnE3Jv+dXIiEXGSdDXCVrHUlhlYZLevWQp0AH
cjADC4s6jHEO9TWtC8/okEpnjFUB9keIjo4ImBAhpsiOdjZuYwLrJQriK3kZJw85
+4bL2HS4DcnRCC6pVjr5KV+jnSWUBbJDfgsrxlbQwaFbssdBz8cTaO1bjf87Xk5p
dhnQuCacvCXGBuZbIq+vhC1vHdmX0FqF0vM28nT5Hs6RYcDqwKNhRnpZpqveCK4B
BcfZtyas3JDLmjhE8OrQPIZ51cmC/dYnz3ngknJEDyeK+0PZLHXdrcG9p5Yexl0J
FRePSOLuGQ7PouAXeITQGMGPOU78dErvzrIpxnZyabN8r7vwkQTXzQZOQV6r3TFJ
46+cuIzD272RJDgSVGhRmKMdnTtISs+yQQCzGt3qD1vafv+lFY6Jyh4gvbTQQljb
LUurebH/Y8YSGqk+pEzjQHN0R/zpZ6K64yH+Qq+Rp22qqBzc/UyhShgR7JdsetWl
/H45XeUMFztiHG9tWYTstvbyXvUDa21IdJgeJy9pqI3Ihym8R9rqZk22zU2pUtrN
cSweptNt8vznFbkv3ctc5sEYF/p31CRp8s3128iSfXEEEyIsZLOIySQ7YEy8LRtA
XE40QiymJ6Il/cRpr0MHNy0Y0X8uFYuFwRo5k157H4+3oVEoWc26dVGnqvwxxDqg
2BtVLYhRz/Sb1Xoj4mFIa6nZpqGZzTMoiefg5ttlzIqVuebR3XyrSg78kpVfEPjV
0fmXFoov2OgGzChAy8qSwmO9zxM51Ngm+D91BewtM6ldyVa6T6pUdvQr5Gan2ps0
s3g+J3ACmXT38/Vbp7TEQLUdZVEsXkH5yngKCOdT6eNRh1QSHoIpxaQVPd6/qGb6
2/4H9WdQnH5rty9oMiqV7wSguN3ZM/yZdO2+B6h0+8irOjjrY1RV4sidEakvBd/k
P10uXvGRvtcBbScREU65FuLx9j2AXoJm27VQZpmFRSR7FkrSA9FU/AQ1gVfU72RE
AuAlPV7oBOGgM+Xz0ZXiwPb1ebrdPzeBwqHbGR9HiUreVPlN3FOS2dGFjLuy3kLa
mXs97g1twB/RUdHu9dPYhxqBSVXa4iBaKieceVKrloYiSnyBoM4idjAn7Fy8RfaB
e/W/UeFb9Z/5PDm4gvpzZCAWLK4nqy/3Z8232e/8GioCB9J3bif/VB/iv+uB0s/r
dh+26kvpZSAMFF9EQ9bXxKgOkWHc38ppuVLx7+LnQrGgpS2mqhCKAHnrAfOMeQMF
bzJEzZvFXdp1yrBC57AGLMejrFNWG29g7YG2Xwiy2OIpshf6wA6VrQN20UB8a2vb
4GDk6nMtDHH1EknYHambkpQyGxHVQA3HRUkpyasr9P/R3KXVITzIYpNLCFozwrrC
vD4d4oYtXJcaWkOq0Lm33X0krn60HNVxgq7PCyvEyaBIlAGC2Ko3XVmHplLmUrCX
Tb9kY7siTIuRmj5D01VS3/nr+EGmuLiM0aJGjImErRWkoqNBdLzeTITVNl8rfVub
DJkmJDo71si1njq7/jTZ0rBolBB4NuXTJeGc6F46vciqvrW8kQi9GVQoz3X6jPMr
VvbRluixhkoW7+tWpT3dAF9ZxvazbgWDwEz+wHwaKwUrDkFvgsVndiUHt0oVpQxr
VYZDDZGyuJG1GY27kzhm+NPrOrg35h5UKqpxG9n83ovuzOqgkBy9RkOaheRCiazM
hqNifQkHjWH33wujEp6AaZwuEi5cFIOmKrCYvugVMg2JPfy9W3WYq+9JPi68eQTD
r6Ae+MgXMqghQYkgAiQQWrDxh1P1WWfEjXhDa4YWyicYbrSgMJl/P8naKUmEij/f
GdnlKiFZ4TUqu49odOWyxL/GC3U/A8qW1EoOevtye3QNfLP9bZ113hYYrVXl594c
YzSOQPQ38qMIqDsir1GRsyJhk8TI+bOWO5K1VquYgWV10BYMSp98aZyodZWoVD1y
1japN825iMSGtKzk5GA64E6fhqQidH4/Xd39egcNvxwKr1HGmiNnrW23gi/ybst6
L0FQnRZS9MxotJLjw8riWCCXvH2NQNmN1T17xIh/fAmcrXRAOLYr7f2BlgONHDfh
EnwpKmec0YSYBwPs0yRhn8x9Pbh6jsDWF8hP4imeczZbjYcAbXyBJeJtbI1AHa6t
lvzre/9P+hInTaXBGFaHM0+yxPKAw/0RC5VEO0O00U1s9i164Rk0nOR+FyZiUt7V
sz6Xj1kb6n4SxgPLykXNcBQrosODwcDQLzp32j6ScPL9qXQ8i5484GznOM87Dw5V
raCTitYYRb+nVjH6CoZZZfRrDMZ/udrbRwA5JelEy5iw5YZSfDfQq53cTa1few87
6jl4RZW6GWez22fKx1U1o4Z52TeqgdmxRIOyunaDRuApcgIT8+/rPNaiYFtoIHuO
HpP/3UA2K2PjHDa+GLijFv2VRmIpNQYMKIL4wTZnjMrROmbWw/AlECt/MV7SNYUV
UH0yG6/t3QQ7c6rb+Ml9WoZGex5TVnB43yHe9Z8+/F5EPhmcpiSM+3iQDtQiGpBh
8JGOWWhow9xC20vvINzb0Kb19Xm2ZFcKuq4xzO8i5DNS+QU5052ag3Ub+OgCab1v
bpI3x3q/9452q25ocik0pI4XL7kwsNy2hyEB9e/Pm56MAhMEB56FqTaJDHcGcVpU
qrRWSb6qPj196vusFsLH7jtXe6nhNgGobP/pAMTVK5lrlFoEeIC0RktyqyjPRv9d
7yAshi8qPDXTARufVrZzbW33JoCDlXrn+KHRveF6y3S3j14GdiQmvL9JhP7bGpxI
XzdhBxvmyPkQhZV3l6z5W19fdlDctKbTFu9xBBL7GiVsFQq6lJX4ZbpJX301Xp23
GD7DlERszQHSxRhJYwZyZ0/ofUfA9yb7afXq8tbspu8G2rzD1PI8gujGCCL1IAZy
pTttWkm3cgFiBtIqLhmomeDx2XmVa7Ueo4P+6oBw2pt3NjPw7NT1Pdtsc+ltBC6z
qhVYjR7a1tVxE6jt7vnvpJ0jL80A2aoPYifLjW2hyyPcw7SOGTmt7blbkRGq6zPN
k6v0Vq7AuklJSLn1EVVVEKyzR0OPBuJoMUwffgciBkq+Xyp6PGslAVw1iC9l1oMB
AcuPMiYhYmkjB7zbZjq3fLgVfyHwvRP12qc4Oj9sVJgwuh/cVjwQWj8nU40MzFFB
Cgx/sfByaLcmiVEEwpeOQWvtltU2ooqBvEAK1OKVDWSpmgNm8RrjhyIT7y7jvusp
mYyv+eOYUqhU4PItGe5DDQa4wgoWGLkCUcvvEn8IIrl1V3/HrgotY0lQPqn4Ejfr
NL0NaFEUL5q9OJQHsLDljoouZyapvq2YPpPaiDpE51HLgk0eEFZffdKz6D0gq0LF
kWqAp5tVC+9JmrVflWjRfGduh4IUoRRpn0k6Tj6AGAiAsCPBB7NWmRF0yNOp35xm
DqLDTRpbZXt65N7ee3Fj4hMDPHzxmcr4Ap6a8tfebq+F31MIo9DLeQqZTal0zCoF
ySIXbfESP3xXjYpYhbDeZ9FFwyl8FpU8DV8jvPqzw5xqMZZslIIPsNx+2qdcgMoX
ajq922LnPmkt0uzroUp1v5HWulQZrNspv2Q47qpSPD3oL5OsKtckMP78m8IRoUAM
de1+iYKSK0cNKXHjwBodOVgLDmoKChlEHVzU0CXbe9jplRjQ1aUSIGegLr8+JKnU
q5d1m7dya7iptUqCWBwRIa/6MSkvi9SSEy2vm14f11uAVI/SUjlxrRZbjunPaiFQ
WyAfR3MG4DM5cMBaCojUiN5KsVAvCfkhKK6xrYRy0P1kxIqF0lIfbdbtVXRf9i6w
slNN1AiX8V8hqMoNTLfh0iwC0+QR8XMWEZPPAtVDFYQrwW1f4pl0iYBdR41gBq8I
xnIex/h2oAoKtnK9JUmwwRZUgnIuBa1Y7FYS2zln0pbwcc13EwcPIFJfpu3838Ty
UgVDeuLb8WX7QbtTb+o5CIAXwhqbTexl/raJRawZuHwvBsPrt9XPcSxfKyqZzvqq
9Q2TPtKf5d9MtzKbk7fqOZpcviI6C3V4E8XcMksg+Nnn35X/xk9vbJ3vBttC7CYR
PJBsw612HVVAAn50IBbKqO2c/V//9+t/KJFlSEhubWqm4++534RBFs2HruRZY24p
oku+yUgeFVGqgmEZExDrTPOQWXKcZrqh3fkQKYaP9DFmtnBB7Knv/4tsioDjuI84
10pGUYe0/DhciHl0hvKUCWjF7NMukAChPEQ9S1EqztCjq1RalLreLUVPxoaOI3qY
b13d8YJWDJwSmacZyb9UYcQh7Cr6AFqA3/r4I4Fb/8JZLoW9kzbfZyijXOcuzZ0o
uDKcD6haf3DrqQoN8Ayn1bIzxNY838mebkrJp0xZ2QmCHNMiO4oxpU1P9ndB/b2P
IwjTRxUg6sqUXsF9bkhz4ftsfNCv34zO06mkaQu6O0wl/pOxIuqfA507ypfoQten
9TqqCQWl79V1St76UNBux16MlSvOzyx2VopeOU4QrWU3M6bllET9G8FGVvzQzh26
5FCn889fN29ca8Axf2cNUdHz2OU/MRUI3ZmgQpshgcJwAfL5y3e2k22PDAV2GjKu
LO3TyEmv9FL7F4xQfeFaLOSqXnORZkTltqt2fJHRrjM5IGJc/H3trM6zDMiCI6Kc
oxUyz6XaE9wswUA7U+U9hnI2Yp8PrZg5Ec7BFKi8vcvccDjk2wdbz3NBfHihuw+q
tJvGfYWE2hoY1iKDNha9j5WRh2AsZCC6u6HfeFcR9K7sXodo+tQYWiknRNVC4Wn/
dsfV/uBjiCMAfvodJGABLA03nnUFpbLwl8gem9LSaoFHwL++xvX8WVZeIBBY60bX
SNpQjzesi97gBblS0/7hJMa6CXeU6dj+96T5Od9jlb4wJT7Z6doiSuYOhNhQci2A
2mSyAEfimT+Y3UEIIhvMjmJP8cfZ8xTVbOxrMkgRmj+kdGBmIB9Lp5+7HKgnfCoA
GeYq3OBSRZ0mm+U/+I/algJKmCTweo96I2n4KZV07fqCOIfBoVOj89mP3vH7d7bv
/cfrVkFg6DeVCtlW+V4fHMpwSGOw3gWnMIfDZlP44Id0TJO+8qKgV3bgp2Wd56My
H3FhFnJ8y5FLIdAaBIoD1Jw479+SXRayAaT4HgG+LKhgKfNtphgLAh1sHlgXK1d5
yT+HAV+kXeEj3GlUWSNxooZ89T1hi2G4rgzNZbsPsIxuc5m4qJb0Uc4Q6Si+7NQA
VGKIojY2nnU35jK0A0FFA7QZJouUAdGfKrZTbct+E0y1wmff0OBFci7vbD4PEQqt
6MeY5HEccSObksL9y4dqqrQF2RrYu6mo4BaIIaPuGAgkZUKTWMk3mfEosDb+iA2e
zC8KIBn7P/1dP9VCgco89K3W9izSWXkTfeyCoIshUgUxJeFXW6gu4v8C6R8n8c8a
3+lj+K+W0x90L9JNPwE1J21CvClgobw/4xfYQ4RYAXImC4yfDb+tMN8OywDBTrpi
Qoquv1dB9sEgW920AFyy5Vprm8UJ0uZiVb23HZVDIAzojT5Bsn9/nQOPwQvhnejY
r+ozWHkrsRxMb8F5qQ3Xy7PwB+rO5Ych8FW3gw+zGYl9kW/vLM/Kwrmy1q62Tcsl
GveWAlU67JQAbBMh93+2egOU59WcQ6UC9iZ5w/3yR/s0CHjRJWolVO+kc+xGD4Ez
6X8WOznd+F/VOSZtEYHXvVmQslX+yeL3i8SHzjovrw7IwImDAitS/CmgqBbntMWt
3+o3kK0k/8gvVjRHPVniYCG53uPdSiLELKii2Wq/KDPFKnU35K7rPw3Y+H9nF5F0
VmaummdBNlyW3hebVTdLYKBkm4Bkf9dGH6Nv5ksXUuUIPaCz9oZWLqcRpjXombgG
sZ4mItrQt/9rsGw86NaeexJmPfwejT1vuUdyliiCpOcD/RcGCUF3PMudZdQ9h+X0
2ugH2A4Yy1OV6spdLU3piP+VRS48P5KU168VwTLzomOhlaLngLcwa28I4dHhndpA
TnIEx1TtQdWDwJa4rOSrHZBfNQ3odPZCRMU5ifmMOphYxXjLGVg6luUAQ8q4n08E
c4L1a1TDmbB+78xAegxER+j8ZFUJDDeBk+2qeEawKUWg7+22/TI6Q2cIsf5Yrkit
TqZ7JQfhOOdIUQLDeYAjowagZ8Qn/NLtnxvkumNXvgsNaXL0Z4nMOfAPMZxznl/h
PemPepBKX53CcLx7UkKth2cSLG/SmKiyjjyl9FmyHzfWRhufjw4SNEyW0/Yty4Eo
PAfBB6WCmxSA9MNOCK2APnsMzFHI6IY1JIWJpR3sOZeLd2kvCQqJD51bJWQWNNk3
CYNtJ91Rr8+dUhyTGaGOU1EeAis1YddaSNAhX61PcyBM6FQhK/rZQN5jx0irgKRf
7rk7Qr31hWeCiB0QPwT9/2fnnWrTqBFdLcdCYYXUQhYvtiXlvyKbXo6x74EabDO+
GwEWXiRBhhYUyReNhQUs7a0hfzGSiIpcjsXqTXwhMlFjUAHpawmcszuT/x1iwxg9
SmbOqnOUAKhEzuV1TDo7AlcAEiGW6r26VZyCKSCtgnFP+LZs2i0OXKWsE80019UU
+ZpQcncbxVYrFjEdaFZkd/qDy8G4O/aI2vDmdJckUxQUj67Xe4LNzxNhrADuWynv
ZvBwo9vpLLVS5SfUIzvLRH4SVvL/DVrB+HMUbnhoI9hVqjYezhnGTIassb11byhR
wisKngxZx8vBBxiZukhgqFE3ttItSxg2SVdzhM/d40VTSHd+Zu4df3LR7ip4g1C4
ucA7i/c8BoP7xObcl6fnPcAc3mBjN9BgsF/38/2nGKbxlw6rT3yKgDNVUazHlTN7
/G8iySUfWsIbc/s+CRvGi1UWvZqOJ7U08zgO33rtYmOeNVB1JblpgDTg/C6Yn1aX
qTCfH9vTOvPDqs/+NvPQMfAamQ7hDjkO9RpLGTpJ/XMgiiV+bTJZA4lgZNQrAACo
kmf/rg7gkPpFD1fEMH+RKMuC7xlvYXGs3Gp2ef5fDgAZQ3hVKrEJMBqTdpPbpmbg
TuhfkMIf8ssjEvzp3bZum4iLHK4izZ/IknWOiEg1MhAQLP5+82fhOSHHkuOOzzPU
YPHP9taU0nnSB5nhUK0HenzXtlC9YOLAowJr26pz1QQjf6fAjy92z6IgKB2CV5hD
9PhLIxDhPZM9N9vwb9TtJkONRz/Jh5Z9gAIb0L7wiMYM0eOk4sW2wuGKCcQc//eA
enwaTVtyDyymfqLQLiQ+3rYZEPwnljdMNFrcW8oVUMEXuE+awrcuIvvgJP1ujRxU
N8p8C8JssShsNFZ+d+xS+7YYKT7kn5zv0QFMgE3dqlajV/zO79uLjw9ey2sTC2Q7
PM6K/onVMoM0RaphqHUFP6AJW3C7n1FuG0J94sOPP2PBKkWxquSNPt9ObjDY6VM1
FOPZDnYFV5R8FL5/EDdaQgUV5MaLZP+jOArkoB/OhOeCTaGs3wpWiOcc7VSXyai3
000pzHOeBmJJDbREybxLHh+NCCO+zqpSJ+6M0HtXPP07dJnePOJoRs1cZn3L1nXe
XK5VRe1vmxBJUtxf8aMELecEtu7YNDiEX2T2w1egpNbgq7xlK1bp95wJr7F0B1qy
UMk7VMp+o/XgoYjVQyhXHmyXXsLTRYYbckan7JV7aM5TsPqlc90dy6nghm55sxrL
R9PlHi3b8MQQBpqCIcgzgGHDE/5FHWobHsZ/D3edRkJuABY1/KJ01VXr5SBFneiM
u8p3VjFsP4afY4fRjWpr2YGLU/gUVEVhvzyfewZd8vAIyuz5CrU1T/rtsGwvn0aH
+3dfKJuPGmqX9XPfIBhnI0ZSFtrPGGTY531FYIHZ95NkQ2ai1Q4HGiSygWFX1T7J
vXG+JSxp4Tb47pFZEkGLU3NSbbj5zifoK0A2dGcpYDuu2oMKHzXAPRY7iJwCZvm6
mV+P9zeweFRpyvnOPni2H266eUeZGkq3xKkJn1i23sXdxGSIdIgDRW4JA2NzMeeM
0t9JsjVGiHheoBSwMIzMfCtOKAeGaP7oBjM/Y5GjcDEolGlhvo/Oun7EGen9UZ4v
vQVUxGFhSd+Sx1gJT8mQdF1eEj7eYq4UtGeyKkUukodF2ZNY1sbsfpKhuPqwDECy
R3PvR2PRAaCanIPNsE37R/IWXSDdEtgNlrqY4lfYNwkKPSk9b5Ip+0x95+l99Hdv
7+150FdHfsgwkkvBtXvNXi3Ebr3AcxKc4g4AgGp1TB1JwVmtPCddqO1cbHXoWQoU
jh1kkd7mkWNNC5wOBuBvLKjvQ+3u4l3f4vbhGFhEK/rIDgF0xszCvoEKu+CEf3ZD
/ljtu2ZuYB1K2jxuOS53JAaG+VqdpO5TWVQKDMEMmnZ/ux4wcCW3QEZ9FxRZ9zu/
fXXPOQwjG2zzRfGpSaPFHUhjcdH9h9n9yHiGdr4t+O3vIVTzjhbnjB48SINFkcLV
dJqQTUQ34CmGRzf4PDtAkiljTDb3r4GSBwNI4o8u7zHKwjq5eth2+kNOSIqwb+fm
UE+Mh41axPGW3DDl5uvorQgTaWYF6a+6XvGDZH4o89IcYGzvDz44nkX1R3zKkXnY
8YJ1/dwhhmPCkIgAaSQjPxHiwFrtqJaSDAJw7LWLn5WeYfysqxa8+FyIxXPUuZLq
hlmHC2MsB4EH5pMKJ758egXmXsCyLq9teEjmKnvexOTRfGrRDPPqOBXHonUvK8jF
wKjn0DGoca6EhEhnTWLnfMxMdXKyv//6uTiKn8jVDkZjCTsNRwxeLgk5b7p8wj41
wzsR6OfIXk+WpT92r/xceGSiKdVDiWp5bJARWk1TEM3Udwwr13aE7Npm0QuzGysd
ynm6f4F3lEdx/El6VL1GfSsavzwTwUyb9+kHUr1L5Kb/jDtIERF/UoopdWC9XAwF
937Z5B1oa69GCqbQdSIhsfsbdRxC5Z2JlFc4uAIR8vgueqo34CIGaP5BJ/FGseHJ
hPmIOsMwXaP9Qo9m/x3xWNr/pB9R73Gm80QFazLmkRr5exoRpdKV+nnlkocfbMYA
F1E8U0jGaNvG8KPgIEWa63UC+n0K6OEFs8eTyI20f1gz2MXt8oE3RfzlW+6Ojqff
MmxbhgbFamiPMLT0cB9IggPQ6MhD8vj2pRfk554v3UZVYlYscOT9gUi34DXfkQ4I
uvqauw7slQB7ZUEYr/PD7fThmcATxUkraWaZHg3RzWIJ7YOVSWR8OLBvHvK6pWBB
6YyIf41vC5Wy1oZp9jAaZjrndlijp0ZN5dakuZjAkPKuZagABztO07S9WUzJU9r5
HK9lPfFVLVl+EYZRG+7vOZPdKOxn1ahT8R/Kt2Qzyv7yWe8Ln+fomdkzyCkzDiZt
dLfKawVKBvryKgVvH0Id4C0ehvwF6TWnD3mjVt8M7/rF8i9oRKenkIfEzAfgjU4O
6WnDS3rbLpcvgSNSxRtTgoaaHzdDu/H3jEIUVNDqAscP2Ejkt+LvqXylxOcLXHq+
mJToBdsfyrPkTKGU2/00ioUiwOSap8vWOcWyvl0VdhFwIsyAXLN9NldOz9WNQKBO
BtIJIChrWiXo1iEip+Blp3NZRCKr+5lafm+w/Y0HEjHOfIvuqXl/caz8iBlTKIov
uHDdQ/U2Jpe4IAcZ+ThWkriLPabbt1Oi1Ze6OecNTNtNyMGAm2b6YWttNbwSMkQX
DUb+hYJKAtAixSt7JFJ6pKYxYRq2WeUWmPaeLCBpxFEDkDNfqI8OmiWko3Kw8k3j
6w61LKnGx6cc6HlBt0IEMluFIXHeyRfvsigEBF1g8jra2UNNaXMaNvrk7SSNzzvs
G3VB4v2SmUhLMB2TnZZQoM/c+A4pPnp29BXMY76ZTgXPUMvUrjK1gtWB/C6yy7Ri
adIcW/aBV0TBMXjFzL9r2PSsASFgBClI6godm8BBGHaXLZhyhD85AGXsuXB1liDm
fbeZWD57K4Cz4xPA7YjmrmeirGTKmspxYqr8iFiddQPjThbbPB4tXAQzM96RnEnY
BUr/T2mFQisWC/wROXfFV5P9MXn4wuKcl9ZLxRxfXP6xSFb7p0G2GyknmAuxvIJp
od5z8ZBgnKxOBjT6RR8BLGXSNqNYxMVWtiSgsXbojQt7D9rL22lhlOdyjljNCZLE
2FEf7UVv/TMltUA+4odwUrBF6jZJF675LUXQVq5pZf5V8gcI3AC9uv7ci3gEqiH9
4uTp6T9Bg3unl5sVxK3JbnowjJdSCBHwe65N5lWG1fmy5DUmA+h8MZ5WQR2vG/WC
U+vtLlmjHG4NNa8wDOwk9Dmn/Z9MXYoDREDvzGBMgBZDcIiL8IQiCwH1aMYw0jCa
P5SDzRrfD4yk6TxKtCT81LZ/bMP50ke6o3W0q9HHp1WvNHXHlBuFJwetvrOoGqak
U7S8LTF3e5ng6zJurvtjP8VZQERyegFc54xwXlxmTB4d3QPeNofF8ZPU7MWZl9Dr
LJsdyQcPa3rfOb6FSmjdcH2wRm2SDi1KK1YUCXiad+IH94F82/yL8NcuQNr4fZTf
AFEnU4x/oiyMgGeMd6OXRhXqVQ7fj3LbB63KoonMJSGWoLkZnaJHyk6/3YVNG2bA
QHLrZa4ckX2rm635JivWTKClBf8g8liRMLYjYzfRR+j9wdRdOpmLvhzV3F//f3os
GPGmP6QU0BMznNo/qf3Y7K8nwDLvVjS3UALdHw1raIwrJ/HHe2FxJ6jAhjcc3Wjv
mNSUHZJSpRwUR254DBs6kCMBvk6BQymVNHMAh3UMvv4lNFn2T0TVtBeXgsMKwGJc
PnrPf9vZArQrCOvKWDOAXbChhco/sEXjC+TKiV05OTGX7oPdHYqOMYfAAfhyZOsy
hAdb9CsWIAPEtbvrPH6R2DDVIxy1VeGODB9LnSqIFpNzpIGeIQ3kJhLTYttTbses
pZyjMfSdoWewLdFYNd5b1WQkoOuVZ7PS4Ya/6Wpd+/2tIHmAcNmJTncRm7pq4CAE
8fgMtWCG+hFOq8D0oNTJsgBF0guGQ1TCmM8ZUoFtHw7dvqT/77UFoRf5OiQJdzQ+
nRGfPBf2WDS2/3J02TjKxT9tDpdCw/GVUYvDhJWSBUDx3A3YyNuNcWMKzJvAc4Hj
CYYzJEZ3uVEkxr24Wg5crSj/UrcpQf6GHWWW2tb3e7xpyAPBO7OAZllxyHH3rq3U
rLlG3vyoGTlyNXOsVZfJFEK+RIThkajQbGeX5YhUQ9rt0ihVMjWmRCR/z6UJw2Ab
zdWKQh5W9cNznxrN62CodaUY5XhvzTx6l0vk8mZ6oCbMG4aGM3SLVzQ5HEE9Tu8i
xCjpSloBbsCgEpyHW9DCm0+KkhMFTTK6np9Ba2xUb4MJ4+PEKTQn0E88qXQVqlY+
YFXQOaqVDwSfsDs88MK66h8xcdehJsynKrKO/7w4xhA68MPDZMkG6WhfiU2Q0cIH
6cmDX5S6FOZqzeYLoNWbKa3TJPslPoT8KM0hrrOpw0p9pMT+NFz8i6WG3CdsSqJL
uT3hKjNkS5QL7ZdDFjSH6NajDDKmQhzM0fV5fyTQKoIAdGAxE8n3PRmn0oi+eoUr
5RBOOFSRGjA8ELKQ2YB52pLEzljqE6hfC57L6FqFCjpqdxeDZaI23oHxejmkJhah
+thXwm1BI27M2oc2h7OMwQ2ixQ57DzWNq1DQy2G3RpP3jgJK3TZAYgqm4PRti5Hx
dEDRPoQjuo305tTnt0Ui9fcgA2Bco8hz/we+c9yTWZjtMH96zybST5kJo4Gza/sd
zP8XlHFDloAGChtVj1dk5rr+qf79VHW1i+hRrmn8c2xsQEEisA5IM7DCJ7D9XE0+
cHZAq8NG75CJKN9goKiAAUsJU4bz5AjvmH4zSLy/gD7N7MsGA1Y0osPhVHNd41q+
xr8B375W1SyHw4f5KgEqpJKhZuchNZmhRHqkuO1qPwCZ2jmIb6mY7OcBHa8+yMTL
2cWmTSxOYaycogm8j+ZAj6XeFgQCZpvl29y5iIdLncAgHPlmlnBzDqcDeuw2cy7d
UqYd30MswildOvpPDm8Zroq9eUQ9P9O7NixDViGewKSFiVHHMnj0+1S0L6puKVDN
wXy/mBZH8Enc/J7+vlBldeiv1bFy+zEfbpcPE2X12gjQdLmI0uKbjlG4KDUjXmVk
rdWh4GgVsQd59j/a9b4pKM74A/O/LiNlzr6l/OjbcwaM+2Fospvjxha7op3Mp/kM
0AzAp22pu1Q0uAowlT7THatU2x302ZVcEY5KnYDvmZzu3IHGtKU6spAqMIJwr2Al
4LRXBOssZQuV5yGw0TCPSmLNy7uMI5Fabg1MewSeEp4z0M3DExTJdSURFDOSEArX
nwe4/LkGO7z98ozaBoCm3ir+1aBeGlx2TnPQXsWdI8lcNSOcziFG1ypEdLv+7CzE
Y2fT2JkHcKnFYIl9/nnWHllbYotVHf+DCWZMoPsFTgUK/Hn9S0yAnxXCi0Ctlour
9DrkjDCP+Xrdyj3VQ0S3kJ29r8BdLQlFCYXxBuH0mDBPvMJsKkdl65pR0Ig2onB8
xIdCzA/vB9x6e46Rhyvryvj6aTZvYMb8yBuHS+OI8AjvB0S6Lzgqv0t8N13lacRC
kzXgpmzSmvra4ECn06X2OVpl50nBt+z6fIEVhvdUZEdr0Ounzi4bOZGfYXCYtxID
dy2lttwQHM5lOISGxoIe23hGQdkCtmd2jQGYS5Y30WkjDIRk5VEX15zGiRGB6k6Q
/wHpa9sHsk6DeqVR8mgfWLDEHOseh+5OxMO0Aqcph3sv27gRcZC0PIs2Y0iPJ4U5
qRDJb+zSCs2bWTL7vFB29s2MmLrHN7x/iq0pLO/1qp3lpI/tv81/KRKmXu9OOE2z
6t8Bfn94MZBfx4vCbwoWlr5UTZjRn05le6Ffvsz1hSz5KD4Qj42WQhq34EFQgvb+
p1n4RlSH5UJ15l7OO3arMkzoDnrI3EtXDTmb2+cTR5I3XiYaHKcsMHvP5ykg0PE8
YHZBQgAlFjZmAv2ZD1pZwNFwdWug7F5ysg5eWXPODz2gAND5WFEJdlbIX69sE+qm
Wx0dMjz5699vIdVi+LMjoP8r3U1qHb9pDTldaQgbZSV9KDHeOYcnZr0r5j6NXRu7
z5dGA1pWF8G55Z6I9rb1/rc40X8zKJ+jny7/o7KeJn+rKNvRYYspCRFQyosB20th
AXJWZCFheheAANIXeKr+N4Jy82WBIcfxkij8W0c1kl7vUFbGv3Nk5dytp66ccW5o
WNem9G+SDvJTxUJH1VkaFfzjrlF7ftWw9OzjxerzUjhXi/GJTew6qGcsj1oe/mac
ZakAbMCMx1ajVvGz8k52RG34aGb7EBDSwGOTry21jUfPqmMQU7cE9htQvFTGfFja
ep8v1NYbM53oADt8+W+A2G1COfoP1jOuoW7W9De4n1m3FMcq+il26X9NLyuxnAwR
CTFTRsja4eShS/mYawm+I99YoEzqr1Ee5rHlsyrfpe0iDTahHcxQ+cEMXeJko2p1
JJEDRIO4/JuRsK7kjLt90IeInZoMjizXGobBvUtnWpewy9dZijZYQwMShjGdv0e7
BxTDVTpNLE7TSSgtsqr0TlUFqDliCy4nQKEZlZeCKPVRLG5KfJcxi+yaJ7pHrm+j
BnJTCLwSoZYbUOJTNh0+uHnIYErrCwC2Xhg6t8Jq3xzW2uW4CL5xCdDNFewuFLH2
MpjAPnHeZD/fJX6ga5Ycf5IBtHDzYr5f8yBsnohDiqwsPlCtAcFgz4WWLoCSGeSK
OTGqsqvKyCi0jwVHiR12s2y+DfeerkeSll8AI7AcwPfn1tKVOsnL70oI1c5RG0+M
VUlDYYypV/DVcqRnMVk/fQdHfMa28qaBggcz7qPXoI50HcJYaCazPCOh6n2qlwGU
PYT1oaDOmbvjH0FXXL12KCDoTiF4ck3G/O2g2m26dmcjNjZQAvjwAn/Oun178Q8W
vKPrpWN3f1QBIHaN3ZgmfaVVM2pYi5bwSUIHd6c+Dwn1XNGkGjHq/wspFwv5xePx
ovXbqKR5pl61zgXmAszu1CTkqAEN6LtEfwwIvJWQkK7t0T73oyvRV9WwZRnlMSj3
fZTvSoU5OaP2+aHLN05PNi3xh/RSvqv5Akq+Lhe79ngeCiqN+ccN15ClAgILQwzb
ev2hHj4Y4zFMGFcgaSuihLX9vDz6Nw+/66+GcvnpK6TXjWMdOZCA9LnhXPlguAJT
r4JSnU4KAhSNXEmY4XigQHHhjvMQRZsYpiayFLVfbpZaLdZW3l2oSYf8Jj8Rv+hQ
GoUImC7F+w1NBEu/GBCz8FfKQ3dMUONMTzLQl/WwKmcoLmvgcB+19smzS05AW5Np
SZjYbd1Y1T7pJlO2rBkLTzliB959QmaC0TUnGx8gAI04wxjy962UDQOLO5f6Ff9J
Ba8KBveG5sv+Dia7LwzXjLjQu9vpZ/PwcJOiEwoStuNJE/mM8/zmbaToHr76N3nC
hsbsRvTThxU2t0fWsSv+JgMh7HOnaLz/Lm6MV/j+nk6S0PZiUpdkBXPgFe2Szb/g
8iaOJtSR0lvUMecOIlyUlizTlu2bEj0GEztod06knsM5xuYobMCg/rtNNyJrLC9K
oZ+zxPYnpOE8oU0Qt1Jc6+a3nGE3CgYYGNBB6qKmtq95kA0hrlSlUYMg8yrNs/xO
34WDK4FL/b4MWNHRb76prMd+1hhONRMeYjwdQeKn/wKHhCwUWuu+mwXTcvyLMU2h
Xb4iDUeK8Ps+zpXad4LLoH6+gzOs6x0k2+ckbTIHWxkd3GGJ485n6Z32OxqaIeix
FIEHQuuYIb7bGttVYNrLKl6gt+7IOgqn3B5n7TNhKsgcBtw3BR+YPMxeQfAgNd7Q
jrCxnxQ5TQXj3axi+QiUpO+prrcX8B4dumRL3kB7+lNMYMM1tT4OSoGnjSHLH2aC
8fDZ2CT4p6smNXL51OAgu8dCJeJA5Fkx3nAj61opJjMCii5XVri9eJTYjhZ0/FPq
MhgguMBimz8OHwh2+Tx7VoLdc3cKafG3KAZDIeChxXeyXxmf3nzy2URUiomsrgyH
Oh8xBlkexmKSMq4C78Iow01sq9WeMf062bU0WtoGttG6CRGeuTgCuUuajbwfjGib
kU6AMVPiY3+UlK5B2ZpZnbZFpqlaZTJD8QNtwgpGRiJGJ3VI5I4ruSd0aJgNZ49X
5rAMumfYQUU2HE0S6KhdGSIDFORb7eO5v9LVI0oAjkP2YiHPX7iM1fTq/6L2u4CU
q7M8iAT7BuSBnQHXf4aWUkT6pLyjsPcOe6YsZy9SYWpdAKD1ZgAx+t7Wm7NFjJlg
MWgSmWR0/vaJxcOlZc/P3eWNcreRkmQDPRRSaTFt8bQkO0Qox3P3bmpUROGvOdSK
wX3FdE9YWuyrTyrZRof6nrZAv/xHkV/J57+eSk80Xz66I191SwC+a8FNTQ/Cnl0s
IgVsubIMEqlSRVtds9dBqTCw/F2Mos+JQnENX3/lwbBdyxMqy5oX9qMK6GiXtwen
y0wcmdPtM328uez45CJD0EWubrmO9PgpNvTI8scWKExfNuoS5vZvmcmlUqQz9df4
viKhejXzqJDXpwAk9GarGtRSsF7r7YNcwrX3JlykojCu1G4xYy6+mBT27wBR31Pf
SnRuEv6dUCwayDE+qlKowl3kKJ4u83LY3D0Tgh1y7mch0aJmKp8+CfUVMcf7TS4u
r6VlrGVbp+BVs/6n0vCy3aVO7AOtGAtA+pxUsvWZgQW/zSL4ACSBqafgr3wKFBV4
c0sXlHcMtRyV0z/SDOzverMr/MK5GZ719TTvowREyc7iUb5cm2rq8kuvhhvLlUr2
5TRUsdz3A4nZRPRIScewwghctS/SyFSPNy3WYChZWZFGsTjUggh6hI7WG3R4h7tz
6uXXY388u6hPBo2M+FlTZQDYdxtELMNmkFOasIFh60hYTVP4VtI558HugEdzSxM1
7Y30xQqN+srOwsLEJu3g4Tl+7UaEpxtHrq0nzsKU/QdHpVmrdz5HfiXZ48bYYR1O
Rh4uHqoOsoJDRDWKzt2hHFuwoVRSKdaJPh9eyXFPjZO/cc/BT6liOVJfZnDIaNml
IKyXrUahSmMlJ0DTyIIesfxXkorwn9Z4TMps3np31LuH53w5kkc4OqgyZtyKSUl+
JXAmiYYDAGIddmCGsXCsBPEirHIy6ltfvIrgVZwDE4Q/oihe5hD5lZ0LbQw1mHg4
M/grJviSWAydxV82uptnzKNloUgZJ8MVCNuJFKS/gE5VL7vDTZU2uOZU9TfbzGUk
VvEZ26hh7MamdwmY8JhbNDR3WUXKLPYMOwXdS5olTvEjFuorGfc53c1AQ0yN1smU
YxZ2Ou6NA4ozr+JSh9bn5J4EMHZXpZzIPpPPf7dEZA9TVcPEU5tJlEWDMQL5NXjr
kqxK3zfP3d55UUxMV44W8kccTFodVq/GoTT1CkvUsoyQRCz/Boa33nF8tJ7g+j0E
2HDg0s0jDpmQiGxuv4yK0L4capv5bQ3V6ZEhZMlsGADcwu9BtuFxD/GuUi7NUN4M
HpIOF9iHxGNrG13umd3cDJ3CkloSutZ6Y2nNuKMQBbjrAIvgUkXSB6LUOPQEztTP
98YcWw5MVUjswj2C3VtQwRZL6R9efDMwl7/88yTYJ3WPRdS1uJKPsOT22QFZ4Z7q
2c0IQV6gxq2wq7NcVNHkIIVMcyb1tnSMKzOr8MiJYqBSsXEvGR2YKGytXr5arYlD
u3zLf2v2n3YXSdIfZps1e/lBEba5kKe7X+ciyGCF2Cxa7WMJ2UaS9lUtwymR9j+C
D9INTcYz9YsGJW+RK6wddfI4ld0qExfMaFhD+V9P1AXZtXLSDYM5qnygv+9JOXnx
3sjKjGcvuyQIUSjexZLaheA06YOgq7HcJNfuysuKQ9SnDVkRX9YqyLVm7rtKxFH5
jhNmyvg0CQq0ICCXLtSm1q1aV7mK7MqC0GMKFx4PPiaA5JDde4cCDwhtwA9jDMct
J5ZIpO2F/YuCa2Ftu+ea45pKejVE5OJuaAvmP25vJghqXXPA7muVLHvFbGk7KpWZ
UCt2Ns9A877RI3lLjlPBozhEo2GWx9b6MdZK3pnqtC9fmSycRU+jCzerOzPJ9mYd
8mRvcxO0vWdgH0lxmekgxaNpvJY78csu6pCZNlKaUEYTSmYMWAczLNRl1q6nk6Bb
7uJniyT5SMu+JC0EErq0Qp9pkYfkbSVLl2IsEaDjv9y7XGJpIXNsH8TxbeV5YEoY
GLscPS2dKzsgt2n9wXOL2OqoMltOIYQHE3+UF4ShCBG4n7V+7M5Wv6viUlL6ZbwD
qvyvzRJxaHaO0dBJMvXZBtDXpoK1xC1I7TiRzVxmVc5uvvp4ho+UGFZSDBjH+1Bn
YTBKrKf10yDhfw2TLFBI8tGfHJba+MC6D7OKKQGLn1KFuCkPpMIfTqwK+em1sJrh
OmEDaLoJHdWpOEmEXZZ7604iQq8XIQWxiIm3VwWDA1XL6gb69KsqITrAllaNPyJN
Ycb7MKdm/0aUGczzoO0GeSQhS7AhfC6+AzbiFdA6XOg9AosFAQMobw3EzpZC3zhh
3sNPU/xBzoGd89MiaoZD0aQC+24n+NteGcaixH1r7kBiJJZtgZkHzZuXa/Zgwa8x
93lg7GfFP2AI2ERoA/cT1wlcGIB9jphAJMIuiOCFAkU4Ypu1qyYn797YMje8N/xo
vMb6tICivcb7qOaFUPQxZRhdCtTFJJj3fRCBgQer0Ij6fGvo8NBOLiYvRsuGjhZQ
q3NNpPATj4AjsnjBwjNwuSPZbT35lzT3mzbhtiWFgPWIL8T5/RvkZK/901JifeiI
nan444RQmulBzt1pBqixIFRHdO9RT2+33M/6cnQf+U1E9iwWrKeNLDjnagSkFqm7
3cOxr+cIfPuBdvarUhl2MYgIL9eQtck6u/L8g9Vk87Z/bFiKBpZ3+n4/Qw4ZOEnA
zZDtgEiM0pyARP3Xx5osrydBdwMmBiY0XVDaR0XqsPPFIJb5JzVeoqAbrmPeJ63F
eSaNNBuns3fjorBl68gAOvLSkLnd+HL71BmwBagPLScfQuE/NpGFY6ad1uNeyMPr
qshm0WPmCVTB0Jcz8qgArEh0ep0D4Zdp9V4nDb0cPpdkTKffGCYgF6JZ10lCCCQh
iUgCH+f5wUPFwFs6D6bA/Pv/q/1pFQ5oOmQox+zHSRClCNlwghm4foZXAGjH/hiS
cPVedwljhLIafYmRQO/en40N/bPHKOvmWZVWRZdB8/EyffwD3zmeBFHL4NhiPYXc
7reFHyjvG2WdXeZcVKD8/PY1tbTbSzA6VQ+1MwI5Rn8L9hz4HVxLOpv+hhMawy7F
m0X4Z8PKY1EYQ06jaFdKAsNGJ6SKKk/EIzHdzXmPr3qib0FSLyFy6XovmxNv/T98
7TCJKRkSd2wPxgd7SoPjGhShcGUUZEU9LKAPfPwgjgPL34N8RHx0QfmY2/h1FXzB
Uc1nt4S2fMAxTmQbfkl/Twt4C4oJ7+l8d6cwzCov+ndpBYUhhGtqYuxb6se8nyXS
R0/NPQU8vmh5N5Ab4NZ9lpMQkpvA87VgEFRseZ4Ib0ncVHbXBkspT3aJc2oqe4R8
/A4H7Ra9UxVpKm59TvN7DOnz5PoX2HIbTsH7SB6j8ogbFSEI8t5JmPDeLp/8VeLt
79Nr0WSh02q+kkU8wWoLnL70XC3cw5BSyg0PTb2a3S9UeWErg8k12KRT+5qvjOlI
8vkzPNX7Sd/wwlHFkME5SU+xibMujHRv42xVIV/EnJ7GX2uJmjJrjzpAkNs0rcp7
6a2CKdUy1Ib9+LOYY5vbDFbW8gnbdExAG7XC/iH60n8WRSVxbwDTe/hrOQbtbDzv
6eq2a21MU2D00NbJpNHZO+3n3766U15aVeWhI1+Xlu+osSIIOMk1KKn4POPySXww
4kTJi9Qz374jzuFH3Clz0d+xfH0BGhCNSmdTHHnHaT5+ASFNtYGiIqvD0sCp2qkb
PffcbuVOziDAibx+jeyoZzlYntva8Aa995xN8/ikBhI0ho+6WBFTjuG0v2hDffF/
XxE6f9DKXmFFDP5OJKxdDTQzZY+X5q2jvklSOWKa07nmskM6hjjEhbzxftxoRHFF
Yr2cnM+4vs9IIaY1XobQ4MJ7m4jzM4pevyH7g76VusKgczbmCwJoI7DcDvgyi0DS
lRNkGQQJfqXK1FrkUQqDqy0lS/h6dNxyy77upadYbCCv3FEcC1HwdOrW7ze7x+hO
lQlzW3iRTX835uDMgbKNyOJAeXkMeU/yv+baUfWystP0Wd6sI1enxeyav87gefYh
YTA9NYkviou1SDNJBE3NV3QoqYhna0iEx6mtVutH2gpS/38uhJwV3ZeXMr/FRB+A
71uhoSeosgRf1Sb7j56ArWv6Fp81eQBii1BD3+44z6M9YVoXxpQtQVt2xjRhkrBG
rd4GvLCvKqlUVJOyfONcrGc89LDtphxKNw8KNBNifYj+J4hKWhgvR3DoY2mP2Mtu
t4eH7Cuw0TTkHU19GyLVRVok0GdLkrYlqe13W25RawOEVusBswS+bt3Qgj4Elkk6
IPbfS2KO3Qn1QgyqOuwnFxtX1ZixAwnM80or4OLcjJDW8DY7dtDV6NJOqOGukHvt
OqjCN2Q6vqODs+uff5XhwjWiMhtINLymqMPZq8tCduE2F/9eSmYmz/v3dtT5LQRY
S/QNW1h0HmuWQ2pzPfjf/O9vlu9xumwHk1S/I6Udplmm69902Y7VlthjHhctLBYk
4bsN9ikmu1MlzL/ErIcohn36laNthn51kVmwJidtKbWfFuoS6CDvNRrQzuU/uJSX
WhQBmB5uCDIGdP/e5ASrTQN5pnBPhP2b4ji6mn+kiE8OIrwgV0/pC3rJhydp0CAk
iFZppa7qtFD5bGVwEnJh2RKqSLAaj7BDWgxzMCKxtJExyMtVAnRH4aDp0ttOOt5j
2pjxmwsrTAcl6kSb49ebDNyKnqUbJyHMZJdHMq72HzeFPL6ZUlcCOMzudnJaKrKt
KK/8FS7SQDuKBuBS7WSUMzDzlqP2kxoh25x9T8RcEpvs7WsvUEmOJhRK+nxI8EMg
wfig8UaOILXswT7biXMmoeEuv1x/K6E0yseLb5nSss/h16Sxw4R3UB6qRL7Aovnz
oXA1jg83/b3k6NGdRuSjwQB9YbJyxxJW9yYL0g7oaQtebmG2pOE2H059AX/3lXSM
R7o3BXXurvObXenIxAcuCZq/U4bxDmzI2WnWU50P7r6QQAAeYwzeus45S79E80CC
WoIcnLJTFybJiHloK7iKq9p8q9mfKzatEIjPzF4ojlzWuskhg2AlGM40CsbLBitu
6H7yxDiWuxLC/p29BJHrp4WdwbxrLWKZ+o2+J6EnXMT7ZbUZtb+ei3Sg9DgotLrJ
ptMj6Z80yh7RH+0cjf0F9KTPlou8LXA3TS4yAen8sS9NayW9+RHm3rDhFjFt4PEH
ePWHSQbG2jyPbR93d3K7zAUjUtP0MSAEUoO+0cBp8b3BKpIg4oaGFnJl6vyIOeJc
sK6Gx1ETy1IRcbjabpl5H12Gi9wOZuHq8M623hDIPNAthOOlqdsDqOYuYn9if3bk
3+QFB5XZfZl2UEEuRciQH/On3VSiuqOyFkcfnb3toNcqWeoea1V5HJ55qK/4kV/B
919A5Q5XQ8T9pOHP5J8vtOz4/3r1MsoSvp464QQdLlpGabVbXFY1aE2eagyYDA1Q
Ed8klLBkeqt4vkdw+L8Wpy+M7BBaxss6sV01U5AHxJ7K5e4cXwE4yLfnXVv+Y4BR
Y9SbAL8+IPPqK5W69IDbGt9HYZ5BtohnNuXVYXmK7sjM93T/4XuCAeY04vy78S3A
AqmzqsNJRZq0z3lKB3C8oqonvINFwWd0FPReg7uq1K4Sr99wWQLVQAJtUyyxqvIu
QdHraYexe0OVavNnBkMUkgeQnUVf6RbaGH4pJZLmUqhftMm88OqiNDR6uUUDegIV
hphvxYf9IwkNe7tNTZfBifIqcgKjneKvYcTqtur0oppaay4F1z00kYlWnPrhtsiJ
YLZk99eoldogkAFzewwdGJbMk0mCLboBX/NRC63jxJrLOLif2I8XBwUCrOzc0Or+
VVJLlKU3Q0AvF67hM0RTtzYhZZib2BPAsl9iBwiAWIWOD1WyiaPSLvSdQPG27V/b
OxexMK8BepjtiopIHFWWKLYie/mjsPYCjoOhwWvehv+uUVFAWxW03G7XpgGxL8Zo
SrGtRHhhywEfbJxQ9JtZMo+PR/gfF1fFM3BIOCRYb5i8+X4EW38V/uT1sN2E68S8
aBvB8gi9c6O3kpE/AJwF4aurFgG8XRNqd+8XISM9FUtaO6BN/xc3Fmwx0tMteDao
7hB7k6tmLPULfYknL8nPriRHJECvlc5uTK1r1uGRd5lssdnY0i0UeLyTmPXg1vH8
8HMpPN71EKt9ZVySdGqtLUE2TFqCXsyheS73+tgdHLJdRDq24tXdUTpvGztKPr6N
InZykiUYEs6wPYuMrjJKC5oZe2OogvKjcwHbRZYYoLWuPpHSv8FhOnfdAILKQFSm
/pCHtwF+bQtz7rDkS/ByZ7qD08j6b4MzsbSTBTTmBa34rWdkFrOQfAX0mVpqTvKL
d0iCLmY36Kosxsk/kPY5qVzqClCFdLUQjZUHMA46G1+ZEdK2iqFn01vDMYlE5HHy
IyYktJxGVnPXCW7W52seUcAFaA6Ei+4CWrKN2ozVMyzAVN6bMsRpDR6x4Xevn7yY
WqLTTVKMIjAfccYG+9delxqAK8wJuWXVwZoLdJD3mEwcIVEKtMKjWQgWOo30kzV7
YUQv7qJw5zHyB1Z2reLepwdTPR33940H20GLWjEzvFCAIr9wki75SScYSppS0PZ8
wEcp3m6mMDUNGM/XiadPhCYUcIkfs6NP2nhw5OzkYNU2ZYs9iXX64E8XlT/F3h0I
1eUh3xMnix+KGW9imC3wma3xWfAWNB9EHGp9jy3VcBKiZA2wUQhD4lrmEjWN4HbB
bB566EDFvYCTJq4u84UaB5JFkAz85faWQT/8cfloXLYX1SOUjCitob+M+SEenyU7
iZ+VJ3XfmK8gYAA8BbFuu6r0eA/ktrCQkA0nOBp9ohWY6DJxlsIBNswocWkPbDbD
c+Ued3hwSle1CtBjiPz10yHDYRoNvbBM99aQO7uCnq4Tl14KXqmPofVaYS4IspLV
Hmn+X7nDYv4blY5E0XIee/6xRI3wbnXzGO28H2qg/9povy4fZUpPfNMN6MkRnCYV
hmVBeuiXz9GkxqmFULUyZExFNWWqrE1HxojYYrRuOwsQG1kQxu9MKlcSFeQzv2CV
ol91MWeYZvUTgg/xvDuSX8ZbFRlfy8RCAHOiFLFmKn+enFVHvSGE3uKQ25rZ9Q4m
RVmQWZ4yESjukqIIptDY8/V7CYWzPKekuS5y2uqrC93G52iRXs++amKSUXWk8/3f
8P69RXCJ6Bg7uo5/mHlbitcu3W3cI9+oPU8CteFgH1dfgzT10eU3WzqM5KBezRQZ
4CtcRsRD6cbzioNOXCgcocDwAbHw8M0k8ZykygXLOE8hAyKZ6DmHXJG80b85rcft
kGgjMg5iND3+NX97NzfhDoFBT1vah8fkLuts2gxTXqpu/IU0zABT2PRESyU5IANQ
plRHOwlAZowGUxLtmMEoPm47/4qLBlm0fCIt1JsTP7d8bu6/s8QyZxsaEXHJLMQG
Up8XF51aLtgDcuNSq9fexZLK9wEwJMADrP3zFNnhZu/OAq7Ayv5tmU87Oa/AgG+y
R0lXGJD5Ud3VKIFUFNMiGadCcQQJNhYbHof02aIaE+KAuxE7aSOAi6HmRm8eyNI2
y4rykrZJsu7MWnxhviqsF9r2mY0366yyKTrpxS0ZeYgmfWkxWstO7DF4NrmdjL3o
9zdiZhkJFRGkGVFlSpvljt52fIroBL+aKUrVs7p3vF3puvQK5WN5mFGR4/tvWqJS
Zc9+JpsGF8cTLtRTN6K+tS9l5cM0Gw1ZIy9EEJCgaoVhN14Jl0thTx6CzcS5Jefo
vsc/6HPmx/OmFNzt3xh1fq9/9+9NDnwN1ltmnWiFnpAK+QC+FH7FmyTM/Hw/6c5c
/sLx5AJNtxMqm4IFjp8mrYZkDTc+eogB/gdwSgpfaBsakjIKZlRzKQRO3nCCWFa1
CrBAGupXj9UtjyxAYqs6V4LFiDLa7URRbNbIW4fCWGFdpqTKCIfUqA7OGoAFwekD
i0QqYEPLJS57xIkTwYpuSePJMGwyijc9oW1Cd6KhysY2Wk4+HCFqZLxLj0x/y3+q
+qUiWVDePpydr1DRJhKo0e/tH+8P9TVRoWB3hsPs1hZKMHP+4FaP1VNua6vbKUgV
IOsBKtrRd+ky6d7zp7Xq4uhDOntVbtgMk9a9hyWSwBEPvrsLahhk0nFOgiA2zB6t
eRHcElsWUKbG7HQDyZioYKuqg1tyWzloC2eQPEQE9/EHLSYgQfyOdmey466YMN4z
SqxyeLZZP27tjMjcx9CRULnInyV03CoiwCrEjq1esDtZ1vRD1bIjZZ2KLzoZERci
3xhLE/I9yprr0sQ+A84zda+sKSPYDPqk0e98iMEpr1eJP3MS/2yJMvQ2VSxXHcEK
L/EUw5P3pQzGJI9kuiWpJoe0SRVu/VNx4f2usjYTHMoH+GB+0Z0v9A+Vk5XsxGwU
rYc92RnH/oJn34BIsX2BbCOIgyLjhJOh5jAcUeMJ1VlvRtlKC7tpgKH5HzKsR54U
7DL+oWPalQfmwxEB3ArDFEQ9htbY6p5HbfFPjXOJf4bljfNLf+26zNwQXiiVDq1W
jOA0M3I2Gx8eD76MBavk6MmG1XyAcatyTJHCMA5RvpL+5mLwqVx2w6wMWKhf60KC
XIRKjCWzie+i4iV17q2QoHtIozgXpP7E5A//c+mlqkP/L0m0R2fCFPOYyucio95y
P87O48LDCVLdk0mO9w6fR6v6e03e/OHn6D1PbYrHO3nCPBZrg59sQEmKiOhpJ/2U
R3cr7COFhwmFEj/VpuBGQDho/A7RkBYsitaBw7bGJsIkA7lp+z+MJg1aWsXUrQkR
/mfit3/HOMlI4Tr4dMTncZdlicznQIhXPKLCBS1MgUtR7E9vZeYOlGi9S4d+0XUr
OeDHSxpVhssXwhm3SC7Wjk4fSJWrXo66ZEZYac53+6B2W3NWJKQzQSVPH+7iA2sR
ThN/kMclXxdy7hqxrghU99dLsr6yJNEBq2bTlmiMfrrScHe1oID0bcr5+oC+EkoH
+94I2IrxsLY3gHtKHA5QHvQqH/2q93xeYRysvpfI/p8rqJcVSbahkI4aQQHuQuEz
Cv8uC1UMw0yJykIET7PUJ91zcc4gRUPZoD5rSKk1EHCbF5UbuLVLD0BYk474FoFo
yoCWuZO0+bOpS8PsuItn28zToRqQ4KgBrYPi59peF6U626t2SwfD5Q2gEePTgE5e
9jB2ID9i56fFGDhp5FNNN/LChxWV4ahpUDgAL+t4WcxZn/EGz41EA7MSf21GJqDO
XXnRewuI2RuzQ2XicmNrsgpf0Qii362JgOJfVOLnjxUojs9LQ2ZFT+OLP2ryTbmD
sdhwWLWGM50bv14sNV2Tc/vdqdMbKO7XcrnE7j8FetgDRJy/AV6TBCR1eeQfVjDP
nKlB4jtCg9+HQ0fFY7NxUXhTAgzyFoXWmajEMwUSQooxxHER4LyhisqyjNrJ2rE/
Z3E1Y1G0chmHLSZZQueBN8oXcJ9F8myH+JPYAl2FPSEasW7bevOO0E9llmi+mCTZ
nWcL+SpJGtYFZYPIKIeT7qAdJ65zEg+zJzmzN8mOHziYEB6griwwV7mpP4C4G5iL
bEfYgyLqlwfXR2VVIhr3oXEcy9XgLGsF4SM/rRQQddE9173F7HbrAjtNWtQ63DvI
z/pgXHjWWznHCvC0Cf5Ks4ayVazbYLcjxYSuCkDuVzQv1qMB5lz3cJQcnewKdVlC
kmmAW3EFjCetwYVfC0rNHkWzSNUwchvUzQWuKUrVZ+zIDG9vQStUIIzgJsgXzfnS
N3Uykad0h7Pa9hlx2w6os0JLOgUdZMnFgLRb0SAUyn72mlWrNBILbUMXI2Td5fPO
l6Rv1wunWpk8di5J1OMRTfnI4HnsVWM/bohrGiaHtZbUcn6u/yssOoepHt/o0aJk
NDIp8+df5Ist1KKbCSClbTqA61wowW70tHCzBnSYOHaG0dIyPSG+MxZkHUBBnD/N
oN7I3E2qMQN1fvMt81VJMNKCPTO804kvSeGoLTcr5g4DMVHqgkCzfcLWOJHcB1xt
E7yOXQgWEncyNwbfoel3870cCKw8jdiNkzII2aq8dvP5YRP0bKhlrvvIuoi7fPec
ap+/I8SdI4GUiN2DudVILC84+h4PrK+TC0932NeqIHclEVMgBWGalKtnK4gfM8R+
toZmwUbRvdkQ6FPQDmaBqr1Xr3jmK61YWLduZOSC5860o3wRQnNa8nla29gp9qqZ
dPH2VqqChyn4wdhXC9WD0HNNaG5X0EyWrgPzamnWqzcU822rKR+rDCaDFl9PaWYX
MCtHEGt2j0pY4/oFTiMbx+y5wba+thqfaLO1VBxMxEFBE8pwQ8SvMUIFPf6Z55i6
a/hYuBr1qNWeOiCxtUY2w65auqaaAuUhf+Am6bMtNrqGKC64vN8+tBO6h0QHdUbt
c/wKeEViGFZc8pl/aYec2I3LhqNChtXx8LNLuj3DyOXJ6/JIREEhov7YQsYNQmX/
BXngImJisDrUld9Rp4C0vCnRrjR3fxSyrjq0D0EdkVD5WRNTn6dXVQMZemR7HofW
LrI8iqasVLGYEIVd2fTNjko54LyRe1gQFAdLTgqAlzjtPLDaj3j9MXhZIVOmT3Wo
dycHDWHEud/0/Z+mkHZn64aiYCuQltWndAp/Vv8IXr447BAVFAxaEdIXecY3m2FG
CNfUPLCodUBsbVbqW5nJq4NwTooNUb0WqMiGHOFgCJdvyUEDhUT+EmYQdGZyiJ4V
tgA9Ck2IPbd2JzPQLDzAB0l/I0tCI4yfg2jG5usMSqbtrHdI51b1JOGubjlEXE9S
1gzbC/WyetZd6mxj/7/4o8i8Z0s+m4tR7W0zc3TJm74jE7p7XS7gFd6krX2lYzn6
jCyYRXlxIua+NXSNcy1Oi7Uxm6zjPe584wdgzPmr0b4Uu7pqd8FxRdSZKNSiR3LZ
XamIA3YBrpJO9Ie/xcqhOCxM6hDKc5cZfCAwWKXTqBhU4WyHUMOQM0VFRRT7DXAM
/yXRKAQ2DHrGbp1FvMm/VdzIWu62nxmcLGv+yny6nYkgJ4q5zlc01TBzqemFdy1A
uVknaaC2JPRpTcgj4Q9Z1hL2q3KPFM6nFvmqIkGkuBRY0NPxK4Ia5x6yJ3FWU3+C
89bo0mQmoyvKh7vG+Fv0lAEsQF4hzIH1/CtcK2bod71ViyUpwSL36MNAju/UCr8P
XVdBoj83kZo5An+qGyhfqMgiGoA2xYEzrqoXw3uCdFouPEdfN5Qec6PF4k1cXsda
0nxbZ8hqqjebr/1iech10gbGjRezFQUKaaV+NX6rKimJvRW2lgNrIdofw4XHP4Sx
kuZddbi73eHQRJbJubI1t0dO6fJ87ckl8Kuzr5UD/8X9lDo1NNxxeMCQBzi42Mna
+HFABK8e1mx/p5ZNQe0rvP2pp2hLIgDZQdVwnPGLU5IfDgNlAX4VUs5O+mStIz+h
0KpTt/japlPcoSNiBTUuht5XGP4mnPrlnzBNq/uV1tBBDfPAesF7T16FjfDmoGY/
H0sgA3SSc2JtAgihxJD1uW9Oo4qCl9NBEj1ov1MF/wTV5P4KJaPlk18t0SQBscDp
dBU1Ppr6lyfNrMCsxxldFpZXXQt01VOIGi7eC8rDsmyk4lYoWCKLcA66m0InjmPF
oWMukwIY9QjRP+DmyKPuEO+Ancxmxek9tMfglvPqg/kZ8jhTZ1UdxaTyNSMJUcvj
EMDFI6KcmGLXvdf7xpJWqRHf9XXsjfgMVfvvkJcJMD8QvItjtYqEa5yEMg1bA8w7
q3FAkrP19KgWjNzayWUHsH6Bc7q57gf4uibMtWEYMWFHV4o2YrsOGy+eq7zWIVmC
HbzjNbevJthzTEhqEdVTvaU7f0/BkuqgVFPKywdaM7f1B/gbYjuLGiXnbRs0mY07
Awv7DtC2cKZPZYyEItOrsCloyRW9Uq5KgCmpvFiafbY4uQICYc4vzKFMA0TSHQlk
55D2Hy+1PFdSRxiHPdPphlQe97AA1kAmbR4S72t3DO33CS/mOWevCSFXMjIZSkUP
1sCPCJaPH/C7rA4apHM4FTg5dtZil9jRgz8LLT4I8waRbowen59tJ6jkv6LmuVlE
lLSQfKivwKk9IDhXc8uB+kBwrlap/u3ARye0wtTmejVdP/4Oo1gJEWAZ2+af2UW4
EOotOZ0CGWYjTrBZFHT/U4CnHVHZ/xqkJ1GmQIr04oklc8V8AGsIwjxp0saNY2hu
50hqssKNv43Vi20brUDsa84cU7+wFCUkXDfZZxYFlXxjVSwoxIab6gPST9I1hdsN
ChfZ5kSI38eomNMtIDPv+D9MaHqbBYofazwXeeS8ht+XHShjebuZ+zokAuCXYf6x
Cm66EmuYc3JluyqxpRCcQMgLReTv3QPHPTIVbF8lGdVjVVt4rdqx8I4kOh1Upw0H
EK6L/6ZQ0lT0ccTimT8/vNNf/XVFmfuaUEbU+7vShnVxC6jtQJ0wgvJK8EVjxqzR
LQaxd0Ww/KxPLNTSqmZPPuaAA3zFKlXql3QIxNRk09R9R56jmGIohRcrf8dFdeJg
fyeGpQZzea3b2up0wrJSCtAfUdm8ZrRyMGI6b+a+410CrspvgOQL7lAxDKBJM71L
CO8GbFiBSxtol5Js1vklCpxovcG3kY9BnNpo5SqYFF06yxUsmCwdeke4mDyfyS7/
cVlaFccUt2ulMnPZFvQFE9AxkmzJFDxCBX8ybTApQigfZr1sNO2Vez4HappXLPBn
srlCz9juQ5KWGAeTlVs8eV2LNwXKHqpDEchhsLf9ZhiIKye2/1K3Z7fKlnb8JsqJ
yfjyXHl8RjlESaP5Lh0WxYWkW49HUroGB3UPZSK75+BojuULi0YfxZTg6ENsUyhN
+aL68x3Ua3OK5yfd5bPFl4iTsKIIcqAvtyLXz212WgbvpYkxA93EGeGdtyrzH4Wy
zyFZWmk5kWNRlamxGsNCDnVUX+mpZdTUlOhFS1l+lc09eVJdRQaIzGxFwzXxM8QV
zHtiq7tEuWcWejvEvbdRGVXyQGNCD42dcHeZ3nixMVbLJJrM6WgQ/JJfPKyGyNvp
WoHI/wogl7Z3uvjQci1csJG4U7Wn33peYVXCSJYwMpuO97GALWsCkQrxDkoeZJr8
kZK187uRDOJEjH59FojOaI6kvNdx3n9MZbSu4C7MdxwoFjVr0kFCDsP3ZcQmnB+d
LNTORiX2O7Oaoiykr7GbjfyqZRHSLRTISqNdEkAVZ3zTmZagsImWn8GFMZBVVnTC
AA6NYK8YGWGHuBmgOE+wrubMfQ0T63S3+Bels17Zhj0a8Tx1lA+W0GJ1Ssv7goib
2mBVTzzpOf5KJSmsquBFir//CKGBgmmnRHJlbeNeUi5b8ts2LC/XmOl9+LnNVoQ8
snCFhTUc2Gue6+Atgc/+BKCPiZz6EJmRsLiTqSLpFxmps/SOx3G5IeU1FWtNXVQd
DEoUlSr1bpw14IwJqMELWxzOhvjvMrgFFZgUqC4TS01DxM3Gm56l/nJjArQzWuGL
sufcK0OTISf9NofJnxkilP+vnUWEQy0E5jfTlDA+NXDWLfp9/QmBppSS5NOmw38S
qs6GPpZBsbfgyeGthpMDO/kDgUDDDyChaKvgtivgp+LHcH09M/lq2qBkzleq+XQ7
/CWtPTokpnUuB6aUraTEn7UDEGShNu4xi/Ulqv1mZk8ELMsmiWsytN8IdHa7ERM4
lkkKtIuc1+xofU8wGe6O5MDMnbnibRWaNLGG4bf/GwX9Ro4+LeNbdDyfcN7S9Byw
LRwfhQSOQpfQl1UNG4oNSO9vzIXiEWQ+9GvQJB4OyE+NjuHZS2+AkkOevvlbRC8P
+N7xxkPqaQYhUJuLQy+IkAKVtUteIypv5/hG8c+Eze306x+KuvKjLqcH/y5N5MtX
Hdrn5fZIlYK52rUV+fJpDaxMxlGlrI+J63OSDiLn7b0IC2RUkuIiLUhoVeS4l/bC
k4lgeENUAFYNFN94WfBYTNGyEuBAOBUIKwdSZdGa6kZtzXQcCT4/H+4hDdC9vfxN
CkWkAw9aHFtnfgA9AcaV9/yTW+1+OfdyuATGPrOeM3/yy3xEPFRRML4pn/X02eWf
XdEYBv/qqjzbPrCJN/L91HXjPPFjvQXpL7DqB1Bns00+C3s9DPTycQ4YDQca5DRq
mrLUjNglKuTZXabwIE2eBrMIabfEVYmwnfmbc3jqBMG5J3Osa1l6XaZ7nIuL5rWz
CWk1+ODifpttNDM1WGybbefPev1waUYd5RYa8I6BRajQgdNUZaxWICnjyq0yaeju
/8NtcyiWTWPLsHFjtWabH/AvjH6yu2SebxcNnQo88k0O9akR+h+ut9wq3J7jio2Q
TtyV34+vXB13xM7qtesRzhk11/b+wOM4ZpM5wQmzwFWnaJjZx3qPTxk//NNjYdnX
NxYdqdeXBTmzQmhVULgDjJTHkVAvrtPSG/NRVjgMd/YEdVPAcN3D0eibWzJuHj8p
3t8UJ/n/t7hjbqwkhGUaFtB7rQ++83irRSUDwa+ku5AwkZzFg0oesJK0g3INbnQQ
4hDUHA0F2QhllWQsUkaDBQHGCgEljTtTkqOuS57XI4eeQZ8DpgvrXgo1bOpFEmiz
aYB0K86aLOqwH7ymv168bWRMeeImdRwBu+QIrx2YYjyfkc2FO5gyDItyTK//yzr5
ktpTwexD57zUDeazGF8Q5t8478X2G8hnaP5v2spexleLX3HVSwGi17yVVxKnftnf
7eFqYgdD/w66corbHjZrp+u1qGUPzcH8JbeTix7uMFBOEhX95T+DDr0mcGrjxfXc
S9C4+hhbRlUBgPwp/Jdw28zTC8mAFCq8OzLt2TYmRtRUs8A8sO0ReTt4ccd9xMm5
uQ2MDZlEp5CISQlcDUv9Zm7WCGgQvxk6vxowZhit6nFaYClh0zsZYlVjvSNOqp1n
op9IFH+xGnrte9YYNpG46gIwOnf8PzS9Xbbrhx8CPUAQeGYu8QfX8I8mGi34z0wJ
vxE7bsML2SN8+sEQwGdDOGpxBJRLiWhijJY+8hmXqiq80x2Sa5x7t5qd77gGrdpF
sQLdUVyENNKBxl4NzDlKKIbIc4zmimXqMiyzOn5JHKaL8r4E6MsVrrCjyS6I1b1Q
jRKlE2uBGn+6vF8tYYLxklW8WWB3q/Ob1hCMv1YxtnWOuA0rH58TkPvUtbNqZtEY
kQ/MjOcDg/BXNThnVnJJapzK9v5SstxM/QAd5tpybhWxwpLyKahjMjI5XCIlmZET
oR7JDXI+st9YI1yc9Y7MDpefKCriaNE+ynURBonikklYPG81qegZO1Zn0kAhWsE+
nDGigs5xs946t4X62iCQndcUGBki9Yy28RvvP4N6h24CtiWSZQWeNAPQJtQfflV4
5QGDCAZWboObFHYjj1wH98ciJXzSqATrjLCelFRjh7QCqxriKEN8bObOZqmcWErw
AgMlq2cgEb2+hG8pjM0u/aZoMDqXCTG9zpptC0F7ZfiwmyZCD8TvESxakxNrV5Ri
hW7Ix3tuFtqAuGJAbkne9891/s+TN9PJRrb4LbgOn5BD+6pWUU6WrGYjzMPo9Z/p
3g5CFERZgnN9FzWzangS0eSUKqpfWItJlRuaE8jpcRV1CZ6rPGbsm6ELFXFbDP/L
JuWv/wE8cYV8Hq3ARWYzR+w719hvtCH14Ig/XH4kGr7CA95MijmPkGYyH+5YWVOQ
yzWLjXlmgerzWtxyqS7TUe4IlAqJH55mWi4m1J18BZN22mcQgiKoyZXpmVwO9ogT
BpR70KEkmI+YA5tAClZ3NXmWzVEVkHFCmkdC1ZjwmRkKdBi1j5Kte9L0qjtIr/dl
9ltd3Yl7MWRFBib4LBS2A+yw2B2AoEOte05XZ2DR2omhI7rCCdMYv3iu1pB2AIK0
/MuQdEU+4I4nsLbHuQznB+Yf4YjfcgIv6ie7BdXLrcvm31Nn9caYkn2okjFRuvJE
365uAuBjMvsrQEGsE9YvpD07xneYkc9Wy1HOeRRqEP1KocvkZn+LLjSoREcJTIX/
tP4UAVrVzsedBzHfe8tF+C48+VDTiRHrFRyphlMMYr6eUdvh4P9X+TI4Q0YXFm1F
O3+0kAMBR3UOIVUfNVfk856izenxbPkqWuZK7FHvr12FegTHwCIjoSp5avsxDfjb
p1tH3ok7ufsplY+gXLrhC0O22AG02lykuZ0bBt5+gVbpVN/3oY4JWr619DKEYvws
jjPcJaL4les28SgutgHegMkzggOefdUyC8MIORRv/mqLEcFWA28JdIUp1/cwLBgS
xSn4+rrGtCgqkEUKfxHkYhZAxwrqi8qzzGQ2faPYp+mnW+N5H69ToOg2SgB6whtt
fvD2lN+Bz2PLTSyECiGueT6Q+3X9WRtbnn43IdfftHF5CYcLZOneQEpMbj5WkCiV
kvFE1Kyiuog8sYUPChot1L6pIy9+Jc8hMy3c3RlYmyKx/rySwBlyZnJrJypYVjaB
2b0MNFQsAFM4DXoalRS/Q5u0zvuuHK5QPZsj3UbfRs0YfIXHCKJIOJ++mo7t2U4A
X79GltKtu32l/ZO+I1Fl9A4+IruyF1OwAnP1+PI0LNDubVRvLpyGO7DvkkGJ6+dV
sz4KRu2Z0RozBwvXT+KXbfRBHwdV4klWi+13XI4j8gyZRBQ6IPMDV4H2mkzZMYGr
d9KPcgjFB6ch0BHKUdKgJkAMJ4r3K0FIS8SC11n65VuqjAgZnNtyvV4k3kG+ssOX
eFhaDB+0UHlyymrtc7Y5Jx63FJl9OVqtiI7EieAc7U9FndfqEVWQ0Mg712Xdgx85
1jIInMQVORXsWCT/h9H5wnVaTpCTzZel9ZZhSKnJ/VOYwkExVbf6BOQ+4T2Jb6Zc
O5oLZdS8wPaXj5vJGGFNFe90S1P+2pdDjYpYjIN0RtVAT4HmoaDQNGmhqC9Bjl6Y
GkO4wtaZN2WdK0R5R16zm67UVu4U2jkjGphMMwT6hR233jC9UhHPJJVOEoE+zh9P
TIyJbKIiDWkiOo2ixgUf1zLnD9F4Jgoiqd0tG8V+vfloLOFPRqlXlCaIVu1Nffj2
QzdpzL3LrRiYjmTSHy8pcorD9vj6MSVMHjBgqJP42Z6mrOH45S14iy7ydX7fHF2Z
wCKjg5aOsiPs0HEDhG1+AbSGv/G1hH9efimnHUA6DmIqyQ5Aoa3XESaPp0EZfku4
vG8k4Lrp48m79wZPDHllYvylxMvG4leYu0boG7smBGYD1uSKoequM08NRf+H7QqW
TgNBau6xzN5em9bInQejol4G7j88JihKwyz4sKW5AE/HL0+OxgjG7ar2emWWY55c
wXHWlaN0igSQiNyJKDYs9Lm75pN/vaoxN4G8sMxnVfLeGrhQDdxoXuGBqwk2mb8b
Hdywpx0VmN6QiQZNiE1cD0njlNiMxxTl5hOaFsMh9cITy0MYZM5Jo+spLJm0tvhj
X9aUFtlA2P4WOkO5wcPA4wA8sk+mO5BYENzogDyv4hcRFj+xMdtm5DHgbbFuRYal
kPKEkNHnTte3GyyihzgAMV8oZQ2H5xNQIOy5jKhZ5RyH8HguDEYNpceTZoAT3gEK
Xg31bearKb/lglbpuXu3tqzwbwnT3/Zv3MSetU6iEXKXCD5tniH1nBv8J12T+iT6
KvDZfnhxkOUX0rHJ3zgJ40iMZZZ5OE896mSwbEWi0W8Hnr34qzqtvbZWo9jn5xF5
Rfwv35n8D8JPRvCQrdBztaSuYIm/m6FzkcUtaU0Akg/ZAJi7FkqQEt63+/irmF5K
F+ofWuDTUK7t1Dw3trTz1JtaeauD6dpVes9PdqVnaXtPLEvKGbGf0XN7zNUvD169
Qlio+eLw/EnyWRar26MA5IxC3uhPBngQIPJLTI3B786cOei9qX5CGt0eSEsUnpii
2pkEQdywjKhj/wfns72yh4epfoDIRWog1beOIctWtmCSzZPIDhxB1hk8zDwhVvxR
IUFJITTb/E7PZekBi7I7BOGKR5DmPFM1c+at2LRV/+Gb+uUfO9ECp3vVZxHYrU0z
IKGiZiaW8uluVVk5g65OLSoGIRMOUMktTL5cExlgIXeeKo2dtuQyZlmw/oiXUQAW
OWau874kwHwTjbh5k/I27VFG6j0+Pm/00qv1QE3f921g4QXmker79cNVwZiWpzWB
DWXk3g0aFBmpADntFqhH2HJwuhuOC5KVqIl7qjqrwTIsFp2kmhqJB9krCjp//qF8
6oci0ND4ZZ/xV6kxusHRgXrojmZA/wU8NrYm9nM9465TqsfkLtxROf5R+QVkgTu3
06cUZ0IZzow4LdI9nXUCya16Z09BbmMxD1eMKylilvLRW3K+k+shqKITSRJTqN3E
wAaFCN8cY9YKsFmaunz1wEgk+PKTjWP9isdytfFaE8pXT4MGSjki0TcqlCcc5x8A
YR/fPBGyFxHvhrMeX+R98t3PjhIekAyaypUuda3S4U9nsyg0TeVNL4VzwjSNtQD1
L6SF7dTSktrHdoGHKBV1oOnl1qgz1qXpsLLpCgqp1LSfo1QJPP+ta9KAB0PMP71q
1fEmqPlYVZHncN6KAy2cnqCm2Yx2gUE8qr8PcZzv1OTaqyuQmsLiDj+p2rIEYRZZ
cp9EuDcQ9R/kYUKQXiLs0iK1sLpn8ppsE7mSdxcvHEw55c7bwkggMVduo873zqS1
SdSUMSZ/eqGBuYjK6ZQvy1RGCKMEIJc0IM9rm5T0CRjy8B4eT384RZX98BPiPmKV
l0L/c4umnxMQH+b0UFOSBTEINqzuaNIe5atuKims90DJdf4LTO60hp52NDGOeBup
G9jpzBpHpmw15BS74goVSzRWkRxeCiGOJiARV//9cD8mCXzV1J4JhYM5qywhSS2w
Jz9edNenhvGUr+55WA/1M2hW8rYWVGCXJ9GuBUQDxuUEel9nQu0S/s9cmu4hQn8M
IyCrUUdxN0oWZwwG0/16ejLhnZFNG1JxYj5G4KQ6bPAnL37xkip+jyLVwpQlEGR8
J1FrX6LxtCSQ8ZamJFJmWdRLrOx22iz+LGSAtAaD0bXGIcZ/+jeiU4c9eRSYzw5a
U1t9WEdmKbL8qd/Yf6vKvQSiWvOfpz+SXZPA/HhXmzy1moybhlcMsRxuohFWkSv9
CQcAYx7RLBthO4yIa+QblFNFKkJFjCa7hGAEo+QKpy4rbDdXKOUB5Sr/WRiV099+
4GFEfdAAfvQqLQHfsHciQRYdC1e257i9Oz6OwBd5tK2AXFxR53IpufaTTUWYewAW
nMoD3EOZqxZ+OgW6VEfErNgX+nYnSDizmc9FVdBoCmh7gShpwiaywm0fuKYvciG6
L0dF4MssZ1CAGgTsHsm73o8lBwOedH94GM0n/xmRsrezFPoz/PIdUZ+H/VZp559A
MZ1QJe0MrbjtejaPIdrJOP/VSpKAXgZPznTj0fBrQa8oW5xK7OEd7dE7v7OG4bIA
BpIdTkqpDQ7z4abAi9tiIK0UsndVb5sHpHHQdm4FyKn8Mg2fLfS90fvD3jMfBtnv
1l3MCj3Su6hX5b3P8IvhvbNd+6mzHdWxOn0XQomHxNTtVAiTt9Y0bqeno8MDflxb
kATXrHt42nrE2Fl1qgXxF0R5AxLAGcsXPVwC4+3Fy7k+6HxVoB2IV5zEqYT8pKL4
NBd+XtFJV3Z0nu011HmmcW87NMLo5DoAuSyKU7SNh/AE7U7BuUP/4/YBcpvOsL+d
hEhLlmSevdyURixLLvAwuNTQpI18Qp5Zz3MJck1dDRg9ss/sIJjeQTunjqFHs43p
2EbRzKnKag1k/E8lncFqbbVMJPCNrdU1ayGvGaLyEUYbmqfcc8eWnS+OADos60b/
8FsWc3Bx6JqFGpY7+XY7qw==

`pragma protect end_protected
