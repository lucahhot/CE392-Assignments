`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z30XgOK4EnpVImD6yTc7eeR9dW+F5Sjwqk8qWkZ/1FxgYIYya5QeUwm58LXVS/y6
hFk3TreN1SlxreLV9IuS+CPSoQbVF6JY+jD4U07JAoImAjDLgunz0999ZShxXVfQ
efi3GCE2GguzGw4s04BnvaxYf6eGsDIsMMze98n480c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24384)
HosKeq3ByI6W7rfif54mDaXOw5yxHzwkCrtQOr8RJ9Z4djr4DF9zDC9z4A5ZtiFM
Vk9lyeVZLpPIrfu0yECbr7uwK03NeBUhudj8whMT3i2ytl51oeLYKh2GATKNgw3e
wjCJL64PAAIRAyiup046F4kyBN2YAa2bzpu8ybvpy0XbjVYeWfSEUSWOGkXiwhdu
Z28t1sUV5HmoWlUK2jrk9gvTAOdM+NHs8L/3h+5jLOycRZdcm4qC/n1EGIBFlGN/
lxrrjOKgzgKItqZvNoBE3Js9U2HUCv5SS0BftKVc9Y0lXhOS4Bab+OSOcPWlnsCR
ENjck6vr/dwIG1PslGBhYaE5DRB2DKYd7eFwaW1UWfTLFdwOSoxyiE9Q7WjYZN8/
R74HL0eUl/dhC/ozzX1qJicOBQYF+BLreeO6MZhSo61DlMXXy8ldNHoXiPHfUkgm
LCvwTebS9IML0ibUzSBu8jQmTG6mkz44VQvb5p55UMmfWWEZ5iC2OhDLYL4DFpC1
nsnLznt0dmyeofq0AxFr7Jw7+Tpi/mMplitvjiGg4yq7kxTNj9wWt2mjhYNYjNjn
ndXmFQKGfWK/UF0DrR5lDbIG8vggWt8KoSXOWFmRBjulLuOeN6+oPLAGuqTKngPC
LFokxq/KN7GxSHQnfb+oXM98bOBtq2Avu4nwHkZ0r47hmrchyUHXgAbNQEK2uIs6
4W+5USTnYvnp703Ywhh5L10ISzfDwvNG6sUkDjJjQZ5FWtTP9q1spbIrApq/113C
hMKwvy4pLVYf7k2mYJG5eb1OrrSiBkSXjvSopI12cIqZZ/UFLH0S9s9sYmlgGZgs
GjqzHeixMPa6AGs9sCNyOyUayEZxPnFiARZd5TpFkKoKIQC+4j7PH17b0nY9/Ae+
Lb6N/Az0x/ip/Q0cShBnv0syJgqbpZcGDoGfUKA5D8EJHP+kRCRZUjWJtNoYje5S
/kAu2QLxor8E6HWeS5i1/gWjh/FbkWRgs4GtFyXc8yjRhTTIqkI8dhyjJFX4P4EJ
90E1UrRBrYZyKVp624SEp05xQ9sV4tiFkU9fdVv5P8wdmto4iIfYTPpO/fcsYhHi
yZR92izRuJrNSR30m7ZWvBIoLNbBbO7IdP6yQau5PFfwdUOAdjKsGAHlCkP8YgZv
CSK8z54i/zBwpfUpQcZdyLoXPgPQHEIukum7qsXvCpNy+AGtd9H8isEQrjxL4/0I
NQiJ0zUYpRjNS5VtJ2dtyhih/In1rJnYuJopndeUe6tJyklbcuCem94w+Zj9wmbH
eDBKT7FrSOIeQ9o2wOPFUBAoAD20SB2OE+pMk34x9/P39vjF5i2Rh0A74NMADRl7
H/1f3e/yNFjNPVHjE9+/Sx+ZZrUk88+N6daH9aEAG+4SObhWFIWCvXU1f04nx4sO
f1yN/2g7Wy0nPIAGmtFQqwZ7TwgSHhOyFuk0Gc+mpOYDjWJs4FmUaKO0zcwkdXAK
MUBsv00rjYkmL+iMvqPU4uFm5cKdRGK9EvX2ZCc4IF/AdPSlwVMWDcc3qRO6i0lO
SeMG6L5wUnWazI0Vp4D6GdRBaRDJLxK26D/rQ8rq8fb7kNJXD9y+DC9mQboCr6K9
cjOImSrPejZ4WM0R8mUUUO/XtVnRGmc+JaLwVbhINbl98pxWFXF0taTcb337+J4Q
rvqqWLltUMClal5c1GgSUwUa026tQRyLOOnViVquuZ4qF7OnFrSQUqjxUmMwMJPg
Fs4mXWdzPanXMduy53PvGfplninxsAKawBP1Ee2gwlhZBWWa95uWfozLu2KSif7h
3VcBK74SEd7isJZk4FHhNw6HHH03XcZSbOyXo1c7gwJ48pOl0yI3C0ahohRZdlIw
CLvv6tR8M+tiUZdm+VHPzFlf0mteQdldrqi7apF0pOGll+dFuiCNVduwXosmGmHL
IS6VY++BxhqIAgBB4jKTPUbhCj/8hKEdA2Xccazi+INHUjUgVDSEbRESgl2G4zni
r6RyP/7/qFbOcVQ9UZJ+2CqX6PqUE2DofQiweUlRs9+Xhb8rmMa/eXBqtpvRweqo
Itc5XtUuNXwYdwezCaS3uSs6tdwYgE3Omgp/CHJ3gkb1BgFG8c8+sS8Gz1btAjTY
3XkW8R19NVHoMLQd3qbbwsZZ8hOR571HxG1Qe/hXKVf71pQhYxPTGYKMJVej3kH4
N5W0TBOqq5ZRw2X1OGDus85l+5+fmizM0HhRPikofczx6cNMvIbisxJk+8psMVCC
RSwG67CBaQ+BEdGwAJsmz29RsSfgsE8dz4lkKCPvuAD8IiKWfEymHSc/mbvFLKFH
dANVbbaDoBOaHn+0G9zx0FieWYorJ9H4h3sFHN9aStSyW0Z1SU/6Mvly23rVXqoJ
QVBJfNKPW2Un7+NyHHlkNpSb8E81UrqVmeHLFwqy/idIc9dIeGHix0pmKUMsvoIs
fniFI/AwR2wPb8m9Ux0iDFp36Bxc7ZC8YqqA930+e8E+F8fAJQylDS2XwTPzdol7
VmTp1KS/qcndamfbUFmqSMFVSFezqqzab26AI1bYiNoVpPUKu1SKpq7Jqzy2cASQ
tV2Fe/z6hlW5vlEW8GrXsYWJ2jr4jV2Bsnl16Ex89btU7TbaTWPWOtTCeGLIFH0X
YXBhx/WSNi0ykrWZpL/d5dwI8r1KMj98seG/NzC90Lu3k7coIqvrscDJ3QK3Yeav
eHXGh6yv84CX3CmSVnso/RuXZjxHrQDodgVeiUfB9e90UNnH29yh/8mZmAZdIw0g
1k+08AZc4ITNBkq6GcQgxeuQRMIC50F36cN2+N1ptr0rosUlBbcFcL9fwg+YaGLk
j8emUht/4oHDoVhvbj6yLDCQ7iQOEWpyQtveZJA9hcICV4/B9jys6hRcTiLMoTZL
KWNX7RuJilFKAn4mg1a1UT/4z29x7VlNtxVWzs8GgkcZUfsAD9CkhMuWrWsxzMQs
KubflEHbwpz/8ypgh9yHWaUR7zYRcbHaOsRB1AfTcXRqKP8NbsUrhjZ2aswuexo2
P06nFYnWg5de4U9gTPE2JFpbhD2gMB2veSDrNx55VUMm5L4VfYA29IrVyKuHadDH
+JjJOc7B6aSm+WoGjafHYM3S74miAbLtb43Bolc+hSejI7zsKCN9dBexoRq3co2L
Zb9J/6YxhlGtyvG1k6xImppBssEvaVXVCnuaSGJzS3nbcfc/L2wJ+v1fLJ0gqe+s
bvB5nRCmzvDFZ4e8h5D9AV+gYOteYCx+iL7suuxnPFuR6J6gugMCRhDr6vp7McWc
iGWdbqNlZMWdRUBLkPm5LKYBp0acPi+e44zaXUCyR0z4Ccf0fFE5Nklu66yog/Bo
wpMGOhhJpWBIGEpNMBP0yQ7ybpW/IICWSe89xROD7DAkTWZV3FaM5I46/fovAciM
j6aImlW/dEZnkzRKE+sBWpwoZ4FbkHAEuNhFsB0yM0NTePG2k07vsHWab2ggO2XG
9J5uQZrNLBvkuXStSLZ6NMMog+grEy5QvPdciRHHw4gpUBHa5g6AfRGIvf98u6FP
ad5LZ8i2+cgAcipq7WqG9DIPbHFmWBTTmzbDEKCRxaTmA2gbodpfg+HZYgeFGeG4
ftnSBXpiRhzV+rx+pA8Fz9Nq5v4A//RSU+n2wvRL6t/QVmxhTNBG75kml3KEksFh
EhH6ShgYLevbIvCYy6W0Or1bfZRj0qQrMyMM64b35NrAO/kTHf17ebfT06vws92A
By5f6oxl4GIudBwoElbV4Gp1JpdVb3KIIKQfPBihqQ9Pczt7ltvaj3DCZHfiQkyY
qf9d4UvpClUiuC7I9kMciv7OtLyvUpzb6sBKG5UcPNgB7mtByYpKz3CINO8BFT32
TCidAJiS1oRDhcr2P573OykfxYWhin+Ip+WUcq4tnFeJ9DpNT8F4TyaA/xAFeYoR
lsMEQ7nox6W/skUlyozxGVG0rUiNRluteAB/zFZ87L9OW/eGjRxt8FIFEf/vth+s
D6Lf9x+3m7sn4eTRQTiwK3Tu7fEk+DXIgieBKj+eHrfbK4nOjSWBVetZoFHkgRtV
Hiyw1drLUBfj/FVej2e1m2zpIXBufZJvuVf/il7/sZSQpS3PIZ/TLBlR9aDMwu2c
iYkX/CL1+tUsSMmeOl0Gc4/KMtGjauN7abHt0+so/h1qqfcx4fLWbE4aYnvKh6J4
jaIqdZ/YaeQvzGhOcNFutxAHALN7fVkLdj3LmmCIDV7GXyMVAab0r7lF3LSEPVQJ
zlnRgL18BE9VDGmCtkzRit+CKx8O0U3MmtLLmv1x6thX42enJKjFyBDyRts8K33W
8xnhV7qn8m/L+zObftgv6z5fPx8usGz97FXkcaJgfHslUyPvFVO/I07Dp0pP5Ecx
5EmgN5KYWv1MDA1gijX2M1CgEAzF3v9y9eUXFXcgXCvxqHvLrm/K7Ku1aM+UP++q
DSpDEcxgwx3KaFRF/5/esmW1mLimUY3GruBiHdEGq2acPoeEMnbTB185PZ+Qj7BZ
qUyyhVOcSIbN6vxp/Eq6iIwr/xR0yucJjPmE8l4mk2oTTnluQD3Ku2Jr9jf142rt
vpBecl24kJzJJh2aZdSmJGt1DAk9rUo4Y/sQHxKUBik+S7aZlA+iCk8qRSEgWGuU
1KJPv8asrlnzTwv25TVM6UURsYfPGDu41mw5G8n5AGAAsRe3V6K5dIsJxtCkgSqP
20j0FGWoMWYsaH9TG2/z7MPLw7bZ5+c3N3EX99lRxF2eLl+yHd8IxXLdW1oO3mUC
pDCKTUy8TpiM9Vk9M3KJgR5tJw6owDqQdDSi5krXTM8eONszjiazqeRamQ8HN5lY
2iOyiaPvh9lzPv5xOxYSvPeh+pUGVzKOv9kUsq0wkDgaDVgs4xYnIxmQWy2pF7xV
EjprXGMhcriqDPcdv2sh3eIQDCSf9eC2NhSZC+fuYyNHnUN1Y7/S2S+m56chbY0N
Z64lf/Ta3qt0OXo8TaLXSWKPYmWCqHybfIAGr3fucNLG/QG02XO14ws6XdxfoSfn
3HSSVx0RtL44m0RpQS9O6hLxT2eiV5lAMXY9VCy24juVZlLKFufl3HtiipQORe0w
EwVBe/8/k2aWXdPL1MiJF8tJ9w23yxdnSisaTEW6R4U46JiPXW300rz1f2J0GLBw
rS1VQdkIhQYNR7+ZWMqOkrwdPDqTfAEpXtz4fs2cnJ2yP82gTpqp3zXy9u7F1olQ
TI0fWqBmJh22CCpP8ia+v29mqhJkvMMofuFDdkTPUjTzJDU23GQZe1PFNfAUuipE
OGvI/m7aSA4pNlO4W5cHq63qu0ui0VLg4JOn8J+QP6tLYgb8EA6atVoTcetAvGVi
8Dm1qajyMo7Wmd7qMIe+djcOFS0YGdwo7yVAmij3hGrPTLBZePbR+CvYoQ16BPsK
YzqzPKYCdapb8BJMmBKPdOp5x1Sb2OrBxXtFwy3j5X/S5mJwsmZ6KkUfPRRjY4DF
Xlw5k09BC4g82cGK4N4ujBuUQ/0WjQ1+sjytPOI76fTZDwhOQHNyjbXrEUXiJykE
dl5K2dZH7UFg6s2mbpT/LHzkZQ9SwMRe6IW/SqizKMFS+6yl6dZr74qf2vKL0Obm
nzIRZmKO9OXHhM9cDojYRFSCSmKDH7ieaUd9nMyE+rQFNZKz/gxGVVi3BDF3og12
R6fJIXuFMvo2K8qAOBgcFbbhfTXNftJdm/BKXu8rn8msC2LVxM05MqCxjO56/lA6
+ZojF0zu5d8vNIKQ/SI8UW5KjzTu4OU9K0T7j7EmU65Mdlnz4cjfaOsl+3A7Ol3l
uf3f8W8XpjyEakAVl7m2QT4TELZkFrZGjQkWthd6OYIr37cqraQ+JtuummrSuN2m
teduedlVJq+ySshCig1aj1r6EjmOdpZ5U/hm2YVCfeMLvxHqepvr6+QUWAVIMdKJ
3xQBef+LBsclQgGUbcJWvY/okvTtjHTy1+4q0woNmVPK60hm+/IwVAuRvcmC17Nl
T+qz8few7egtMLKK21xaaRv95PSwcOeURL++sDs4sGWLbY6tSzLa0nIDCvOebr+B
TUivwMWB3yXkataMP+E0EraKGrWtgxBM+/60gk2vQ+Gn9b5fnosF/HXf7ny2AQfo
s41fQE+VIrefL48q8H1SFIv9nhBx/vFJXEYCpjZX0xXasodg1C9KkMDhUptLhLK1
hLJAz2HChOtYhA3/3M1p7RUIN6VHzL/4P23sXz+/NcG4GkCob5yF3D3/xLAl01kc
7L3zwmC7KPoW7vEZTCfHGCfgrqGeWFkBFED9KlmxBX0wMJYxrTExjtn0+GcAIq5J
qLR6ghnRvftgTU2q4/Ah4ByqrlOn/vrlB3WFsZxsoWE9RHHnnlojRQpaINL933Cl
sx7W5tBYhXqc7hRQwieIH3eT3HZPw+dF/AghVHnSyrHgh/E5/Sr5pJJIVPcAjqQE
qei2nHHXm4qmv6SXxUGkuXSYOzU2V6DS59sI6cVw34vNvfsgk+jWQQqqDE1GvCH/
tYLVAewwYanJF87Bg+TvfF6VYxP/vw/RbX+gy5FKs6Bb1JlVnOzSVUJSg5NmGOAc
U0ghXgTKSHSBbKg/r4uI6zCWkkBmVAy+azpIbov57WOM71Lyf43LuX2KmuSgfqYM
rZxZE7ukAqzApu29MGSmmKpHqIirvPs1IOq2/prS+8lQEYILnZ9vAigRsQdZNq+U
KX2w8akmZcNDY+wJoj2o+THBy38aWoJWfmvuWc0Znvcby0qqFMdbysXS4E486zOK
maUeAt07wyJmX2BUWrZ/1kmJUtLc1dJanhX2WdVQhabUqz2eJLvzcG9Vccg+27bV
WgqNFXIjjwBjSDE+YxjxmsG2g/IEHbsjWgcs6UHjw1XqyDo7mFz64ZE0rdfNIVPr
KZk5ymiUol6hCgh9HuvFxiugq0HNnh2diUmTe3B9epf0JylQWOkg05lMytQuIe88
Py2PkGFMSF2+t7yka69qHhJ/FpnWIl2qnz1VgIeFxZXs2bcj2MML2IZSEzTxdpmq
K8q1ITwM2t3fkm+DB1YyBgm9EoQAmhQ1mRrk1o/C5y27RaMs1tdtMz11L5bX4FD5
+nfdsKxa8vWJuEVumqM9eXkvJzbBYu45cGeQ+s0bdQ9ZST0mUI27ueGEv6uavgXg
QMubg0MMYB/rDSPtsO6yz4GlmB8EJTtqkewdrQSkW0oKKi4zoTo/vOVONf/fdXfs
bHF8WyFWhZHbLzHmMB2jFRROecnjmNdLsfQcKdQgp+6Wz696brU0F4z/oIDChAyx
O1VxeZaVdoVAtLmxckfyn5fRFar4Rwgw5K6pVj+bf262ZJF4uPv2yIt2u8es2FCc
XF6z3vtDnDpCWWC7hRO8HTnvGlXRTpAmEFoLJHlzdkTW/UOwvxnEZwpGw3IvaijR
gBh1q4zSTym+kvE37P2b4b02V8d342KLKIUyi188yFVgEZKgjlE3FdJj0yuKetlL
fAl/PE6+d+8R9FmGMbzAtcaG0jIXslv0k02yDFISFM2Kdh6Fb6oVSECizY+wcf2G
5bdS/Zqt5OqynUn8i+S9DTID6fVIeahvVav77JsM/x00WO2hu8GI2+DB4xL1YbIu
zyJpYNz/cY1NKe2POo5n+BGz3snSEGcDB4RcTn23u7ceiTz/jiJMG7Ha4b9Dd5C6
o5M9EO7RnHivj3xBDfwN4YWeu9a1cWwMxviQdRZj+9yWkD5Ioyt9JDV9Fisw7yY2
qYiiGCiSlARb8cMskfHDko0YbafD38vRk8E9AAa1ooLb2TOn+RLhxgSYu3JdfH3w
GnvKh6MNsfIV4veLxotAixQMIQ5bjRdI6baJGK4GvTaNXkcVi7gTe4ogvhE35bVF
7tuJLPsDk9l5e9A9qSAlN1IVC0vgIdJ6QTR0B01CF8NgeKGwmZR4tKfny1fm/8rv
xQM5GK6LiXI8MPlqYxNvuamf3dmZTTpNxqpCGhGQwCrJtGx8gONMJ8xgHkCRW+Aw
YKnHcQO1yH3yFxuREWemNvZ1DEOONHyIphZlIjFEBEHMDUk7DzHn4adUm1BG14ZO
i5en1hlD5WLDzbRPXld+3ByE4mXnxeDXJnqMl+jj3RLMMlERsWR0h4tB58U4KHrT
dY3Th5O5GQCPIbZospi1XQoHDDFIibuQckwTM+6B0ZnUdZ/MH8xJzOFg5dQ3bGHz
DcNbBHfPuIT6ZzgUxE15OfpJ2L+/imL4jXdt4a0pfTzJ3EBjCiZBuzF7bQ7KChhw
JY2wuxsmpvrPz/hJbM7zLROayPqNB8iaj3RPO4JYy4nDy7mCQUqiLk1FoliaawZ7
Bmc1WDHhF9mduxxEZgNqRueA+1u69hNS+PaHmDV/98Qk+2a8FdbZ5b7dboC8/xGN
TNR9LoYRZO05oeqccy3tKFQOn3TkbuJpIA5x2tdwDPGc2KbB7dMjMUL1qpVWXvbN
0d3CWX2ZL2EFcAQtGeKOUqrS1eiyoYGPbH5gDLgqN8I0g6UM4mj/4STW+daYvu0k
FE1ALFdx3vGrAiK6omrEgyiUYxSV8GTsGRai41/7MQLRLBckmYEizFZqORa3GVOE
/JPR7A5Ra3gMzgsWRKkHjXqsqTCqhi0oEBvGbYJAbN159/HNR+a/Y3IUm2BVCoLw
jpnYJl78cgjwYDpCQ/w6smBNIR449ythK2TQv+mUhr1GaBV6NpRwIdqsLu8H5RML
vUnDi511cvucoy1kM8zv5t5r7uSJ4VKRB4YCBYxAyqUINZBxG961koEtVLN0kSKG
RJGpOcYy6i9XWaCLkqdis6Umjg5d2veb26aJgt9QaGQAACSWoHzpGvM1aAcnfg4H
Ale60qVUD8admi0MtiLHJAF64k9hJsI2/2GnSSN0tv6VLViOZe4lIP/UVPviP4AZ
FAqQB1SQVM922b1KxPK/9SWLtscR4AyAHu/yvpy04xsLYGf8kVGDL7TciwibKVG0
5eGv7zixlQMq6nuAsKZY6JUg2B17se1JB+L8qHjEHH8EbOaJ7ybFqVqHpKNRYxL/
NqJRfhPLTNQctQc2rgAX9WoG0gevpckFOD2fpT/akA7nYYDQKNHgkvKo5jOpu+s5
otLvuGX2lFstaC8WkX/XLPot0XUOJjPQmU20UP0p9t0OoX1Z8czdMWtMm0zL2R+t
xFGQb9A1zj4vbNec2gl0qWWr27RLqQL2WzQH7R/CQ0koTm6KX4D3gPfU0irFVl1P
/vBuAh9q0wH5RGmKiE3mbEvUz+JCgswu8ehcseG5xPxxM25Y9l2KAq5S2j+V76Xi
Fspsf15wZZUWDYkSXeScJDelA+xXybYrEir7C6upUO0ihbRtQFDQHaHIXui3JCCM
EC6qrtATrybvb3AkjGPrTdAefoSxc88Ltsbl3LsRcDFSVtOIJTWuiveJfB1nmrIn
OGphMfEOblpR++BkK/qj4zsOODKd84JAK+ug8BwK/wvn/pm9+20EKnoTLkOp3TJh
qUGg4MsPheMAbba1GJkqQLyKC84WoofLFmOwsILJZzyoMbl5AAb/gIhDqKpOxzpp
GsYe7kSG2G1CJmG7QUVzKRtnnylbW1sLfY8X0VDbBQO0s9oGpO1cS68TuBgShHfT
3PB2bfQI54g42xZoPMWQPK77L07ojCu07lcAgUj7PU4oTLxCAUdzfIcNVdEhwjb/
n7QMXTOfa6u5QaBzqgVxGW2IVAQCYZsdgY7cKCK3HrR39Ku6x+W6xqaEUCVNe7ig
3ORDvdqf60kuZ6tU5H9UfEW5OIwryNIwULgbx40zkJ083c9M8l4kQS/mWXNTj/CG
QfrAPNIZ39Ynfw8f2N+lI480qIKU5picevFA+ah6Fixl0PZGhVKZZGkhp4jflCiv
3LTotJv2MOlSmdVujIxWLzxKA43TZIQSMSBAlbctWAMcZjBMJXuEkfGwBqi6ieEz
Gl24XCzN44YHWVB2rOjCw6VTSuoemo7GR2VFFQLgWAD89ygXoNhPlVwkwJiqnW74
53QrjBOU28Y2vR7dRJoDO5JtmxSICzX/NmlDTbKuMrK0LKCo2RionJOqBI2IRLGn
Ka/GQXD2wUBaIkKSYbrwTUGr9bmoy7QvmY9hBPKvxqYtoxlilD05E04aZ207GfiV
BD2KqhUxfTAC68/UFqNMVINp5ESEFmETLO/jwpjStd8swtQ6J/YW2Ak3KiBl7fmy
LbovdWzLE3AznlpKUG3GKU9K4y0I7i4kfPrwOq0O5UAIUovJu3EaNVf6t/FTupYa
PdePs9vu+Ri3QRrWslzRARuGnqq2aD2QUsA9EWgYHxN+P4YLCYW7bR4SGEeMi7rS
zOGqyJ2rAnXS+mixAVu3EfYRR5ChTzG8LFP6r44+5Ka6jTSscMfpB3VUs5X1fLXW
JyVQAz/jis9czx6WCdfBCkDzqNcjvUmHCwcChMYtzGz+LGASILxjDvVvi/RYNRfh
3JaQx2KOyIRkNUOdSBkWqu5yn2LMVittLmu7130yRCTgxdCS3rzkWjfKE/I8cFRA
ndwvfF9qMLvF1FwPeg3OdTbTSvaQ8oBEmygOQd8LpY36pVGq3jbBQ/+3LIcmiseX
9Suoc/A/jnCDAF9Z5wyYRxdIGMtR3LbUhnV6uuL7TxxWmyTGsi9oaU14gaUDDHb8
TD3gsXJ61tCxZD0bILgxQ1ySMe9FADSce4uXScimViCeXxRb4bYHMX5e5iEsTXLI
xkMd3JUhNsJuwCEHo31OaMpn1PdkoJ1I9k1Rf+ahxXyTT/5iqenwIeJqE2NfGYlK
gjrHUo9m4PdGyQwubfsWKVprPEY5mrAKP0jusXLbiPyFnLwa4wzPv1C972w0+zrG
w+eqzwBOKxseBv009QvJVmOGOkk0HAfjHEcvXEdF1mHLGYzQCu32YrhGbWeAtnu8
sBoYM5mKf7Z8t+WuCPctOP0O1YQunTIh1i0OydyG65SQWNM6cvlliVPijHml23CY
Ts6qoBW1q87DufnzUwjseMKu9COwm6bItE6zcrLsJijxSBsgE0x1XIaVuDbt2OgX
abMN2rm0yHFklhCUaOxhHrMR4EurglFBC9BF+AQrvFn1S0ZqCjznGWTNcjRJR4Vg
6YNA3duzAyHXuPA2Q8RmJlDMlcYQH3pUxzFCWeo9DZB9sqAu7vdhvMvEa0RSfz15
jQsE6Bv4IYafNTSCo+LgksJL1OTroGVLpIyVcm6W2VeQEZzjX7U7CJaKJzLKqsWz
3OyvZ+Ty7F6XCsJJntdxQ4u1k7nA42mdJZhRMzr1xJzw3uJtMoym2ScRMUPyREHl
5kWuHZ8ZiOW1VyCUAjEoRX8oDHedFDM7flWxhIAeDI59CXBKJ5mF7R6ncX8vL18c
g6Lhw9tndpaXSkymObCnfHoumPiiA1XgtZuqDZLREJ5QEjScaWxi/pF01+q49j6L
cRSuaRxXDS47TLopw82piAuxjLY3TkYmEvb4IgLeHi+3AE0VtDp7mRWxhCD+F2Dm
V0QiR+5+0jiyqIP80t7RQak2dd+eWpFcaE1IvOGhf9svZP/L1OF/4xPqFGXfdGiU
14Pnuvf3anWkbnXYp08fUA3U8brlEENmVst/ohLf1PbIXBBPjdIjUY65tpDi+qVf
2sOPb9XPIM2dpWD3y4m2FGuf7x4bzD+lNJZtqnorQcRvpkp9RqcO2kX+nKl4tU8s
D2K68UOAXCcytsaV1vBCtk/O73Y2olpMwd9HAJwTW3URcpT39V6IYR0LEk0MJ49l
e2c2Ai7+r2cdz60WP7NO3ltAGy6/oXzZcPOErzatskloonXJljeZ6EbBy9DvK2Ba
FXCZ44clI+NB1tDivlB9jEougyBdvlCYv5tBXR9r0rKXqGUWv1G7vKsThmNzkedm
dMq88C7yAaRoBMdJWl1fEKWVKWEIsaknqeEOs3X40aRovFJuKdzqyYWlWV/lPX2l
b/qZKYWNm6ONAoaqqBoavBXN6A9cV//a/G2Axufr/AFUdyWSljMv2PPobQmy+aMz
qaTOKHQJoWbBnk/D8Ylv5Mi2IMJYCWFur24AzQp0uDm5ugCzov0l7Wf5pStJPyrK
LD6oNZidu/w2RtfvYW7eprtMmj44e6QUuxpJ4PXTwJLTjGy90uLx/OZ/4rc9L8E5
7YABgwj/sH+E5fB3lHQtu35ZZNSzoOJpwfcpIf8JckFZ5+I/MzF8OuMNOy0iSIEG
yFwTqYXfd+esNBwb+wES3LbUiETjHNoz1s2rZuaQ1somFSyW3X/DoxYoOJzXYhy3
bfB3vcNHTWHoblK78HxKHxy/Cw00u3sqEzk62J1mE2oAWRgJ8Th8+HL+fhfkwtMn
jM7Wqv3/GHl/QTJT48wl8+Ux8wvjtQl04SohsUaCuPVOITZ5Mw3W6ugbeAd/SJcV
t9ourQ44wWdo35SJp/xvd7fk2y/QbfcO0xECJnHU5TeWg8w3do+koCpPnt8eQmaY
au5HIOteD3+UwRom4xvpa9wJdHvMww4HB90zaK93jWY9NQZ3M9oHpjAR1Xub6UTx
1TWyx00jYFC/8WcG7KmJnVYMtLxIc7AjkZHhxgIdjn6OA+14u1fFoxyW7vGVTLdd
Sc8IcPmrLJM8m1pwRTP+ntD1rlNNNWztmywJ1v3QgUNhVnCWLQgOWKmq+JzzW+V4
fHsI65mNE7qbTJaGpt5ia9okhYZyOHrti4U+mHDzbL18KFMvYN2EidbJjepCdQhK
qQgFYHXWZbfBTdOe+Bz5aVhD0cu2sZlv6c/fcIR7IbY8x5tOEXSWVhsV+SrDLrlb
9r2eDSUVUJA4/lwzAAY6GWKXZpOc907h+JrhhM5GDvXMZK7DHinYvtcR17ZmcClm
Cycn44ZalNaKFSGNLLYsRAZu3l0YiLUwOU8ICbOQ8xR2f0ZsPmwRKyNgnM99f/8P
LLh25WlrC3AiuA9GY6zxQqvVN5VHGagWrD6nHn3HQGb2aRU8y81eMLODHWyQ9S+P
iPKG83+0Ky5QYOTnXJUp2xnrqp+uO9Myt2HfHOOF3qz3hqy+MhEB2XmfwnTLpsyS
fh5WVSHJt/BmqR8741D6dJck5ULhbgQ8cfBupkX6P4hILOV8B0zbHj9P/KPYPt+G
lu3D07l3rjAiglm8CsatRwNZg0NzOn4T+rRdwjqz3ysLttYeem9fiz2g33MH+RZc
NkDUl6qi69v7oOEIbB9AOt/EVKZ4Z4oQbuTjGNtM9PjU3/Szd+e3QT/9GB8mAGzu
i3w0TpeneC84p7Ycb4W7/3Dyqu8GRt+MEsT2BZwnIDoneYMNTdLoj3yazh80JtvN
2z/L5KXWGOtlOgnE5nz74sGlTWPUYdUzd8b+u5VETbVcxLQgx7+VWFkacyXNfJET
x92fZklDIxYbMyBZLqmLi6/hFhUPnZeuKCG9VQye1uUSkZtPU7+Bb3+fJxVSF99e
fAEWmMpMWSmZbVn8cSjEL1dZZKan4fN1up6MO/glQ6Eq2QNeMw8RiFJFPG+9r5SG
rJfP5At3rBnbaYZ9ANtXD5bhqJfjR7+TH4c9Hx50F7mWdnQfrczLFXJm0pShBbm4
YaEsA9/PwfJA9NiQd3IWn9ImlC3JyMBgv1FaxGiCQzA9XPNeo5OhqqZmVGGsPSyw
3q4dWm8SWZfe+NSFJKPLYRCWyagx2CB85kTmYTFXTav0n2EP4bhxYicKi021YbFq
Ec2u//9RzqrZY923zS5hgHmiQ9Yt8yTBsA94P3W45ANhpgiOd7iKd73wb1lXTtM6
EmdVhobtvyfTiaZIutwCPrB78N0QG5c4JF8Cq8ULj9b0XbqI6nN0JFw5DDcG4MQs
61S+kwGbsgf7foj2F+Q+2E8b46erbcy5GOEcZh4fGnEEB3fN5pZg6Hs+6s7rL0lb
k7cvs9gpafRX4mheCVcYd5fyMieOb3m0yGijyRmB8LxPCYa8n0uA5mATfZGGTSt5
qjgSuVZ71M8DwryXErKJebEpx4dIp01EBnwk/UhAdlSoP9n05GP1H2hls2QJUCMx
exlNx3S48WwSuzSCkg8X2qwpyKijaHDmwVltusWSwEUQPrn4byzcoY6uiDRtWKXc
xtMjfrQojnqP7sAXG5ukeuYa8s7MVnUfqxiAtV6/Mhof/zw/00zo4I40jII541xF
0IMthbMXKZ0X6dsn2alpJHZwy8K5dL5UZxfKDYQahL+6X9pRNuonF8coY9Mba82p
2XDphwQGcqPx0lmxoRFk6+YXxbAXC7QXwC5YaVek4FYOuHKMRqGOBKp/469yO+0M
rkHv2fIcTmtgCwh785u17QWJLKY7lsqnHY1wbsXcBT28GvxaXXeJ77yDhI/G78Bn
Wxgy9TWRbNz11ClD2kyITYMtVgWV+dcAYDBSI9N+UFneDenVgmY5cbWJS+b0ZwVF
SIG5KG3MiV7SMAGN4ThnYMieZtnk+915PMUUoRwhNSQFjSM6KTmc7FzBqVpv9Kgn
WfftidDA6dEymRibOM/Lalixh4OlJEQUcAPHpAhzcMLCc1LZYDmDdCorCPr5cayn
HF0f8fHRTHdsvaxxWFUc3X+BTcxAVoLpCcI35wY8FrIxtzBJfjw6Fb99PjxlG2pE
bbrN8va5BhLjAYPDwnLv7fHeS0If6xmgc7K5a8yfH+iLny9IsVwBFJ0jA1DvcxXM
kjGOCqfBEt5WRxaFL/4imPPaG0iz6kpz7/iewZX6UhTdA2FwckcEpLLxn8apg23g
5WgAg0EFCsilHSnXsZ8WQEgD5WIaOVeHS930+Ld0aGaYBPjzCW4ZczfPLJied4Ju
DNNxaS8rLTpxY+4b/SvgcJKbaHy602QbSm7rqyD/jG+ik3fiSMtQxyMVaTF3wRf1
FQ4zWhrKfHirbEI8j+WenFasgqbDA7cLXb/zgpEPMRifnCmtnbsGLDY4EvDHUqFf
YOcAskd+LplVZQTUasNKake0Gvg8Fk9q1oVpqgVBU0iFA6jI1kBNPlgtFSfvb0A9
YZH2QuSEeao9t952UOu4Tnf9hDQx9tH3V58Y7o39FiqnuA8XKBWBlbMIOne84ia0
l3wQipnNDjfvoEkJ2MGcjAehq+VW+0/QWKqldYV3ssTGummRIO+M4ArBLePR5lQs
NDC+Ge6RttkIqKgunJgPU8qjlKTbEiabbRPw4yHXqXcxvqYNZXXzsPIwIn28Npi/
Ol72XQ5jWDqm8/iavBN1J4WQZQ6Av0pHx681c1hoLR5v8iggliCa8BlYY7oXAKVk
4G6Lc+CDF14DhKvv4GF7QdWcaWelRDsJBwZ6OrN+EOoB3LfmyXVIX9tn4yUCGQPH
ZbscQqe8b2/CtZPpOTRjiYF5s5cciRK7EpTkQDsS/p49EatVaEoHqVoIgcSY+m0V
yO9WYyYRXiOINHFsYoVnuSamR9muyIFOfrJGmQaiOof5HYtxHOMVqkgO4ZgGrOj6
qpjGkt9Ma2wjsNfvfmz1TCtz8TY6NfGYT8IXQRk1xboZJEBZ1hl2qpt5kk7r3D1c
Zdrjbwa2l8ykRpCnvRFh/pAXNXU25T6qe+IYWolCmcEXjAjFVN+t4uJLQTql62si
JgQ8i0S/vZDcmzg1Tn0EP1rDJCi23bwT3XPrcu2djBVX02rX4rK+LHcmMgWKhhFn
GxIHmTo1qOFiNWltofjzT4fX+5D9v6wrlhiO1JbXN3jf+XCnzchwhMtWKI14WeNk
CJiXFfO1bjKNw4zrQiPDcClxs9ARbMGNDdWwu5upigtn7f0fvGjplIq0q0ad6eM0
jIAGKNFEnFrFPni3WoGTNUkct8YU1Z8/vcPamwR5qQTB3LX0yhQP1M8NZjytOPjU
k8aIkHBkvMLW5cT/NpIEJtkLm53lNufRmgmMXwnpHqB0VTopGrlhQ/RA4eilFVic
LPGig/v4JEHCzHYutuuYQBoloigo7vG5Uptbyxjasz7s1akQxdv7ee9n5OnwA+/V
dzPnU9PfX9J8RQmuZoIbO5Nd58qSGOL3voPFVtkFjVOmQcHMY+kSnb/b3J7DLuIn
heGUFjorI3KqjRUQ/9JiC6n3Zkad0G80oK8pkgwC0lVHlYl+x8MTzyozwQBFQcGQ
TttilgyKGlktctnR8CAyMNA0NdxSPNY6KOed0uWDWbs44b48v/Z1itdfPjBe5eC4
TNdijn0fx+UKQvrgVouVMgwo/bYjrWsSeTKToPL/TI1W4wZzdzyMn756z2aoveLg
UA+AAte0kNTQxbzYkKKrPOErrSn+EX4H90JksAHzhgbRYr6hiiDyNoATWlbMQvJd
BcSFh6LfEbUD4ZPXfsBZqCRgaHfAYOONg0usuzEhblziHcPUlC2qmoU5tvGQBbsT
46WUk7+78xZjNzkYabw0m94kxCxhWzP+coZ+4qCLZbOgnBvmbyN+Auq1ztY88i1O
oGbX/e+jWWIktdCp/R1CCYjT+DqxsjG87A/tycgScdHai97t4HqeXyh0tQXl6jor
n7eNGaz4TBLl/8ulIET0a9mcmY6PiPugsXLpmJFsShdILi1PZ4SIr016mFJmUz6P
kSP0Q0lMcXJDL1/wGkAmtdhQMhwOXJsG4Elh7vZN30dKGM7+Emyl0T3OMAY/aMX2
mpOphOEkUdSWq1fAZ8j2wMDE5l+6yFb7ZtcwGvhmr3W2wxxKsWKDGzr2ba9Rgqwx
o0EjnLbMLWgrq54oZIna8/U8dvcKqG3wD4Ek3feFcNd8tGxMfMF0Nhd8OmHy9rgL
1Xw39JJWrUIbLaDnFU78tReHmykCgnYENAh6jQAFyCCB916SY9Dp6orjqgsisndW
yUxq0M3EiHlavoMHjWhYkTlH1QzqSL6H0D5D90gOEQsjC5egkcmNkMT+YagoDN4L
L24rawoZAl2v+aOq+C2ZYWcxnvHdcbNIsxh+1UnrlfHKYSrvB9jKsM2D1gAlleRs
2jpUpYUf92JxOOv61nLIR3J/6h1g6CX6HIChCglxsiBkqLbbxA4oRf5nsHqH1Cmz
+2rXlN+npoSaL0n4xjT0o1mXCwOKm6SlypbV67LTQFzaivHD8Iabxf59ykrIs+ex
ZQPWMNGE6/i+XuoLV1xBnSGjWgOZUh6rX3Lye6tFHNouGdhRVQJGGyJcHDlmauYs
nOtSRdt+I3mtE6qtcKTJfMOUDyRWPVrnmQAHqNc8uAEwiILuKZDd8osZmWzE5KZL
FXWVPrYdf0UIN3EowhitIQLCHUffSeI3AixkYQzqlSq2wSezufhZFKa/nYxM0NOv
MfEsuu//dQLISVuyc5ne/M9CJ+aHRmW5zMKPTEQqMnvYD3a1Gjw81lh4HBD3HVKp
WjC6YLKlL26rBynHV+dwjk8893iejHRqJan0yjIbKQdAuE8K/jHBVBc0n+FTv3jE
ldMdmFEe8t7lnKWUN0KDL2c5jbOsE97Kq0bueXM2+dxj+/FTdNaIeYNMtjjtsY8n
Jj+iswpqsZyxuwQi/HUBNtJuKuAoTiQhsbVeBo4Vtv1Oh6nxZxLq9+y3ohGuaKTm
DcIyiC94SXXWppaYbgtMz2Y0gG/M3zoyHVkBp50ItROuwN3M+dEpPHdg75IsJOfk
L18jCGlORJq0XlsUHiYWjFXLc3n4bRlRlXI+RvK+dUs1YZQLZ0d9ICOfYvN7WpRs
q/hTaddnwM42Iz0szN/bCFcdqoTyDP62+BIH0bo3FQ8McR5KR6tWlloQDiSvtVAr
xE2HClUmkOOYT+4ZFq2w89nXVSlBaYL2GfrfEhZMzfKlSxNKMI3xrBHPJEwQdHmA
DQYpR5n+RuVIfLYaXIRi+oaoEp49tDCYkIOZfwr415szVo0pbQ/ZgBrz3/UcIJFt
A5Zi0PwpVtN18cxuEzrO6HMXDrI3l1HWUpoBqLD3b56D487alSkD0bh4Jq6Tv25j
eVIz20mjS1Aa76+nTwJhnuXthnlvkLtL6TparQxUgT+Z6srWrBH9HxgAj2M6rg8A
5xGzJMPb7LhOZJUNOGiYDun2gYrQz8AulCYWC+MtAyk65qgd7PDWwJrEzJ2kXMUV
a3eM1HBrVCnhewnT7OWkWTcZZpNFLSx6C3g0fPP9K7Ipe3FXROdwJtIn/ZiYrCjw
65hvxDBABB8edTzzEeZ3RVfm2HCHiuFuFqkG26NbUJQ+0sCQoe9hDjgGtIP0CbxV
1ozUr3ynJirUtch2t8N+UXrLUhQNvAWhXiAol7crUZJ2iOGYoKuhYI1aJ6CHNDBw
asFmgDhMGmfM/2zuZwwBJYMiCAjSJg0soF49vHPgdkSf7Xs6YeyHU5hBApx/0jJl
IiEXP/ap5zmezHdyBmKwyTgPWLZvWMjBmzbPnZIJmorQJryfIzRAPvXk6IOlAhYq
1CASqqAg7RudfM4400txUZSd9MIBlGICgYGmzRLvrz5lSphr9Y/7Gj/iVsJOJOjo
iVjP2srTtjoQ2X+4I6i8G2xakV7o1SdtBcGA6Y8Pk5e7RUBJYODqNlCbnYsRjpTV
9cVfksds8QMZdas2db3J6LLLR8MhUFHFoJCYIAJZEva1CFAbOYTHNNtbPsbYKe7S
h4rHFDEqyiAJffP+tHqVitVGgRiMMG5qrxpoGgDB1NWe3XhAhhnPQf1C3NIOFfeH
L4ruZwtetO9sp+7X1BBQOle79+0qY8rTQzYhAhjqcw9CKX5dSUtBq/vm+83ENdkb
9gaTnMMJPhMpy+WksdyVQURQHHBeAGIV0S8k0qUnBFfdJ0XVjIAGAFcYKEKm1Ah/
wXmgQctbv6G28NO4asHflt9fnJJ3YgEnAF5XbGLL4AxYZMbl9CPdOMa6eUK+IyYx
OOWGT5uQc7wx3dETZXj40E/wkjeusCBLPzboyqL/7URLGnhjL5sIpiWgtESUKwyb
0AL9yaIQlwM4Ms9SN/vZHjeBKIVrmlOFtpb1SwPgVGtTwi0n47re9dt3ztehk9NK
4WfI7ZyN/z1dNU4JWmIkj2T1sZLWBz1aCXCP3XBnniJk9BiKRHr8Krcd6PFIXLpH
q/ZIWGCOzR5GJu+qHW+ujmoygtwEpcxtnO3aFa0HQd8Q8brM8r6+HnCtO2dqhRIO
j/Q9/rTsFTi26i4cg5fSp1aXTN8I7F5hn7wLdhzCbaImpeCYGh+OzTI/ou3Fd66j
W5LGggoxOH0hanXcnixvsa4aiVdfYmbtkVPgFmo1c4pSrCg7w6WMZ9/K/CBys4ey
KURFJWs7XqHm7KoUOt1aqmj3idxt/wfqEeYudLWBk/rG9c0X6Xux7730VM9cSlyk
WJs1HD3+DVeMl3Hd5B11vjNc4UbmYSG2Yy89df9ji/YAx4f7b7mrwgvRoiuRkd56
isBTdzJkswukkEfzIUY0bkASTrJLQFC2hxCN9qFPQWOn9c29UjlENUZGPbfVF3L2
hofUkSQn4gyhW7QKTOMUC2AFfE/q+dOgBstaL6jelSnNST6wyr+R1IkCuXdEaKvv
AFIKhhghbjRqC3phikuBrVZ++ag9Ml14ZQuihyBnOWylrDNxmzVYfwB45W4W5FUg
DBs651KM8zOOxvKNtj1fvzVwd5kd7sru+9fjTPKzg+ZOy+jhVprpkc2eh0V8a7HA
5OwLfDBs/bf+wbbhJht4cRAu0c+oqCzckCaEuFt+gM65683g0KcMY60Nia4q+i0O
xGhMO/8n+Yk9TZx4AxYRmsIujHJZlYjl6BMHgrIN9BKwbwjx0Q3bY/KxwUcClQdF
goTnj/fMAaAOdBt6Ooh23rsHPijrqn6+s+NHwjBNEGKSP9WaICqyKpmBXgzyiJNR
SgSXE5ynmcPeQJsIEeUEILC2y0n0Dm0zgSIEd42KXRJ0dRqfq+QUabxF/LtlJ9/t
S96ZTyePTF28qmSBKDi6gcSMQk02COy93xDvZlY8mzikvrJh3GBZ/QHAsWHAA2GZ
LDlEGMDj6j3d5hnuHLcUB0u0pbf3naTAH45p9dex/HYopYGQkRZN6VyFM2I2IqO0
VKAdH9OLuMIkS/WeVvAG2pnzu0vPkJ6MWHpG9UiRcCYR8KrvkqCM8fjqGl+GsZIn
UpE4PeuDg+DESGSWl6Dzldfk4flO2QIekM4/hcevAUm8cJ4JNKW/2Oi2EqOTWFbr
jXbMSSXQO1sPxXhYQQ9orXsIbc67DRuQITFW8LOWfWplCM3UiHrmas3rKCR/McSc
odhJSryqCWWgwFHtB0Om4Oem4rXo50XzLUQJS3hlDF6e32Kv5ANJkRNLBTLZX9E6
KaKJbxCcHveIf+pcxSWtHnphdOosm3UPSY9g6uyW/CfSWa6nph+5og8CmW8KP42I
8DCoODSsoyYllCLI0HA8Vkc3HhtcjYUHuZWwU9jt5ssLp30ylH8qJk+MaWUWp+ZC
2aYVqUJd3rYL4VCx5zTul6wvU0BUugWu4gRXELZbF5CEXGfu7Y707WEBRl+ZYoJQ
QpAReqr9+NOI7higSQfTSr8aeVjzIr6Q/hLf9fYdCW8QhaooRuVui31hXO6f2ijZ
TiERsIpEJ5QwPg+6Vr8koDLdibD1H2NcvU4v8xqjMQuGAvDCqDvwGbghfH2lRfgD
iZKrUGJHJeSP1zL6cDBPCeEqK+U4VKG+V733KQs856+LsmwtI6wqhgaCzh8T/eqy
0dFaFOQyUEQk27VqHnT4Q115OJvqAFUOp8Pa6JC4m+DqNJYA02Fk2oTxb7qrhIgB
45MV8XXPBbBZGd+MjQBlfOaPREWoL+2clgsq9p8kfFpmQAQwaBc6B6WeLIgUpygP
hkGwA9D/EBi0qYNOneKTOL9AV1o32xkJh4FhrugmSyJxB+ajgPYiTyGkh1Y2Gvs0
P/TjHX16eh1dhYeMfARGunZ1TorraDPKGZ3jAbRwdDVIL0R1cO3M10CHgc3Z5Inp
c59/lDd07jVtl3gpEmhfts6BZHbZzs4RxC4mEa/nVv/1pAtszb2nCBitYmkeUfje
Vl87SzRaEr7kXjlFRmGcuh5vXiUNjvjIZnRqpzoOItxPM/gztqkFn8FzjtDZehvG
hEPW4U7RH2Gim/+HdM86lnUkSnT1dq6eTtpAf+WEieJgixSsv3uNnp8zCv76CIAX
liGmLufLtcSUNryYCbgNyVYbICEMf4MPy+pSO9REBYrHFiI6djUdld1wj6Sa71eT
C8seTSkHvOW2Ye9oziUnqnv/JIsjP/BVz6rxPBWJ+gfxSyRgiVoz4x89Fxce+glT
pFno6DD51zKl+XCo0ledquK/7tZ9xhGCPFa9oIO8ev9SnKwthoJeboEmrIFoUgXF
EpOScuC2XqGoVFoT4K3JVCT2X7WIcpQQ2eZv3OlPMjHWlFEPnTynEttUJ815mefz
T83xvppAax+Nbxi5cPI+O4WtymT+aQNXexhXtIctEm/7fqpOjoL73WIK5lvkDQIG
mRbHLqag3VtuRsvbHSpS4BHJcHi2BjuSeDByA2FGSdLjiCNkK/JFi6g5A7WnREvb
meXx04KkBIWci4nCnaL/qpicd8BJ1JWch9s4nqls1A41VLN7kG5+f9NEsbWwp1gg
2HZtMUnSKlthJdWiHtc8hwtVPCVxKc09qmd998IIWKq3RS6vNWABXBmra737IqMx
7+fIeVdFtsux9dqYVDxrrKFMkHJnpU+NaICK086hz7/asknGIj3Y2v6IWiBzKOf3
3njMXtSsaVK7N0ril56Tv+Os+BfQvDU8iegq3Ppl10eZSLrysJk4E1ROtvigyXho
5DeN6i9MnAsApHiJkic5mTLfvu5KxNaCeoAVswCCol0tK+COtnt4skhowc5btzjV
JtsxgiCNNx7O0GDoa16ogO3EAar+oJu6ZsrPSHoxFHV0zkrKzxH3DdVIiaH7QRF6
+TL+vCp9st7O74ThuyMzET6VkdNpkTcGgvRGl/d6yacpBHQ7x/0lByT9JLlN4igS
k/aUNuYcM70TwmAJ/7Wne1ZUjUTBx/9WN5nBPxE3kA+leZrspCcVY8eGD4TuKq0D
rJ4sEZ65UUZe+6r3nE7vRiapVvqF89lpYPfnc46UnTnQx6fplmanIieaYCnawJqU
OkW+UOtPf3iYajGJaYmt2o3loBIfTiwNRW56UZQlXfXFiCehhSnOyJDKhbXVKoqT
Q0imadmOINMIEcKSARWNjZMvHVkqQupm60WkVRWF+qLzilWgy1b6tW2nH9e9MzpF
sjqy2jbDvSN/lSY6aKWGTPCNptQD+G/oQPZtKsh/Uwn3OBSB9urYns8P59rH4hLP
pQoHFhopLVxsiIBzdgrbtVuPCM0d8WWtKIM7ihNn2LI0E/YyCfKQXA5Q/KrtmGMt
bCw6+dy71suyKff65LMxJJT821GQZw5UAix3va36Hf5Ro4CfHLiDm7sMO99yMcPJ
HX9wUFSDx2rXdl2xV7HRxrdfyzCsUJzzUaEc24Du6kKhCC+qG7dTJS5UBtlbcJyq
03P45ys282l63OEftCzCaURNLUTNqW8JoGjxQQjPlfQ3Q4kukXUc5vbf+QHja9Er
b5kyf3dD8aXwsY+x+nXBPt88BSK2hxG0stSMmO8e7e4IkfQwVM9q9iv5L5ynyFhd
WIk2U3aEo22RN8I9sbiYufxdVH61uF4vj6hkv9lNyWX627LmlEk1Oexu4/baPEt9
mWJ0l4zhFCRbD15h03RayOEIwCbngRH0CFbwT44hYf1PhwVtnzPMZAqUMIv4kITF
fQH2eLcGhaLj7UXiMabEb3XUh83QuLfgRtlPN7wx1dwcRREGfz7OAPL4CSwrYbQy
ywikvaxkH5EDQ+9Bh7yx/EC0fXrMKZNNmcqoPDsOiDw34i+tdoEGPCIrVGPjG7IS
YSMtK8mVShxm4wXb27BDshooy8kRrGUIu2VnokUbkWJNi2MW/aph8qJCA/u+hE6x
L/BK4ZOGoCLjvEhq98fvoo53UUEy1GLeoUKQhJXfkRIESjbZy+yhrBl9vvnNzBU8
/XqFOhcy5sHQy8eIlzfAZM0n0I5fEYn99zypIavMtUVMVAJyEN/H2l2ivWMY00b0
kPiakzAeyM+iy6PZaZsYgGPvRqA74z1yfn7mtKahsZ9lurR9S+C0gjfDH0oREqiB
1viyoA7venlSyojEzBdGNBOyPd70mu4saU4z3536SzM5GnaTAFD6Nyz3Impdf3Zd
7smUS+nIiSBJeFlWZBszWIqJmIKWJrE5KpHFsVpa+G0lLm01v3SX4rC2rWDncrnX
DaQuwBclKzGLB9Om8K9/ugfoQ9ENBcr1Te+gG31SuOIfkV90n+V3+sTusKDdIex8
Xek1cnjqf3obxV6e8w9cKgEBprKG9Iq234RyP91QUG6IduiiMf5pEWJFqFpaxZ2H
2kfzucmMxNzzzztGjhSdvIx0Hk4J+v7x/D1ak/B5/OY8Jb0o1DG/EUMoV+WYORNy
MckKrg3ZVwBTKCCUohXwKG6pW1QcKMgeYovdD0m2Ps8sMSqWkREI78UbqDMLUkxL
WSRUS1u+4Lk2KANxPKWMtXqmLUglU6LQqJt4n/XyTBNc2UEj4QhME849GCZQCYlj
EzDASCoWFTzTTcarl44+wX4xY3JrufaC4NOrpNIWroAGiMs7TVUHxsI4t7j98Z4/
7uLJLHOTh9iR5J23BDASZ/VeeBHv53Oe4zwU461OqbC2x9D18FxmIqGvF0vu/Ywz
td1ZFIy6I/s13ziNrPY6M11968d3Vf8Nt2hqfjcFLuOZP6OTAsASrSUlZPrqh2Ff
x9L95G3OE2rpF/TFrDJmosXt7h2jgoiIjXSkLwG/dVn6PPjdylX7+RfEXa/8z6R9
XP1gO2Mu7n7l2tm4TKYfKAp1yFVpV2/O1M61SMkCzWyB5n8wrPOQqDTvB9jnqZgy
41xlXHuU48tScUTijHaCcDfmLu7uSXKeu7aAXkm35pIXf56geRkDRLPhnMcwCxmw
2cWVA5/XJnKhFKHO74v0AnMZA3d/SbPLFXWPwuiDmUb05CyVhorGgmiKzqax1GH5
98cjKZ/PyFwVMxb2GVG6v5jleabdE5g0N6jpasOJmc3IpoXmkrP2qLMyIVaZf4Py
I/A2zonNpQ4ApZsDf9yxGZbIFm41z9iPxgWUj107kVf+j2ngkgFXKlE31VfvEbmx
VVQ4m788MangwzLxd91ppA4LZMr0tQxtawvc5UnxYkNyMIx1y6zJykwDedIE5MsX
vm3axUffFQTya7cPTaNIR9eYknre6dkXK5ltUNIn2tiifRd3gAKFIbmQaXogmJs8
06UKQxyXPwHcsv/9ZkXn16cEapTwMc4hvTXO73H2QXB2GrCfvO4yVKXa5D5DaHol
g1A2H1WH8QYZ1NHNm0vjhd8AhsyJMgLIcLCfXdeKt5dyTS7sWx6XdEdqzXK3/79d
3sIPRCZjBziYLqCZiEk/G5hS+Z4Tm5Ofgk2lDmDr9RKGz9oBNClN37Hw9nufiC/X
MsOI4bSIQcUAGSAGd1IT7VBGbDXuVQHZk0X0tMiewuXDCKBJSk4qHEYL837v/kDi
PrQOtrakKU0DVCBBPIHJGFksTSFS/JpqjLoOkHcc303pExmmIqH/VkA83UjUTgd7
DbjqWNFfgRRokN55O6psQd5W0+bCLBxKAbPAnJ2fefWfkc+YJeQhNuD31NUI5T+m
SLj8yQBJswR+sUjhkmxHGguaaYJ+/Sq+UHTLbK/9nEBaJVyTcWilIexcm2tkkifC
KVJyWakSYryW7wED4b82PhovK5DDduHYBGuo8M/PUuRQtGshF2fddRnnMfvgBOfg
3zvNnknc8WqfZc5f8fKcgf8Y3TAJBUaNhmTQnBoinFE+nQBc9qVGz5zsyrkJI9+O
XaFe0FQar4TkgkHt5UDS7LgEHwD9bP/T2EqiVH92pjcM+7hr+RMUB0ajndlQ/HGp
KMkKSCQG4lspHZ/4ODq5413Z1qb4Q/JhyUNhEaQCHrBTdPTy8wrWk9mCD8s19AGq
rpR7JoJ5Z+9aDjIWUolnuPbCIMN0Xayr9++ZfAIyJtSsjPzONHr5+q+ahbEMnoBh
u0y7+56z5HS5biIiZvR2RXv4mphw3opvJUhytCP1Ls6fd9XFB95WHxPIp9mA6bYk
jIjlXiHOgfxT4Q5fGIrMTyT0ypBqdVeYAB6efUgj49byRZZh8WIxThQvKmV2/7cQ
s8X44haIkAi3/tjFiYykldNobR/nWOSVkBr2yUUCo8iJYMEWKIIDxxIrq7OUFgzl
rnQDCPDOPeh+N0+tlgHZPT8CvOFXegLT3tBsRAzS20o2ioiIggQj4DAKK2ryX6XU
hRUdfxaIDf4yfvPfH6wQ+bg6KKsnQHd157s664pJcA2qzEo6NUP9H56MxnkS7u0K
mjNWucR3R8uK5OTvr4h/KiW1RauH244k48fRGjun1wNZ/vmu0CRqRYDTrPqBDepr
ZgNYDfxh2ktu/tTn1TbhHaLHrGk++9C2LdgVTeBe5Y6AQhgPWNYATd4ogyNRroLh
+H9uemBX1BZFk8TYmhRy2KQGj+txuwMFECMHP9rkV/PEkzWJlDJkRQRyqR/WuTNM
yNjUQDs/tBhqrBVh8PoHXk0JXcy5YkeUEcZAjAC2Haibvc8xGZvS0yd6iCbqfrXw
UEt6YtzKanGijLTp470+MO/s0YDqKuwPxbIZSglvc87Iq/ljMaimu78enKZx+v9x
irKn2OZgYd6xZ9iJ2bHpYmlLeJRXh1LVl017cVumOD0yd4PoiVZjSNNdOWmbRDlr
VvznNJ973lryKIyVg7vP71osEy3mSV4i0zw3lW0SwEfPBGUkmPd8VBEinyqU+dKD
W/E1iQ27yeuEhmQ3fneRPhV8Hu2UqsiKqflZLMHYxob7DdI7yjfsO2ZqEP0s1E2S
pdWVRA+K/CLwtIwZG7gE9rIZNhkA+FTwaUYDQP8tNJiuR2Z3/kwVpuq1Xfo5W9MU
31B4awaSs7dyWijVHFVjV1fiYFvY7Nh9sc28nSK9tU7lGQKo5ZnihqIwIIamKIUz
yPThRZn8eEsMwPd5bEbRAAF74+iq2k91XwDnI+Jr7U1BrlluyHJIM8nOKQ3bHbzJ
XKix+ih4OlUbx4MGqktcrDfRF7PROa77S5cNQgY7Dr9kM+bJR5auV/pPgS0T0OvP
vZSehYhymE2a0NFEoeBhW0skfmP+xwUUH1l4BLkcn91wL6ljUfKk3ZWCdjX7FePm
ff8K1VYjp7dNcsen+DwrtJi0qPXhCF0v9qjm72v7MwgWAK28puPM6x83yMBoEr5+
KqeyIJWNYashP1XYsrYpJQm0vZtdbQnMHHQ/K0PtdTFos7n9fIo6l/Sztp7roKcV
y4tBzKMEFi6YmMM8RehK+BkmsWHU0wIrkKTpOFs0VbaT2BWiyrEVDFGZSFWhhSdp
lzqjl+zDF/DGSkEVze073PWrlLTpCXCx/kCgkZq0Fq89/eleUsGx4215+Cvcxy21
2lJD8UMx8ZzI1bxEhHjgdO/XkQcquTJMhDkkqTibDadLsebKFU+xfKxR39RXbphu
Iy/oClwQaFfv+Y5YY9nAFju30zsqvzwCi98FK6NexABmO67ofia8Mhp/37C/AA+F
jbeOqSBaBAYN8f6n/NBfAQM7ldmwEN0QoeUyrsiNm5SMsGJkrAjS4/29eZp9cCry
p9j6twnbhyI5QSjyRRIoEupV1wNMXGgrEacN6GJ/K2n01gxLfQQDePnVCM+tEpyo
OVVaH2eBaVhW3QCs/UbpUUhnMLXF6eRngtD0Gv9TYeWupGOf8gUS8KwhLaY8CO0P
iWEQ3Xkj11KvYdnxPR3x9A+JZgFsM3fl/nLv1hKKLIkul02opuU8BdnblW3y573l
aQ3WLu/L19ifYNh2zXmlWkMxULvzAmUvDREg2an/OHSJpD3MUBD8Loi4OVrdduVC
KqOo8IL4FvQXWlorz5k8s37TL44If+KpcDE4dnRkgNoL3VvX0O6d1UudMjjG34WI
N27LI0b23pMAmnW0xeVAZghEVo5fSuEBEGZOdUrAY+VbXMoY1t3dWIbBE8599ldC
cmg5HmN5GrEQPxwEHl0RqR14a1jedIBNB0knW6tL9EaGhN15gPKEIK4ey1JNEdPC
2SB6Uh3SxYI4DQ03MBprH1+VnvD3I47+klbUlqLIDcZaVL3SxFRBs9KTC85lYg+1
1fWdLBXdYe7wjYDrYI6Jtb3GYRQ87gmzuBg0CUBfwrNNPVd7VrK0Ao2tcivrX0ZK
GmMAsVWFLepYRouRE5fjwY7MrWOMma99fK9SOpdR+ymirny4686RfzJp1CCILw1F
zdAIrnkGAGurf/oqa9LSIHo8CSMJuvLDrXIXuMOv2iXOO6df0s3KK0e6L6RrVtOk
aZ9iKN09i01U6DSxKztAg3myadpZ8T4R/LhyjLtaetIqGo2U47OrbmGMoTVLmWAZ
pk0ew7onW5vuvdWhun5vpeGXWaigYrcj6F5tQftx/wVvngyBsJyZfJSeUL34OyeP
wDPjhYdXbx3D5OIpQSvEfCxqLGMmCG9+R5LfZ7xzAp0kaoznh3W++2016kU8vz9O
MGE+ptcTFhz3MIIALzvL4v/YE2nw251PljRPPVnZfQscojtqpWGZBHi1guODFPyB
RIOpsozXJAqhX3nDEoXxuf4O0GFBWYG7yKsqTWH6HdRRrn7FRcmswcxUQE0DrIXB
9w+Tt4IufyoFdyDrqoQDv75IX9w3JGfuP6uadfnQjXGOL6a0ZQceFA5uOblsdzU4
cPswyGayS9mEHaIlHg8dpQ84/d5D8++UtH3Nb9YTn1gjW8ws7zMT/uZ/s7CPQ7jT
XvxZNI6K+NgVNJWSm0vdiZ1NFW7WeCqgqgJNOAZF65XP/9HkN/5x4vk1vYFLlbig
6EVEs1yaYszk4fFqGN+3Wjz9dorOfClmktlFCnyvY57DhWTEJlDxVI1Mst+S1RtC
FJ/XZs6SyT/bsExXSwk8ASP1IJNV0X2W74Gd9tAmNL4J1SOfAt99EntHh5X+8bxD
HOWjdUB2o97RsTLZRa07rQCBCJATwnhDghc+BgXO97/tP2vKo9XwXv3y2ttdJNlo
B8mOB3qyxthE838KO9mj+kJu6OLmQ1Rk0GHfH0t4IBW5ynwZXKPt8tiifhTCN+uP
H+dIeawmnJVvVNz8pkkl9V6LrY8HMuFfhSe/AGQ1NpE3VqlIGMCFggR40dJoJfz0
f8dJii90ihK6tTbxR9bhnqjSm3wznN1Edanu0F9Wphzte/4BWEjRbjVafIAI+8PK
yvizWG4ZC2+zf6FUtDtwcs6A9UMXwDpc2X4K+YRlr6sx8PoB7yotcrNeSEJiCYOD
XaLwKEVQxiRYQ9Nte/J8Rtcg4sG4F/ifqnB8f8EWRN1za8ojlfwi2et+48S97vK+
5rxOm1rK4M2cdaJhBhcdE1WnQb3yT0Q6Ec5zdGPBazJNtWKzaMhMwd30WGNUgJYG
iVO2tJIWzks7yLr6ewOg6pOUXice4e/rgC9b1VBPPVI0lJDNI+1Um/BifDmbZQZY
qsAK6RV58GgSZpjCskUryy9zE0kHDazBuroClLz8U6hCKhuq5PYZIhsaiLsOtHND
ME2A71ul+/Ovc/d425UhjKTw24PsUIpfBgbPkwGwDDBeLa/MCon2KSYhio5kDSsT
5JLq12gfmreqLMiWVlGJBB4Jua0REX2h0roiK4qYrqV78ZOWzPiFpr/Mj8W1hk7A
AIoEaHC6arso8MHtfX8o+xORuXcB8hy3y6ra05/zGq8vIz6rak57e5QdyRXkTkRN
uZFV7rdDO97PAjoUKoKTFU5HO0kXUQj/15BOzgP5mcAC+NtNaF73DmDwpH3dn6lK
RQtSeS98d0+2HSZEkVdByv1VLEGb6A47Cl797qwCBysGqaBqSKTi3/H+9VX9LV4Q
xuX+Mmf+TCwf0rEYnjlEP8IrmJgyyPsY0zUdVQ/KVOGKbOaXbpoJOdt7Pxfv8/8f
0mxnNjkWYBs2UPaMn4ZWuxUL8WkD7D1kmxlN7MmQQm7HY68BK4cWKl9xGBO0og/9
GNep0bj6jl/HR/Ac6ploMfQgq88QYFZLwkqYLpuOCReM8u3jZODe0Uh0RsLJ5CRC
0fXLhXFMtMAbk89ywnwLSTixSi7RMdWtTlWZf3P0KV7JRU6izQHlSb4Te+eN/o9t
9esSuKQhcc0mp3Li7bMv5deEjhfyY7V77NNOnhB95NAqznfPi0LoucOKrYCQJqP9
Klu7XA2ZPww41KyiG42dTI61WhkaWMkYdKXGP74Yb/4Bn2uavqj8+0zrqcgkqzJ5
dBtDia+oJB0PpuES2lK5rBX0nYU0u2rjTgk3DwoHDoIXJCFnFws6Ne2TeggU4X3S
jnh7WPI1XcCLADBlE6gher2Xnfds44jIbsnK2m4je/JQNC37TgRItgT1VWbzXVb1
nse4g7n3HlLv42BS1mDF+sBlX8tvvdWcID8sGFcPjPGG+GbS+4qn9xRDTtfBeqKP
MmyOS9dt9XiMJA3Yl075Wi1+uRSrNpX7mf1On/gWsrKpC0z42JF+zobXd+CP1KaY
0vU+zR+W6wDm2nVY2qZTWNjEPffhGmAHOogeGa9GquVzj/JV0Th+mXuXnBmNEYXh
a6U2/XqCwuLq+chnmbg9pZUERpQh6mwMg6M3apn0pYDu0bBSG7BGltvpZeGMqMOs
LODBH2K7MgIOUHjJYPJgr6l13bpagu+XcdIn1tECS+nuCrjprfTkR5Ecoft35w53
5DGTaKvG6kHrjIbp7Z8OqFvjSwMjm/FM5YLMlsx+WVaRJY5GynPgy/xaQaftP2My
d+PHNhsQo7vn0Mo2NTfB73Ii4iItLsnTqeEsL2bNRfKtWRbrYTfFy1rBFPVWUs2S
cyNLGJaZBOdZZe1jh2tpQ8ZUIeMwlgdur90cwTmr5MqteMMQr8UAA5Rm/WzMDH6f
+awjnr9pijW43UZPPb37BS5Rnt0HWpyyEXtT+VKSSzYajGCIr+IEmqFDVt9w/GQ6
lLt7J6ZSQy09nHHbpZmgagtvffRtAcLBA2LSbWtqj2xy8MUU3eWoP2UCRfhx1t6U
J/l7Oci0Zg8gA2Rh8O+DFudRlzEfyIzcaVFsnSFQ6mR4xPmepTb8KuiHAMru8NYd
cCRPNU1fZWu53WhVgk1dDHyf2NL0sm8GIjc7qmhF0+ZqZ5jW6JQjYz/U01uvtwxt
FQOu+iz51TWrLJ5A7nmI3zBy3RmaKL6B96CMt96OK6fh7/4rpXEDw4W7gHFCEDik
cMJrpi4Qqk70XLZTnxu5poIjNuqfbgwo3xoJ7cPL4O3Hp3wHXXHdiw2UMHBOsnZn
DXRUUuyw5MUiduOagKT0vaVszbTFjCiOLHQq2Rxudp7wXXKDgPpjKZJ/myqLrcPY
Q1MOwPwQx3K2h/saNZz5lJja7KYj257x+Og47/Xbgr85kCouZ4PdSbtYhJjrP043
FuSvB616cCIMhvSEdSs3K8XTLvQgGS/w/b5xiXvC5Qa3T2idm0GyamHbBUdX8qX/
WB1/5tu3YX3GQ5Hp95RCNJbUiRbWZCRLcniq3Y9QT4/gtAt+jdunAalpGsOLJ4pK
CqHqa7W/LRRBlkO687IlHJAx4LPR6a/RnL11O10Mo79OP7yEA1WsCbh72K87vLmc
DDURvz16TYIJtw9uu38i/Hk5lfezox8AQBCy5L4n7jcllhnp+Z12aazH3l89DkrU
vNOSbzzVkJ5Zo885FE7+blcDZ8hbPTc4MPz3ZSb041bMNbi0QiohCxz8d81rrUrg
1CC3rIvVmLOxzXPk+HqASb5Lb85ljV04iEifA7BsyRHU4OzjHlpB8SKQQ2OpRwOf
1NcMH5icua4wSysvhuwj8z1sU0XlgY6wGMUqjrQG4rex6evC/bAQaryEQ/AMlXgI
a+jteB7vYrvWGmyaUOk8dBteKZla4Y48iJjNFXa5YWcT4UDmDub2R9+0y2yyLcaO
iEKel6sJw2x+rFwLtyTZXDhHlztFK9/p8Xw2djkvkB/0YzVULFHIAE08G5wsK43T
ThELfy2bOhy53zthQCwGy8/ICK87dn/gXIMIizr66uIryqS+h97tTv+zcB/dsFfu
WzS+cNmD5CQC0UO9GU/7TWsMc1trnABkZCtXggyPGe19vIl5TLttDYN8IQPhMJXv
px32PFiHGziSKt4cSI4hTlozs6s43SUi/iypuyjQIIHU1oVsofBCBsk+PCNdnCHI
lmq3B58UF+4pmVDi4fK6afSDH4dHmBPqOOJuVG+gQNKX37ZknfeJeoKbsRXp4K98
ITgYWYm88QnTSL2nAFWMeOT/c4Ju4xpV4FbTNVjFycjeLFC2B3OEDU36dOd2u3vn
lHTxkx1imi4+SnEHnh+OZrPiSZcXeRNnDBUR91nV58/DCpGOtHqdOgdkK2ITWOG3
COUiHyyyoUclNJbLEtafm82BrviwOTQz6WNj/slMEjT/uqYeWTfIqmvJjZJawLJ1
+3IJK7QXjASPNWf36NwH1PJmbVw8EqOydKwqA6mu7b8qKz5vCzK2EzQ1kjEohG9P
8WT+0wXoowP3NQCaEhcJZ08fRqWa9PSbjZTQfRV2mo/9tdyJlN5sRhaI7xi3SAtN
Iwn/qdCoORIf7+ZpC/nQz+jN12UjEsly/Y2/4McM3I0jcw/kX+sG3B4YiT7GNdlX
aEVHxmxtQRW1wQvNEVmz/mkF1u89jmAtIov7ML3NXPAPoKsbSw33r/FiYfyiKwD7
/MZmzkKNk5EHBIObWDKot+OtBds+eyBgiSLlsdMcXy0ycZvChjo2kWjCAOKs+xAw
sDmvlh5D3f8SpsOvPf8LfRySsOJCipd79OHf33fmEQCi2q7BjBNJ8zsRUGEyg2Zo
XyPbY5owKzhn30VQasXBr8towYj0ZU1Ew8xTc8XSQJ2XA2eUBgijB36d+K6jhY1N
4GS8XI20SoDAtrgEiA1PSaDuw+yRisHvAUz3tpxM7kE8pe2+kikuuZGyGb3hko1r
y5TdD0IN9sdFe3/DtZIywOxPbKgwB12xWhFdHdUXpjR2yiWKDZ9THqg5yDPc+pmf
pxk2xj6f+bYs+eaRntgiL9nPBKp17cOc867iLXcYi+znegxEs1s0tQC925Z5DMX/
EtRSflvGkPz+QQrq+B0496LCP3LtpdCv/nnare/Suf/vLDfMN1An4b4y7wp41znW
fqeFOGmsYXEC+IdkNKvZp/UUuU6TsHgXllkzfmAZ+QA3tprC+cFzA95ovP6AZ03z
WFvMmJ2pnc0FlrVQ1XRXZ8Q/5sewDgStMu7FqnNiNN8fyU6S7znAfLHaKdNPi//9
bRTAjS2sjhBGjm1zimz6KPdN7vHokFMr9XcKLtDhJ/f3zd7JEDeja8h3Pkh3S349
aIR4jscAvO0NoJYhZ+PLA2cREkq189vV+jZ/Jz+nEKCmjBp9w3q74cIjp32JD3oQ
yIHzbWf96ocpvTVb3FfBPXBaVaSjA1ZwXzXASZ6VHS/YWMRLqOSNjU068V9R5kB0
3YhC3f5NeRFptO3XaK7rKaIkYSqT8r0sWwT9TQjidUy3H9MLJbV0WslQFIgK4Vkg
OGtZJxd41SSdrKkY1tkxVjGl6PfmCdJ9f4/89xOYMHddVL5sn4c2klpORuwPKlAH
RGxHEKSCkQY+jiVHcJrb3EjBXMD37z+1Yzv5nFTdIlMpluX0Mf5UKlf3wn3/aDPj
DB86dK4NjM9Uiz3+1kVIBEA0h8t7mnGNRp2YpRIv4MEk0hU7NJR25OB5CF4Jrn86
nZs8hb6Pbve+ogUJ01W4fj6390jKTvBKBivQLMmgq6YVPtXBITqlcs0KmlCdQUBW
`pragma protect end_protected
