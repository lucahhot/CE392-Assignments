��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_)!{�J���Bh#��\/-�N�}�5f%25:Q��Ȳ����T%I;�x�f���zZjC�њ贠����<G��'N����!���ɫG��K����*Dv�"���ü����P2���-�3,^�ٷ�:�cuݞ��.	�:2f���e)��O���/������e�Gt1���V�a*����!y�D\/J�!$��et���Dn�̈3��5;c��
�[>�����ؕ9�~�Gf���V�����S�ڃ�V,!*'���w��#\U�S��6�6�{|�eܦ|�~�y`ʡl�_4��9���?K�ڠI�~�|~���\���7�U��9=ś,H�/�AW'v�����>�nJSU�n��mN#�K_u������^���:Kq�[V�Ղm�x�������Lɝ���iC��r�V������BP_�cө\揤���k��Ԅ��!�mɞ�_���T�.7�/#��������g�G$�L�mB�`��Q��>��@?�'N`�g��7\�$0���A��jđQ��I0?�����09��Q�V\�Ql�����'4xc�t�$��V�6�'5"\)�o�;��7gҦ�	���DL1��ȇXz��܅�G�+5��Z��#D��6���D��P"��]���p��4R}�%��+��Exa?��ݛ3�e�V�pi��{R��̈���Ͼ���w��f�I{57*����kZ�W��c�n�x�L����R���yh�J��C�f?�B�Qf��g�#ؿc�>�A�j�*�K���Xa�&D��-�Koh���>ll��]�[添6��'da��@������wsR#(�KP����9<q��qmmKE�;��f�� �6�Ն?hlp<��ջ�}46�v�l�����$5�/�fc.���>���<��"�+�z���N��|B�|ː��fP*���"��G��<�6{ZK����������e!�.i�5�;�I������	,�o����[KZJ�;�m����/����.6��I5�		�X�퓘dOE�gG���A�����8q���`��e��6Q�$4ɤ�[�h%��3�}��\��e�%�tJ����m`~��s}���@5|�H�tM����w��I�����E_t}PJ��6#�I	ynG�3��o���*n���j1JBx�({��A�M�r���l��������!�ێ���F�yD���*i�x��y������ �J!,q�y����=E�Q�w��md��i_���dh��7|�eW��S��l�pc7��)����us���첐�x�����>�s��=�7�`|�����?�/7������_���0	�X���p���u��z�>F��k4ﭯ��G��"�y%Y����1�d�3��N��+�*�f׶ay"��<;�R������Jd��Z�(��k$��ʉ}�υV4�
�1v�p6؎�(��t� \Y(V^)��*����������Y�o�v�����)O�U	�\¯!T��'�5�p��u�Ty[S�7zm��o�Z��^�g���$���>Ք�Wy�eTu�Y�foz+�"�f���G�*lr�� e8w��6���㮞�5F}���<��N��[�q�O乍l�#*�e�4u;��Ã:�P� +7��®�~4�*2���p�B-qHL���]�����^DXd�Wr�e��ť�����}�98��Y�c>@����3�0�o5�?3����럯x�P�7��<N�ZB�����¸�PAlEJ��Rk::�p�e]=J|ܞ_T��%�=9�~ �4Eg�ڇ ���/�_�����K.��HE�~��K�講o(�vg�ڷ�V�.�������O�'wL4�S**���.�)����d=k�}? �:'�P#8��(Q.���I�������Eၹ&?���f��xՑi�Ψv����36:��Q�}GP�����UB�6p�N`�R��gx�V�C�e�;�6�}�n��O���ʹw q���_�Eԥi1oK4�1�Dpy�bX�vYCUv���JO�P5����`^^�d��8�U6&9� �Uه��'p������\�/O$�mZ�$S�ML��%@�ow�Y��s0v8A�p�v��r	������1�.���ۼY��,I6m3�^w��J��=����{�L��9�s�S�pG}�c��ʆ2��2�}�B疂�S��@������;��hy2�{ k�`g64y�p���bv���{�]M �`1���T@���6\�ή�{fd'1}�f��Y�F����6��|��:�}��}&�Y�i5�U�5,K�IwL=�b!�ƳL�[�^�X=�*���^<U���䖬����R_����*�B�%��mOIF7�X�@J�ґ�*FF��\��½m�U��i}��o��aA�m�����ɇ�3�Ө�?P��0|TP�*�p����2�i��{�b�#L
ʊ�K��U��nq�z%qF��|/J1t����+��*4��R�$G�.���Ɏ`�nt��3  �r
����`��_c�4	�s�ha^�y N1�x@!f�B��.�
�,����� �U�ވׄ��N�y(7˞�mꂻ�����!�j�W���ȁE`���7��'��@T�φ�/�φ�	��fs$�b�b�铝vv�?��.�KE�>��(k������?�:۩���N���a7�f]���3��Е�ӓ��|qX�@�fKb�E0��XL���:�ПhI�*k*�Y&j.�|ꦜ�z���R|o#SZsF���B��7���O!�a���)e���k��В-s�]\�}����QR������DL���;E��3�!KR�~ϣ�r�ss�WB6�mQ�ZL��� ��\�h=��K�W�i�D)�Y��en����:�/�)�N�sƿꅢ����V�4�Ѯ�X:u�/ۨkj������Fp>��ޚH6�mZ���0Ϛ@+f�F����uHCU]��b���I�2 �����XC�T��t[���RP���Ѥ����o���#��؅�$���m������oN�V	[�ǈ��	�>��Wݫ<�E>�Y(�?����4��љx)�H��*�>�>
���m0ܡ�3�G��ߣ��#��\���'����A�����ǋ��ȨI�^	��t��5&ɑ�1�R�i��F1�]Ֆ�� 5�2�8����+j	�s"h���t�a|���eҫ@2�ġR����v��F�zWg{现b�ϼ�)*@@6z=�-�a<lR�ԇ�+ix$|A�X)�$x�|O�HRVa	Q'�$m�GѪK��g��A��r��Ql�������r�P  �V��3��Ket� ��i���FXX���5v�NQ��O��������:Kr�X��lk�Ќ1�%���ϙ�:���e� �<�?�%���;��e�x�TR�<����E�%�r���?����@�Z�i<��l��Y��'�C��8�0R�M�K,���٪�H���Q�uJi;��l�%�s1��L'�:�����x�^��k�O$�ߣ��G�ӊ
7C�j4%�N�+����EFZG�š��zwK���P;}"�$��8��)$�����#C��7��½�X	?x����tB����B^_������TȰ�mӡĜ�0�]���4-�s�~�	����e6�e��W��X�K�'�E�Oº�f��m���>WH�<S?	e\ai�Z���E�XW�{
R ������s��"2��d�}�MUٔ�q@�@\�a�uj��Y��k���T���ܮU)�}� >��;4�os�SE�oq�vU.̰Fn��A<�q���@>Q{�$���J-0il�]�٪�U]J�+Ӊ�|�ys<���5��U?+S	S7>�]�fy�@��EW�TZA��a�S�k�EZ�}���:��^�%̉��܁#�x�c�:�j� �Om���Ʈ��פ��!�p�
_�E+=���L�w�$�lh�pp,w���:�5�7�kOF3��U�h�9=}����q��l��~^_�I�5΀{Ҕశ���Z���l`��8�������vA�v�FZB�b�ƙ��GWsScj�r�O9/�{����,�~ԧ��/+�S%�pZ��Z�G�Ԟ�)�  p��`�x������jH)���h�Y���th�r9ٻ�4L���a��)�o�T@���;L�z�p�g�߆ZdrI��	�FKOB�ϡ���q"{:1�s��mr]�,�Y~���ؙN�z��=�s��qqI����d{����f�mM�̏i�e&;�$C�?M�0��W��m���eP>f��t����(�0$T+; �KJ.cL���pxFXs�w�{m����$6��0���X�똽�o�oA�I��=��R��b�����F�����4��c�P����\�R��;�
{����ǅ,<t�>����c�ɶ�>��ԗ��9ˆ\~$R��.a��0��Ļ�7q�k$���c��oZ#d���.G����]�w��n�'�L8���9�TA�-�սm�Tv�Ud,S��	w�C��������o�8�����eo�$�WPnԀA�^(�[�;�����^.�h������FFu��#u�|�S.r�wDU��'�c\N�׳rP�$=G�\�M�=+��ěB+���c��8�����ʆ����Ն�R$ p���ߘ?{.L��t��o,�[SA�֝{.��5��gdn�}���3>���"�X��X�&��\�S����]o3fю��%k�����"��������wFU���
����J]X�D�1
�Ƭ�꫆&W!�`.UŤpX���GI#�8*�O�]�E��v.B�W�S.�V���N�&N�C�~\��L���U�:����xl�x�VN;Po���˂���D���'ʖk��8��LYϼ��R?'��Fe�������6�� V��ǩ6~�Qc�����u2�6�彯�U�v��H�Pb��J���4�駃���yk@��l��������LO�WV�M�mF��������*���
-U�̸d��4�m2��.d��h������G������d�@��C�
nO�)v݃�)t�@er�:{A��!��y䖶f#�?I�_}����F��.5~Y�<������HС(�2ն��q�GW%>�wZ�νED��"��ӄ^�/wx)�����M�N��-�}������`�Y�bAO�	h�#4��?n4�%���3FM�x�#T���]���4��!	{��g�rs��ڥTv}��W%4�c��<9n����|ڰ7qQ��3�*��|�������=�@���{�k0x[��������1m��i�����m���:׭^�e��i��Cu���4�v�!'a�ɉӛ�)7�G�����+��`� 	��%�k�[6�������e愯16�D5�i�%����6����*oo��ba���N�+ǖj����z�`HT
��?W{F#���Ji^���^El��h��1�.����b��`v}Z:O��ُ�C�m��	ʩ

�7�4�
����1�����nG���?�O}r�����
�Ϫ���1/�VGi���=��3���
�jQ�4`$X����>PLHe9�^��xם�����`v-]�{����T8@��a�]���h���U�Po"�Ӆ6�P(��s���|������1f���:B�3������\fW�{ANR���tR�+��Z���c��6�G�AN��F>Dw���fu���ߒC�kUw��jx3�����M/�@���|cS�l���۔©�B�hD����!B��
KU�DyP��}Tζ'�������sw��ec(j�Y0�pUNh�q�L5�Eb!�+S��uG��� 1��O��/�\�n�׍�4MI�a�Qʇe'!a*}�,[rS�Pk���fhE��ks}'e"�:�P,� ��i���T`K��M
�3�mw*2�. ��ӣm�I	��$�����9�h�������@��h��!u��,3�+�%I��DR���[���y����?�2�Kz.����s�݂ 9H��eP+���_��Sk�$�g0�N�� �Ӎ=��y��Xb���!w�2���)1��#�JfB���$ ����gB�՗�6�&�n��YxU� }F9���a~� �������d����Pт���o�-ܯ��'�*�]=�dv���Dx)�ź(�pf#���F���	h�S��p�TF��
2��;��2�f5�b�yW�_#3K�u$�4�枅 �$�&=L"�qk�E߃L>ms����3��c�Z�%6}���D��Cݭ�t��UU�;�P��K�,�@��_~5�򃫾_����P�e���5�����wc���AQl9�< ����k�W^���j��"����C��9�!2i�NLy<?�9���(j�?���ZK1�5�^���y���ȇ_�3��6"̌��4�c�G�sdAQ8��M4��B�t�W�"�v�(gw)��C�4c%�PZ�w��C�0/9��@<��p�S�w_�v�n�����]c]���&+7�<��T����ؕP�(��H�RG��M=��˵��~�ڪ��[B�=���,�+��ϼL� �
�%��%ɐ'O��lm/�&ݍ���N�"X�%���.���;����V@xR0�Q::�-���~����:��B=�ꎘ�s���L#�Kdt�G\)	�妰���l�{�R����e�m�ݝM��Rׂ�Į-O�@o��P�Z�Xv�L�@&�%~���`�C��pˡ�룞���H�
{|);�	�KD�Ú��֛S�H�@d������LK�/�Aɻ��v��C�P&�[�>;��Fl��ǜм��K5zz��{M
J�?4���>4��l��l��)|f�tga��{w[#�[]���zZ��.c���RW6�Д����=�+�~��W�U��D鬆�;��������I꓍�c�g����Q�b69,p:��ա���A��<G�I{��L��SSB�3$^�/W�:�fy��!��!an��o.����q���8sny9���
5�K�'�_̲Nd�;\��K�\�Z���X�P��k@�D�lZ$Zw$��0C��0���F�t?�8�u����Y5���!��aL��a]�-�l�W��2�m3lS��o����=��+�O���G�.ߡ���?i4���8�B@��\`>��PJ���=�nG<d ����s�,��(/�� B�C�>��K%�s+�#�L�?fN}/���;��=��{��G�;4/N=���[�QmՕ���2�"�u�MZB����OaH\