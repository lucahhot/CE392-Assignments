// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
C4sIcZRv8uzFhQFvltycdNrZdRhSNRURb9F5u64IhKnEs409aMWeXN4YRPYnlIQp
IYD94DhjVhBvm0l7tDZljXMFwjcYhjBOu8GLnzxiP+ctR9k/GOs5yF5eBYVWCmGO
N7paKwJHn0Lp0QfjlUT876qlfBJAWfvzwYS0u/Fj3uk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 12992 )
`pragma protect data_block
4Uz/QqMnhl2aQ8PdlCGZziELiipqzL40Z2WSvQXKXnoJl3plMpv7lQREAmCr3xRk
j4MhhcB1+AQeEjEKw2WHTDxRYWTAMv9xkXUHDHQJVmD0mua7YPSMUYXy2bWBCrAN
GkGB0gljtkSuUlXb2kVexeLONh4NPfcBiryLL91wsCrKbD/kbm/ssAvRxGXJJQC+
LMf1Im6Dr9zyj32MWuVilrkFaCZFM/XE5dLkIOF634qYwDZd5o82ujchFHGjs+rf
hOokJA559dqCikTLRrIzIQ6KR/coPvtdI0FNa5pU6qbB0ikDq7qto+5xrbHM/3s8
WW5nzylzuWTykVggZIcpEhKOkmhFQQkKsA4+986lyAFsT4emCdb6r3FjkB/IyzFv
6lmQgTW4rlw0tMV+qHSDoxjcp7l2NwxNNQBLYC/zFf6l3UWro4Hy2nyQxl+IaVq4
hTN/9+YnBgTSNjgoPwn8E5exYhPk8w0Xi4NOD2Ad9EmNpQ0AvXPup8mIIYnq2F8z
tLhtxl7LgFHrk0p7/pIg/TnAhJHQNNCFsTL/nZqnDtuw9XV9HWUKoU3gZS1BRyG1
M1DC53CtlozZLLAlY3QzaU3BXTTXBHcpLe8f3MrS95ro5FeZ2p6AFcf9qbQP+48i
skOT+AtY/Hob76RW292k231gqAvM/r9wrCksYnnGI4FgRfvxb3quQa5KhwXJl5/M
YB7DEQWNvcu+koyBKZf4FqRQ6iWVVHRYpapI69rhPA2dN3tUbCf9TiQ2SJJOLzRx
Bm8mL8r/UIT0I5En58w/yAh5Jgz7aRpIfZN4hmgH8eVkj6iAoVy7c7DNJp3p18fN
9SW9HvgVokPETIwTZ2b5elty1KFGYIvjWtmjG7+SU6tNnmEHyM96lUfyTMiYAhyH
ORQbML/diBYhDlHM/HbiadBLkIQTKRrcEm0ALpwFtU1B/mKyK0RMTvGd0Q4fWEzd
FVCuLcdM09AngQtWak8G5qKdo9uIcRcZzeEUr9w1cIuLd261S750h4gBdwWNjXgG
JyTUpmhfUsyxVXwl87svKH/Bw3oojSlTD+8bKSZnFcP8J/4qba0nn7DCBG6OGXT+
K8PX23K2uLx9t3l22WqDHlhzcfZg/VVVfeTjMcu4l6hXDJ8nMRQ/21s4hA7OlLGD
Bpqc0xOeOONi9GQpbUC2eQuN0LanTtNZc/jL/O1CLOJq1ZQfDvDXRHvW4W39HV43
RSc6Bpss5cpCXb4HRXB53ZWcZaC0iaycBJunndkcKLDLiqSYxit/jkdV79vilNjX
AjixLDueV1Cjz6RxY76KnYHaeaulxflqImkz4Ltuwh6q1+dz9bwVGGYpunVzwB8q
vvqJfs93lhhnbVBI48P6JqT5h8ZwG18XHGyhuiO0QznDIQQecxViU5vQDs55DYoY
3liNI0OJK0wTfSmjVcT4qDC5eWZK+nlAdThPVy0+xdTuov5pO0M24Fu6iUsEBUFf
5GhKBwRIaNka2FPXJBOoFpyBM+gGGMQnRHbCKgQVUPhJTZNvkEQ/Zb2Wi4DjzQlw
NM3KWBXw76sDYwpx3UEVEykJNwxRtExiDrXLwwNFtqcyazljz1PCnJPe9zvZ/1Yh
F9LjMJkkpvFEzmI0Jf2xpvUsk96sNgVnBvXFdj4CR3fI55OqcH/MI4w3rdiY/w55
Qnj3VKvf7jt8gobvxFdkn+tzr4HtwaKkLFu/OnJ/+F3D4na2AzTZef5GSovA174s
F+xlKBPXnOCXoFVJZSnCWKObQQ2pi9t7gyPsVqGWwTulYYYmcC5HOdb1c5a7ZCoc
0evySaXMQAh+a3tZ2aZuXfQJacH9iFy8AtaM40FjAwPpiMxJ99Q4ixK4thoLdiKs
XHHHjpFGMrpOeAz11zeWsO7rekfVNzsJEPbcfevMc3rNnJYONlZuv46QqUHyAIN7
/XxUlOQCLkbnL90e+4PQhDlzp+gwfG209b5M1M12MmYWjiQssDSfvsqBofFG1bt1
ryMNcNFpr79XmbauNWqLyGOjCS4XHh6s1WSaNvJT0GVRNhyJkfwkc3OTAttPTqhU
yBrhWWRw2tdzaMCdWWWOyMOjgVQ+FferDjvOfKF4DXUzOzQzVMy31/T9biNL9wjY
jHZurlHxxIaUcuTai97ID1vf7VSOGyX/DlK4Dq+FQcooiZtxeRSOmI3WdYUvB4d3
FvzPHYEN6fgcfBWAW8tRe78rhcyIGmPoW3lMZYHXulDRQQ/G/hdhOVqRHAksjAl9
hBHkeYwxUQo/5jvbDtL5AeYrUZEpTRHSnGRu+wmvQWPj73KuRilqTPe9W6XlX7I5
QtSWxLKYmfKlQhDxl0kFMOq4dI3ERw3gb4OioEOiUDrfxzWTq+lP6A/pOznYCiCl
rrDgPjCbpJ1AhyRo6jvHod7BRZdB6BWK1RuD7Xz+qEjFngAgeKH1NoHSkg/xeVmZ
q9ykTJQz8pTcjKtUl2+muO7eDZZVEGrvg0l2M7xLg0InDMV7mPBF30t8A190n0Rv
wpGiIh13MVh7MMvY4LDTIQ51odgqnHF0xmSfHPjlCamMgZhwUpMPs//8pjdXpwZT
5SNyf2FwWtRc141cz5cb7BuHEF/p8N0Csr0o1AmRpkbV/+XqCW9zFVlahKcmh5wE
2PERsROxQHjfNzSDVXkXQfBFcs4KvuHOgM9s5qY+Fl8QKh9+s4M7Q4Rz1ArYZPrg
0Vh1fGvaTGIhHtWJTLI/NMGwJ81d2YyNzINv6BTp3Cvh0q0N3yAsBurMwQ5T7GEq
LDvczhFshl1+MDCfIQBHb6snTHgyc4rrdwtnJu6lk+PekxPfeDy69qXtzKj5kM24
AqUGvzUMybYXoU52G+kugKjK+LwtW54XCE8BdPf0qcLAqzsIRnQJK8SOYr0GMLrm
YbnjTmw8n4F3hqXBhgYe+bT27MHqKpdY4MNbGLvizl6yq19L87DbTZESxgfLCG9e
1QtaRjruf9lbpYnitCKM+xu+37sw0zGq7bre4aiPudTd+zPAanszFzo0c2SdLSFq
oUIGmZbnW+jxZSIdJKv+HOWPlzUdZ5C9BpTGRTNduIYjLeSefYsc+mgr7/lUlIxJ
hf5PPZ/17M4tznJvfOH4K5eS1fgG3n9XBvxziIepS0xdxE7IE9ifSWnUNf8H92oX
MiXThyuNAb//0rCxc1Id5rOKBehQ9I3Gs2co6K2MvwMhx6GIp2LbGK3F4N1oCjUp
OywPfCzbsMK9CHaxJbFueNCHDNQW8SrTVLnXaS2luIhwsBUDHUg90dk3aQkTeyD+
J297qloKn3RZAqufrcNYV3YgDhbq0rvHSiWXEzNlE+pGH3j6qiNqNZzlS4H7Msom
LFRud+KIeeY1/meDPuKRfok+LVEuZpblTQIlWVKLyYRWxlu0q/d5Z+RqZtGVMlnN
DEHf2QfQDXLXRVRCquurFOzezihk+2TEHKeOicyTA8/aAOPMYmQhOfeBqB86wP4W
4qwXAQPNlmMZClfiFnmuriXOalT1YVaDbHaKMFj6jqgLOqcREi/S8c5VarqxLbCH
HVgasWIytJwa6jtppO/cE0bryAp8Cr3gG6f6XVUk0cVH1E6hZvRN+/58eLPzS6TV
TzUeUynp0lHC5V5VKwpblgbGINGGCc2yqIVGvAvLyYEHLTBc2LZyxunXXIZJINUR
8nUjloMNoTyMUJAwrI6Pcc7TD61+KUkSDLGYRcKVb/GSepfQAMNdXTBhpycG3lsq
oteM/O1Ur6UZrXKA07CSjvKLu5m7AvN3B8vwipI8OOhN8hGqzBkBgdh5GfVM/evL
4BIqH+ZK3TDIct1CvLG632pp/b6hTjyyNrGc3bnQ+z1/Gup67i6xEcmB+9NSbQKo
rW10qaim3IFWhaWo+FD03MgBUtJJIYRqsS9m759aSiqSGY9ax/MhgjZvLNvfiQ3P
7FMXqWGC7kbsY1CyUa8oEvv7HbBg7zOWbB2iPBc884MH9DHsS9ev7DZdnq4LST6K
LcdXnNRQ3HYzsAuszQMg9F8Q2aQf+Mc0W6NHuBEXXN98hxuMcD7O2sad7jFfI7Ld
y45LInKuJ+uSscMWELmlnSKajxm1tFfhEcV6UadvXEV/QJHzYt9dDQtrloYnL4m1
93w09j3NRtFx6/8A7wvm07FbWFP6zBGpn88hIohLIhFBH8TtTlwlKQmuUF7HUeyj
xJO8ObheHWsMywdw998PWOgZKYO/mUOeHpFM2hAZALSnW5IK6ZE0QVNY7OlqY26h
yhuYsaMKBV4iABAA91jUYgLjslH+hSLrhCSsCVF7VfUunjyY/fvudcx1Wckc9/ux
Ea9Y5qBpAAkrwPYsa3xbeCXcVBLIaeovfKlUNF4y6pfZlorb/g7oFt+CD0+KKxzB
mlfRm56W93Wpy/kyX3AAw02M39jiUoUb4NGV/kXV8NbmAmG+tVDlh1j+97rlhwpG
GTh3IjK/jJ9eXprU94HVQCUHYwkRx5dVgs14zALcwvTMnF+9Hv32yy0vyzXae2ub
fxo9Dv1nlg7O4NWB/lQwwuRQcIMxryvADzKzBpCJDrMSGDo9ltyF/fE3wv2wWwJV
YMPlIaENahGAS6KCuUBEah/dxEOD6I+d4fLnaS7Ozr0x1JTjHeVthZ+lWL4D07ZV
BNX6GFQVNiPX5e7G2Wymsq1DETNAwHfqdz9yG1pbK1DDnsYyAlF/ZizEOM2S5v80
rSZWGQsjjB8AI56lnOyR1KIEPVbumzS4uv6Ns9kb0nFssbpyt3+aSXBpY0LgzqWa
oZDBfG1vpgCdsmdRZg/YH8Px9g7J7BWpYBnEPH8cvR5nBoITGp/F7K625+hcaZaI
sES8o8+sh800Qt734uWsr2qhB2pBNkaqyIMP26tuHlg9V9xyVWsqIYANh6/4t8iz
NzsgLjET6CKcjjOaPWwHyX4Gd1EfwoMjln7QPY8zxPax+ZHqkhgo7U5om1IBygCo
9e2kpo5EMFuqEXHgvBFFmYRTUuxHVo/PpBkRfjegtSEBybBapwEx08G+2II/zG0V
MXacJCu3jZXHW1WOvUheG3X8xNNY92tjVzEcyxxsPDKx5W1Em0vYCQBy2+LrdcII
ajNHd2kBr7DqOSjIMRxfU75E1ur2RXZCxcR5iG5pEjcI02/PBLVXxQ8XZa2hAEBz
xUVEOcnZ44WgJRAGOc99+5/c8uFXt6mGMpuqUCW0yC+d67tYJj5SqdQ52R7Umuvz
aQmEcZi7LmErJe0txqZ+NzhEbE5KeNDodDCGCL/gnPUUdEjBErLZjFQdgubj89Dz
5OQO9bau1CvQ9IPRBtf2ktc0R5B71f8Tq4xYXUn3XzUaBP6daXbmSMVu/3DcNOeP
Q6Dv2PUr9F5x5Co5mFISry2u5MGPuImbuHNvWpPDFC19/vWFlEWieEx1QUquZIEu
Vxtj1NEIa2UsEjy3tE2aZuxp+/DtFlRMoYOudCzNi0laEIIUKxtc5bgQgs32Qn7F
TjhAaMQfS9bKdIt1KdM2+MCYqX9skCc2gYwUsh2ifarq83j2843R3AeD9AYQ/3S2
TCts3OH+YFSxyqPZ2OeGn0iZs7v8/baFWG9difd0+AnUkqTPY7/S8X5ZdG8RqOcy
CqX0/bEyFtuwOLzlz32wiECXD285y4KgsOysiTfTw4UiWWqIj/WT6q9fZNKFQ0K3
TxchDZ+UaZOCg21DY6SgXypt/cmV2+UBbqenC5uHFMr84wOJHtEgVSsjOybnm0Nu
mycOvptR3YIcvTLc3i12ygsi9TXnPmHb7Ah9WXLBXx5s9hNnx6vOECnCeZ/9RlQb
+Reyi1hZW/yLQDLpLXEfwZeAFxaWxLUfnNQN7b6pO84iLfWbWe4E0f5tdYn0Z4oS
QIsISpxYbbZmz4r9PweOS3t3AChRjydybGmkJ4SwZvoawtoIsTwN7ETZrOiLF87j
RQ9ltb7PNzDJio4ZT3H2R/7AezPA/xyy3givfjHs02gQ91AuSQ5f2SxWMI7ODK5I
j+rwwd4YOGfsmevzdBOyywvNowvnH4TwtNUZQpKeZURWYygJEs+qNVYaZawO+EDt
+LUJXbPTg2X/q5kr6d9ATLYI6VRk9JTrC0wRAw10TCItcgXaOeo/i+Z6vx352Exa
TlE6WMU6yX2GjCdFuunxOquo+++zjZ9llCUaFsRexzudXpJnTh99v/cbEccIPIO+
eI5qCFGTE7D8kw0+naBRu9y/cpwRwFawosiPfehXohcY2X16TRFDQutD5/ml4FzJ
whYOfXL34J4JLSTziOXNb7PBmBM3sYYsCvZczZ7Pb47fsXA40+MOan6nir0jLm+G
qXzdKRpbC50gw6ZjMdHNmBQ02aR42EYoUOiqU0rqvv8C83QKXR+sxnhmeHLoboZy
amg6zCsAfqk8cR+VXOlw8yVo2ePyC6K5p2wJ0oLdOFNhnrTjPxepn5gJa1f7ltvL
WeztDFBaRkdzLjvjfLuDz1f1VKiF5JxTtah6tUVzUbQ9vLq0UZBIfJtcha3cHeT3
GM91PhvyjDMJQ70nKhoxGCx0MnvIWdC4Y+jeImeSp4OkVzavceGGVcG+SiZ2gWmB
MK/7QshTTaZYmE9F4xbTELrMYoW4MfbMJuUTQg6QWXL8Lv0NjwswQSbAHZ6AwRJH
wNY07WcX5D592qMT/VsAUx++gBlNtec9/7C8y8s7/hMatLYKWD7nfWxvgfzFmgmF
LqR0EsrcnHgJ5jX+9/S4ZP3qM9bQnLV9qCkrXKhSKcOfjCBbS0Wm9aftmqc095R6
nS+feJpquKSFCDInWme5zqnWTFvqFUNV8OWgRkF+cRHl8wBvj3KEZW7tCeJ+KTum
b2VRI/g/nIKZZvvavGq7KVk/a1qRfZg+HoKHT/Go+gFOn0F5n7hLLipMAY5D0tyD
flgGXTbZ0zHZeKGLwyN5gVpBd1bUnedWHAPADPZG+EM5wN/ovr0ZabawmbNNYP3w
lO8nPB+jf68Ff90Su0ty9IYeSL/iFnHXrfq+G45TvEmno+QojX/LxnAqMNlOLroC
GQfzqLU0qXFXSqNTKQLc8rdbD0tUTczQdTSmAKWSjJGJVY/bZryI2rvZ3Gw16nqn
vhDTKtC3rY0kzBmVh9G3QFLNMBSTUUVYn1Te4IY+mVDj5KXWxTkkpGHFs+7Z5QEz
8MqpDsh1gZOSf7v2VrZGG23q6tGrP5ArZoMSbDJxDZG5Ti4B/DoJiA1aAhHFKCbq
Oda27dTC14oQKZ0f2gtqrkzGuid19ngrwpikU8CAsSifKxdZq7eequjjfMmHZ0o2
B0Wn7iALIJI3+2IA6gMUXfyqGo8Cy0sExCBuUqsQjDI9wJE55NVHsoqyRC4KUy0X
R31CW3KUZ6HuQ6Ye74/dGeE1fDXpw5ueCC8MG9c8o/i4nrEXyeDnGIOEXwazvn0+
27UlRs8IW3I4YyxorJaDvEx6dkowH277Nc6MMtV3iEFzNQ9VcyDTLtzS7xQTzlLR
l4p9w5VkL3yhj6JPCJi6uADKyXzeRFNW4CqhPwJHPyqH2uq5QQdFpGRgMWeHDbcn
s08cYrf1A6Ydrvyj1dvFBbsNkyocfaq7Lui9HhNL+JVmRall602uCTVShtimAOZE
uKZ96A+gNK5qBzTrGGhFKEr6eDKDzyQO42nOZqxRrLK8wOCTxo5/up+4R+fHjRhZ
vYGZ4XbOEQHkGOkaVRftuP9nW63fyziQh3wbQNhUF71OC8fd++oQHSL3agogp7Vi
ezJUm3VH/2LIEY7mBbXXz83FpUvN7uZatLdv0Fxzmpuua1vCEosobc6EFAMXwIie
qvaUOg/Ur22tbGc4ChhpQXs1PwKrVj0v6rC3Ekbyvtn4OQWjWUrzIN7Ff2gZPgx4
JAt2xxJxQ6kwkNLL21czZKNJKXGnb5Cv+p/eJCxa/D/3RCsrjfx40k28pi7SpJjs
vUdK5aGmgQRUeGyynG7LlpMNMtddwDDWKmFK9jl5rhuVpoSsnwNGi+qGGP0l7og8
JxuRH8YAkxJZisTjSZE6RPiwKXPYCrAAHaaWKtRMSYCInmw3jSVDi+EDXw/dhndr
bQQxROaG2GuIU4MAUQ6pvx/+jX6YcPuTj3CwVxYclDQyNsOpNU3tRrFck4dp9JbR
VUuTOP2x0AM2pRIsqkL6RBVAaGNRn/gFTDdE7xOUhef6Jf9lGQdDvayH+0vQvKxQ
SsA2pelVKVqy/al3e1SfkixMqSAnKj2h/JgNEplx5c4djO8VFiVf5CZ1Cua7sTeF
ZFt2/o7E2JBmj6QGPuX7arXluireOr1Xvh9ekQPzvmkC2TqVJcYWJCDzqOUMSbzD
TuXCFZy//J16MCRq2iAyclNyE9q+KRKxp3JJnxLq98GcWscCcI59Xb6+EqCH5sxz
ysjdpmOhCGtQiWyg7PBzN4ETRUzeiBuKTYkn8HpyMfuprpDbiUHgbYgACQd4jB9B
KJMgKSY0DnwMVj/5EOahjX/4jdfR39f2IE88f3ZFdQGaLGnkbJMpbG9o80V0L+bC
Kq5ZlR6Zm+lSw6b0gUQHatnGzEsNOKYPi+Q0GB2lV19nCKrHLJWlOKFGezJfjf/V
OpdqeWjWuEsBgz1rWYOKpLpdfEZhq7WadiTsLM5PilkLjj1QWEhM3klbvYanVUOZ
LwRBEcRzepT0pkgbjMZISZ66Ed/rjTYKZQgxksrxkiApckIw0fhUS8LDY14MRIZD
9m0hIS697XN8E/2DM0rW0I+pyhislJxEQYnHTFvjiDutq4sm3gBFlt5wtHEuKUPA
DdPbi72Lc46MKoPPHI6ZLtUUUkcbcv6zObV72XYGj1F6MFKCbZii/36Q9he5iZex
XDZrX3tKcs04k7gN1X6xywVHK0sQQKhb+DTzHLVzzDEHW9kOeM3dYbas6IsiKH4c
v1DHcPvM9dsktLCMJTBu5OkpaF0PIM3UMvjOpS0rqi9G2vgYQPFnV5+0MdxB+wCB
EksqrZ6JWxplT407AmbKZO02XjEHrw27yfkWe9844N8Ga84GKqggo3iZ9u5fxeUl
tZ4uh2TKqjBDkrpA5m1+dfv0iHcQn56lFGFS0oLmYEO93Lz3CnNvM4Ow/dpnWlqk
4Lm1MwzmIWyevZ8vblnYomuhcD3uqt32oxX3ZzV+Jw1E4aNbQnSdCqHW+twNc2nh
cXcHEPQ/f7mMLqqVF0X5tbhRy9Y2fizBsx9D8dxyS732TmpANJQw1A/giqSY2uyJ
a9vRHiPkmzXRmNKzn07qbUSON8dr907v00RwJ2iLqjDsUZCEJzdFxzEVttET8eBO
HTYPJQNQCFT3UH3SMCpRIumDgNP/KlwZszYVzXVjUQvuw55uHxi+YRcC0YeQwGFK
VY6SP/9UHMYTn+73NyTJhOJimD/BAApKWqo3UaSsR27tDGTfG3wppqYLLxFDkO0u
JlUJekeDEctgF2YhxmyCZq7RwGU/kmbh4PNujUk9J8WiXVPVZ8JybhCMCYyriU32
DyVL38oQC+WuW/znqVN/jHWfSFfnKbtKHWL7+ZKXVlrAxk2AsNWRfQ0Fi27lXsqh
FWSQxRd4tbc6dnGVv6mTcXdrjTAiKV1QrL66AvrbIjLnSnsAJF6hbqo3axLuF/Qa
hq5vB6RxFycVePMCW4tsWUX/6r/btSfzTm8iHT2TxwO/wqa6jOoyEDheVSqjWcg4
LEq2tgVhIc/VthFmic8WGw4LAg1q0u2+ARMLjF0DgAAlxSnZd294vX/2aA4UMEk8
N111NZeol6P2REEhHs3vwe36AZq4vMqh0VzyDY8SfYsoSS2nFIfBXIjZ/5uyUhUU
KOcv5QSJYDrRfrztx2xc8c0AKOEJjzLIv5hKvHtGdJZvcmrTW8gW1Mfc6YZI/BSp
xav6WtgUdRsRFvduSJxqQhfftQZw3Od0Q2pzL5RKu6bfSKwOjKDQjS7Lx0b5PbvE
ESYooBml0zNfQ7QtsYgR0HPQOVjMHSIKZPPAHddir8KhlRagBOfTSzVNZIei9+Bp
DjqdqTd+74JFqRsNvnBdemv+FrGFzaKKhg1IImnIoqxd3VcWe9CQ5fHiEsQwcQTU
EMSGJhCynampY0NA37HDzXmlgYFNtr49mM48/oY3S4bw7ZBooNJxLw6zPRFXUU45
gegContXxtkjjA0A/FWYI6qvGOk4fNmub/3/ShKuxX9fCNMKJpalETOfsoXLfBxK
gnCr0O++tjJvnHYMdPUe4WCjkayNmYhY8KaYBvFoP6L40a23VLCSJKFDqiSYXqok
j6neYBObtrWIF16g5tBH+hdTD0+XIzrCI2rvVbuvzz3BYcgkmuYMGEFpLTiOkdGN
576mfuZF2R89d18MEhsmq0EOfjgTi+ZIsFFOECkPaGp+MrUIMxBI9s9XEfIXZa8A
2uVtcpibvwE5dl16PBmdNwlN0Z2DT6mHI3tv87sTpbcoyhbt1Ot0wilWRChkv1Fm
7Tz9Be9X+PfnMNvzqK8+NDIdQx17GYrh+Doxxjf5ut4x5UzLK3t9osM7q+KCs3r6
n6QN/hghvXko+Hu0qE8QimQHqVDP/JTM7fipQ+Tdbvfo+qHDY0jqc4MyIw67Z576
7oA9Jv9Ko7Jr0YTgHWmB8bGA+QFlE7Sg/6UET4S6ccK/vg4y6dRSR1Sy1KKzLS9u
w8wDEilinaD6MP9uCXuzcFIV7Ald25EsLabhYbnFzaUvzimz5SfiGtnj80OPIMf4
3LpPgucgXy28uapi+4+Hy913tSdn6Mfo7BMCoGo2gi6LtEIDgwDrrCggo/+14dhh
euJ+14Rh3/glzi0fRx9ITx1sOk/YchV4jD68Av9v5qCZPkQKhNYkq1t35AKT72pP
rluTFJKSrO73dK3UX1zoU0FWeq4X5+yWQjrtODge4vzX5Nveyz5eE2KneUzIvS72
/cjiNIv3GgqnIPZbngtGibI8+m93TUKrOigr1pifciIcUYOGNUX4i6JONHFt16dX
dYmomY7ZXu3z8wmtn6Q27oqSkRY9bvpKjVT8Lvpt2Hd2I6bwADtWkIZ+ZeZfeqNn
HTNkm2u0vTHRlK/DPmDf4Nu6xcGcuT+/zAr2aefk2TpNa+xsFX+9HtIvHx6aO8Bs
aIB6vL+GLi61la18Ctov6pzyCQFj1A2yvwD59wPPR5tFehEBgxcLkEN84L+8y1zz
RLhgM/v26Y1S4/d4im23Ymi7Z1qYZ/ZL4riqYllJBVdqqNMEwD+SaOuxfQGGL4Vv
LUdJvplFf8EqEwIMAxb0NVCStxSx643+bCmrwcjtKXL3lr2G5FxMeD/8cNJ/mNOC
LPIVo8iSI6/cNtiRVEe7XXAO1vLQ0ltwXETqXXNtrIqvgdc9RWrmtHR1doievqn4
LqWMcNx38EPCkBlfm4x72aobpYLNedf2b7R1LqgqMC0h/ATwLUa6zkt2BZSGyHZl
OAGRIDBjnSAabq7x5ptYLpmQUuDMIcQa+up6FCeDaoZx2aZMEU/D4iHcgk2BtEJd
kBtWK3qK4G86DKQLqmvq9DmPlT6K0iDycxwDP3FXofLtL9vR8dABTkqmpFTL8qO4
XNcb8Cj3peCa4CIHf+16ZUihrOb05BwFey13iCcSXUUUtOJfGyyuvHHrZs72pDS9
FwZGbSAY5hhvN/w5mdXq8fJRqsscU8CM1NmgRxhnAIP03dgx7q43UZDvORDOyPwI
UHhHXeLbJzj+n65AazHcWrXx7kQUH8RQLtMy0W02GExuNF7wMI/xuiy6risDOkM3
ygqVooEoTNyK+oJUvfYrXedpfKbSVvMzhqz73WaVPniOPj7WyjA7FlQt/mthovqg
3l/TnT9Io1CVsWMnhTuGA1GxZF61wM+4/VHRYaely2cC7+Rg29uyszQb7p3vDY3P
9ELCCnBEXoSfmze2muYJJmvP6JV/h7F5DoSm6Ar/XOvKMZldxmM8pqwobL/j7O6k
c6C7Y67QbmIxc1dgi1Gmri2zRqQWHUrHOj9Xt/dOzgdxmgKZtvXDPGinFyAVt8O8
5uSv+TWGSQSJN2xkk8QIwwoP6ebVUg1VTVP3nD8+/kQ7yesRI3KO4QV5RzCG84f9
JXieElojkaZ0PadJkhqsenKogoQ9hJnbiY6ih2ZsVkA+QR2vOJwRsxTBISvC+s0c
tw/vvtDZFe3UJQex1wf74fxWSCMxVeGX/lyUj5kbsnFvCHnbeaCltU8P5S+hEQNu
TYYxCNCGnQTZSQM+McgL71WIJssJlP6+4Ce4KvLVpsBtzFTYdYE3UFUMmBmncvdn
f73XKCz+p1FX9SjfzifeBhnF900/3/QMa8HA8xoT/5B1pOjcXTgbm7vQTCDQmXI2
CfOorHdBo7G3H3Tx4Bfh7vI2mb+EgyXIavzkOqUy/2sUvOJCFAEbKNQk+7Psiekk
7zD4r5gscr655HxxS2/PsVhnWU88qBwc1mclqCBvWt2qWCyJycIS3v5ByR5TRsdz
7zHM9ojIXUGZguRnTSU7+o1F1XxNi3RWfdeUiXJYDxDTNyOKboPMiaIsOg0a5nE7
bcxhPLPXsUM5bdUpyXPpx7b0CQoswYMY3UqMaZcjLXJMg0Stuzg+4plgRVyNhDOE
YAIfV5jAUWUB6HbikXrRdxrPfq/erPK6MezIZV4I1S8Y1MbreHB3HLb8NmirydsT
k5Rp9WP0rmnBiV4RWbHqP9AdglWbQ1z5biGDqS/11GYpAZ/tT2GDss/FzYAEIass
qia4FGxgwPeCQiZGKlcyVFh9FBWhQ5jO8ZEwP1XDq8R857LBDR3EwK/adNGIyvtb
Kc35dGc6ODe0lV9cUfV/CufF+J4zCGRZbfbSb21QbTMO0bbbnPHRGH9MPlxmXi6a
mHhmdgZf2e0g2MQDJ2qKwxSRmrt0Ewn8HXtJkje89A+u4BhfRxIZnGRVpz/Sur4P
gNkPt3I3p0xZLkiQ4W8sPhyjiaKgEWz6O3rlby+5NYJ/t8Q7EjImfzCPGarX9Rf2
VHtHeDPoR1FMBNtzrR4xUO8vNOWojPiW94O3LflsdOelvxauRurrkSrQTaVprFgU
WBosWCVA2/jJu4vnc9D7Kx5scxTkIswh1VLFpb19eRmC4ny+JG3ECaXrcYsVUcgv
eYe9FlS4wwrfyDCiJHYOCuPNVJ4vJU2gBX1CuK4vLAVRdR6VLXn9SDF4/hoU033o
vzVehzdE7Agixq33A9opKYz7g8z9EFOk1O5pLJ9sSypt1nQXlOO5evdGrrPpkW8H
U0c93jWBsZOP1aeqgEmCw+3xNEHs7Z8GjbMvDcK7tfZkI0oP2rdpVXSkB9XgtCwE
pyY7W7IIlT7K8UVlhcq9r3hyyYL5Buo/LDPe0/r2lUGTPQEfDjZfku5R+r43NO2E
O2yn42c51Su5jmmt4766RaAUI4Z/ujpwndj8h+w1W0SCe0h9zw+JIpEBx1tcFCkl
ynRAZPxcr/uZBGfniHLPMMT2O4Ud8Jd32Ky3kB3aCTk9vdt5AQdNgwiViLt6o0ad
6+KB8fZmzVAhHJEEZ1YbfEJz0ogYK3b4fOHn4MwZAEToKtXMXwvoBkDnXosasvPN
AddZXBzJ0jONPDkUwXjnTKCrTaE+qWlBGafrOT3TIAK32cCh7kMmJTYHzO4ivLzF
fqucOUDL9dBJOWiFWy8qwOIO4+5jSHavKp3Q6ZykB5miM3BOxAVYg4RBP484CYPU
Tdo4KD9KRHdxvFQaL0sErMhSCLvAIKsDxoi+BeHic7TrpB5VO8CRHi5IFZckwI/1
akga0iTknUCSITZFSsVeglYuIXfqqRcU4jF10U12njGN5o8ryDz8HQzpnyjGp4Ei
AJsoVj7SKz20tQ97xhCngtymd/jrxju4Va9S3vBagaS2qpK8cCY4QdBKc0Ur3ibm
rggj8PK8CD8zG+Y/jc+Td8StZbFj7KEyri1KdskHQqLsqFaukzGp2Ijzb81FXaks
rcdOF/gJncFS63tXAk1pxIXAMPjv+1gESW++ywwOURSiILu3nHfL0LWifAzAogO3
ArvJW89fStB676uUm2Wi69dKKLH4BcODjVaESOeUJsfu1j0q0VIRYDsDdPxJ/gkF
KaYutzQYB0/qj3zrRB8L48j/wx0TrjhB+BoquBOGkSy1hJG8rncVPRQ5Q4eNlmGw
HVYp/iNNpq8VbfeeeUVFSIgdHOWjA26IiTMsHmNkk+baXxANDtDud8v2tTRhuUFq
vf9D+m61wE0JKenXteLVMPboTwX6lYJTTaNlJt5rjyjJ9yXHzN0SPLEWTyhST7td
TJaaROBcGVPJFHcgBwOq+Da8fCl+XomMrIwPRGiRalhSyr8nhfOGxmdTSypRzHFy
l1xNEfodOH1xUEW8yVeANsVzY0US60HiPygSBEYHyIaazUz17+P+clHQo1f/DMnC
h0vXlcJGWY/B2uln/8rUF7M+JZL8tHHE2oJ4rRNGOUgyuew/1aYCpFKwalPENkQn
9RwHlMRoCMHM9h6CjS48GVJCQHslcunToJq65j9aWY/kOAZ6RT/gMKVkD2TMxeUy
WnKXdjaguj34pZRS7vJsQXN/FD+iQ+q2Klp7HlpK8utXGjbuu40ANYjel831konj
oiO2w3kJuxZUGjhg7HV2Lt23gP/Z5ah603uYL/I+80eV1MQIo7EPB/16Dua8Jql7
Z2rpLsqyunAwMy+o0wEpyJ5wddLl9nk79kEdN3Fodc+oQ1fclFEHJAIiLgpS4MCB
Yz4sxC0PZG9CDShX32Jo63Fum8gtzvVP2vUJxwiCzGjMrJ6RsbStYwZmgPE56sBn
P6x52olDflTbr9gEuiqjf/1J+c3/ucpWqNpK1K9uMSs06DdSssg0k1eY/vUIFUdi
QLlLVwvOMfK+tmHQR0DJMHR+cuu9O+oWA2hVBUmRQXlfKze3uE5R+tNRb/O739kY
QFalvfwcfCI7LauorKn31R5H622NAf+63EZTIuihrRJ3idtNZcNKoj3RzDyM35GF
Gczvyc2wI5RXBVqhZk0YfpuQDii+JdgrIGwr/TRFUDN4cbDUJRAvFKFq86yxwizY
wJ8i/S3EPO0NUjDan0SC1l5aLq80Fp6Kb0H8m21WUOXlyxE2Vf2F/VmFXB5X5ShX
8sjOa0s9zrX8xqJhUKhBvoMhWgB9FiSsRcYv9bdT3Ut4JNjdW03TFKL6HlQt6BB/
uvesTUMje8aZFpWUWU2oOB+F86XG3r29cixP1CUPZtBLn5d9Dy1RumrSJK+1XrgM
Jv1E8MJiua9u7XKWFYZ1ci+m6nWoksBB4pWYv7u/mG66yZv4o7IGRlT5e2wGcxT/
yucZCSMQRsUzV/ODy8Ahd+9mQRUB4CGZEjJFJ6/lAW4sOnkUaitcqOjNVTLKsF0l
nXwVMs4l7Tc7koASYGJ+NtAI8XUNIaovnsbPmZLmagk+QQv5BGBC3hXQ1oPeWc+f
cqV/EwKXJ1553STFRYrtd0pcqB0cCer2pzH52YXtAcCNhx13Zl9jeDqKt/bGwl/L
9wTdKvihwO70ceIgB4EkWetZg1ZeL9qmPxPmGD9mgtPckfFLuf/pI1/3voBmav+P
KyBBMk4CReClkHrwAmRixH43gkJ4nooQq3VS4v0bdlmYwG9cGs/V57r6vRwQXjPJ
qxzXmtvCyaDLOGX3uAm2kOfqCxf+yJiAbew2JjDhATl+7NlOlhWHTnraNX7lg6n8
nAkqgArb8QwwWcCumG3TKhvcv47v/KpguKlv6TRBn7923M7CYFC9IBAD7VHhjTrt
/HJql7HvSBFhSMoNKjR6SJY8GhzZZccqJkhfZqzpqRRO6g8rn4x8z3qR6kAuqXpM
Hifd/d55lDO/+4AEob+OXe7DuMHgAuHby8trHDBJXParwutv68A6kyQA8bIkxYzT
zEa+sq92v/2cL7Vop3O3mgPVauE3NFfyaoHUiWjXBVOVtW/qWszSt+AdfvHOHQiI
xOd4rRTP+4YVzD74J544/NQe97wksVKeJ4fT33WYxTpQEAcNeAJNuYhLSGirLaKk
aiIU4gh9XCJRudLabTD+rxE1zt+WiP66ViNoiyE/l9lNKCpBEBNgrWXHQfOBU4yx
HNSXdK+1V42WVnNRJeneTHNTGxWm9U96mpCsDPlVdYh1zLwUwHjcCImnJmVlgn1k
yo2n3m99ftFumBpUgcK492kxsVt+mPAnMWf0Ykqlb27jMRQdQRjGlQEBfDniLxHA
TFDMGFXX7UwNc0R2+OMRlYI/HzAfSqjuJc2JBNgVdUHZkCxHXq901l5ziIJR6GZr
C6RYnIC+Y6X50XzPpRg+fEMBh0vUVC9egdC1cxp8r7/5wPYYSxzgVVybdGeaZcxz
TQgEfUTVIDXpEpn5aFnUpAs4jSNWeAcJ/L945zymgF4C3VEDwcEK29TgxcMc07/1
07aa4QCaoQR+dI7iPUb2lZ6g38YNAaEw1GDPjnjz8ZhJj6kPyCXvAq3h1AfkhEtj
o1/Swbh/Y2zwlUQoz6KVQ1kIAdpwncrOIoB4jmrS93HRw38y9ief5Us77ym9I2zx
DCymb9E/z9x6UIu3dzHYpWDDgE2D+RcZxGQcNezw39xgPc6zVE61Dp1AZmDsy/vx
V1rhsuf0iCwhsxEJhG2iCPFKvgsgMDreMN+MHjh/swaotOMZTIY/N92a0goGSSbs
VtbELS1lvlxzLT8xl1e1oHHSlaVXryan6onx0A6sMNYoEhGhH0fpzQuKrEF5y1lK
4Eam39jMZyfLUmwLVGiQmQ4KTz9Od3AS/Yq/bqEZV4mwf0Rl8DTX7boMA1wcJnvk
573k77bXErGLSXjIMgUcntjQ5iTXTatq8RNSUMg9SkEfj5CI0pBmXCqjG0bM562U
GFbUtXiM4l7yE+ezIGPtyKWaoYCZu7AFY8yjRSOlEXZ6rvl6rCAVsiCulDPCpiV0
+8rgiy3ZRGXF6gOV20Woxns9RKD6KPMhzddtm2nGVAT/2Js1YCwMvY11OI0Ph3ph
TCkIOt11wSjDeP+ZdMn0Fh4oxeC59LQWv1USSG8E0GRX/d2jhayWv2IBG0D9ZTMh
e1QWWk17LvXTS+ydg84KuPTsJoV6xBU8SoaCeDLTUaaPUm6IQ2odDMYGYE3T3Ir9
tp0bn3Eeoyt5sVQaHYlyK/acAEN08bd6Xv7mUU4l9oIpqBsp3CLymtS8ZFr1Cb72
OYG5z5UfTLWoXEgmlpfaY0H7StHmux1GRKgSHcYjjymniBdRuDbVs3e1RvyzeMkI
aL55huhsjcM+d3Ui6NaGx1jyg0N7c+P7P86kpcGIzp8cebTdn1tKKpm19wnDy52K
btAM5ddZOCD1slLkdW59Ix1Zv0fSDXXZtbj0sJwYBsRU0Cqohfl8li5h9qDYB/0h
9B/bikmi7SafHmetvgJw7nn6R2IONQCv49KkMegQrwpRxJmEowEJTuG11BIkgAS5
Rcg8rswoMeh3qMVlPE3YZ4KrzFBbl0Pwqk32MNQ4+jU=

`pragma protect end_protected
