`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iJ/jisXI2QBsSTd7xGrgzcYkLREwkywwmJK+AzXOV+oDMDfi3vCpb2inqmJKFgaE
rzTyOdyiooXAkSK9zCweY7+00zdZKKtwl//MN6yn/IVwDsd+BNAFOjN/VHJ5yNHV
2vG0+KT4nzCafuGJoDWpHctnB1cnnSbe6sEA47ykCwo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25312)
SPlp4AM9JjKgwPP6El90c2tGFKAp8k1einhDeC29B61B0RczyhepX04FiCrB+wTl
QG4BBQl86qQoWCOFRW1Lii8cHkqA7hZlXPErXuN5iAXpH7bEo/6FsjU+SDjG3/1t
S1KsXoENBgzIXEF8jakeglw8RXYU5olM/YNWIIotI/EHpp10xhgpRTWAKsVLfBmJ
v7aJ1la3AdgVm59hHJJjHCcgdHnk09mpim+shtr1xWoEGz9+CLIra0xpZv6NwC54
dBLBzxhnpPrPPZmmM3TuOPmRRHhbFc305rrwZo0KOanwYBRf2A6+2i8CQ+U9bq5z
bS4I/kHjdPdW5CiUeFyZ0EyQy8Njcsdt4y3vPlCPTkzvd3juv8bcd07yMrznm3AM
vVJbt/SxmdvpGgcou3SpO3pvwlhQQBd54bYwC2YnyNowrauo2hfiaALP3f/aeo0b
6KESxHN/J61H/JLvhn2jIK/f1ForcTeBgH+d5Ec3pJ47FFN+GbpkopL+/gAnLuBM
1b6Cfa+vbwg4peqQZ0nWOOEHEYlJPjVGUbeMRnsmMMZDvkhQCBjfsNyLPZRbDWVW
sVGDYnbqOC6wCWWwT3kxveqoBBlNRSREGUoettEuq1PxIgq3svM4w8aJug3FDbNe
WOEzeX6/y9r1taWJ0YyK4ssxH5WSS6zPox3iQvFjG2m9zJCq8XtsFAVzWqfS47ry
9DtIklEquotvj30d83L0kFTJAQHPPotaz5FYp4rSnIbxV9hGSw3YRjY0eGiUmyxa
CYHdY9bKZyFtBajSaQXKc45MElUx7pq5zmL2ubV08cWbUvH0VciHjaD+1kNI4zc6
xLX0pSga8FMzHQu5PHSu643hw4elDWsR/hJ+gNJ2Q3G8rm/8WkU+DFGr7da/i+hu
/75LQP7UoNiujQV0cfsOlGGEOx3Aj2aDobAgTUTXUJWH10YhhbB+EV8aegpk3h3o
ot76j4DmQXvrs+xa0cCpMKFN63VucMESzRYVKJcGwJKwDrwZQ7itRZNfoCnu7y/+
OzkFbQX2qclt4au/9hqZSvobX0+fxkJIOoc+OJ5EL/xR868LLkNoKlFI2636UCLb
lfMCXbtVLyNDllQbwbwQAQgNZnJHIOsiEDhexWm2ulgAzir9iQoBzge3QRgamCyo
VJ3meAjYr/JIvXQo1ziO74v/WmbMd0Z9//By173XspOnfYTinFmb1JIM7H1fvb4b
CeACIRLEYHwgiU9VrnADmCTjauL2pHzGOQDzYcEZlgHD82Fxo0Z3ztDKFCG4SprA
t9jcFT4GWo87Ww4frR4OktHzOH6BtzfMtJ1SUz54IhAYyjuU/BZeAdSzGFKgAQuf
SCZXSZO/mHjzE2SoBQngtmKZf3kxZ9qrqHdsmPj8GG85zSnV3d6o5b40lw/XlQUo
HvWU9tQ6tUmpkB5X87E2//231PDMvJzVVInFincz87k8l6WvcG6NEwPK+QIcuKwk
EIPreG8g0AMacWy6eJPuonQ/m7oPtYMr6W3/Pi0nvOwm9Mzx9EovH3jvkM6YWULf
92z6Zk5x5N4tHuRV6uge1AkvrVnI5FB3z8V3f+4EZzesLbcDDN9N/5RzZR1m7bzS
t040ibHhKFwet3wXYsnJ1m2kSmOpyaIywunF4KL1aqvr7TjFHcRkGKZrLBW0w0v7
M8l5n8Q8tYFJ/Ct39qEFEDT4HxRhOa1NV2zqCZG+WZMyb2QIErTGAg+Wl8YtHWgh
3AyVkMqI+++XR7eSdqUhtfN+t3hDAQ2nNr/cltARPByvItUfoE7lr9+B7JgyD8Y9
i5H0Vdo3MmQJNw7IYa94FhFo6I7XifZ91kZ30YxajyppEjyqUEYssemf91kr93Wx
mcAbHSwx5wuxXJ2qoB9d6B9KqGh1pWCHYF8/fhim46Qs/T8OG4l0n75nC84jsq+S
8Gk6Y3AoQX4+9VjcLzUT7E+JwY2bydkp90ZnyCF7PNx46aFbOOiFR+grC8KPP+u6
uTgzf3nWgXRhJPiRzZvCmpH748U5g8dKL5M3wEP2uznG5K6TdwgO8F504D5bXKQx
dSu1yjsxCaeerdJj1Itfh+SVuWHLDnH2VBOu06d6AXHHVaSqmT+VV27s+4rsaDCN
1sUx5YCoPhaA6kNwinnKKdzgS5t1fXRt5UptfTdYWvolvCwp2k0+mMR853sz+IAG
NlG2Nkv+Pji1d+xa/HpuzJReRQNr/G8lzJ3AbcM1UkTLORtN625Fb8HhyezwOBoM
5DdUlRNMaCtQOYtZTqxCYkJB2lZnHhbgELG7NpKMSiXnuheMWaSBJNjMnGoOu3ow
WeXGjIySPwE3b3zayidrIzuHQmd1q/Gz9iKHHzwJ9Kfwy0oUEb3DibDxAncb9HRk
h09bhzmqyeBeAGwtIs8tK8BtM5a99+lILDN86BPJpF2T698YJouVp5GNmphS/6ug
g2zpUncmude5BqrgPQqukOmQQt6y4qLttHOMvuXNNVurQKJK93E210D/gPGvzcpa
W+kD27rjwL4lKJrKqvgAJlblCVctC/VRAv5kHGExET6TiaRy18sC48HvfP6+bq6k
RARHAMIfrQFUu/tHLk4uLzfyQwpLiQ1EWrVDY49cfAXiuHhyy0Cn2tZDnKKENMto
6dC7OdHkl8MuCo1DjVRZSSd7wUYxyW2Ca7YOKtwi7o8RIAmn7A5+nviu0lxpQ+Hy
fLe/SnF0p9sMdPia9v4pLfdhQ/PFXmIACod9/4w34gz/HT6sHfLD+5/bUkbr6ZY1
RkaXCTOaCqduomRyAlzMoe4BtXhBXH1WJOQ16q4FzbERBqVPTY8G39/ZpikK8BV4
D5UCtm1D807Po5woL2MoRnHPRWWI6HFwxxKEhXU9gB/whLm8UVGEaNg3GXzLeIVu
54xY2Qvga9ud/Ec3DrRn8jIPuEXel+HtLAkaUnh9YHnYplj5+8Pr4XnO+U3s6jlC
0JRQypzLcxDy+2K+o1RGozNsbmC/X9I/v+H2LEZjYQh2PgFuu4EnDiRNO/kIpmFU
s8uHZjWKz27ioAo+QAjGDBb7V6aOkQ2d5MaanrNBxfPTZi0XeVCw1GkOt0ucGoao
cXI13tu3xT6iLzul4puPu5lvtkTuQPF1hEpJI1Sd6TjxrQrgjFG/sr2TMuVQA8Y6
9I0rvcKyAbOg0sNXcV7aepaKGmtG5AN8ADCc2gtsap53CpCrKnsMitEdtX6tsVGb
62M1sQc/jUKuQxRps4JheypWWgHa2p5XzblH7NOHRIbo8/2zJbFsVAA8NTYOT5fZ
POBszwz9AQuGyWwlA97e+aDigzj4VJZHZhQmGyAheCF0jNjFUcVxtSJlclLOdUDg
ipgU1NWL6s0C4K5Zo+V8M4zm17ilr5WlC7rczzW08iFh+5GP18B2FgUZPSEAlz5s
5oA29nCy9RZUEQ/4mJ8LrdFSxKdqiw3uwxz9wXRA1d/QDrFOZMy6K5i3gHXI9/bn
4+l/qagaeCqJHqEosb7W1D9DC4GWHxzD/qq/z/CatoYN+708SxIJOpwWG29iSpDb
RZQzqtuO/PXxCpf8rM3g+OpDId2hAHWu1kpXX67PL1teJCyfhvw48p6x01nlZQ1F
cEwmowwRvO1uhNM9paAQ8cI0nsyk9+vHrtOTbjiLujslc2MeW7RVLJoV16CmhVT7
8AKBPcopFcK4kLejPV3Uv0oXI7F2GaRgw21ZVMOiUqJ6nwZRJLKzH/ChJZhWMZgI
tspTn1JsViGtsAgYeUhe8l7W39XraBJM25AgRgNsK3ERx64mBwzo66ufoHrp9bWt
xhFuT1OOZ8L6QDlVVwJBKSudM7srfGc8l3LPQVg7I9X328XgiPXiHUhqUZQm7Ttm
wdQvlF/UuhXwwGOE5RIYPVXy4jEtXZWRFUXdbNCg1pXFe8IfUpKUdL/Iaz/UA2XN
NeUAFRxeZPYKXtpIUysjKWbE6VEMIeMFDkgQI2QpML5ltEpSqSAgELYBbQ/Ugrx9
IoZsyas+ukOSguOSxYVPLTl85138tP76iA36tfUAMI9BuRjfL7+1Fy4stLvNOnXm
sNC1H/mSnxzHN7OOUGD1fwSzrHxqufNpThwS5DlpialqK7t0BqbcuUQCVgdjz2Dp
34A2SxdoePYrXxvuNMr6l+RKnd1GcsWdR/utofqOx/zMGdo2p2oZNvmecm4/R7DD
TSjKXFz/RudfU7zq2wIsLOgeqwtsqOPBJTW+3QOi8J61vSqKmGETRgUC7LBXHW79
lem5mtdEQZVCYKIX6RQqoMXqCKD6Au0R/zTS9zzRbKnXsHJwWFfaLCt9DSYqEWPA
xxXJtWEpm+8XTa2csJBu2wNd5TsUXjyQ8TWp1VDbS8z06UrDutGfAwpQF1ChYRoG
PT5Q4d0mFCDG10WEm37bkFNQaowUAgsi3tj5TnFb2LoXNsAXXZZ/m8jFqAmB/VQR
gHVdQaL2FW0HR8rrc/tYP+U8m3rl81Fbtlo86oTyiyLHyYiSKM4Br/A+JIu25zlr
+sVX3KrLdGsHOenTlJntx/b80NrJ+JabkB/F7w5LKHWSEYpK6tQ9/BIzlmOxkrpw
Ymh2N+OU/48Y9Z9c6+2/sCP179XSpPLEBi0nlaldTViF+5fGR+W0efS4Fi/zaE7P
z6lUVZK20jp6Bv2/5ezRbjhaAZGKdIHy9Lebowzt53kXZ/xwwl++rNIQq4KuVsaT
DiqtQyrDm0vgUHT9An00kCFTVHHnHRWQV1DLxFEeT4wHHXxjzsEsPwnmL4EWaS7q
jBYu6sBmXU4BfsXKrobsGqXbPhMvL1kB74R8E4F5VqdzCaKEvT4XUIkW5ew0NBHH
g8VJ6PSaoJpxAGenI1NxNin4HBPbZNpi8ZO/xrHw2v2nBTsEPwAffBOYfWRdVrSU
6x3SQnsUllqsAjDge8tTPC8OVPBjMhOYrBqrrd6SDGy/b76Fz0g8d6UIyliR4KgZ
/M4N+WoqVH1IjNSpvl83e9LMZOv2XdVJSTgMRteKZTU4Bl0mGVjmrYVBOETTzOrN
iqvISkyIdXcPWnUgI5bsXaQipz4zrtkuC84nBDe/g6GLIg4v6bHYr7EE2eB/DYDK
ehtcaxbAHIKfVt3n+PWSPxo7wBv1fBY+tRYDlazl75IcCpodEFl4kFlSB3SQvhi0
+NgCg5lNGEm5O/4eP8x60ARTLNZ6KtHnyEsSRbTWrXEOOp7gKzYpAbEHZCOZx0mm
3dCJU8fxZbkewQqldT8ZBr/BclJ9kV4rIg5JTNJrL3RGiQ0xM4Y9p2FHig2iAUwA
djGitbLF/U2rxASuiOGNgc7CtCYFh35A8xewjipSiUVdm0VFJp36spcvinc77l6w
g6lqfmlr0L+V2XoeklIXFIRe+rYgaOZmJ5yvQPJMVJARY1Q9LkACJFDOyk0cF4vp
PXVCwqYQLrrj+3Jbd5rMfN/CyGWPSPq7532kqZYAO/byXQyjx5jLKsvduCfqU6zC
ramQQHUozqcjqCWaymYdKyzFsYWDV2kjAaEUjg4kwVcqLzHGDU6nm2L6OTCbZ+dU
wx/g3OYptwDo4z1LweEY3g5ihzhDkyRFUMlTslmPt/el15Kt1a06a67dcPD74QJU
A0IsmynqVI3F/m7109KJ/VdhcwpbtKL+mJDiPBSQOCAT+nTcdeoE+sB4Gu42sV2X
mjMn+8eFKbzHARq23hisI5AkT/gug5Ia7haabVZ3q6rJ8QJTW1qEPeDY5qtTan/P
zqfdiRDhe1DT7qDJKj6m35xCiOyJtG9a1HF+b95Ux42B52UaBHZBLrsG66Pw1le1
NmQrzdDvniBR/BnXjNAVLFs+LaJZMlXUq0SLp83/IuYKWku2+g+wEknbuBaHXs/o
uDaQMhXenIohYMnrXz/fyLN9EUBrIiDDFVHoilbAt9BqK6Ctm2uIy391SfCGSLOO
G5XFHLdYZMgkTl9BGfmK3vLP8cIyTpvibEX89VaHsvXY0ntrPC2tpV85p7rZ0KYs
chIQsU6zJ/u9ykqlnA6eQ2t9ErSI2BIOpxuUUxqEeyxu4PHMhnjpDgnWWj2qVuVB
xb5mNPD9xyWHl5J05Wfplc3kpVK3quIvQFeIChJZFeKcLpcxZoKcGyjSAI7yVVKB
O4Rkc4i8atcKkQF0vqYMvofHz5RnYakK44tPdgVdH28mrrl+OLqlZMFEl8qxaAot
z6KapM4pWNmeloddSsotXx6NBHKry6Lh3hswZstwTZHYQEVdIvRNti1TZHSGmN1c
U3QDq2JVsui9/BdRwvoQs74VqWTmsa8/rBaMGIZRPnbYOccLIzzz3q/w6apHCTkR
P7mf6by/nSBoeO34XEpgXEET6wcWR/6QgDHKXduXP1Cs7Uio9sRoFLTduuFtJEsK
c2t4nKDdjBw4ddBR6Qs4Gi2+aBxDAEeKUbJU1JafrXc0AYDRVIzloEJiRFTnptUP
gxvGeaTd3JNHPxGbp3aU6vcODvOdRVaZR+UY5es6+OO2mn1Ldd0k2SAy4EbKfKug
n9PddpXr4+zi6FnzyYCDNvXG5qMnL+kvQrRNctwBCXj+vxlCNh/VVblIvT70qsxY
U/fa7bGxD1yq8ICdmYZJPCrQftjj3bEVkzv7a7ZE2o65hM368uYICaEwKx9FZB3c
jQ48UlEqc9I5o09OlEzeQXE7VdFcjc4jzdrvv2InEKx2FDRwgLmbtsdOlLCAZqz7
3EBTreYVvq9GEydf0rlZGfa1OvQ8kVy+4LiCZEPvv0JGTFOPB0YO28XsF6In8dI4
0rzS6RzVgCJse1H9IVKLVfuSwwtHOj5HkDDwf6DKPUvMr8k0EXyvVbjHKMorj5p1
FxVUva05yP5n81YMZFj5+/2PxzyyOUJ+U00MN1vqBrpFqmAuyO+2efd0svyeqSxb
bF9otJMForFLnA6L/YQcjGrb8uGKAhY7KizdsAJ2J92GKwcyKwu8oF263s581WKY
l8c/UHuMmJodEx438eNzHwvZ/Rzqf6Ahbv7RLclcp4LdDjyD2KrnYwSk0WpTtaPa
hvRXiVedlRYoZmBoPL4wgr5IWIJkdBKpKrZPIWN5MrF10omzfqRrHeU3wSwoaF4K
mWiNt+dalk8RjwpC9epaWmh6ccvQRqZ6mqehcz6q/YSSc54yqng2fcHOMgowi4zR
REvCH8pnFLgWSOR5udLRIeUujl5d9EmzNyFeFV6USynhjygB90xF7nQr08wj2vza
S5PAk29KEuQhifti2IckhDlHm0XjJQEgAax8caUJHvx1BLHAHJGt83eF5P4bscyp
2mt6RuYtopQFzA4yfUXMCPNCHyP3RbOKWLFGm2D0juKNOpbOBGJhxEaXOjHWEPh+
4BYUYB9s+XfOtOjnsMmChArbemq2i5htAEl9zw/ZOjtsGzFvDLFyppLTVEYGP47q
kFNTWu46jrcAaFSMQFkpidES8KVb5oGGb6BgHu2lCF7IQzyeMWFmzpvIa4DZF62y
pouMdWDLf5mIssMD2ciRcZ4Ci1TKajvBhnm9Zv4T09wBTCGL7ns4Fn37q7QGzW18
fWBzMk+/eVnCWL6J+rhhf+Snv6CGJeNy2q1FRY59E101wXkAKohmPouvu8ZvkQlF
aoVoNJvSYT7ac1JHeSIDLNmfdDdGuUsN8RdgSkvEqRZCYurXfcVcq7h5Kg6q3yX6
e9KzzRRr6L/QeN29rHVDBbf3CiqzxkpviklEtCJn1iZnBOvY0M9MlGqeaz9r41W5
FtpD2t5NZS3zI64OztlfaA/IF9uIwPSNJWA7lUXi0bLRqhuuUyxr2NVSLzsrGeyn
2n/tAPUck1H2KN5gZFSfM6SRkH4W+nnw+Bv74sWPMHPSJgCV5NgOmpraUAsqlFRX
J/EvmJMbEQrKaU+zL/vzTX1ipKb4uF2v9WW0chxonEVOXM0JV4/KNE2qIbSwM1Or
nW7kVzsctMJ2ItAOALc/fS/K+LE89rqGI+1eEYyCjTMtouGg1/JpIJ+CQkpF8hkb
zFKtxOjZg15nXHgqmQmPVYK3TS6Ir8Qvsl8VRCQXQP6S91NX11q+DktDwrskskeD
bk1/oJgF1nlrkZosAHe/mdonl5FuzU/jt8Eb/SJPzqUYgrZe9V64fkX6mlaAjHw0
aNRGT0Xr35oaoM1jDIUWA+gr+jgzxtw+qdlkWNAOfBbNtl+Q/JVuFCVjn/4YYWtV
liRSbjpplLDHFcS6tcvoHiHjRYRKKtxmEYlagNOxXr2pPwVxevhWYh/ntXLtsCC2
UjiUygpGokv5WfpiBgmoFZZOtb9kksMjeCOMKTwwQRgvraAMpg1LampLj2UgPgC/
XrcL/U5YdDr4DsDazqD7Fi4Cnb7EYFVoSfqweeDlvwSM81DLeOQMLDtryeR4KEbT
8W+fK/4yq3nh4B3sc3WtRZCFcqFUkeaV00XIYqEphbusWq9vluVRLofwl5uxaVmz
PWswC6OdC72zie0HQpWmOLsCQ5iQM8fv8CG9aq7M9Bp41HCTJyrzEC9alfzDsoqA
WpMpxt7wgmZUV5GiFeHOLJKEXaw7tkLPN+M3nDapfDbdabt7Bxx6fLvG96HhlzVm
9SY6VnKMwOMYFZVcaRRnfWd2LqcdxZc1KLoWSRKIiMMUsYCrRDaGGtnPa760FoS3
9QLrn9ocpABgHOci/L4KQVm1ue8pmpxOdV9aL9uwtq5u99HZaGi8NbF1SO5is9Pw
7lKuaMFJI3cafzWhkLwAsS+oykUVtvc5wyMNhJOk4T0IPQC8CM5cMfcBxbkmBOjq
xLwvqKldZXmcVH4Qj4YG1LaswPQlXgUk++nH+duJzb5gxnMxy5vodfFwG8W2fVhX
W8aT5P4ZVPvXz4F+UDN5qXDUjIbtijqUdna9UlGFg2V5q3I883ycvC+AVEBmtQYQ
UvAy5LnijmideyyROZ8sTz75MgdYU/KujXRtyfirOzad5iZqyLly6rLfXuHoW5sw
snVh7FGXQWTw3DTqdalIxe/CasK71BvEgASPK0t7n076r3pknzA3X6gdpBYfKoNC
GW0D2D5AQZk7mjDfTT3Nr3xzzWQmJ585y61RPq8qPBboh8KMNI3dldjhDvQy3OlI
e6MfmzD9A2JiJxNcn2H5zG5qLxr3vACeIgmsWnSfWnnZY1l5k3D/P65ynxKu6XQs
gkSsPpr2aGKXwIoEEhnyHidj1p7kwtWXs1aDtTzs7XmNtRAANh5EahCXXAg5jJPu
XNkk2AjpvBfzvlm7paj8iHtMZ/cD5uB5AYDZ6fPfTIdAYOA3nblk57OPz1HP4yU9
YuIU8xUBwtMHB31ThJwRuMteMHrRh4kAkCGdoFDhPqQ4zLHlUEtIjKJvWmMLRLzb
7b2I3LBTS48Snn1ElFvYmqr7i20hkCTQdcCJHcZm4paiVYNdoL37SZmH1GqGp0rK
ehVqWYD/qZLJ9mcvONeiGFJ9qizaQpKPTKvvbaSs7iTDH3nyH4OFUwWSIXSlvV7r
cOHYhKWVWVmcZVPZIoC32boMFB9bQLr45qyqAfzmNwO7aMTG7fRXtRcnA4h83v1H
mFBEV/MVfEeaETbET/Ec+1x/oLEsoZ91p+lHgHfImz0Qs1eh3D2J1X0+HRRIRCLM
3ShJ5IjNltbS72GuZ/qAyWCh08Yb3BPJ1/iuoGVG7c3koHlpBlufMMCwdYEX8laC
O2ucuD6GPCr6pPP0TlUZlNnGtsNF9eUA2U6kVvEk+87k1+X66WFHw2ROH6I9GOXJ
+9hh7hwXAbJ/VkXeIJkPYDiNJtTvTEhA3AYgqZxbEiL3Oy4ocLZM2p/iAz0rbrbl
pxNdzD1SCiI9c+bvvlLSYFgRtnW5Imp++4Ug7Ojc+EKhWilCxGgxeBAG/CYRxrEU
Og3ZoJCg+RvfV4k5bMGTOCZ3Qdz08BGIssRqPJYZVYxnEp4gw50fBzUB6HkIMPB9
wJyu4k9t4ZyH+Hz5s3GOTxOYzSA6fxUzv6bsaOxVBrFakiVgwnuHRSSPlYBdE2Q5
0tMdEsBj0nY8JXRRvqRec523mo4SwP2vDD2vYJLeWhs+i5Cg1rBSL9vt1WvaHapy
+YP48aSZ8mofpvbOKzWbxNcSvdRBdSISC12ponzL3kyhH6jOVLXhRYfnPD8OCbvF
EvbyDeYjaqa7kwH15LuxwhPXNr+HY2CjqvFrhru/MqVcUqvOdrI21tz3FhmutvKk
iN7Y0x7QVPhGwLFLcsO2jR2ILjU/RaroJ2EU2hIefNURy3WLzMbCZSIZq4/01/St
eQIgu4/1PHDYQ4C/DsVfcflNe6DRL+zcMKxE7n7KMcXKTm+3eLAMvXjC1gkttDUT
oO+gARJ/nKTZGitq16MY5HoWFgHTs3efdV9ZFJApbyPgm+2zF+14VKJvZodWWlyP
USb9Sxrp5wppUuAsRA2xuH7ClucNqRAYIMZ0u1QXVsXaK+dNUBUK0eOuudFrzTLl
vu0mkh2d67S2PLCZQHd1QHizgNMdasMjVHhLN0OSLr7gPt062p/T0EaKMiMCU3+A
ghrZmf+1dUXrUugddxqxOCQrTtCkVltjXLQ+qdmKIwM5ETOR+tl+cmx02LZod9JK
V6Wjjf550wSgDdGtOVtV87up0A+SlAL+O3l4WUYxkXYWl0BJpQy+Zd9n2FCD0Q2q
7t9i6Dl+0H0b2ral1Th0oipHGjjNldFbwMrw/G2lUVx4jZ30ajHtJcly65qip1xT
+03X6P+oUKCnzNRGxIZeeEb8Oi/bSzB3qdMRbKQwO8MhWkEeqQgpoCE5yzSpjidq
abpMmMMGM4EoqQFDI30QwENRlX668OTHtDJ1E/6XJmOTxPdJI4fQ/NFf7lyYWR25
kcxK2Ve3613TpULXCquF4SBAjrTv76iqGkHjJ1WexC2+2R9OsWqOHJTDkIeAY7QN
Ja59vFp5e/d4E+kdi2kj59ZLtiOIjlqvs/Zr2dtnHGN4QSe2pbxLYlRGNL58HXJ8
JBh+f/8QT0JvJV+rZ0xsmlwj5jja7qLx5xF2eFxrJmodKWSbXOcVJLpIUC2W5Wn4
JXr5rAxsGJRWxBIZGTyR+ImzFFtz72tyUZKdZ/CzBQUSapwXedu6eNTiCE0gKI+d
kJVLtCZIDmCi6DFt1bhX+m4ejpoeLsJF7UOSy3ZGNjj3DCdgnAVo6ZD/72Z3WNKu
Rz/am/TfhqIOSDryAVE0Jix4a1ok3WPikcXv8scbxKkPrNCzxjsPOisSGrdve03w
bWlG4Bw/aFb7j9yPskTemVD5mQQ+7g71vu18mWtnDL76P5yM95MDkfNzCg2eO+/8
f7bLi2hDffSil5tzd0DDVJdveKOExjRjpZHfxNIGtmBgnr78SEsv2WshipJKY5wi
IaKiP/YDiVSMn/g0c/FVIehE3Y5qEB4WVauzqF/fKoNdc7rOi9w7R/Npijdr4YdQ
Z5Q2OpR1MmJXNypEsTyGq3P0hHWIAK+c6MK+bTRKTUVpS3vkjwM1YPsc5us7IpRW
HiDj+eA/xKX0YYcM0T3Qv7G8miZr0qZF0KjsB/TuSKTCPBL5nIA27Ez7cv9h6Tqv
o7pDOUHqcqGfGAjr9ch3t+xDvVUd3LA0nia9RiU46R/lkWcp8dx5BxEpA6sil4rL
Rx+vIuE9O6H9HoMit1iNw+Zn6NLmEozWh2Km9tlt8ihd+Xbt+ysjSpbmUEeymza8
zWILRvOgdGIb8pnvfnQNuPIevDeIzdzRk9dX6yFiW8EXdE+XVDGd866RsPGjlrW8
WkdBe6wElCx9bt+kSE8ftIaW73uRbgBqbSQ3vJGFclYoQPa3JqAxHjf7hYRFdvct
G91eIiE+M9JTohwhuBrBCueHkn64Xt/mcNvVZBG2RDIVbxwFFOKgDZPWVqPUfC6q
Px3zBEQK162js1dr5QCn0UFDCuWJpul2sJIdb18PlkqdVq5mDa1Ld7488PSO0ig9
jahEoYy4UR9X9kgpubUf10Yd5vqvRux60hsNg/RYgp1/jtY33HSFM4Eh048X/Y6v
sPTatcaZv36mtAa4B436fbNNnUmz7KMd8Xq+J5Fq9FqC4NsjmRWx1HAXbuNmxCXa
Pkh+OoMWtHordbp43DDqKvSqnOA8r67Rk316hjeWU0b1sa3cmrBiEyZnJdDUGmUp
3RqREYJngwO37SQ11kjvWS0VVe7TIePrW11Qfl3VnBjT8eYs57PVA/qS7GW+eKwp
O+6QXin9mh/CQtgd1kzsX7MsyZIGH7taMMwuEwE1DkWWGLlc9dnP7QWJyKUceY8j
qzySQ2oePaZ/ghhg6Nwmaek0PpatRC9BUJSgBU0d4A1/JV+Cy9OED/LzJX9B9KnA
jGs8rw5cVOTKFYUA5Ti4qUimFnt8AvFJgcGh1Yu94897IIpWZMKAcGvh5rqkFy22
921uIFEWd1allC98v9Szib2IGywMHZJlnZAkSH102WuC+/7C2breLM7a4d7mSic2
tfKOoDaZyX3d8kYc+5QU8dZgq6Rdk+ZR06JMOft5TtLLqvAr5BmbreGiDv+JWIaR
mc0mpBfMIKvqVnNmeYHqhJcQxRNuk1s2qWv4UZ33BDLPof6n3cPzqVtQcN/RuLNk
hw2aSMheYEhrKGElnXv0dptN8NM6bdj3fDeOeLj7Ma/47YFTADn8SB1sVFUQj3i6
5rsPnW5WL1i9d9t6y8xWktWiBUmLN4K3r1nKGhJSf4lF9w+IOkLnuZQT/T882B7p
Pdx7OFM7oKYvCFa1eyMt2+jYJ5Qa4i54M6DUjpNdcZeuDCNqWNHKEoq2wMdOjCM8
7vmxfEp4o53jcPLIFPVKhwCnSrMw1Y9D79tJzNCt+kBjOniQd69AarvTfdLbt0MJ
SqHXetTqhL2Ia4FV5JHrlolWfx0Ku6rNnMDv/3NmkhwyV1/e4aZCl2qnK78hboXv
jaJC/H1zNGCTXyQXrrD2RvqvSAGcjjXvXxhidx8hsN8O4+xOn3WHZ7yvj8X/4X/r
13wlMoUuA4rPk7rYLXruEcO3jf9A2q3Ua52q/RTolwcAOnugX/x3GeonbgsprLmI
LR6tQT8YmuSF+/MTVNWcUi/us+xi9fUOAw9jduccKs1d9cDU8jA6gOO6euaTsyIF
D/bFcsZ/JfZu9mzZvkZYzGz3gG5rbfu3KWpZj7dRm0PsdgAMFpm7fDV58t9plHel
042h62UDSLO6qFWXtrKxnezXTntt9sbt2dZXZ0enhUatFgEWYywc39Wgut+wIqy2
OOKdx8RcNEPK4OzN6FRzQwdlzPOa9+WnJ7T2iMsjieVX5veJtXanjh8ZFJuBPbdh
1phjfSl4ybxrkD6SNZPHNr69CuMvy7/im0xNaUjBAe10gRcjk8wH4gEuHapTC3d4
RijnAMO+AqOXh6mFPIH8y1tfY3+Czs4a2m5hHfQHcl7vqyPxYoOqMEM2+5BUds39
H2o8hVpbkz/M/XCvQcT+lBkbEIuJQiaMqG5bpLGl5W6c3sQ7db4fLTrdDhXLGAJU
QEdulktmska36W+1PD2WzKmth2rOGQ4bAAxY7/cQKhQeUlk7i0gj3D6H+gm0WWxJ
37UR68Nl/OdcrzBW5U4e1oHYtIvn98NvgutKC3lOdquN9cRhG+DmwabWc06CMC5H
egPj1ZJMMYv4GIQrpg+aBftcvcF8LeClCjP0knnzuQBYa73ge8kxANNgoWDDxGGl
qXm+ke37ZeaaIn996bjNAJl9GH5aA33lHXYM2XMEaQsK8/Bze0ykFjsno2q90FgR
r9vSJGqGx217VhvETcfNDX4sdw5EAiwG4nvl28VCxok5mheHu05nu8x+wQxk0tAJ
aNONa6fGU8yAPyB7Qa6Tolk/AUiIaPusk3Uuon+pk4IaH+hX4sj3dfSl/wP9ayOZ
6ufgwEGoPyygvd992iCJxui89oC16KHutIKS6Kiv/S2Ep1mBGU1suy6VoSTsLyiw
CZSq8JxA9eVZ6qxxeHj5mq4wIkKzYtafk4j0kyIwdpKjghrl57X/Ja1/wC8rc8PF
rg+wAsGaVYoyWXoWRri6V9omkNeXfuOI4XYUrTi4MpE2r4k7bpTeer4elbwE6Ldx
1Nf2zSGgEUxcCTRCMlD7Q5ydVkQjAXpwgRz4B9EPrlHRJsBH/x+64y9DcrlCQOMj
89/SPYFz9udfPDNKbAZAXbC1ogQyZPDo6AHAbkMnlkKWLtUH+GJpbbCdqyV8iuiq
o/16TGErPOBIc7bVNT6cVq5H2Op2TNsPnFDARLSUfXO8C4uPSzij2qlICES6dgGT
9v3kB3brzQGvoadGC6hZ88INSXssZ1O+IhrhR748vpQyPGYgIUJxBgE0TWcpYhyK
LEmUJ7zx5TgXG0aU3/ezW6Ajx8ty8mS4cT14VrxflF+5cY6C8XY9ZI0h1vaN7cZO
jnMFL2InBrbJJ6YcK3C//1TEibJRspF7s3G54wB+dxXmcfXnYVnCqE150O2VU6tI
jUTvpY0qbty6tDQR7/vJjQlRwixfFcbnYz36wBM99Qzxa9u87Sq6NDGWJDs1wiBx
6xcJPQtluhzwemWHLoxyRVipLW7ZVwNNCtWuJJbtw4ZYLUj3+1cM95IL+gIkGkVF
C14RdnZcPNHXAFWxRsN5GAMBMVFM4bl8rIH7rRRGktBdQ14NYCXKpoX2vo934IOE
kQvDuqbpnVdogzClEyd02LyH7l5Q4CEEVv9ByCRaGnc5rKeO9uVqLprEZ94s76O0
vU9js8DW4wlsqmESNNqqOjZyQTwh7J0WJUjoN7S7Y5taZdC105yG/9owmI2IOMGJ
/ci25azO8l1PYPhooCh8eSfMch6jWuQs54pRCXMCpmVJs8zQblaonplZliOFbTBy
/ueuv7AqiQIGV1p0gK+LuVJojY9g9FddX77iYf14pw6enMkY91HnaqHrQ1Qa2Tm6
SDyrBwZZAq2fIE8LJ98vfZDOkR0K9NtaETx0fxC9ctXUr7+1cwWkiBx+15A1Yl90
4xew6HgFj9xL38L0WPSlDLIDZS04h0OkqPikosv8+TwI/6SfSconruOCnNonm4ph
/Q/Zu7rB1k89YALMvwdLcdq250CfyLC7Onh5KmHU/JhT4n+mrtVHRGWrj3ViyYJd
YViToFDk2bUhpWbBnVFeWJm6fzLHliRf5xN1hj4442VFXtY2K/rEW5d9g65pH+9q
3Q2Zl7VtYbF6vi+EJc1mrye7uOsqbPWWZCrlJI7EkBGxDnqVc0+fdTMZDF4EuF47
3ulNAa2DtF4nWptV0DKotZ0u/aonq107VBFXpWPQ8Oqo+TeZ8rFLZ2rSR9iAJX5p
ctvBnAP0VXJTs+yv0rDNGrA1JW3M35HbyyT0LOyWId8lMWMegLnwCKGolABkaBqZ
duWt8zG4fyaRlUxTO4jMG/4gqU42jnSlJGPf95xnK8AMbpjWFoFqE8KmoYyEsvKP
T3JzNYKr/jDCFEf/eWdNa7JuaqFKsfFjliP4ob1arROi6LaZdoQqPL1RoZQq6p9N
+a+MlvhmPA+PntumwuUWTMm0BgCXxkBa4/4N89d85lfIGMM5FojT4wDwNfEaG2HT
cO3ag0FFUcVjDRIiPGQmmVAPmvKA4ciGv+dW5AVcYHV7PKR7+tBTRtzh5fHNtyG2
AeY3/Clw9bE893sb6vpCjLbj++N8MJ5JylJpvdSEHpTfKbkAWZb+2fIOkW7MZf8V
vIKoM99rOUtDkAGV/lQ7KUp7BWQw2x07irKrvjmlpDTO7Hk1KL1iI87UjA9cbUNt
XTJH6yN1+V1gH/Bd3FKeugl+/9tQmx8ocAnmVcRALENGKZUciI3i6WOwD5+rHEBE
VU/0qesCTFT4HwbjvwMbDOegKwPlgapY3cBtOPfmXo8wY/jfHN33H2YokCih7fNZ
KbjrkUOaM2kXc/nDEuQYwrV5s5qAMWNdNpxN6mnupt06Q5B1P9lepMDdBfnFxS48
8BqJ8b6AtK9Ngf8YdinnBzrdUDGh0FGRGgWiL54/2cXYIy/XeTpi11llpuTDYcCO
e5RZlGGeH/v9Ad3Q3Dx+eU/p04qnF5Ggn8Ky1ERF2f9NFUBTCigKx4HTsLgjX8QS
RujR705mhmGjOhMnBximB87iiWQEHs4pNLKr7Y/VHvCkyHfiUJwN0TiCibeJVym3
owfVuDAkobGkmNR3IUuzGU6ygTWVDeqfWUn+J4tgvkW+tALSuHHP3y98hEl4uyMI
ovoR8+lOo6FOtxh2C4RRfOv1FZ6Z+DfwupPwi7MEtQsTfp7btgYKk5s662h5IZjF
NvJA66h3CeqvVeLL8j+uaa9wWyvsCbs6bxYM7ayzQ+5PuoNPIkNlLQzanLiuLCIa
1y3Qwjnm7KxhqRTaon0UzdUayiqIElBnBkjrNjw1D059NmMntX8T4GL05HuLA7Wh
CNTydLQCsIJdPZrVAVvRXDjPpec8fzalWbhvkE4HoEJ+lphBvIMCyh96+HbYKal5
XTdToXJjF2yocXe+LilriXUr7BHiygy7duXJSLUz/DS9X27RQAM7FCVzvmZA8ETd
Jjs3ub8TSoHcEfgv3M4+nox5IQu86prLICwzEuIr1dcf1j9BdLcpM3x5EFXFjdD7
q03+Y+zmshHf/VbadbTBTngb5+976gGRl5TAukYr98GMTB809eobxpyeJluCYAq6
OSh8vPEkd0ArCrMO7qY6uv5Zc17fJMecchCzL+XjHGlwfjQaDXxLZHExA0ZtKGhs
aWWh+X+ImaWWDaLHvhyL3GvM8L03PelgnOnrGcITw/2N9n4bluJR2dgAtGk5bT3u
Wvx2/dDAF5suVa4DwcI00B4TwlvAhVCm7eS+zwlFtNvIDbduAgIpVCov8JX7ITHo
kKQvKr3che+wpdUGgcni/CaaWw1wjezwh86scpa4iPP6pSN9mbcEkvjb04CXU63o
Ho//dtLrdiw3lkWKWFsIfNhomdvQaBWX5Ilue8kVJ2WBL1efqNEg8wCM7ZAQ3C1o
cTB8qudCu5we7ZUiYROB6U8RSJL1Uq+JUfx4abNtzNWbXTWK95ztt+OYRBwU3ZHb
ozmcEV8km38egAIliq3Cniyyzk33KFuMfAsKX8sjabEmmn/3Yc3ks1/kXh4OGKjT
xguTaBYkvgGky262ND853Tq2jni7owSMmVPfsOXvB3RAmcltJiKltII0hx/ChFjk
JA9KKvAZtc6ekVJIQHDU2YsDloxi61HzcF71HaH55dgBKvnuDwirRbcDLBnaiemO
0GVpmZevF/htFSMo8xbBBB9gE/SokZ70VeKCF/KNti8Oe/jRz4b3MbFzHgLZGEXT
dF9Euj86UhwBoliWgE2Ae6IZ7I0aqIUBXa5vUrozW4jJYU1rpOHIbjEqc+a7puY5
iYkbE/t6qQKbysanGl20ZieYnE9v87qi6tVFfHL/yAXvSnm/YHHkoCbqDU8y0Pry
208hergQ0BYVw3HlVyJv+o+h85w6BdUkKkzlawepb/LSnb5sm5C6nf9kxacUYaDU
AqjYed6dquuZWCJe4tAjzgNQ7BNd0rIvce0St+KfT/tQN5U9+kFYjw1Wj95irhtJ
2TXNHRt0ydWb6iYjXVCo3H398GFdbyoOKasn2sWRL89/c/boAUuJNWwdvjbmzFM0
FIUY0R7rF3FEOmqHZnbn++X+FItWMX9dG/VfhsQGWG7ouAcMZc5JSTxeY3DaNbwf
mw2/Hns+KmI3IykKxTO5XlKDDkXZrnPXYKrHEtWSdaaw2D+tC80Wb1n5M/9oNYFC
sMUoj+8l6jj1FaddS77pc0Cvrkll+kwtvYkSO1JICnxKuYSCqLEuTDLa+aJ/F2ej
1auy5Pm3woaEhzV66Xd7shxuhfoVkvoteT2TDZc1L64/DggWZRprbOfP5xtvTNh+
wx9fJ6ZXCKOK1w1JY9Q/bG8H+TgcYiQA56yG0M2rMzlXLI3v+o5Ol1mQmVwIfJz1
IalZk/UZVd+kK9KN22YMV1NDf2LRmyHHsS4jGrWYxEKEKo218aRSj8hFx85Hrbgm
Ri94G3VqRLS8KG5xyZS7HxDDicI7jYis/KDBSySvMVSJHXp1Cp/K9xOqnzanEdCf
xeaqzJiNkySTQu6E1hNTLy7ZqNVfEMaYe7TGfvCxaCVpJ/FPXg2VKPBpvHf45fsM
aZ17SHLIiMTUEgpeA25AauzWtoZlxfXmlpWi+fVpTZq/WCvRDGdmJajfLw4jG0X/
2haKZfRvWNyZj5fXx4Ppohoy+ebOY/Ze62/wABU4UHvwnopaiD3Mn10H8qAwY2kd
cpZ0TVuJQ4x7eWiZCJKx2IvOP16kf9idczIUPJaw7Gu4+LrO7QDPr8DsP6vocq5D
rSXRRx9ZrBahy2up65tZux/22L0JGQ4+xjzPsIZR4+s3pXjBFFT8sK6haTevd8XC
ZQz6/mXQwI1Ff1ni4IeGX7FIN0XJ1g9Pyjb/wfk4YLUQdrMkU+EOp8K9jOPNugSO
CTb8sk7ypEy0T921m3mfqoZkcfQ6sWaVR2vmz6MFU8Pxnf1hS+uzzVwxCVcJjhW+
/3lzPX23JpNcQw9E9xbFrMsI5WGqVL1l+1bnWvymHwFy6KYGakn/hBWcKvZw6sYi
qPYUCHYU472dI6fSFrqgQLTyEdS2bzPVjcJIoD5wtJ3p2FBVzyZzsVL7H2I3nlRA
k+TpZA35yvs/BpowfZTkDoCfk5quBHEL3N6wAmUGilhX1aqMqTUp4SrrGAvS6ZVq
L1oQET/5bj7AT6HgtlMwqcd/lPid3u+9a7R5Xrvd8yG011Xm+57Xqoobk0KFGhlL
Z4O6Byke8IWFYgZP+0/bqgWSVPAy0AFQdNBaR4kTK0G6CWgTxe1lpfh9JZoRjxzJ
/pjYG6VagFTYcQ5X7ptHkV8fpZ9H86EkKCSco3t+/Us3Dss5ReNV4aePlZZuaz+1
tmvaXqVFiR3E3IbcZuj9cdnFEBfJF4SxOVhrp3R/FB7V3AIRT1pa8qYnYaD2P3Hw
SPJhsRbDWPhxfQT1UNdtRomkX3bioUl2ZKhf2gO14MuAzbZl/fPXjCPubk4nn1RI
/Qg96LP/9mIHDm5taM1DxIUaO7Hx8sQEadjrhf8wPDBjre5eHvf+YMIBhR4mXqfP
U4fH6GRJqwUOPbCRrsMGnnRzDaCzBWX4xFnfNJEVsNtrZjFcClh4evHM1iMaqEzg
pwT585EbqQOjBgV6K/Y/icw6J4WDsmIl6fqGRqOKevRZqnnHSDjphxC898EDkrGu
bzMz62OEGZPbw9z5DFjp0vSY/97UHp6/YUSsoxgclussiZ7lQuv4bFPHeRwMEGZX
AOkZTkPNg5VT7T0PI8gs+e0XyuDkHYePtY2UJI+0D15a+Lv6g/jC5/OAZc29sycE
1RUuhBq0VJPv45z7aEsSnqW3mNJ7DzsjUNySi2MRAo+bkg/6uh+8UpCvl2Cwc/G+
22tBIzTllEoqCF1fRGeQAnaJI2RuX7b48ulhRVsg2I1tLf0M2Fe8+3irOcCMgUXw
q30Qj3MIxA6OgdhZ+ke0Yq2XrdTP3tnUJPVtIJ9qSR/1xD+VP7JM447oMaW004Bo
ceFgz+VO89fUdWdyJu5+QkLkPTrBURA4ZBolyIduGZ+ccAGXMFMXigCOhRXjETW4
nQtwUhEE1e3tYkKKACSZIpovN8K2YvRAQeg5UP92PtXHkWY5utrE5VSGWtbbU18j
/mO58OjuWRuDYi3+8jMgVITIhsMVIrDsQ7JUNqDxtpColNvWzGaMB6sEFpQqYOlB
yhYPWjZuj4vdY2Zsx3KsXXxfACHXIzlO4bwuEu4p+E26y3DvIJugPECraKrCcN+7
ErIG+cLAdLf2Ll9H05pVexmB4U/o4422m1PzDjnYW6O8hoypveACtBo8P3XE5q6r
42Sl0u1t+/BFqsxHwK6aCI0mf/awjyNWYsjKED+HHcxCK7YUgXZQwBt9lIrNspvD
TYCiCl6movWI7DzB08DQsX0JR8t9Cn4vp48YTJb2acgWzYYlihmQWzjeLj/sTswO
e4xz8jHlPLiwE7xNJTi1mLiInbXro1hTVKqNrzLVVjNn/Jx0DG55/FGLMiLZOk4C
1Vd7cGeXkQd3/Ua477yAxXQQ9gyRaMXRTaTFq79xLQGxbXulbiDpRuH816GvN/Al
VPbPyXAYCJIrBppk0hkRrdzjk/eZgypeP+GTLoDt5iuOrSNrAg9xJkInO1qw3SbZ
yEHz1tlWg+wZcEefgdCzzTz7dNAa9qU1o510sNgDp4BCDh2VxMgn13LCxeHbCgcA
2Yxv7kMolUP4BHP84VUICkWufQiEIj2jMOOk2yElEYuyOLyEQWq1w4nKG2d1f+mg
S0xIecyCFAEe9mYTWkUzdhceRmWIRecZlIY8eHOxPfuC4OzwqgzeepAGOFzCiipG
aK9pTtRP/9LKDWb1KcL8NBwrFsO4IUZ05cbPImLPFnZp8gV3mgxLXjmNL1rt/Dcb
aOFWNAyVtO+pA5p4huV1WY7PBCZ70VR2ltS1AR91E4YyKGelsEvOXGKYNTh/Wm8w
w/BM6tzBL7PXWzj9kR0/zVHmNcBUpCWQ3uURqVh4x1As+5mso6YUFcHjcHngIBxo
rb4zntloCgmoXUFv6/OgD5tXVz55mgox5A7W6CpXZ39n6a3UVUjX9aG1RIipJMJG
O1uQ2ZPvjkRhBA/EbJdZTnnxWrQJYwucOYdtHHezc+ibZc0rFPbdmJdOcV+49082
0pcLMcnGqsYF7GuVLeWH0wROtRvPd9HkzOHvUUjVS23jYr1b97puACt58SywF+zr
CzRUi6pmBAbNzr93ferpupj8HL6wkV88H4SARZNdbQMppQrEafNzWvLRgYIPuXtt
5+jaHJtRhISDOVw2oAW9yLuYK76Z/GPFsb47xiTrYDwbd7/aZbwWCthVpyA7swJM
MjISIy/+R6/hCUb8a9WVxk1VL2OqP5SWe8SuEp6kjd1S1p1Tbte7hMA9PMAnA3wy
8VC4FMRhA6N+HAEKbvVVvzU+sUI9+pdXsBw+JkdFt4glc64apNPR851inmDusG4J
MrqlXygxyLFjwWNgXPD2y4Egal6qfHT+CnRl7Wm+ld+viX2p6a+yhB86S8q3jVHl
jFOtSXEamg7DyL0MWgYHggdl/aU3edik6PsJ7pIIZC+IUNXst4B6mWPFn1moNYVd
+6ppeRMgnJBG6wFFvMSxSMrLcJaRuHcb1MofZpX5teT0AvoomRUjbxVW5waHC+UB
JSypekY2gFgkIz8dKc4tb30/Eo0MqRoZVFHgmIx2tvXcVJnE4IK/Ii3S4pOhjtHD
nLGutRHx24/5QXiHjNrDQwsGMr+3JCdF0rKd+em6KaC9rRC6jmFeGJlMKSlTgmgV
RduRC0JtvPNL4J0+Q1UTFhfwk3olYc5iX42Wx28WIgSmwjieKjAkqWSj4DWV2yr9
VpGKH5DKgGATMQP1m2oHtelk12ykjyEdoBYUOtjurbBQT0pkcAmnoQ9ie/SyPNbS
k3uP7kZa/pFV+HwBl1upXgaqTkSGSm3IyUn9heZz/VTLFEjReb/9Twr9mQ92qQQz
ZTtH+nysG3YHlorsgwW+aRee66+Qam0ji+0UGxsMIWpLarSqujvRcDtjG69AFZIG
MLp7e/Rj+n/xuv83LbRO7pcf1kYM1oq8Qa+AmoyI8w4RNsBFPFwm1q8ZwHAufjmz
oQtlqnHd4u2UjRuAxq4fvHuWamN09oagQNZBdWzAdLxnoGVhRrHCYTQxFZDsi6jQ
b6nn54zNVcRbsiicGaZkoLm/yX/5jWdldMsntYgFVn95o065MAfND8ZDcP/6WZDJ
OUc4zxmL7yuOe9SuXZBJVQyDbHOP0k4c5UrsW+FLbUXq83gY5g9kdGSnzr/53i7d
UH4nsg6lK6yM4YbOaUQxpqw343NTilYT+H/M94RgK2OPZcXONepKL4YRuFtRHQFh
qM3F42t9QmOfTa1ejjJ4A0VbCI7svklg8JueNzRXE2nnPEuY5u3hmz1aBgXxPyc2
a5wqtAWQrl94/aug9l8Ku8SgQysjQVbX9V9AWodGfgQOlXXGb+yVysm9XUsYMNIY
F7PS5LZzmGq5wkKtGp/3XZt0XjuTmQX30V5CC9XPE9hRY8l7Lblw9BxRbK3+ebv9
Yo5KqknG7yvxuj2R8QnCsVDJlofXNnXzzdN5eltB7LiFQeh8nKhQAxrUlifcOb1e
TedQ1zqs4NGBOE+zmHnSDSfPlY7F2l6J+O3FvDFIsX5F7U8PF5myAVacGWrlzj5u
l6LPmpBS54vaSLahHY7qsuhJQO7Ww3WtnOqRVwVN8zrwlpQyUkRY/g4g1ppMtFV3
hiXxMb5FUTByppbKCUeEBTOVXj/wJFbN6bjTZZwxpPiJBKNZJmscn32zGpL0b5FR
YynICLzQm7J0jTk1oDy2jtnjYlMZQbjXKTnN87wuceSydSfnE+gOlnrIDi6wHDoA
EqhcGFtW1lc5xz2PtLhG8v65eCR0gRRK9Zmb+uSSTTctZScGYuLRwsneNl5O3EG3
//OL64CdHBbt7PcckYky7wLIAc+NUsbi3ZNykawAgG9hr/32NFCDJov9i8LOS8Qd
vgwFqXgEPXLUI+6Zx5R2azAxzV7mz5LCBYtihYA4lnzuRUK2PmXDx7JcANMOtI85
9YKHuLWcWgd3wheTjAbqNAQXDZoYGdDiarVHk65WqnpM10Actz1yhxaHR4KcGCk/
w4xghPLNESFPu3OaGizZBWwD1BxOQgWsB5ik9jqaCV18RyysBHNU2KSB2ju13Jwj
zFagSf7qggEWvMzaCjvLwyuJyiJkTs8gfROl7+93hqXshN/kCEqOV+6EBplOqKE5
1QU/lHzOce6UBAVO3KTF3wwrjyxbYvKfPO0JpaGrpkxD5fT11lvnaLWf9XqHvk53
gT1vRwxRoCc3J7W71yhE5U1mpuepTZyWxCUZtvER87vfmZGd4vy9Og8bDT0yFSuK
Ilr9tCHJUoJLGuewJ51R1habjURK+vImR4OMeaysq+T4Zlso2xcwqDuLeB4K1gdy
mv7dplipJe406YbYnNExI4popRmlwid4PntsNx9m5U4TUMHUrruVZpQTvqCXMk9Y
zfLRhUoJA+Y73BbJX1lKeva5TpyHyIjBZSt9V9On3+CXgM2lfCh+bleN+7vJBESr
KiLoaNAWuYnwPUU1OtU5L1Po4bcQJOa+GcrgogxbYbpaBVJsTwhd04AJuYtjjTFT
UF3EWQIxPJx35tkXGK19IH6B4XXExTtwwO3uav2l1dqWrLW2yXhOTdxIJX4EIQR1
F2t/N6dEzEwN4ZkzlG8VQZgR8hDDJVH3XKfVzznw6ySO0DVsP3Ugaehh9HMUAr3B
kznhIF8+Pnvm+qE7EQUjZgUOdaexqMw7RwlWSSuTz8rQ4pZnRbw9m6CFsaqNTd2B
I+5ouYDLIMnpRzjkrMq6tGbSysMU8YxnovWMOCs0Nj6GXxLg8aQJPWPlp8fnBXYm
1Z7tpWMHjmBgFWncgunLOOxxTtkw1VozxC8PcD19iji16HELSHbc3+npClAJIZWV
ph3xGjRWq30op4N4fqiVI4ciBb0GAIYdNCCbaEH6Mg3VV7770aCfg1SEyS1BG1sp
74pVTRUtXn/hNScXw/YRjwpikbDcdXONCE5r5Vf7frwBl6/qgTQATcNw1LgEjk8C
XcCQhgYpJ5z+q4Zt+NfAC54bN4dJaycAOrViCOgMd9BjRZyjnCwPrxvz3RP0P3km
jdpMh+Zv4tx1u7M7OKWsrRrGzVr+jrm9/Hjkl/RcDB2TiNkCcLJNKIZub455M8Qs
MZs4LG502amn8F4UXxzX8FLQCTHpWivxrdEigQyCzC6xOD5qyyoKaN+LR7hq8FCM
8byJOybBYGI7nvjt2nkBfnhclBRgd/2YZwjWK2nabqF3tn/qmfm0aVt8Nq88USin
IOmKv5F7UjPNtxMSKVfiV2CVo/D9cLsqofL2cbwQJX+RZLfomua+rTit7eRn75rF
DhrHaKbjCeu07veIhx25ijFxH6mlE6jOSEiGBVJ2gqVfJQOAIZCh6Ah6ytY6U0D5
x7WrrslmqaRBZYAF90LYCcU1l4dNL/X4ktIj5mrLPebcCpXjsKuPAeTwm1hGpkmC
xPeliazhXArokc9vRuUXnndRoFY2853hqB2y8Fx6CRfwzlnt0rV4wU2bdggSpaHO
a+6KLSwcKTjIVvpVrhSWMOZ2bKsYbXbbTlV2kdshTUj63nTC4ee0t0eZiqQomG5g
+IyIZ82E+lqKe+WdknZnP2TH+zeKQBw2w4pkcN6VAHRqGj2H+nJKsZquh98kWSlR
HidPFHAipep5vKzF3tnh2bK64MsEL3lxtSWusg/grUEZjCyhAhRpVgNoGeaHKfrX
dWbZCT1wcBMv+DVHJddDJUTXKp3SkIZ8fysCIrZXfBruvjSRRERR1z1qv3YYzjni
LIaumjBtOikgUCL19YxnWNHIGdHN2ZVVBn2E6bAGGrdGMikqQrxrcCrhsZJBFP26
5x4MwcRrt/KuozYezVaQnjPm0mm9CgpV4TDTXjvn4Bq/toDtg9EKduLAcTZXoDDG
GOF936kmRH6etP4YtA3otBRx/+HmsOs/z0d2qAV1Gxa/8s5OSZQYMMZU1ZRiFTPi
dQtVOoJy3RPlSyNTRGvW/PpFya4UOMttOyvFgf70Wq0RR5xLz/TF1KnLAr4p0TMZ
h8VL/zr6xkLrsu6z7jcB/Jk05d7ptI3Dlq7gTcxCvwsy5A5soOGMQlS0REsqV/rk
OJr1Qhg96SfAa5KHY7bSvvw6LvZdMz76GR7lt1lEudUuSmXqeT8K3YwHPlYo/0jp
3fmBtzR6dxnzkfBWJR9+EhxjrqHEn1cUo3+Kix2YQ6z42u7MaOuuAmz7eu2d2Q85
FOVAmTX/eH4xXGpBSVwT7VRYBWP2mUb2RP2kBSXLy/X5MA9P4to0fnYXUSJasOnw
8aL5/jNeeBCrfqeOTDevTzGfwf7N15+WdbQ12zST8dxsUy4txJx+mjSGQapLXviK
HeFK/CVuSh9+isp55OVWL3TK58B/4llqllWH0l0TYiqVYbOUGvpN6r8IHH4M+Ap9
17xSerays/WkjKU1Xwbv7xbgLIj7AWVD30eTw+c6o99oZ42BuOsjalTnQUmtdI+P
8rh5YScet5YcVjFYr+nal6smoPhOEZrYFtoX/s3hOvEAdkj/EE7nhPNIWN4RWgze
sFvWLTE4mxT+d+/xOFhYCd6hn56sM0+y5574V8cuKkt5+Y2biCgVpCLqBD1P9Z8+
7rjZ6xFT4hY/PQlJUHC1abS5zN5GDlFmXm64/THBZeC6KFNeXM1POVZoxEMzKJcD
eZVaBPMyQbf+/baRrQL9eAAYBYjaIzsXQo4KRdZ76hVcq3XjAv+c/UW8P34aW1nN
4pvVBjRQjPvI1eFNrmxsDS/7tyblQ+xu1+JXHqwOD+/WCjjSPxXi/m4WPLDIDfRc
u8I2ktEpZY2FRs+1ktqzkK1KjcPKy+UfVUWXH8gSYhlLIwDhr4BT00Sw63oBEaFr
a4O2EMqOEwa8ViT3RG/7OlGwjl1xBUNN17d+UFHHXFOmLY2I1CQi/PDRrwIlv3Yj
RAgFHO4EBImNabXo9xs7L1b5Paj0tmo+kCCKz2pFBjKTuIfb9t4t9zhuTXJfWXIl
Mo6g4occB54oEDDXzfsQ6cEfXFUtAyCGZ71NrLfbg5vim1Bbgvb/wQM8xkgkYswR
+A1lMoXJjwemDP77pQg9bz2/XjK7mYj/UR7Wp1FbtZJFq33AZpCD/Nud9z4z+vyd
wGq5IhHWqYYrEQE++QzPTRXSpcIH6mepgjDog00VKM0ZNFHYsH4Isckm9qwoykye
X8muE+nw4mQtVsLnSM45tmyHNwiK2ukYaYdsNjJEljYWjCQZKFkIaDR0patNYqAC
W4o533v8/oSQfyS/FITisiezzROg8ndhQp3ak1K1fOTOmwquXS4/2cozPDj/azT/
2NR50qsuy9KgfRvtFbFBuSIJmqYI3YaYbkR/lxkDM878/EkrGdl/xh2c0q5ToVQT
y2WniZIy1FofRf+qGbKtwIOsibhB3/9SpBBNiow2KJQfzF6orBBmPvp1i0V2+N9Z
ubojrChoS7j9SxwjxM7PCBhhhxOEE/bTfRVg9lJ3egEQ4VI5MpmvARjw9eTyD6xJ
7ipuC1RRdD6Vvci89IRw/QRzlP+T+pm13HHa4hRebcNAXc+Zj96AmsFO3D97S7ZJ
RlVYhKKl5NVjdL3v5fRJrc0V2NWuGovVqqyEq8MyFFLCaBh2QFvnYsweRxx1g5bC
4+YM0JJDG2zahTVRJ/xDqaW0ACRmnHnGGo9sNR0c/j/TiiUH++fuipFtlW0jFElQ
pRRvlsnorrVyl4kUmL9r13g5YeNr3JAka8VWhAWcnC8cA6//mD+0K5KnK9xxGnmU
sdc0+st7gW5jBvKjffTHqcRn1LYJa3EoL7IV2RglaId+sE5YwROc/r1Jd7vnYekg
FfhhA1cQt8gBp/62mSHiQ77ygUSGuK1YEG4N1WGueLdLa8LtjjgUk5yYx27mLrnQ
KHn8k21zFi/zeKdlBbgtRVj4eTfwAdCTzpDKdSDgR777I7LrbKllOcsMfzilUbI1
fKTC5GOTVlOtMBmyJ3hLVXFvJSNd0TYIX6XkK3nWJSoVhOt6PRs+rE8AZbHWzjBR
7HwqIjD821mDDYbyzMiSWNLv2Cet7+jlRyhXhbsZWZc+ZvXnLH+AHLsillXbZVLI
aLDeXlqV+PEbdk7toYb/j1ehgzlVg+5wAuRRWHoQB8/j/XMjQKnY6IY44nQVK+ak
g+eUGuZBR2RLuQe+bLrtHhlOYUyOzQsVT8dPvXAsw1sRI7/cWvnS/m0dAetp/PEs
bI/0c5dMlKZdPNuz8y4FAp33FjFfGh1T8HtpBHfuwdelsXCjn/symk5kgHqiSSB4
nb3Y6Vv4Bpc2kkBr4RBoPfDk25HwlkBy35vTFmyuocXYZjjB5i0CDfDYpqgcLI5Q
fuASnbD20vu0qLvB4vI3q/Ht44KjhmIsTPjq1AY4QY0WLwFcu/1KRXHMxnIkvSmI
ybqPgP1Tucx9VrhTmyPrXQt3ryzehLFi1QhmUiY3E/gNfw08ALRovUij9UTWTqsm
QtNoe/Fl31/5pajd6f3uEtSuSNJkQKK32luMzBP8hF2I/VTTk86RjqBmGbB8vgAe
Ktd5ZIMxbGbeB0sjlZz4w6yUJFuAZzgDdJ4DT9nohXbOj1+NWY/A2tdDsZI7W5Gf
tMQ6kvT4fQItvuOnAjXH4vMADeWmssSjGa2Fo1EDuV5jDleOA+yUeZWGhnNeLUie
g4ObefP1x0KJdC5PxFzcLfzvK1FSLGwAFWEgaVr0FXHU1hTD3XjMD8tq9oilYJyr
u8viL1OfadRl001aztuGsRAh3jGGlKXzOzLCoYeWB/BNaEIHE6fxmf2rQ19ur2Fo
gvevKUxl37iWiWR/sRK7bLKTlNTWcAoN+EP4GMruxqFwIEs3heBHJLDgEIPd9vmr
v06Krn3Il97hpBdiU2a3JeSHbQ+yQYbSBLg6GqbgBR/Z+3S9g0dvbDu8qCdukTg1
qw+tp/BgSQAJL+SuLcTEe1NFo9bqJEjlGXadpEXcDemvICbcdxxyjEztlssMIQnM
lVlj1QKpRaLoVNPjU7SKY1z2ST74dJ+zYSRtnspo9smcsePTFNyJpCuOb74H+tn3
CiXoK3zCvSR6aXojyb5t+YsPdI/N6EomCK8CwLgT1PItpmqHLEwtgoOg4szDpmx/
nrf4NFeCYNVGWPveM8MwYDmiAjCtDmncM1T7QmEX8vhLw2aPr+YnLJfcM4ZQdAna
ki5OCs6JWrrwLxNzpmcMbwv3b4Nl1XChimH0al/G5V8lq6IMHxmq4qaFdTIbIy8p
JQA5HYFcBC6IH8+fl4P+uMN4klbx99oQlLJdM9JuZdRfIqH9teteCcHtiQUKMGTl
bD1F+f3dzmgkMBxA5I9CqKCTkHYoQm8MhdsjsSG9Ja2q8f7k4fDZV4MU63KjDX+B
5Z3kuoyPjxOdmJ8Pr4DA+G2oBvzpBbYKBY1M+HQudrihzZKDZePm8KUmJsoJKmjU
/V5MU06waIX7AjQ2gQ8gJPVCQp6Zykb/OwJCWx57EWf8fo5ZHogZEX3wP+s6BuX+
rYnrOjYZAc6qWjnErJbtmvCfsd/D/zWXv39Tmt5tOWJw5Ot9seYgFjp1HgHJrmgr
KW5jSic0/SXb9VNffnOQzLbSEy1uWa1ayCSF5SFpSBipqi0uV5Ph6OZdwsWABDCa
D/kaGPRZknQ35EDaI4o7ManFq0axOmnHBcRIRoEBr6g0loZEiLvZVTQEcoUGRt5o
UnqwWvAXBWo7In8B11Cp/883TWOjuIB5eRG0I7QUaj1RYmib9yfISafH+F1abxAl
w+wOwoMzDtYsV05cE+h9bOKZSqbGrjlnOPMohbYc16ayALutiKYV8AkzGZA/m/DU
h3nmr8xLevz09x3sS4e+UyodOtEwBHxyOcrAzmnw4Ua1SuOnhh56O5uO1ByTFNkK
etHGSFbCgsCmx3uJ77t7GJXG2VrsEtscrYG9kY5BjjzKL9X6PPHrEfPwH249Fk+z
wFdgtAPPUj0vnAP4UPs86UKhZy9XDiSdggeLe6c+7n/E4NynunEnoyda4F14FQKs
Kg2oR3FEoaXtNthmuDXxz+IbsZoeNtWmvl/WxoQKPGbJQoj4xm58GSkN+zIxHK5M
y9SBT4AUCbHRTp1na2B1IpxMNpKhm0Q6MpD6rpJFKkwM3DjZuMMw99uPaneApB2B
c/7WV8fHH4XntsJ/bT2MNfrKD2fNxGf1RBDhT7hYJIRnNSJDosjhgm9dtoahkV/z
fLZP+UcXc2S2X92sUyxz99Hmx3+xW/amCoSuXc9So9U0gTCGmrDwA9S12fH8vr/8
/3ZG4wewD9nT2glzQa4iTZMxDhHAh1VZfKD+0z+9Kd0dlvRAW80kVj2F3NMtkg6H
VfUCitoGpbPu0lcqKr4IlXdPlG2mzLPAaLse4UjJm+Wt3Zb/Mmouiz8aalnomSvb
LTsDIaGGs3fD6+AYQCvkpCXRTZx6LwrCQX0knWwGvGtYVJBRJ/fSdfgbzk0MIax2
o5wWfeJkucrbGskIB5zl2w5Gy5p8h6OQHF077C1SkfGTBy8kO06WOBZFepW5/vSM
1bYDdf2FH5mEaHb8v7uckDEmrOfibWsurxgWLsBi6lyWXVxqeXMNiQCrec80HAu6
6i7SC/GVo0pCHTzUV/1JZiGW4Lh0BdTmArAwdMBKr2Xbe4vPh8GWb6BLJn+Kvixr
7boXMf2o2mpIyJINYK4HSWbjsdkkSGYfTqqDzmmbs9w/Xfj0MreV3awE1o2afnFj
1MtsZ92lCPRa4Pcr127wogSLfZUfY/0zPghZGWIAtMJD5+NosqxKRtdXSrr+1NFv
xSEO9l1rSKkdP7TmVwp5mtQbk8Sc/fw2vxDp/6wXhUj+EboHkE5Ky89f22A6HTF4
Q/GRxHnOOLJdSNhOkr0+eGhwla6M4esNbQfA8hTU/GnPv0cvSqz+N8pKn2IfTd23
U1XeALOf6S2MNLsaY2/bSxvPbyHTtzk+UBNgFZ0BHZ1UD9hsTzLXD9IJGpWg8I7X
KiK9LKlSVmOD1+vX7l3h27wwkvS6XruoUURefn/kTTLYNzAcDn18PfnupcoRV5nK
LLM8VZm7Xoet3IsAdIVKFAH3aUM63/lT2frWnAoKkA0kh3DlMhA8saDDfbjlK5yb
B0QJYnmXGt3I0cbuMHw2rPVqKE3hcQw5fzSPDBpSIloR2UGjzB+ul2brWnDwhXe4
92pnvCL/78pwcQJsBlL4ZF48d8M79iF6GNMiVB47kkiYcY7MDlt6pni/5aw9L3wY
6aY6+X+6GFG4n+p0K9ySdpnaFxiE+tVsnoUIVvfRci6+54tXLeFYwlYe1fYwn5Tr
K7w2dNRvP0Nbg/8KcmYp9Se0SVCIKvyODhsJ3My8q0UzM2fGvGLjdJH1FBU6nc2G
oZI+hTzPhiWVtTTZD1dEBDefTQ3TwdPgMB8AHMcEdW1Deu9DCGV+h3Iz9XIMw0U2
+fkQ8wI+4pvPkrDomYLA5Ik4KcmWSvfhQ26uYDjqasmJ9fc/k38lHjsyNqrHAEg/
MqaBmqlK26tzNzYo8QtMw602udH/XdQc0kuYbhtEqwGub73oNFjo+djCkCM2NID/
JK0wlLzCCOTF4qsiK5xK4/qjl0OiBi3GLfgFJUPZHl2SxGMEXd/FYQ2KgNRvHOnM
12ly5bTTsBjkMZClxGfHXlnlTFxbN+Bew0+5/6fTD0Q4mOd+jeXEuucUIK6mQynn
4AyI0kqU08EqCLrmlW+lBSIDXHYfGwSEO7r4wg4enj5/wfCpO2G1Eq+QjkBA0hLO
qPeAKhhwqat5/gDzJHUzpjc2S1GY6ywWCxiWr7nWZgyZ+hyb7MFjiP8NmEXHu42f
Dc+wj6xtF0AEqVRihPb27r3nU4j7GN2cebr75MeicxwQQtRllPzOT79SGWBszudK
az3HNEd0DvjOLQUFXzj6Luzs2HgSC0wAXRbHQagwSo+Hlp37nxqkN9ysjgpYleeT
E8HuLLpDtE49lCSsjSqVUEbpVfHdJUN7IxmNL4Z/fhZT4JtGrmTDuQqtRYr0IWZh
mfUGUqkZM0wjxlQV0fHefEFs5RxINQ9dLEtZXRKXPvqIq60FE7KY/+3fEcKT16C5
NLYocd0k7MYhhheu8ArfDbyrRQzwC7s+g3wK44h6NMgM9sdrjolPqWj7bKLhivzt
nxl/iPg31sbzlw8olLuyBpWEv5edqsa89r9DpA+pahW553gHiqLnNiCfWN6fQpxn
LiktRtktVqkJYjaAQOqaQ9QL+mMBxI3sRJYnAo4wRb3OuILv25BpUg2zWeLrvzkU
L+w+R4KIB9natmTxN0sZn8GTuWPiB3qnOyZ564E3uuKLMAxYEE+DlRNVYQ36AmAE
/W6snygp6VxkbpqtNmrvWQivrEn2JkirirKPd9ZqUX3eKvoqTySafo/AAfBozPC0
/nJI7A2g2tMJ9a9wlSSkS+1qxRhgmwU30rnrhegxW7MHXqv0WawIuhbeIMPvptrv
xu3K/B9J05Z1TUGoxLdha9O4NzJpt5dZTBwWLZP5z+pO8MU9BUx1AoyK/dwIYHLo
AFuB6rHbxMOjRKtXVsfxaa7L/nwGLEpQIJIUKvgn9F3DNz8+fC1fWyUpn0hhOrOO
na7o27S6p1tPL5T+sn1RIKLernASe1oRhzkEdDdxCUbViQlVf/F7SUG9shvjNFDV
Nqql9bt3+AosMb3mn0HMiP0jLgbKHMKIYIB1xK0v2IuDPvyqMnSi2jTiR6s62wwO
wMl5Bx4f7923L4IlzNrcrSaAwshxmBXhhJ0SUJuAYddk8y2jISlhhi3+MSsWxQ4T
ZEFXdG6Rs6oIYBh/f7kxvgnRA943Wzd75dpoRmTEBnmCfNpb95muJm5+8+M7V/SW
pYSMSwQDFSyMoij98EIDonb7z6KWickITMNtA1jLdUETbm0sd4Y41m8LSWtbqnB7
s1ayVC0QQEAF7szvAKlEkdMiMNoYEB8uaIy4lommMUpjX77TOR3c95kkKCY3kN/S
qqJcvqKuY9MK4Zepl2jOWoKrCjj/s8VsZ5YqNV2ApRrJDFbwB0WiiqDcdo9tz/ZI
73DkV8vnz0zrYX0buya6Bp09m8Eg2rCcnESTHvHgn/gk1NHqaejhlRrw9lsF0qdb
TqBcQes3FykkMCsZlHceb9YD6Gt5UYvvSQw9w3czxrJFgIft6Plnm7QgqrdwclX3
HSFuUyuHvV2K5Af10b5BMlI3GjyfNpJAIZl/voGvQ4P9LMzk0SLchNfdhkTXse/z
LkZ43f28/LMoYAlYJwhZVxGKrt+BrOmhI8TFEH7SoQo8sxyPTNj7Lk0Rd+WEor/N
e/txHa4P6f6rBVG/P5WbmjVqaMNTq2OfRyPjfK9bkApQb1P4dGdVwMKFeyNkw3ht
qB2esNDEuCAwyL1GZ0I2RRZWPcioSFbO68IctIzDI5/PaADebsGzeWwzp4uc6BgI
zI2er8/9EwTitDpbJWCRgn7vx40oWmCQxyFeg07Tw1rxwM+0U6nccdRir+UMBFVj
jXxC7S+K757w+GeOZBMivRB2K4B1kfnRr4IQAuDaSly2Pvvpb4Lwt4bwMBJD6ISG
e5tcCm8yIp7Y8Xyp14n5j9FwDV3vaHcGSA1sNuHAo/Ds/DoWzb/igKbLL9Xz2MgA
RuoTQmq15zd+raMGZnx9hFCszpEi4mDqEhoqal2zt3oAdFeiyNJAKI51Rl7oYD+3
Z3AV8PrMqwkci+03fyUcvHCWlYLoFn7DwqMRBnpVpsFkraO9CsnCEoj7DEUHhMUT
pmZU1I8NK7atkjuxQtDNjgqgvpmEjmIrDla4mACWNQfLxvaUBqqNVg4MqBiWYx9o
yzNcdiYG5ji8eBXGG4GwQP7eDQ+kJryReNDw+kFAhi2r3Vc3eQKA6srEfUMmRz6c
cuyzOGT1hx48mHNM5NFev8kuZ4e5ktCc6knPSLysYKF4S2EfNo3Fdbdv6hiBr/5N
/7hdyinJM687uan2EtnlUOelBLGOuLc7G8vmUXSa47p+aZJEVpufH+ZQFhfnsN7j
eXsp6TfpmYenAaxymrQCgTq+1UFQFJ+0rdvdFTWzq1LSIrksLMqiby1n+fsKZ7cl
bfzE4TE4u4JXZIbr4Ztm1GWlrvetmvOf5OsowW7wxCjIJJiKjBo0pZsMk7UTCMVe
arzGxl3w3qf3yA7nkttxUQ+i1uhs7R/g5rQ7K0yh5cvWZuh62gmPnyheCi0v5YG8
g1iaOdCf93NES07u8ydE5k1h+FPRVonuziiq/7O6u27KAzm6lODa5AbLXmERIjRc
FjTCKXggKEl7+UaJwxb0a2gWqcjEwIhsXm6v9/5bTTcBs1RyV1R/G176yWi8U0Hn
epl2MKXyUMYuAv9+56YORn2r2BQJyYFrLrK7K5AekZ+q0HFRkshTSADCvnaaYaug
Pn0IjiMOm6jiPJUOaWpOI0IcmZBfcOAvQyvHX0/5xMfqkJTlJ4ykSL1wFC8h5b/o
SJDDjLhda7CEbls85D/MO5FNIWWNlH6QJjs1SFEGNt5Iw8lN2Zcq0sgfJk7OhaRL
4bkqB7CEvOj1siSckr98Oe84t+NVUn9q8eJhNkgTzE7j1EBbxjqNoxjQGDGop8Zo
c+oQIuSC1Leax/CGn8ohTpsg9vzloeDF4CxkvbZniKEJ5z+UAB0ZudtyktG64Qbo
hFqYf+Cw1cYueYOmewkMoqN+5ZI+petFjUYSXuUB7ovWIDhxcWV07LMwL31BEDvj
gE5OvvduC/L4zOQIDWCoIx3/GbVI1KY76260mYBvQ4ONKTqDlRfQ++ham2KN5dIN
LdCYUSPMJJghGD4TP+CLh6eMgziLkDjD9QE7u4Mc0+RkdKhtKvJYVva+/7rSTzBO
QWysnWtTl4c8b1P1zJRuQyrUmhg/auJozp5bUm0MCEaVjyNkBq9QwdWqZ5H9Ldl7
eXTp6CH+EpBDLaabFSZXV31Eb97PWYitqsgSQB+f+/3xjTCtKj9CrpPSbmu+Nt7u
8sCACj7oLhXmDd93Dc9kLc5P645JCdP/4izwc+rsbY6V1TGrR58l3Q2zP9RfXIJT
uDcpcznF4c25brP+RkcY/Ks3uHTKrST8KRdFOSNzJRP1blKNgV1uG24izOFAnYB6
JaVzAsPT8K/Pept4RpmfoDjyqTpZMsdM0pgMuqmjGGLsyHkO49XJzewwg0OibAEd
AP4k1p8Gu8lQWlbKjf+m+JJXv7DdBf15lQ9IA5qfK9V8IgMu3rJ0OditqL7lvFWi
kwAJD/3FEMpx5Hb+tM/K82R+aL4N9rVB2Qm6Mhp+40Dy+znYZNaEyU7OGJPZps1q
XBidczvURHoSOX34vFD+kg==
`pragma protect end_protected
