`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mB3ZYvbmQ6LYDmHIu6S7J0C+pkJl+UVK0BztZ0/Yx8PXUvgK/csdmw2Q3SOwM6qT
ztzOx4C4fPDsV3Yvo+NuqK7WtbYyy4BvGATS9n2hai9cyB4xBXXCPuuKYFX3MEy1
z0mTWl2qWzdOpIs6j7OFotJz7RJ9D0+Ki2pdOksuBMs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34432)
i2iR2UH6549PGfCYv/GN2A5h/fF1jsi++VHeFQqHviGMvoJnwq3lCZOlfrou1k0d
DUHMNvN91fr93uwQicxxTXhmpXQJA9lh1D6tyes90hLPt6krMdUmyRx596P2FzUr
lwFILImJn3js0eITTQtdarYVhM6lz0LgOmk+ZGmgOv9UGf7x1PEqihYqFOXCVn3q
pCVrVMaYHz9FKG2ps7cEUYrLjh1EY61EQsU4irLNkK8lGhkoBaIWaa0/NekAbeiI
JkhZyZEre27kzQs84zBDrFh5a0KatFJQBZaRtxPdkmcP6JVo6a6EVpK1A68JOWhK
PXUzohCo7QBYLnc8/pQYgO8PqSZ5KRI5wF/3lggaiqxjD8qM9KHTJPYzC/iCQdFn
6daYiNwMG6LdA2x5OlPSXF5uDiiJwPKkqDXUrb2OkmJ3wtU/e+FOCWMDPz9aXqwC
UfURzEu+XYcsCE+UMaC7eF+sTmUdA/VEPawu0cODHjci6NLLL+fL7575SzKjDfxz
ET3iu1RhU/P6La6JypTkhk0BCxx09dQYATNlFzSxFWk7JQ4MVoHDEO5gqw/oiIUq
6O16/UTCrKRHMaDIiJt4AGs5P1xrTMXPRPxE4uy+zp49cXBpfRAFGz0gL1v2c5zR
PlWfrC9j+Xq6hx7ZxPc+xs+ebdUVt3n3CmJGJbQzlLjaMZ9DkQHT34iATl0fOEau
WoEro6cqnerxz8iaMJRZ+BTr0sPOYFZRvzuVN0Tb7S0+fP6I8PswePyWdwBuK0mP
GnS1g0URrz48dyaVISCo9kHiGRfn3tV3yXFa0S6iKJD861qYliudd0kMrvYDGWIj
KDWHw07Ev2kFZ+tRVSHen0omFNplM/yt5/gpofA2+vqdmw/GSPoM4IsXtnc04mE9
ANEH9fLheHFVxE+ZIk4bDWqTUMy45FBX4dJZWUJkmO1dfRoC9sXuGKE9GvKmu/S7
gwGrtsBrW+Kkh3sZqrri0wcqoUpNRjlG+9G66TbRhyCEk2TKDu3/3MCfW81ib31b
gBt/oDjwc/ycMdBmhdwtItsYJQuYxKW8xCPS2aZ/naEThtgCU1Kjpd+4lEd3f75w
ZWj0aF00vcwWrOqFd2C3HLruB+YutcfuYV4I6jd75s5VKy+psAvfQWemZFlligKk
7UVD23BXgL/zXkN0bONfPfxAucJUL57QDrKC/wn1UE+HcaDfmXgrvz7t7eGtFeMU
IEutRudJyhTPrbr0HzTB47A7L7VpcEUdGVFiXN/IHkH1lHfoD9E7kT/3g2JltBPn
XDwXxapXk2L5uY6KxS6e5la+icD54Mri6gabr6wALsCVqxE16HNqpYSHT+SL6Yz+
hkdOTEAY4AkQhBDPuHHJhh5TiAQ/fRZx+boLHeXvT+DvLzoRSMoAMkvBKuttvz89
E2pUGg0uHY4hqQunMl3kor1/zK2G/WTCdnM/JpFXvMVDhbIs9MbB70G70B7Pbnb1
UzZZwHfaGm67d8X6597jMCLZJzFgsGwYy6eA4vuHVp8/M4To68DFvqyv5Gh0wU1G
vXGVcsSDZFwZktMt1e0lzdwWW859a6w4JSLIQVHriU0FdP6NspPGne7BD5YAqNYT
xJMPVs+qmSOsMTYplqLpC1zHcjxZ5VUzLuDmD06TWngC6Y4pQupxUG2Gh0gnFYoP
enbpe00AMnk3z/lmvYyvvEZELrTdW+eM0SCJJLowc836HHv5uNc/kXjlf8Cb1GH9
WY5WQ9of+Ci2LrdYaUXCQU0+mnytn5b8SEdgzOZf7D/aYo0X7OYWCdftyizv0jaJ
UCrbfvYT9LK/8tetDxOxHWR/faF+WheqWJdsVtJAKIuypGWa/BBS69FTQaJrsiVx
iksjVQ6J6vt9pX2HqT4CNIeOu/zoNBaTJptDxn8Ht3Jekp691OyWmcaeCp0tZ/4W
std7sfqx1o66CQoLRzwoVJ/jQ5Fia/ge9pQ+Mr40+O2lbKIpo908Fc2so0XEn9F2
WDLNfmndFgiUmNfoHIA/MoE6E5etybX6KEF5+6Q/iAnEmSLL+vjYHQ7rd5AIMqHx
4TBbBTTK0c+i/k9h6342GardJO90ToDeef/Gr+8G6Jixxj3rRghvqDg4Dq/MlWOn
7I3QRdQFk8DvB92Vz3twEC0bkbrbFtRYpR5ubTbeS4MMmqIJtnzZ+17D4w2WBrMh
s0xiBjRoHka3PTd7fR6NHzxwffg55NdZdoe0nLxuo9avObLQrZURA5onfe2CzPUQ
LgeC8O/aajXzM/Fultd7fOV+jgR58z7JdSbKhpLxY4bOzbema8GDpLxcbcMBgQ+F
9liAqkro+BIVwccIaZ1AgaQtEv4n85tOt406qoqv+pLr91YYjE41Sz4QaaRd9tB6
ZlL+hRdgdDghdRH0D3pSwfoE3E6KYAtzfBeYO8NgNBXodghKFDplbx929GuR2wWV
+VZeRHi7rEPiNY9SQRy2qW4syWtgp4ivV2Jay0A0dhhrzeR1Y+84VxJfr6OaE6pz
qkr45DDuCbqSFpzpqbJMSt000QOPQHVCScQQ5QYfPciVTyE6yjlqr5PeS5gJMDyd
de9CJ/VwlPU8qMUNCcGQ77MGCAZTONDs9X1Um66DaRMMjY1h2B/pfMBbQI9+8o1i
i5TjthPNJFe1xQ8Hh3m5P55yQ+YmCsO8CdOb/USI/zkYZyAzSGG7mZMdo8UXNcZg
uMDmoxax1M82ftIdAGDM0m6UilyE47jnseQsFu49zzFRCcfvWeaRRObLaKAZp+va
WgFQHufhp7l3kFa/mhu4i5tBWnRc05oIMubiyGsii7GcOcwo+pB93UG8JIHyipt7
LZQeIBS9jL291a/aKLDzEG+xyRhfT6d1Do4iYAmNKmQLolD5bzUQ2j0WwOSmBZca
rEHJ1uhKOhNp4KMNnqRd4phDz7sj7JxVhqWW10XL+e46I3CkdhHT4m28H4c9ta0u
/zJy5sxpIzok8NZSUk590HvXbtPX/gATW7ug0Kp3Dhjl7WMH5wkxcf5Fp1Du1MPV
Ok1oqVPWk6nyWtES3criNuWG2IukshDjNO9xz50KYb4W3Za6zBt+Ps4FA/CFEid5
/tepgFcshfJQmJz4ckj8OZDcnoqQxDNt375Gqy+8RF629/xpptxbagM66YoTmYil
lxRr3Dk1P80DKwfbbOztG3bf6IEvnCbx6uWxAVD9H8iZITD6vzMjmfaaYSZsgfX9
ncivE8Te6S8Iys+v731xhimQrnUMZpF3rNIVW/Nh0rGQtsYGcDD4V+L/31Qa+UbR
Glu4wbYAT+BhTOlmbIEJyclAVjU+wuuaSy71lnbqqApGUIlOoVa3t/Iv8g+mp6+Y
YjtfY7N7DrkGcOAdltMPSA9iihXUzPRaUxbBLdOQLc3gs51LcNf4iVL/2cFC04EP
+gMovRf3zeYGf1xb0FyePWB+rwWRy6xniwvlNCJ3MCxiIKiN0KfpFdcUkhzLmjSu
y96k3M1IjARVAXrSPPtsYYzQU1Z6egj/V8Rwxx/NA8BClCIfddqcHypPaTQn8avD
DVvkbHffVXeHFNnvdEV1wgbXBfPVYZclW5j6eqvZNoJZ5LOU6tqfToO0KD3irM4G
30rPF4kgf1R5UHm3Gxnm0Ae+vi0cHjvtOF3FUayq+3F1cL3SSEbfaZXDXUS6M0Ag
kthv9pEzRdwwiK0tDpdWJQSqcTncovopJWkDKn893IoeQdhPUgqs32WoKGjHyxvz
Zrv//XgG6Ghe4JbIGTLLon9xj7VJ2Wq6uH0q/91xN7p1a2wJs0yYXhI5RYjtTtYH
SO1h1PJdo+125tyJzrBEdH1GVEpKXD2Sit5M6shGPYpf4pPaxd6Z7wT8M7UHBRqF
cYVahsa1OuS5zDUULc2iqWQcfhpet/aOt//dNwtUhq2JDTcHoqGMiknamCKgS/JR
6q/kHc+QkWIbQcFNpDWXyZKi3t43ltSxzlQEP3VWTrRoD15bBA9b9W88NX9Lv6Dl
/R7+KWgV0/RP9BfOr2Jpevo6VMsfGzoEcqKVF9dsng7Sg78GReVRH6Lr6Skva3I3
zpexpUKtCQRMSTcTjlbs7EXlNwzTXHDhPzdLBduqltyByEH+2Ed5AU/xGkbSJTHz
GzJn0rDm6emFyviTticmdPGvs7siw6CSCdwzCEh17I02rL6E0DNrt1FlGg7xxyvL
5lb19Lfbz4Oe8Z23wNpbdMGrXCr6tzxrD2j8+IKeQw9q+XMpIC9uxo+95I2tjQL3
7OJtdiF5txS/wCFzplLu/VHppU0Mdxbq2e+MRR6btdxjK55vpeQj23R6CKzobr7u
nDBrqzSHAtkTy3XspAeUv/EroepJXaflzbpfdg+JY1gxzlithhXzRG9c8EukDJHn
lMxYv0FV3G8HddFqZXi+qlcwdHTsgMQ2i4YX3CHKo9055VMyEdHd9/6rw7dQMit5
hQL0cIz81ZHBPiC5dz8qL7BoGMiB5HB8FxfTo+bx+TaFHasNQTBv8IKrvBDgRcmY
Azr6mJVT9jpAE3TcKz6y3z5AhxUy8NinI+r7hqxlIvGH7ptcMr9NcN2KwfpotSNi
usssc6vDZQseiR1qCwu+dFEFmeqoakQN8+ze1of/kZSV0gBWWBcvtOokkoJZiy9T
jIZVEg9RU3DaRbUNE6rDZCfJ2jaa+ueg+nOfP4MYFXySjkcSc5cgqYCBvXFbHu4e
/iNKWdKgM/2c9V8YYcwzXZSGSKvGwPWElXENMHuqsNshURWDefP2UHOD2ZEsdSMu
BhIHnpdmK3vIEGQPLeb/m4/DqIDcpWyVACfzp4BO4MkH8Ay+NFm3vKqLW4hwNQi7
OcYxgitGH3B/suAHNx2e+eMH8ny996Hm6C9l9r4QdiLEX/CB1yr04nua48a7tciR
JQnwIERR5AZai4Uo5Vf/WpsZ7PLZUiiPKe5xeS0mAgkHR0mkl0CyrsbUQh9cM/JP
9ir6uwTa2q07V94gpGPFUI8Q6hGMwmJm46UOLQHBXGTTNtnAHBafjVXQMakq5lrN
4HQk9FUVZUTbIGP5/XRwjvTarcGZ2xkRhH4WjC0ZxYeMehfpFkdPxL/uQeUkZqdo
wi3G659wirmUZPvRlcQl6s9w98HvLobOEJevrb5wFnJqtZBqcxqcA0BhXmTheA+n
5RllktOeZ7o+k9cvgD3wELZCMaK/zbrt9dvmSdVtIuiBKkkesIf0s+l+PLGXZuej
ocOnuHbbwDCmxi/XaLKPpL+b9kIX6L+9ML68rEROaYb7ct67SJ/xwt8k55FGOWeK
vW5Tjw9HczVPJf5TXjdhG2CNJgfhBs5mHX1bp/BHew/R/82J15r1cKGuONT7QWdA
N/q/cVXmo4qq0jsoeAg8eBfXUEhM7sP4fYxi08d99eDOkCtAVNKAtrlRUUXcCa48
hyCNMK269nET/R6c4gUAYimzaEm9ixRbHGzKpUPdNN1iAxpqb2HK1B3kgqb6zN6f
+7h0wth0M0aazYxUGUBDpZ53tn3F6cMKqT0jMuUh5l2xOdnnEtSyuBmsV/XMVRTR
cqO+ufHC9eslQRc5HH7mTW/Otfh/nVXjFROdlIx0DwRU2eLpeFpHirwKcikKYxFC
ya4ZGcj2p4tSkG1g7kbnfXuZJXw8zDZBAxHX1AJMmEMthI0XL0kKLyKci08FSYDg
s7/Fx1ghlLoiSL5apRmtgeUljB33nTeG41ojbJgrs8fVEdDF0g/McA0ZhQ9lD4CQ
Fl6xnt1AQPhPdKqOqSgVet1vmzm/gxugR1/1zBPnAzWeo/2pL7KcLbq6hx+rQ3yu
W7thr6w5/YdWj5bcZDRlAT9EUB9NGIwMVkNcjvpiTCcYeWTHqI77vAM+XUQrXz9S
b3o64lawgZbf0tlCvPCy8nicw8rApGpLSsQoZXtnzMOfuWHX0mcj9Nl8A3l4dfqG
/O5KRFJOpbX2ERP7wVWaq7Mkz8pH07sJn/mS1xW+aBrVXMLwYpPUq5kmL1A8ZTHa
kE/o/Mkq9K6Pkyva8Atlam75U2elYUcY+8Qg7RcX2+T/WHdolSh8qBrifj+2tN46
nzXjUNj13TndPtnqzeKIF1bEpF4iarurAhISupHiohwQ2JOFn3x2t+mWQx6iQcXM
o2BswzxEgStRydpEKvxPa1SPczAzkIEVqq1+o0SQzIQ8jmVwt9hlYt0zYbaIrZmW
8kjIpuAuKprir8E6jUK7CaSaLLJxydBIeLjb1FZwMZEdQBV5icT5gkEN5souz7AH
SX2etWIehnQ9lsMF4lcEBiFUbZ/xSCN1CqHu4haz5zr31Itqf3iVlgu0tufg7yWJ
NBru6kRxlC7CL+03NpXjroXD0P1VPyCMVhf8EFlioUF78Rw+ATDoLHDOkxxRr3UU
EDoCFdpwQWxXyxuQ0EmsF+8FhOU6gD0v0vV0UpFj0RFJtpwGmX81WttKAt7nSUGI
Of8mGYcjfV+rkxaA1VZGIOwAvq5NYqz+YZrBz4XTeOmlyEkgkQbj8HL9y8b8rVuN
jsHuIVnm5XB0oy2WNsQAQYf62R9/VvfGcRJ6qvvvioUxGb0/1zDzd2dS2zzewGfP
NGRz0feySIEMntKt/Pm+LFO11Kma0wK9bswqFWVOf7nwZ57o3ew4c8Bu8XzpZ88y
mKxN1/imztxOBgAbhnh2MhoiI9anyLqqKyHdV3CIaqySG5Q01R1IoEveK4nv8THv
c9+qO0tiTqRtpc76c7vYgdfNhywOf8OYsO1XkjHEdQVHlzr9FS8jPHneMk0mhEWn
XMwtla85KAkqo0C9Nv9kGL8vh1NJtUUyWbZxZbojewSP7j539zbiZn4mF1+Dl5kw
dEFSrYlgUrOZWJZGyHu9bB4UDon+FUpxShgoDCUOldRNu17iqPx4ZMNrvnsrx9hz
/iq9v1ex99tVeja2OxB95RkQccs36ih0gT+8eFa+ziEeejusJpwFlIpB+QiJyXyV
wntslYfbyBiSRlX+5X50EyC16Jq2c823QlssbDZAIFqZEskOZpsHFkcpfcwF3lfI
ORET51Aliz5yF8r8lLjJiqzn/agzlQcMELytN1zLJ0QUK19eY6eM37cS9KKepJ+0
j/BzrRI4We1mGuUTraiiVSMYlSvFKiBCdRmsIPlYueKUngGKYaS2YV1HLL4sBMYd
Jwzr5/EEB+TwRiqPYzNnJgCVXlbH8DlRtLtwLr2Edaan54QugZHl2H9B3aFOh9FJ
zktJSapqfhpCaszU9H3ETKhURHyP2yE02GT9EBmjPks+WSo82udMdVteqPJftiyC
V8pbR6o8qZ7nc/pNWqmyp/ZBV1olNTfDaTHAKV5QJQF+Z+bTwXrmEQaGIbfTefzh
+F2SGep1/Ir/lM+Ocm51eQEFRlv6O7uq6KhzWhmL3JK0A4enwLzZQcQy2HwOM444
hG0OI8RlrY1ASQn5u2nuEzXbhPR3NKPbJFPSYFOBfXFe6/fEz3A4aQULqC7uinuO
HW3vRTamdmVvsg5Kjv3WCNK/BS+m5nbT8fMd4V9lBIM7c5y61RC8Seii9M2poSAI
glz2Iox+lroco0sRHzHPRzwN1LjpxwVVPxTN6IoPpbdOnZWgjR3QiL2KIgf6RmBY
wgcwKDqQq73mT3MquvJQGeX4xuDhNpGG1Q6E2QbOd6exGeOLWq4TThzfS1n3wddu
9YZuH+uzd+WCl7u4q2Q2NOMS5yRyVAky4lm3Is6LpVkKAUrVjg1NEivCaqj4gU+Y
XvISYHl51dk0s7qvX9tOVdAyWr/K87UntUkTSwVQ1qtg6tHFHr+Oancl0RFcqz1o
ibGb1G7Ik3FfbxEMKjX9sd/c3UQTIhVQSnHoJ0ZI0CVZaG9/GKvEKg7bj4MXG7rT
uV5UPu2qb43LkSxbWeGiSHLYNwJS6/8dGDVJuber9qQVIMF7n+9rIt5nzEDuFbu6
jWkVjCVwf4S7aPesEoD3AsotdMZ9dleN4W4D3Lrs0vMnHW7JZsH4xFCAESjKgqzV
KslgRMXeqCvYkr0rHlEJkGoSGUwdP9WwUwajYMTEVomv6jQfcy6U06w6eQJ1MdgV
KGSeTWU7SYT7lR2C6KXg7z0OUFhT+8MerAu33FyKh1S3FP1YCQObcXalFyeUPtaJ
Q1p3CCsninrZyfXqIq8vRGke/59oegFwXqnfeSGXk8vV+rCr/uIwIzClp8XdEJXQ
PETZRH7aGCSpbkNTBlz39+o+HG4hF2qBji/BANpbZzTioXwZjySV/GUd0I17bKRr
86pfxnhuAfCiUDmAgPUKnLSALsWgSEGcSAsCEzD84iiEbq+1JCzSPYth5XMZmZst
LlpV8yt5kJFoL2cYgmKUPUAHGR477eQ5UR+zKk/TSRzVCHFPZ4cxa/SSRxE8O9nv
oJrJ1VdujCuNfTc4d8jBHMoj6a62GwwUu6HxbS0YuDFZ3+xaDLTLmpnXG2i1debd
p0mCjfCnhufJjM2jM+6guCW4vDs1rdPDYs5LQYNvNKXe8eXkNoPWdYgblyrXQ4Ky
ul3GT0U9PlevsVyLkHTxU1R80AoQzuM3swWm9Na7rgBE1wim5Mn7+nO5FAxQrCN2
fxHl/ojATlju2rj+LxninCuBGJ5kJX6U6ZWM7HqqOuXoHXfpUakVguo57UYCgia6
HBUZklRA3eOQIcZ+qpNbroKSGIGrRzxxicz8+gaWIvlhXB+zSaMUsngLDbw8H6pH
7+JfByBtrHXc3jQBC+25/DyTG0mf7zbXDrhOhmOdAF9Qfa7u2mgSY+pHF0bXmctc
JB4JWMho1yVWvIPkFl9jLdkHPqsgAJ9OVYkcZjZWnVKq6j05RFRn8oA7EBumF3fN
r6O+UaIYsYhEhtrl3CDNrg7KgiKSljOLettnobN5QVy/rPvIL05syPfF+FXhG2HV
qLtrnb9TBZhjhrSHoJ9dZ3QaDbt2VnWj12VVD+N+agzFKcIAMCrws9eNnA/xwAQw
/qkosRjrFmd55iDQaKbcLgYCZafXT7u+X4rJA5quT9MBBeQOxID2qpo8pycnIK7r
8zZJAM8BIOabJEGPZfK/mVngEdbVXoSHdBPQxCn/geBtThYgdcJWB3U18IXj9/ij
VZPUBILdUDMOcdhS5A2IsVusW7Bl56LrVQ7r8cnPyY9Wm997Lb4+yTIL7Sn3yAth
h+GB5UVkVcC+rJs8fBIGfHU0Zf/Zu2n/81KkK5HSSo/HgkBk3dBe3/qX3pIqNmRs
xCORSok5Ve1qhMRhF4/W6uxwR4hTRtCiL2MMB7M3be3ILbS07EpxpqqdSNjhOJDy
osKrneb3giAfpqNI9q28TDmOE3xoR/QZdU8CFnRLeifySOwurY6PY2gs7s0Inaht
ATrpgBXE0qyHE23FrLls3uMxy4pJn8HUKPP/2qWD3c4KpEMtOcz9oQsf4lebjztn
qpmuLpJi5dBvtIRRFrWC60lNobYpJuG38dBj5vyIRzYuCTeMIvEdH/y3zY9lYJAD
PG4DmwcJAzmAGdhdYxwTvH/hB3F10UqGXd2/vpbEvXe7rFRLGKqiQIcF4xm/m1FB
ZSYkAwxV1lE0r7sME/rk2KN9MGGvZmMSCdnmaRyDCBz8YEJUwPxBL2ubPrxUMbji
iuUEwSah7pZxusbkXOf5I8UPA8Ii4UAh7gQKCaE6Lb6vgv79Xwjp8CTinrCuNHJd
JNaDkfm1cgMw4lIfMRvCKLQr1QkSVG6KooG/WpUaumxkW2q/plXefFe/QIsBU1K3
sWAVsUY7VJ5XXP1CHx9lZIkBQBre5zjYNNRajpeonyK2YQqlvB42coX/b/+FLs3w
VQx8Bw6risiAEXC6SmgcaeotpxfWcs41KC3ugFPe2sRO//vAy2BHY+gHfePMguNh
vsJTRrJnocdrPxIp4L6zv/GNUwP9yiozcC1xk4V7RYbXm/BKGu0gAXJDYSqh7tnd
qbw6xv4uiFOhJMgI3Gwzs8bXCqXgcD3GyYHQJV47rOLVFtGwjeUPG0uP5FfPlS3+
znvXELS4k7YMVbLKVSFYx3GUGpgbjV0b9IUHCag9DTrL6hJtcEXRfX1fb7FW62ME
t6LUOowLPESizTjOC92ctHLRjHvH4enEITDPsJctiMR5jNvKUCBh3kN8qrzX3yVD
sgyuhlmPykA920ypNN5hYzbwcPN98/NuGZdb/TeXkExNdKX53MFjDx6Hj+HzFu0F
t0nrQlD2MnYfa3IHzWXQZZBgg4IQf315nsjyf3stI6k2cCS9Ket52upU/3miEn2E
QuNZvFuDMgGagAHXIUrVO/dkLhAyxSG2IxWJx1pv2ho2AWnUFZPjWmIoOZq4OIxU
/KI4s1lNtUioVCs8KOMwjBd2LaUZV4K8yFRhxdO7V9ZwpLi3xFK0AzGgy1qnTRCp
LtY44NpZ2KBX8ff5LOwZKCRCVd2xIruXc+Xub+dnydf/1WUmSCXuKIKh4NloCEGY
h4LoOHTno76+laqBVJVKc7iOnhgbl20W3gFHBHwLxKOMocyPRGoxICk9G/uCSZdh
miZ7rQUAMPXBvPtGkJ0N2dJr8M20nM0VbJPSoT++sT87R0kNFFhoWx/UYCJ3Qzp3
jkt37qYA9fteAe6yDvBPBscj3NmPcQFh8o6zZ+q/H10FHoROTFSi/EDiHbpf04tg
V9+vQ74dNqGAxkyrpHR4pdoI+1dz3boJ7WSciV60eh15zOLHLZLg8E0L63knKoIh
dsL8eyuVl3ec4QPHE8HflMMFBDhmWHKyk5UsX7fAH+jUTP38EtV7AhTc5e1LGwel
ntV3ETDV7Ex3vXbB7qXIn7II72mslxrU9q/vsAoeF+N/+sEzf0dRopuLmNhSInKw
5Et/qe/K9e9h16np30nJzBBDFz+fi1U9IECaS99N1kM357zlhLsOqRqN/DD6Tfh4
e+am1XaMtmqNn6assl56YujPM1jFhLj/flNN9eW+X25RDR3oJeC2frXJMUkBkD5G
z8Pvej1M/Fdl1LN5rtp8PAmIApAYbKld3/On+DG8Bcji2PJnMJjFO/4WgwYHaFtO
JKCr2MtFIlphEkJ5eHAv05AaG3XLn76qJMCu72Xy7Oxz42LhlSbsSlizRO4F9EmR
m/KSgyL8yg3jmuBfSN1hWcOKm+anMmktmn7wTbgQ0b/Unfw1JmZPvRILvsZvX3Aw
hz1Rr0aUT+IYJT5woPr4xcHZfOnosvRypgoyCT6fKjE+m4d/XcIMNWLZX1diTvbd
9fS07Ns+/gAXdnk9UTY6Mgghzop44J8FjJUYEReWgvXbGDR56YFXQoLDhWKqge74
HnWeH5OkXUTXLNBzbL44RyYLp7OP/Zq5hGeLQFSuOyuNY+GMEbYJ8fqtP+8jF/VL
ZGwEXkPEzmStqnxW7CSlRpsxv3pK0DjRPAGubDP1NRLAY5ppnbEPyAQ6uQo203am
I6eFOhB7Hcap5KqEhWx6Vh8oVh2wSkMULqjHjRYgOkDODBKFgjmIUtZjFLVea/bz
yF6Sw6gwgjdX0noAcCrrcUFUHruDmGTlWWq4pgGZ3Wr7PgkNhuWHNquNJIBzgShQ
OoGqrH/+SRoU2y+krTaxezArGGPx3AC8whB5lrph8BIgguzP4+udZRR5V+Ry/HFj
MjyTmsEMkEHJBCpFrknV6qT9gHxSCs69UqqrbjyuohpAvL4i3Oie7pvf4uA/bbm2
XVyjCe+Jf8yBK00AXGSVOmxIp4p8g0gMO8N/fOO10Q2nMeh45Z20tn1GWvfgUnN8
AyVBzOLTIWsKgDcc5p6TPbZypfkPnqncTARQz/00YXGW5PtN8eJps7CTxVYUTRgw
mVlXUfbKiCREy19iSOrM1qlKXxl5FuTK3UvPrdsGWFbNw437wMZbI5KQdkDsugWb
q/gt2VAX7FysEeGBbN1Zn/buFmFtOmnfUDQY9NcjhuyqXJsqxiH2utLWYfos03XB
MqnIlswTNy7IMrtv3gnIT4mgArcvB8B0HNoVWU48vSYuV0BSfpNb0kqw4+6yH881
FVhZBOEJn4qhslNOk2JWtZFqW3YlOFBj+lXgiEo5tuH9BwW20+lKtuoa6r/4lnd1
avqDUySkapn+gQaOzMA7PWEY6t6a9RqJFQh6vWWsVAhhoOYcfYro9KZlrcP657C/
AnmYLmJXTVE2QzFrGo3CByqTV018bWBxVqNq9lYCWDjYXMpWGVQz7u1fwaqV0fAI
EZYnPFiVxVowCiSE7nMK6JS2lM1VWigsJjNRgucCLNGH4Dtb7R7BwGhGuDIJrkC6
YmzzSB1EmfaHKkXk5q8wYsBENeGj2DvZ0+1nY2iNv4Etxo8cl4u1OB9lz5BxeE2K
6u0H0eiw+pN9ikg6C8zlx/ONy2rTTONBcKB9+kA0wSNjj/7LenRz+44wLGlAhRgq
Y/Q/pUeL09xwJrdJmuOrJ9OhRWN/tqQKLHVb5Rtkszl01jqHbqv2aZnzYDx1MLzX
YJU73hJ9LmErxU77yIaCB4Zl64b5w44znOTUSmgEGLpwLh2E+ET3S3w3ldUyxj0R
aTBnK+lgp3PkPqZeyl4rM2raM0rVxkc8ps/4ZI5U2qvI1r3NV/Yjf6GDlnmSCANH
qFSwmwmt5rFo4VgTrFLjrwRXwvcjPFfFGTLcyKW5YVhPlG7baUwHuO/MXBRsl3Q3
Q+kbrSISl628sFDqbIvue6T5c7HmHUaAoba7iSDFzKfkOzbEfrmljQaLo9gtJ7a5
kHJiJH9N/Dn9RdREdkwWq6hzs4w6Yeh4SCRjU1BEExC4OxXWvT/IVsU3jhl8khoM
fLvv8CyS2cyoH3y4aEkOjlzbwYvLywrhmFL2AIpHPU7pWPNn+qbnOoM5BYDKXH9+
Qur9SeIL8tWscF+i5AGipcXCLqgxZ63lI+/kwdilRC6ZrcJfL3PdtRw0X6GYPhjt
PBJYyf2/6bGXdM/uX5tOxU4lhyHG1WoAlrSjbE/5XVxAfUBChwwx/ZB4o4obk6/1
IZUEAKA8qLQoMm+O7pAyXULXcyu95/frDAtn2seE6Em464wss18NBEs2/GqwvrwC
LEQaqqTdNx0VP4CImPR+mskxlcQleuVtR0KB9iiJ7KeChqZSJp9TiWUbaUNxYlNF
avPHWhnZ41hCwnGfLDTGiCAfPdklYablB0S+tNUR07pBSD1ynY2xVfwScdgWGBos
jcJFprNTKqsEk2EzXeQGznz01jBcb4NKHyZt2QXgsidLdIpIs7mgkqddJnYQSGvF
sw3znHnIBDTR6bf3w0C0LdrUZKPxjvUy/aZuL+LZcWzCOWn3zipkvhVkcTTo5wZo
Qr5G0qTqvXcQO2IhqEGUFgN5CVF1UYCrHISb8v8twOszaBRt96gd+x8ljUVqb7uZ
t8+JtUEyt+uLi5/SjrRgjQxSlR5q/2czz0MxvtbVzQcymSGneUoxz/xbIlR74jgY
Dp6fAJtFMWEyUmeKcNb1XYmvZzke3s7Ty1HZq63yTpniICbh7M04v+BHyv90ixLL
qz7DxMju9ewEzRV9fVuQ/2VwygM5+6c5Yr5aNpqAcXnKRUKjDmV97krOQ6tx4kqt
wH3CS12/Sf1L+z0/y4xGPEYcAGQBfc7/87eWmIOOAl6hYfN24VnTKEDFSFPda/L/
F3DsjzdOn4gtScvM/Ou0SpBsu4iHs0XxvMGRjYN9/huueKqHocQ38gXd+L/1TVEe
i5kU/R2y6SjsgOsuB5SYQnkDamVcWCzQdOP0aDCGU6gkAvG2CvOv8XFYBEgya5RP
LYbjNLPqauckUcoLPmDEfcgZGTYah8dIlIn3Xrf9LNbCeSSarqqih3RmqmQu2VBz
ZzYRvy0dLFKnq1XDdOr5FkVE6JhK5rWb5zzsvUYZIeDaqVq5HCvBEVdX0eL7BoN0
eyf1fNKdJ8r//ik422KM1pwhkRpzK62d/6ol/hTEc60Jstu+D8mpOL8peyprd3mq
hbcyP7vUVujjKhvodDwE57l2rJTfFqpDOvFmRpFQ451Z3FRxFAzi9D3PDJKFVJOi
VUtmtAMFyPH6/rMpY7jg6J3KnIrPMY5qlQA5X9ouTjJpSXAsSeKXGTUp/IA/CQva
LV8clt+i5YKpZBw8LRfPbdwy3RiPvTxpGTtwy3ONHjKMNBgA1CR3tHsYZB+AHCNi
CR63T3PGze5NNtYucKgalaROHm0jekfx64Xf44xve2U1OLMB4Vs0acdLsla55c4P
JnxSENPCxtx1Zl3zKH+1kuRHfCm/iGqVts4++BWsC9vn38xwYcUmUdePQ7knf0SX
P9SQkrEkBtbPMSimJsi4IL+W29a8ptkoNpVXcZzshvDW3V9TyWbzRrIsyW3G8TLd
SSOl15I+YvPDBNNCvwIYxZHDvoIMMrQ9OC9pNurDxzyI1fFz+mAlGUk4F2uGB7DJ
f8NWyJ1ed61QUNtsdonhIa4a7Ld6F8v5Bt6bRaVaF6yTSp1olx7FjWczix9PwFUj
w9W3rLWLM3yQL5PUF41gFzbucY8iGluoiPcifoqVNuzLo8+zKfh+waNUr/iLvM+J
5a1IkIalRZhnlLsZKF7ooJjPg7LkDKr0VSTgnJ5H6vMhccxeAK35k4tEG9HF8V0M
qlFwwHpjstJyarT/4dvmShU0pVPiumEQQhWFjbFVPzS4OwOF5qcVN6VoA3PkiyfX
10z0uzhDsfrL4De5l2YzcxL3m0hvA0EVPuBbxMKpUCWwo/6zwZGN5prwgd1x9G8F
/Ah5IpgptXKvlOiHTle9bJMIgEtVr665M79eI88IBQx4NBhnOgqveMBr8O326UPo
O39VsK8PX5LOg3ODh1goT6HNgf26VYVf+2HdZNzzZkdeLzf3dLeLBUummHCg7wAO
RwBVfzaXqefU9KgxMXpm9R592l36jZlp9QZzmslXFU+5FiJ+Kvr+Rm1ijDijVC23
0J3FQv5TkDkmB3V6TxMZNhwSnjKD9uSON4K8ilxPyR6lmPYdjGkZ65gYlK1z1QU0
AAkBjO0N2owcWKW1olyKgkpTLBfrVj71iLIJWIyc5jxsST20yaBcxrKzSO1zA13r
UIfpAxTtf8HWtt4pIRqPBX8BbaR0omaII6l3h6gO0JrC8tnkNsAk6m3Bzw77AbqF
0QNtoh+wnLZcwCY5cQDl9gLE85lLm+Hz19H58Zl+MQDpqDMK3HXSUf8WdreiUA6M
OVP6nMachUq/vLvvJmtzVyYvI+jQptg5ob7VAzwqevaSEvGGgZWFdVvrFwjGh68x
Q7oFQjvGvpYglHlTPTFfXiu91Lz5M5qL5C2YXy/PnGRMadCfmmQT8NyHmFt3QaSI
Cpic7EcFqPf/fa7U8X11odzneP43uj2GyWtSukloBmFgqZ0l8bAczJHYdAOuKq1t
A5uf53oCwmgrevYOuGQ0TjUy0JBrBpUZDig5/cp8nW4A3+PjJLXJxUiRy639WaRn
0QzE9zEyB9HeXTA9gLQIBdqBt+WJeNu9bB876nGJqzmD7IrkK9LPuL3wVwNmdhKZ
gaJQeWplqbRgHn//kDS3qWAAv+WNUkSRt5OcMoOIUtqpFx6nitaLV5O18blC6LOx
xDomzAqACw2071HT8XAWEwhvdc/p3q49mOlPVPzc/huYB4EBQqtdpolaEQwjxQni
Dp8U+BcnCIPX1fOwLchnJ8QxiL3lSY0JDFtifRI5Y10AY3X0mc/xwBddQt18SgbM
U/LNHr1sjif1+oKzzg3rHuOhxJNZ/xc7Y+Gpoa3IcuuVkPKTZLQFZnvdygxwqDuA
QOLV1LLsCpSinrQoN2IoKNQtTl4MWxvq9IuqLJIu4vI+S0CYMlC3z5KWtS7bmlQv
woaULfH0p6FEG4Dv2lKQtENbpQHup9A2qY5T4wsUWr04cu6UqvKhtch62Cfjmxjy
yUU4E3J93xiWMsmMMnf6tdLsoctVvVFYjbPRUqFwP0iVN8JTIt43cTMNUUrMefmi
KIIlC+IN0JvhJCvFCbfkNUMT/FZ6aFvUveYDiDtuPDsQI1hBr9iv/WYhoekqHp99
sVx2H6Q0ub5x5HhXLCDUMZSXJlOD1KRU1Cl6KPQRoUcBVKJNFH3Z/VGw/kBFwO5B
WCT8qHQQEX4JfAmieSxM9Ii1TFrJY6DFkIxnhApSs3KEMTqnxMPeW0Ch4xzVMddy
HUT5AT5rTFjfBwiccFdf68NCluTqQR5b+GkGmZ5OwiPa4ESnJu+MIRxNn3HdZ0C4
Ss2b4aFNlqfQfjB/HzL4yxipqXamgnFlHL7Ig7++GGOjSL4tqLfVhtWJNUSu89p+
H39MLj39Z2dZG3d7kcwOTIbxDmY62fQjLc2olJ0iK0ofeOBkcDaLJ1A5CjaeMOpn
2VAaqT3biwCiOrNA763OjOTiHjxE8E47Bmy2w4n3UHypHu6VbyXQcgEWKQPAZdS9
vuJgk9bEtB15ENottQeQBzA9CnPcEQoXjvGdsyd3DgoY38aDrD0G+sdXyYDeKXwG
qWhKnr1/UctrOnuw80FGdZAmXjvIVkNILUysWtUXd1SgyQqkfn4Kg2A8Xy9S1kfN
gBurVDZcoaCmLh9lgZVKXAzPvrPt2Coh5sxizGJZXU3QqfTkXgXlfCr96/BI6A/6
T/BrgHElXkin8gMvNeSx5vwNUsNSDbbsVu8CmA+PCLNA/wt43wpP1onX0F4zhDP4
K3T8BnD3gJm8wVYGC2y7LRJkZYgOeHGDabHjLa5Xkvvgqwd9H1AtFO5tlx1wt02q
PJ08tLhJNxXxYhhjqNbgbd7QYiY3BLPGx/9tH4kgtddUMqI6PZlgBQ1Tl33BQWrX
n50uYuUS73CGGhg4vHfSqerv8jtMngGSW52NZXOxBIIKZjdrI4b6FqCh/YIu/czP
D2Z+v0vzSDUXwJmV61w+aAN5DjMzfvgA723uhHdesu4gV4+pq8OeW1lC91E1VYCf
z1TLu++iOIkqnjb9MUclRjPMVbe+dNeLD5sOk5wYipw/4xnzqpfczVj7Kb/ERTCm
okwvrggfPzz4LmWpRZRHy70NuNc3o64i6sKhzslxhrSKx7z75t6Xa8LGr1qxRQCD
49iBgN3ebXs31aERJ9UMTBjEpj/00KqCIuh8e8wJubXXA/WU4/1fl6bJX/NSgGBA
eO/fPgeiKUiwzxMEZ/VJq0C7XiwYrLazbuALNesEVdGjHoHXDMnTU/mBjwXBd1vt
Ld5sP8tji/F1UVM/qZFW8HWRVYYks6/w2lm+s146Lp1HDpP7TDsx0aLoDRhAhEhc
vjQ2qSCuzhbVTGcQGU+1R7N+E6tF5KRtgW4TvmcXJfMqbrzR6E/36ObD2J6uEJSb
/37jtZyYEfzyhlBpZhAWQWZw3y5ubFYQVtkEfivXTl47tqetbn1Jm4kxKq1duHhB
EFB5Qk+xrQ61sHC7Q9bVbSHYyg4uIPQbgAoE0OsBW/HkWk31WHXuoxzlJl/7FWwO
AA20FN+4qy7IKcOBf+A6QE8mSchqrY0JCWp91m/b/NbXehHLHPIODgRnuamAi3Ji
y4Gam8zlJNdwbyfCFSBUz6AOVlz7xFIHe729E0QUDstMHeJba5MR5KaDTEosqdkt
J6BX5sg/Ie02HJuFCeFKkXNelw/p8gMkoxYVtV8tWM8LmrB5XWmaeYha8xjamExZ
clLbHg1f14PcYgJzIUTkXQcwYOflTBiLu/mstvUdbJqaeOsbW6i5ar7R4tF7WotJ
2o1wmOYja2ZowymS5bxHvnA0QIwLe9P17RF5nsyDlQ8KcSs8cSykKYpD9AEY0N2d
6OVBpphAfV0nprrtZGA/n96x7AU5l1o4Bqwv6wDh3MLj7UsvknyHfY9ZL3xNG/Ok
vLHafwslAJ1peXy5OjUdFf1IuXdFnLMnzbjED6FZWnABfLY/4q0bKBb8VsqC4nPt
ixSXvMuQb3wPmMnalWycSASQsTWLH6vfwaxcValn9A/iHt0VJYRKbH4gVloPHVzy
m5w9WvPoQJe1KL2JnVEVHwutD3+fDZYNN4RIlqYxFjymbZ+6Z0t3IYcbKkI1zRc+
Iqo8OrFPHitnWxIZ5wA8W4qGJ5Z8j8gogH2XwTrZP55IjgbhNxoI0Lk3me2kM+ny
rlrz90kvKq8fmxW98pQRZpyROX136luzg1OJ/sGRraHJ5a9Vao8FqTbY5vBd5YbP
QyM2aFx/QyA/VNfM2u8SCQZoxLzhwkeDrhXx60mB1fU7k49kk0mmo57SYlGaqpTE
XDS0HYIIVIX5+eALGwhXTgPMxbD5OfiWAib4PIjee3hd47mEUPBed8+BnJJ36Hkr
144dO/MFkF9UsE+JVgAxdgQLC6mKO80uF1cQ3+f4sN4XA0mVUdpKHcPKyjUT7tio
wBj0VAjCigqgKaidXMjP2QK/QZSL5sdys7EbSyAbc4KP9TzIXTUeHyunlemZlDMR
PduXojTn8YGp9v9LQejE0kIBWUnezwEAKXchxM9gx5KvfNuMOxIcqz2smZ+4SNwu
LbNS/1ZEXOcLXMgNdeRVzuuLXE6qlZoqMekoM7jYQf5D9eJl2dlOm0B8UqpLsyRO
+ODVA/uduwBKhetuQ/bGADZ0KQOKexKRZ6se9pZoSRRXIgZiVjtXsLsThkMimReE
YNiQ05EPXAibfw6njME279IxpxG1VLKY894LSeInQY3QV5fkULjsAD3QrONcQ5Dm
btdWH2av7v66iknI5YwOcJACoN8bvkwiI+lm/Kb1nPk2DnGRe2STE2cSqDpLC6OW
DoeUhi+7DaO3s6Yk/0e3ou7ssBNCUc5M40krmoXWE9OJMyCt7gPdzTXQ0h4Eg4GV
b7dyjkZ1/vCLlDBJObWcvfMYlz4awGF5u4bLA2WqEkMbXb2McIWbozm2UGRkBNQ+
Q6le40t6rCWLtjKhk8Hx3l6/MnoT+CXAFRiFvAytyyu/uC2FW+yzIo4InkJUhQwn
i7hBpXnwb0Pyt3nWhv126unXqzJl/k5UX7zWuJscdSQFVznt2nXlMUdIU/dd3hgo
tw2uBi7XjiCJFDLBWd0OaFXMnmQCAEOQz+Zs1pPQyQwM7dxgKBmOq2dF5A9N5Xdq
U5SeD9Ck9v0sWm4bcD1XAA6DalYvl12axeU3tr2dO1sZLTECbkp728tI07wPT9b0
vqAe+MWxuE+FjD+BoAdKURKjuIj8ea4SMDHv9ZPZjgHj+gK5wW/5uXqMukDD7p1G
AZkQ+GknHKEm+LIN2N71VlxMewDLkEmSrvGYPzY2qIGVjI/ehFdRl6goAWmbgK08
19PFItP4MZFQWf7oNEYKW/UAekyWtMM0/9trhgNefcr+ve+KjgeZKh1KIdZNb8sc
VGGJlmZUYjF75HxBL49Sktcgh6gzzRjUifri0GPOGEapf6aNjzwOGd5CVpk0kFan
Bay/lCGqlq3/uQ7U/8cZYC47u5KtzINmwFhfedthQRe36ZRXtdQqcb3pIxaRi7QC
Qa+PmOSl6xL1H9R83+uGzxViS2RI3eAz00NLaKYprzx1NxsQvZ9dwowXSYidBxp7
S/UMJFznLF6TXVD6FaWOO51JW8wdMKwogjcwZJ0f146TgGCoaImhKgyp9ecnUyDT
f8NsCS2/jxmjncR6+kEdnTR/BpCt4KJbQhP8Nhi6yRoTuTfqw8HEWUReDdcub/bm
aWvq0QSBrZCyNcjIxU59TL75Km64TMDnHjHGkwSNZ86aQyH5IYChhSwlH6GLlEEP
qzfzWmGwacD0ix6l1iJ7nYojjZO6Y1WGBSmBLoalHMphLVZv6UbDtw7aWvDL2krH
3ymMDd4zNrQyD73BRSaBntnVa2uJA0GytqU6lXA3lgpV4PCQX+sXUm9xHMAH1loq
KUAzzreNYz5esM7YaQGMxSKOtcmQOePICwkKxKiFR3EF46wfKWbsSugkM90+apRs
886KSdjALZ7eQQOY6AUpB/21CAs7d996O3pzt/M5CJFaB98m07GOUpnkaqspIi/T
qdJ3mHq9TqxbARNjwx4EOQHZoA1UqdtDomPLXyxfMhqHnDgXVwiSEY1ty/lyTkvg
sNVfSCpOfSHwiljr7HaichpoEZQF7td+GSgff1/Z+sbMzN6JHwlZQv1tfqLEq50U
3JNgL2Q9JqHFML1MvDGGy3NWbmG9T8FWqc7eGmx9mc0NZH698ZFpg7FSGhaPg+tY
OmlvdZcHoUoL+pILJaySBpPJbHaHs2gEDb+p3HdunQJZf2C9VwXqFWQHUUU9n8g0
RFxwjsI1Ckog+L8VVQfFTASUtt2n2Pn+57y9GrOeoFCQp0pMvEIe8OH7yuzGKjhJ
Iq1uFkC52GN7EZ8rQ/9MFXJ/vILjUX3nSv1oJZNqcVpc4Fgi1A3qG5buxMjt1euz
4Ep8H4fpdOqAduSELdJOq09JJBOBtP6ELrHEd6EdKKxGa67/vkRYzPnfx0Y0+3cy
zf+0laN55mcj0vappmBI2SGGwWPQYE661lhftyEV8pN7cznV/m5toM9wmSC9h7lr
rb2uwblvgGgZWwI9/hqT8K944zEbogoIGW1cnqSLdZcjlIkZ9rR+AjVsrCsza2f2
999iOIfzg8s1pSh2an5T3GkmbMCyF8a0a6nFjnltootzVVIHDuAD8GwVB6LSdsU6
ocveUC95oM5jo0IKa34LvjuMkZKQMG6xLRCHBiCD3yi6w5V8aZq48RojVxkTlu/L
g3MK5QQGZqKTbdC0qtkbKlYYjnYWie+1TyKVrdO77ziPqXLl8wRIdxjCMo+n7/5d
j7t4J3VQ/8zocbyWR/YrEuLgyYabtQw8E8E71oD8aLWbM4tIITlgs+ouu57nsJek
CvxKbbR9unNGcMCo+dQQqgPNddoSDQqhMPiKlXpikLQQyKwzGVMrgx/t93FHFnJW
UKa0wffv1sDUU9OjRWAahVouxxcS97HjQVH2KecK5aWkDTE64zXdvYyk4IEhaIOz
RripylbMXw8tG+RYNQUSCqYZ8z6zlfs9Wuokaan6y3/ii7SUTmq+tpHmQCWsZMjS
rDPdshxt/S4v8IbHHemAM2FxglMfjsLxMSqq70AFsXwleSIvUgiScn6+ffCmcXDY
SZUXWitXDmNjNg3qKNr4oqk49JZc/62kSvkMwj9hgnkJWnL1EN5lau9efPok4eWP
7gtqDn8W5bccldqIYBhRJDtO1WDlEyd+ct1xgtxo3Acqb7bSsSRgM0a+rlHMPgBa
wnR+R7ylNBQLBwIX4Pae3qzRURL1OqTYFMF0v0IzgDLUqlLFcPfqctEzP1yHFeoG
1hOIWk1T20OPDcsTsW/cjVwc9zsoFIiiZ62cNoXgDEDZnE713bdgCtp/IQ8o5Hld
LgtfBEjE9fu7WEyIdTHBqCr3xVXKSkZ4xzhNfdEsktCIAGikXPDO9UISS2EoEmFH
TpMGsq/AlS4x3bxmzvlBmYTADZI+cpQbpJMGtmLviQUHnng2QApH+LEiBYh+vOV4
FkTLdrS/iUX+2jqdTQZl0Txe18gI/G1EroknPU3ORo11e3kUu4EyGiA123f3ueJQ
uJk3QbiKU1TGCR5a3zwEvXw2Y4Cd/L7ZnWKNVVZrBdoDmpyVpURdgAw0ouomOtpJ
R7AiyQe8B6I4anRc3UbyXdipfUi2kzvmDehQXeAzmYIUBzFtTd0C0vq7RND+LINM
Dn+3HH+rghe/i5t40rDiYLtl52JajzNO7oUYAkG3wZqJF95/izWuYMP+uyEdSXii
Rym9q2yYnu6oelp1EEEC01/UrzYTdR/mEuiaayocMP9RibWdAh67cvzzdtzv3XeS
hrFXCrKDHgu8Z0fWVMOBFu9acWV1coCUDerEoEacvaIosO4FVdUknhTKKOYPcR3h
W1Atsuv7eBFwrpKs5Hvnw+GMaYyx/Pcc5S+ct4ExLAnZdEHdKDKfBUjq4ySzu1//
83HmTM9sM7omsCXCyGD07OTQSMX0BxZ7FluyP8IpjOFDG2MuRXvyz+fqKn8RgQOq
QKsttJV7J1qcWha/DQA/SZrIE/m8OUHJDwmyUF8qg4jbV3QyVlz4sbNivdSvzoHe
pQBN85S2Xt8CcYZVVzrscoTSI3ulwbMSGy2IOH39QzPk80QzrhyFxbYp5OAmAUtc
wmKYCsqurPPvk1AUIcluH6YN7pdFvEqB+z8yLU52JLcZT7D55kIvWMo6uoFKlDE4
LMouCcksGaY+k4/z4HQZROVyfhll+qNnqcSIYyjsu2uFdRKObWvq6gTd0FmmRfD4
Ld0XgN8MpxrQafzAJETVvD4t211m68E3i2Di7mpqX3K4w21LQHiDZAuI7+pRmxNe
2DO5bsPbK22YPN3KCM5yO+df7SST3SQ0bY5VxGzAeh+GjwAanENKvq/BawaFJQcu
tOxCI2uHV7UKI7917BdI42XkECTeQFJbjXZfzywUep/JPil+awglkxiKwf4iseFg
LMil5iDembz+mjznRr/3dQbzXRK/MFezEmc44wd3eChPHdTKpUVL8JP3uMLwx1sH
d6GWOzozZ3Dm0udD6VjIZXlQp7nhwZxavz+QvqYw75zT08eRDHnAINWidNuit8VO
6PMdEZRb1XPAutrixAChFpvGMPouvU4DeRpOofFFv//doZJJhRIyHPnsA93sUbgD
bGJ0HKdIny4QJg7UKAxSHmCHlQSs7wRG4+y2XoZkbS8DEjyEe4o0aTzCOc6xqmeN
C1CBKxA23tVGTtjv6XnUfBR4LyrupOVNFbGGXn013wzz83CAFKf+TK9HPGKvnHzY
pzzuR5jh8h1p5cR0hBYRcrbaBZwISKlQHxEOQhNbLbqWWoJ/ar33chXRRJQ0Bulp
bYaGxebVbpp7Rt5ll4EPtpkXc2824+fiBoPmpqdqu6mEw3JtK0YERpBaMwtyJc5B
AggPzF0UyPtYj1yGhaDfJjOhwXUafssEpNPyD8qxkULJE4P6YvDUq4eZsy7HwRnk
JRKK6EFut940Sk/xXSIHN7uAQacgMFjf+z+1becAXDV0ZDjOs+pUKWpAWkNNMtGf
vUHrA29ehSN3p7ujpKZ5hq6oJWFZ0+lhtKpeScKKtHbon50X1H7av5TPGSvYDC8+
vzIVtWe10d7cTBl2CV9uzSBZ3rJ3cFpQXmgMS5J9pd6ZEf/KudCmTNJsLnjc190S
oaW5kU0/zH6d3qaaAIj0kTuKcJoqghhvCGOQ9L80C3ogv5NFlAsgoOx65mZ+vFyU
eao2r+YLWabI1524A31ZKxquIRpxWYKd3N8cEpvhRr6ywBboCbD8UfgaIJIi6Db1
n8oz7bRNq7uE+PVYNo6O/wC9yBdujtt0tk2V/Tjaj1ppPjs99cuk3FfovJ9geT9f
rii5u+dj/D0GCYyrXKt43+jLu+97wzzeXFANT/w0Ebc4tYsH+ThOhXL4+GrtqL2B
/QwJyMVrFpqgRNgDowh3pZJJgJZnMWUai5wMr4D1CJ7ySPsAe6oEv0tDJKIoyykd
7hJ2aOOlpuuI5FsIQo/M9LdIuSpzWETlO8XACQ0EfbVkkhz6rI4P17BuQIRMiSEL
awH3caNx8Pk+PZ7K5ywBUvP0mM4L06n0KOamQU1V02mcpt+5+OWl0rq5AZxLvaiS
ogxnrDZkYFJ6ruE/Oimik/EITgQxR2z22s24Vo1JanrLQOpOPFxONKAhO9JYWnVn
BYpPFBTfO7WiJNUZAE5hp4zxXHxZQCcMM3fmCAtFqNDLTHOrX2MsZ7WNIKNGf+6V
2UIHBrEdPRFLPjMay4jXyP7bv8i/Z2y51cKumVJNQQ9BUmMI+2LJMklshi0v1Onz
V12Rn8H1Bz+XxeC3KKxNDNmplr0uwA+9QxLjpgyXew1UjdCXHy9sC1IWca9NBd6h
BTd0FuWj1QfRxmoYdB7vdO09HQfGF79LiiqQ4keZc1WZuH4EqDPo8W/pNccrkW5O
IxM0n+tECRLxemWB7oEsl32ynq6bdgqONqrmfpI3qwXvckqOev/daho10LGaKHcV
QDs6ITV1aP409/K1C2jQHC768kX2LZxYntIcehejpQHJP3bdNym40mc1vMsPVRJc
Ifn/ZWvpB0Qf5JDPP+S4zWh8OKAbFw04J4WwmG7MDWO9t31I+OnfhLG6ndsw0I69
AylisNy2FfFYbgKpR8nK/jsLg7Jwt23qTmJTrgw7KQ67cTSonFNoEay2c61Qs0q/
NbE7NcloRwCfGSavrRH87Z2ufBsGMp2pWrCracFXkcEw7yjsmysMDfDfw2GQKb5b
aUEnlzoyL+0FcWoUy0w1Oj+x6EADseWiZwyBzUMiQUZzf+gdP4hChgReGKpma/Uh
jfxDsy5JuMNCL+olj/rC+D+ji8uBzi8Jcvru5i5M6SKeeJvCE4cMQZB4tyG37ANr
zh90dPPEMtP07YUQFodPS3rNeWj+5m9HpR01F/FzZpyGDH3O07LtOq4faSCHc7ZK
gynU7dw6nACQ7RdVKSMWqE3GRPND9Wt35qJT8L1ce/rejkQ4vn0xkWlARoxfLXe6
2KWj29NMXA+biEh03Xm6g0mCCxQAPfe3QjssdPnwpKrYfQt5qwqOdcEhu0iLEjYI
0pMwiot6+7g4wLaMsuV//koBDwVmqD3wy3Vlb2FhYg3tt+fQaT85fcaBR333sanf
RdVjAz/gxUfvk9tivWjzTLqSXVRIvBNdWJfPHt/vWm/KnBRg/ZTB5nXogSjebqQQ
kYd+zGUDChYAmdWUKrBzbJQatkq4h7FH0WMGrY6vi5eilHqgFpmqvL9xhXONo0zZ
2m+GASMiAbQYIoevOAhFuRkOqh4MeFeKPESQ2UeHfQP2SlQy9PTX3NL5taof5HQd
MZgajaLMaZ5qjvurArLLAM5DAG8VPcofhG/Y7Z9LjegDgAb9r20nhjCelf2TDWvx
d/CnBR3iwFLOYBY8UocIkaNJrjs/NHi3oQbDzy5NUf4OU7izkTpNP8K6PXHwE/Gl
NVMjOnbhSWlywqrwrljHNAvoIOMVAC58zszfm8tJaaoZWU8vOJLkvTr01gItk328
BsihBTK3kno040Eb/lfaY5YIPQts75+LziLd9RVBD9NLeMdRPRhqfEOxwQtTV9yr
9Kjygg9x9F84yknD4m1XJhDO0UX23nGTqEiaZY2eMfjf7DIuMWNtJYpXLjf9OCbf
1jh8XTnms4yopuNEx1WfXGAqER1Nl1zEUzpULpzXF4jODaj9yvctTPtkXFLprqSk
ZkjzWBHT39QlpZsbd7dRcPmSFJXCPx33wVZiES4Okj79+3ymxX61H08YWb9m29qJ
kq8m/WBh/o8kJJrs1I8qfW3txM2M83wQ0e/76mFp+0/EVbkiDu1/p0K1y9wPiw+9
jOeRWEW9uOY+losV00qUdyw5hqJHeUnL7MDOrGwPwxJEbvTXCu/oinBjjLzvSed6
BQUVEeOzunEJUCY14IriOXJweyN0/0H5uEz8tizTKWMKHro4NiZdFKCTTQM9RDMl
jbdwolVlWG/czQHwdwGtXvFol+Ks9ZiuVpG3mFbwmXMUEiR1/+jctaHLo78qreJU
Z2reVlSoVnXJ0XE1+iBEc5tiTWuEdzX5PDXJKv2MTObz6rUz/6iSzDkFDkNu8GH/
zAorFLDgydmGUvYWGECW3X6HHrsCixUTrsHS4V0s2nJL4u6Vm6f8hztZ8lLWynNY
Nz4h1i/SgDDT15xSRs/VnMU/NP0o5r49WRep6sSWrfurxCiPoYRthYTl5XCGcuHF
dmTIo7uDwn1dWOAbNhjpKakuh2FQpY1fc3YG3cbewTAG3reB92ZPTHthtLq1mNbA
SQMiYS+mmWLFfjKi1DNXE1/NYkSlUBOyUIhHr280B/TLawsv7j7Dabs0nF1l2hzy
WJS90QOBqemXw4rHQAqj7e59t30myQjripnd5hfdtSKsge5F3qxxQFtyQ52z8wVz
Wvx3rdbVb6dHi5mgwl3+reCMprPNN66d0/s7W2GasqgPT0CU8OIioW1r9ZYLA21N
7et/IM0DauLqUcP22kNunlEcALqgsW1vmDL36+LCPEOJdwJdKvt5So1yd9Q58Nxy
93kqYQDPz/TYHhW+hwAU8v4/uQwbDlwstiyAlmhREBW8q+w2+HupJAbOQHndzBBQ
DDUSVdwgR015mSkYtR+OR51gJGD3gN5qI17VzkAHtKCQ5pTZ2ScZlCMKkQB4h4D5
vh05eUgc7xD0RtQIjLb6S8/eYi80sQq0qq55GEJ+HealnnVnMcKg1liFVda3edOC
OYXGbftbOilXXIeouQfcaG/G7QzOEMSKmyyEV4PY+4JLLAvcfFi9WyM1ol+a1KXh
eB9K237vDBWnLxNHbjNRENplXYRM8dmRQUJCf1Pcdf6M7UVqtXLEIotbUj+JzcMk
+ZAJ8+qhNUhwkZm+JUOmCXYCVmhotW/5Ee7mxNx5ZmLVI1qNUpRdZpQFZppptMjY
eOYvxV6Hh3Sm6Pqpf6cVXuX95CjwWncSArqEBS6IZrdP45dWfTQbBqd4O2bA5wDr
/SBmXifSecmVfHsMgtrPsOPilQQoi+rcJMurd5k/0A1JJk8/eNie2TU3sAJkaCFY
7zf8gDWdeQdWF3zm6dyIwwrrrnDisiWrYJwCU3T3v6NT77BcBj9HRrkTGSlQkhUi
CtTXZzd1IpMznYFSvttpA2i9buJbsnzTbfPpfABlhB6KfOsx6T/l7ALpM4PZAdjm
uXtS5XuZYycJENymTlYTLVt5s+sinBAzLNP7GV8Zz6Q0AeohMNBQee54WGoJpDO5
11kp+oc/MOUoJ0Gs2wE/LD5o53RwukgLNUbZgocEKRHEHPMQS5qTLU6xm5zdKQHX
FcWE0aXJUOFLCxYrFQPhSvCzva+Mmre9JRB93q22qfSiBKyx1gMDEtwt8L2WOFfB
I8HpdUYp1mYnkxc0/kwBABBsKVlv4iG4fFSmZuiL3hth68Y0xjrT+YXRftMznNcz
2cZWGFYaO2XqVMRCiLx3Q5ItjiGxi1ESAyhw3JcVxBtJZ3tStWrzJA3i+3lVbJx9
EAELWkK2wteRUNzCkbruiaKw8GYNRNn8Ufra5Zg2DsoTll5/tmBY1LIwdvQCGG83
LNePpTIlbWsKkD+xZBKizn1jFMeCEIStnKT9lysGVHKKc2lBuKArZdUERMNGOUQk
NCR3IPQGtk1Tcz2aJuNfvTHpMR1JhrlU0dbMiTiZYuB3741grT7EPan1goErKWiK
rYIM7Sq6ss636p9Opr5LiEM94rI77I/oSoUSGKOLphSoTFXiH/0aDbZKYt9vOozb
2m72cxeHJCmebW+0WH1P89ypMPaWlSDpPpDyPi79KPBx7MDHOCLpn5Rar9TPM8NI
KLUpDaLlAPfVr2zFt7TPaTvNhrXQwWln5o0Tdc9sZAIb/VemRBAldYekz9A1+euf
gk+8eklXtFpaAsBeAb3bmBctYk3rAuSVbu6v8uZ4NoILW6GFsC8SpJ5upLpzI8Oc
RaaUoq7DJDp2h5FYA9/e1EoxOjP+xkjE0BOpsKuAfAJgTY+Qor7/yMODRUO/UYnP
/gluIzv3w9y0quxMxSZ7bHb3YYk7vvbdvkD/KI6dEEpOrz4aFPeNS/zGUcePMcvC
4VirPS0mkMm4me6jIT6OpR/nA7s8ph08ZBW3gUn1IpR5mU8CGJssXwkfp12g+hlU
9f41jJli5Xs/RkNJUWGTgUjzUAiYc/o9QJjATA0RU5LsRD3UHCp1qDmmpoOfzpc7
bpSdL1fF5jnJ+KNYl/q91IKu/JPEUDQL4Zf/sd9BILtd33R1+uwSwjw8LNeFBmfa
x7pVBdIOoBkQtxYI+PUU3Gopx9lMGEWfEPBEqBD+NDqPA6xGwtOYr8I+62KMYvjj
kEpigP4KuYVrdHQY7tyy82uII1V712zW2JvqSQjlxQ+QB+SHMzyGagNvRzSbV7oM
1RfOpJoJ//r9c0JNJiipHoqpLV4nsLED6+U/tqYk/9m7jpQCqrnLTc58DedEN5SJ
DMrDHcGOl08RLZOcP8ZMTfwck3fKpJb3F6QslzzA3yfpqDJIv5t3kFF3PRvEgw/F
m2AdCE1zk/UoR2nwZrvR0HDXYoP4d852V672rLqTomKnC8W5ekPEp0dOkiPAQQk2
DQQvcezbpLrw9YD/Ie4LA05pvQGgWNzCE0+1g8DqXJqC2CbtnnDuabG2WYb6Ssw6
D0EjD/cdrgNdpRysUbWr22Yl7FC4jxd8hEMaYSjNrlAzeg8dtzl1BV4nir++rZ5v
A56PJ/ED6kedG31WB9sNl9HV9kK8paJQvQgAVentUbZ0eKzwBjiCoEeql1OyLICY
BDvv9Va3QODTzju741EjJe7Sg4RDydLF4GbkdhW8xyqLba781UpxLgLOLn9MlzVA
D3qNXQvc9iVUMXG7i4u95bQc0ZoH3MpuMqWNtmzgynAHjfMYViOJBTauYK235APM
pM17DUDc3xCfy/qdHo5zx+91xjoQ282mxu9GNK9RdhRzyd9YdqHpo43FjBTQY2YY
ufDg3Tdjgzd4knTYVCPga2qPpySd0KXeGaR2PBuGIveb8nxamu3dvMgMAHTTwsaQ
xHFJ6k/c728W3Tr0HLYnAk2DpMYFnfzbYS4lpaMHAhwhbe8nmlEMcfc6olelRCby
xprmxzVUEvxe5H7XVnyMO82rEvzPidGrRFzJ/UnUbNhAOAOFGu71URgtVAR+pIYX
I17d5i3PiOQGZ82q4ggn0s7jN+MvEWrNG1w282j0aBdMK/BZqOZB+N5yY2V5x3WR
wpcdy52JWasyLpmWQY4GgbSEfuUdYjU1pC93A2+wrLrOc7eIERWzVF+fr3THXZCg
9cU4e9htVcmMWco+GxHcoEnEthCY4yZlX7Mw1UjvH+ZLQHWZMBrPHz09Ognu+DIg
GBIs4IX1ZX2tyZYPxN1+TSaFfTeY3iaV5FZZY1DI6/ZDd8Q+LmGDrLOMF/W5hRol
L0AEeR54S/Q+1SN1UJXIjlalTlrVpMokusknQS88My1PtoQELQZmvEFdKhbGZSv2
zCJW/jR/+69PFMVCn1C3TYM7StZoTxDqp9Ggd4wEoXGa8bAMKgp+nZHFXiOYZUd8
nV8F1qU4ZBWYHggkRXPJ8J5WnA8L1QMOKmibxS4Md7IMQkVHsprXuFXl7d49t+WX
bW0pMs2tk5hyl/P2AUiA9h462zsZHACV2ATfyeOvvCnvkxSS16tGAwVG1Ij4nA8m
7AcDKazIEG57fZ2cDvuN+leoXbufhoOO0tWqJJl50BsYCQuDvz+m49PGTTWuCIF2
bdyKUY0nQQQvAsYxrxCI5//DVFkPc2icxyprfI3TewX8EaCcx8St/J8ZT1n/1xg3
sKgCLvu+17M3Q3XDCkDQaNwap5q6sS9AirQcILceVTkImfHXuLXrOhsTC1m/ZveM
hC3kmfTMbNBbDIkJqk74tjTyL7V+nX0XR9Nbtsf03bT+nTjCdRssHwZqtxh8vyWo
rgLQQBImQFntOkZTxnfhTWULAHENppgTvQjwKSMEGRgepqxQ5Wgg/dIkalC2Vohd
JepVRdSRTaIdl+JtO6VhpRdEgw2bNLx+H9oc2qT3PaUmMewfMFIU4jBdqDXFftnF
xTXruiDIdR28iQp4ChgMMO+YwzFb2RTns12wSF2trJN+EPZMyhVd8IEhGHgt/INB
w6KnGUoiHAAin4xHdfHUJHSxo+nR1SOvfkimfR5yFSFTsA/ydj7Byn5PR1wtHOUl
d2pe7lzY0aVSrtuGemDPoJaRESnUwTbhPz+u9akA4Ll96WTpzYCgkkqutOJOeb+g
GySleN5EeEAUt91OdAUYWsoxAQdrEt7QJa03sZZF/KnzLNSfer/RWgi/un5bBUT/
Nj+pGFPGd31s9zkaWt8jq/27HQ3NHZze7RDh5DfYoU2tNrT4EkMh2kluwIVMdCRD
AR+S1vvS2asT899u+Lf2owZycuuax93gpPz4DFxyDk3zzBAB9CuyxGyMm6W9fbiH
2bhBks7ivEqIU5XZsAgWks5cu4qRzp/3A4Fk04u4GsfM/u4B1M7W2S7qTNCqMS+7
CQoTd8x1UiEOmq7Fe6SKYCXmXfd/91/cIFV89wupiuVN6EN/5JvUJCgmVvetnY5Q
QC/y4JE/YePt+HgMpvGU6b64gcKralo4Ku5IIk6hWXdZDrjp+23PygHRDqsfWgkV
ABBWvtHKbpPHV1E2r5wyUaKXwTYCBnfab4PpSS6wDzGV7N518/BVFek1HNv4pg3H
GZnChXzIRfE8eml9kSPQM7A+KvVPnmi6corUVY0Z5m9PaPBCrB3Q6s6lHZLrPszD
fGUV4vvVoRafu8hROGPwnebmTS09zld+616nxl9Dw7FoB2HUj72O/I7gUllF3w3O
0a3SFWlGN8L5j3pHYKJfCSIBZod2n1f0hsPLg7FsOCP9L3OlF7748e5JhdA5sB8/
tFz5HP4qL50diftobNGvhHV2GyvdfznOWnNH0W+6exzZ1fNo6sMphOR3yhpKEC5E
VJ7cwvR/1ABf69Eep/gVvnNeSJ/lJ8KMuvwwpeialuBlLpNI07Bp8hXtPvTbfZDi
aF7b+fXVG9f0kF5bqHismUrsbf+vksYKg8+D+wP3yTI1A80/QCbl3HrlGwZRkPjG
BXa66O+n4DnDa56wxfzUIpZwJYBMiYi5nNQRlk0ZkDnfzGPoappIWjHkILAnDpB6
jwBhFBRPfaiiJTcLKUN3tJxs34AXztAXQlOO/RIWjPV2Ybz+qxPr7K8ScGzyS29c
4YkJ2BvXisHiVbbut3LhWYUxLQVhnD0P+d/3kB4KvOEgD58pnyv7BZELyG6/Wtkc
lbMO/hlzu3f/3SFjuzHNmppcQ/sDvHL66v6jJZUQXvnTA34fWXTQrEHZk5XwDbZ2
voN5e43llbnJQPsgQiSMiJgeqVITESz905od1ZbNZGnIejwhqpWQlGwnKDSynGLB
1Nl1RGii4gfjZpsqboSggzSksvJ0UAotUZKGJztCMi2U6s/rsIbIrB9dnU4Zw1tE
DVRZd55KEftySLTsRiSUPnBt3hAGpOwPuVDyOvjJKw5D503YCpaemSi+Lck7AD7k
kVR6Z1QoCs8CxIZD0RME6TFbPZaCyrgkB0MX6Btz4MYxV2ET2fzJqktu922MQEZt
V8gicl5Yb0Ersfmei4JlDekiMymvGkfbh7EfDBSmTdXMzmiPQ+hHT+Z2DD5a0s7r
dKXz3M+t4il7MCRXNzKFJheSE1kVE5diu+47kFgxARCTwh9k+tfRkrWY7sbBY8w9
st0bdAghaRyODujyligxjKytt45gT5pe/2tF0scBv844SN5rM6TTTwEkDLGylrUX
URewN09ZWjIsljowfpkH33a3Jk3kmkuZ2eUUNBy6Z6waBVYgf1fEP7PBJ9i8s1jM
C2vS9JdkdnYlYdFw+qboODMB7h3BRzusohJptmPFVd2cgIsjuo93A0USnrNwGiQA
dVeWX9COR1ucirJpEOJBVHdmb74HQ6rEYxcQB9ApnIujmKZbuIrYTk7oOVnQoS6+
pwuVf/R9PKB3UlWmi9x/KBbPUrVeHyVOTDTOp8jEo9grVNgXruc/MBF5WrVvzR3Z
qNYo2Cwg8klrzaueP4j4wbOenelO8DsdAzWTEN31mLgWuowsZ4SPZ9cl0+zPOYTE
j6+o9f7kXXSHybXU591TxH5MsKYrFoOIMs+arDnBGbSyewy2UdJLXrD0gMXUjyyV
Bqw8orc/jYJDb9AIYc0EaMegnMpfwXGPEfod9tH0IyQwUpnzrr8NL2JtEI5CzTP6
v4IIk1Pp7pTH5NCRJ46VK78GVdpHQviGMcNSxEuHLKqLYmlAq1T+6Esgu60JO6KQ
BSK+NuzdSI9bJ3xiLrijjBk5jlB/aC1Qo8+DS4EqNVaX2uoCCyz8HHuo8Gy91ehl
3VbE2DRbuHZgLjqYUnCWn4iciNYfZINz64VS7LEtGa7stxMqMhT/XCNkYaMk43m2
Qj+GD//Gnau5D8gAIsxBbvtvxLHUjrDodgDeIWKuZFa6VIK1REl3r6QACZu5SBe4
RB/OSuh/UEr5wQCANcGrBbxzuppPfPsrITgsHUV1T0ZTCMXx5o3/0swRA0nr18rV
YfGGKo8qKTArW4gjmd2d4S2P7bLAq3i+wJkHEloUH62ZGACnAaJPUyIvSt6yWh6F
p13oLd1rP8tGKyroa/xUSm29gdh0KGmmAn+tzHMGKSRw8L07RBD+2CoLCWy/ZdV3
XCZTX+Eep4OOfJoPekqD9Q8DPTAPlKAI/bVH9N618akCpAzS5MChP+kqXbKomxyJ
lAfk49N3eUH2BBzSMdqWc2wjy0+BV2qhzFuIQM3o3Gf5jMSt87n0IZYow/4fZoF9
3xgkJNspP2SZwgICAbizuA+00hoBIaSn+9XczHOs4SBgFisBkHrbUJwI2l4ZJoqD
7tgdEdo2cp+0hSYUsGyv1VuCfarTx18ATyqHHwtv4VVZnhnlq2nA+C6nF3UCTMt6
b0rNl8uIe22BNK8BpM14GVS/gHtAbaKvAc+LSCObMwocL6iBbxaf7f2ZTg9dFm72
I/Pq2Pcxdxf1fAruFEeyKzxagWxuLtpUyubGD1ttz33TmhlI5bPsE/v9stcHQOy1
ntY/+IilfL6ULF0utDbgnAnrWqhz5uGbYqb6UNsg/+JCAKcWUM4YKTmz8W08Tn2/
Qz8SqcdcIbxIbIcPsMqpakhqw5ia5GAw0pdBkzBS998Zw88vyHcxxYlHRNZLS2WQ
hA3LIyYPvFMavzazSXvB0cV+wuFvgNj+PN+IifZ67z6meC4MIWQpLgPh8I9/XvnJ
p59TTax40EX07zRhqN30frrPNXn7/Vvsch0x0Ad6BaGjDcIIhsm68oWnRA9gKXjL
vP1E6vDVQ+syflDsj1E8LOiM7Fl+us+OMFFpD2e/wQFYrNKvD97NV1dAMjmL9osn
rtJojhow2H5E5uinRVOBRCyhLgQtynXqqVQNyMGW5b0klsYqtrBKMJi6ScTYCOqU
FBm96nxO+TjuzkXe7THkkzCGTB84IZzOw4wop5oTAg3IXM7HJjZGVnkMVIgv+GWr
Jq/L30ffDSV47mZ+OqTC0hTa3djY2U/N/FSdtZCNvCP3ib5qCfgkNRmVKyWOi8tQ
WrfbPF0ulqbmvvmcInsPW3oTC2szw7y12aInYRzDw0fwGeyKmW84yO6TXEwAHC/k
L2aQVG6fDGwvJkDrlM1pgLtrm5HhScmzDVBY6Qq3q7WTcPwrxmOKtTJR/qI2lBGf
JHat2m7EvDvhGFA4ypOp38FtvbaUMSbzRKmqjuJ8dIJoO23vrQ0tUkA/VWZkF1xl
OhQ+2xqdYDicnDzhIRnKg7c7ZoiaSkTNGevY4/zc68O0I8NNManulqZef/uyn9Ef
LNr7wojyTbuh8z5IzunUeq3Nnu8J2zVmoc9z213KFNajOLVitYlEk18vslxOltZL
TVoOSwh7oHJWDo0ZhA3hnGP2QJIl3/bEcWosG2o694N/ZfP+3zNNmY5i9sfFPuBV
b4986AVBt5RaoD+vB+m+3CLVGSffbF1TDul7VkYO40f04uyBt+9rP17cpzkD103r
YGI5ORwSNsng5S5YvZl+DUYYSzfxrb0IwelE6CKeZ4vJyZRH6DVuN2svLE2ANySv
Jhtq+IHZfSNycth7WaRwlT2CS+f9TVSY6tlDxKTwFcEwZ3H6of0UuJKN9jHHFlpc
XPpyodq3mPjd7L2rul6jZzm481MnksBqpda1sRSLQFviq6gc6PuqFYsjZLFJqBrw
0Nc4DE/2xe55rQqNee+FKzkBTPqXPrC/u3xol+1ovgmODs4EcDF7r4hLcpiwC4Fs
RnjJUG835KDe0V/+jN3O/Y/A5+o7t3erqE/yLndTQFkYjphI3U1RAV1cKE6jFCA/
ZiZj6gls3KafCDTYcozjWUdwCiznLrQv3qGmmHvApqfj1JaavXwn0+Z0aSaLVHXt
micnbv/XrVPbkWn1b6jo1EVKM6SHKlnOmSx2oheJe7JffzcFsEgFdoLzxCj4/Ifn
VRRICttpcvdpVREuX2+WmC9hT6H4iovY2seUW1KQOSBy0WnUYzLz1+6WMl5dlcJe
ToHfFr6vSedewt7yXXKlnJGDTAW5NGSP2jSTrfgL/6g3cvRDfq9aNW4LJS5K0hnU
AAHl/ly1QTHppi0KZCZLvhADyVI0AHoZreAUAXADtwO6SONpMEqLdtVr3wIPa5J/
ton0B7Z/e6DqpgXKDV60aj64a4NBbs4AUeqk+5jGSe+jVGp9DQx9d1uCFQlBXS4e
xxaATFz51wjJmwMM4Ce/zXxkmFClrjQblbevae7gqYt+rwHsiS3tEALYCn75iW8d
fiCbKv8VfG3mT/CfmZt+3u611Qzhw4kh2Q54B2lyYSve1ue/a4Lzl2OcSO5hKo8D
9F3MoR8JRnUczntaaUws8pjqjV/SOAN+EN4u4PVq3bWSpdKTe8TT9ANJf59ZMMWZ
pLk5juDIvwmXeyO5F13a2nKHaHR+JW0jhejKqvrg1GQkx3TRg2oC2VU3iAXqSvaN
aW8jIP2iU2zt2AsmKx4Owripe7XSsuiCIM0iqjoWgRGWUOkyJ1U0t1Gn02UKhdEv
cCGNhyANGqbyiJ1+zlJIBTA7gxtYf73mjQt6aglfvrKcMGUSmTXQWdICWTAXVV3v
cY/Fvc1yZ5DeDGfkM7/5hEh1dedvzNz1/ONlzDR4efSVdDejtUxgcfIZTPLNHDYE
7xDW0yaYZBeVtIjYIrUjeng4ZUehRyi1BEFNMk5lpOJ4A9Ix7GVBEaORBiwnnHN9
+utbT152o6gky55QRFMI1/zdmC3O1cTrTtKpHbPHVbbGA+aiG03/tx6qzIWw9RpR
J3dE9isGwuDIY457f+Pp1PGF1Ql+pvD84fmyqiuPv5az2ooeX98zLFtTwSdakojf
bYJbGfSxsWJu3BdjPyNvaeoHux2r2F9bJJXZPLd28qNgJbn7anQWChT7Zbd1KPb6
Z8BqzgqVHXShpwnFDmynCLTYORKsxoX6F1EOpYEpMX13hC5VCBcuZs5ZytAUfi8N
cLKzyLV9T7MFW7QMFV4HH9D172YUdUxct53nJhl7pQUs6WgAF/NN/H791Qg3P7s4
Iu1oqJAqPa1R+tfpOwgkDMom4vp+CGqszXciQGVZ6QTpfQCUcCfHJs5+CjS8iG5a
mrDLEMmFQG8CseeG3Ukb++XbGfbBE0WOm/XZvbwTzLoXCsajeDvW5tU+JraNPPaT
YXa0SapmiVQZjPu4E0tNh1kZK7sMCXAOuTdD9MLPf4ksuslJwEcLjNoagJqMpTjF
ZmHr8JOiVoMwkUnPAZrtMqiW/F1c2sIFbaQVQJ4w4WNfLexYbkqDubvaXey1EVjH
qmfd0BBT6WkwB3oM/BAHsJMpHL07L8TXKTrxRx944aI/iCaWMwRA+dBVmMUF09PG
TX2fklEbJ6inaYhibuCGrNEtkvtjIq+c7PHUB/t4SRW8G+df5cdBW2Juo/r3bjyq
ocZ3Lm1B9M9KIdQjQ/PnWo097DPBMRFLNSF8ZdaZ/wdWJAwgDBJR0QX3UKGZRMax
9w8dP/7z91EZ1/W5f94y2nMADuIKN6eyabe2MuY7UsVZSxaHY7XBZ1w7avPoo3tJ
c/lLVVs9K+LRGqfTl1Igq1RizsoiavLhUY3mgzkQdm2hW5bSTEji2grvjy6v+0lU
5wSyRJuiihCKd8To1g/6XtJfNVmQ2xDGyxKXX8QfJr1XqX7S+JPTO9zgHs8yC36G
HkJekFA6j7COap/k3Tq1VHKKt6j7xS+eqr9TpvHmbkq7NUW8/krtoqlUsno27coo
UbFAnWJk2zQC2I7EGf5ios1QUR5AQ7uXpQSjg0OZsw8wEhqEtwYgkK8RORV/P7j9
xQbFIKhXFSOFIQX35Hjehurp92CZym2MyJ2KIn+cNDP8p5EZYxdQ7mxdknfwXse8
XlayTB1udUx3Y5XjFl8s+NMZ1ppeMtjRWgx9xjQLbCDFgne6snKn+oAu/H5oXR28
xZJmVK8/i5EUNkxQPEquNlGDbMTdJvYlS3msONjpFSk8lmfmeD8AJAQM5HZc7XRd
S6JrdwGw6/mrh5PVgumnksK7pGlLcx97PUuk4f3U5NEAH7nQUAVUm02MepyXtHw4
ZM1q9bFW64XhoOM4gqg7bK0RC/YCFbBmxXnMJlz4AfPmvOY0H2KCEmLxH97uM0B+
/Gp6KrBKzBrhZYCN8ietQdwfcwkj2itb9d1ha6af8ICdQMIuz7ZcBnieJfAM1FW1
11Wm/jFwpGeUaeiNQFxQJumVVYOR6UNfOcq2xr9RVeVu5qYhDB6JXCIXKagPHiXR
CKMh5AzMGDgTEgsn3RucXK5MUEoF89uv8DQiETCKYY1Ezk1B3oeOtZe1eVbSdqVg
SC9u7R1h021/slq6tUQSDDDqZSa5I8qJVM6IsRGJw51IMwBeNNbRpGwpMe4JRdFt
+HV5Au03RMMvYA7d/QC6PtmlX2VZEXj3w29T28mJzFOli3se4VeCY0BImilCD8LJ
sS/nmZXZco9uSglkTp6T+7HOa2gnisK3gyo1bfkOrT9bBtIDi1EWIc3D4rkmlPBw
nzcJONg5SQXrIpa/tD37ttFXw58buSoUMbCmeFIGhaWy3gNW9OVOAwrg5aDWgpIX
rRo7sGFEtHj5lHAKoyQjXp46Io0hmf/YltRn4U0rVUAe5A19N8SidNGU4wMZVj1f
M8/bd8B6xwgLeTolzmZNHSBtJ7F8pthkDa2EZBdyo4/X4q0hq0LkmtD/nCb+YJ20
tPnl/9klibGX8rEh0EsryVeo+AkCLP600ey9hDpFMU/DGDXi5YQP0HJl3Sh9Kxm9
+ATZ3VOyjfl9+LcCQPxKIPfDwrc9h/RSXLdjX/cNZL3aqQahT6g5gTlZV/kYSAB7
r/tXYRxiC/k6FVQ+TfKdaQKI3dP5PeuM7NrKMtuI4DnroKksK+Bgupw2gGd/trED
UhJdUJuzkpbDkJO4A8fXsDN93xyLItNrgyWm9rTJ4/RQD06KHyr0BzuF6CNux18E
tkxiTPuzhnz6FWdtsvmxjKEDA5NxC96VsMmTN/yM/HEhGUpwHD4bTUEGmPcrQNkp
hPvcDv3xsYrV2ukKZi0EP6te7QB/HEjnzmP+mhfdp0C7adERgLjms1Rd1v0+G2CF
9ZjXY/c8qYqLI6igBDc+9Z3T+4liwDgb3XsKLVxWXYuhZQRqTLZ2sKr2Ch6ercNN
3mlCbd0ZMx5c/s1NSszd4CAb2bX+vmWkCZktw+ieRZue1XAweZgJ3vMZeMGbaLxA
xw6GhL5WbZ/uHmSHTebqf6SFHyTsPyE5fjvpYBK8OR5qSffvAm+KAKnuAxnCJArG
Q/qoCgwB3c2KXqNMLG49B5K5JAKq8Sx+8gSq2TT7lKo+WxAj6RZRdU125h1BVADa
lmDSbUCnfy6OmMS3aJpH3jQ2Y5H+TMmPffMOBEzWEVo/PzetGr8xI58H3Rh0Sbg3
aOR1/II72kStcd0HC0lCxCB4XzLdeZIPMW2eFSPZ3um9MubTH7eP8ikXuD55Zid3
NSeaCXav0xy73BI+ozT91LWy7sWzkpf3wh0dNdYBSr/5kD02lcIjOra3EtrXWOz2
XenFTvbI8jp/fq6jC2Wl124atyYlaWKnT2n3z7GBsYsZfmR9Wsi9wcBy5wtUnK+m
M7pmoQrrIXAsuLq3YMswzwcEbmNsQwD+jdRqYPJQO5aSNE91b6CIfQqy42nGX6PJ
KcXcSBXQ7rHSytLCaGu/e2olNECg5ASLvacH2EkZCTJxXzNYCqJI3R4kfh+Us63D
nPmKk7a3dbMlkaoOsUfZvieIf2oPoYoZx9fBjLPP7nOeT80c0I/KD3taiefrZzkS
xAOjW0xwmMJE7ivYzs6VZdGIMkDIpBlM1YlR62B+GfMzgWkcCzIUXJWmSGRyGlUW
f9DO1j6ooIdkS2fFicy2vREJImzbc1TePXY/+5V/+Z561CgBi3EPl0REE+rOMQf5
PHMCC8fSnsSULZdmFmGu4AW755bSi0ZOgXycx5v1hp4SA9TakTwJ3IF/FP7rEiWl
ksOmlPxKR1JObjmNGRq9JxE9nxzluUn8P5tPLbJKA7KlwZso66kXgCQbU5M1wQVW
2VC41cXNgJh2AEPFhiZu+jKduVmpQGYziXOZKJEjn0JeZkxVidLJDfYNFl8c1z0J
oSNQpeknWsBzD7bu1teHyon4l8xRxxAEMtfYLdmUfg/BzoZ4hPL+w6Fc7aQ8G4cu
4v7KwZSBwdc8y51/2nIpisGNoDQwGVCMK3/kYlgd5OjPEzz8sYGph3rvXZbZAqGH
+H+Jyiin8qGOHJQle3xaGQcROQoDhuksIaed4IvGfR4L7KfFSG2Nksec4qeTIIIq
JebHf61FzK4/+5t0sUPZL1V5m5bl5npWYN4Rw4uvabi+zS7jYimaIGwClY6OwsnO
17hxRcK3EV84B1g6mROZ8FSsxT+oc16mlgtIxRsO2d4xgLvN9nwaraIdJm1wbOvq
Y2yzIaa+GgcuQi1RizJwhys5hoxdERXyILVee0XwQITRqX1D1XOnErIOT+zOpUFj
gBh2cToH3ldqc6lN6Rlq9/kC/mX1DODgY8o7XfoU7ecSNSiP6vp9hnkE0Zp7oPzF
xxkiHM9TXuCFZPlGZXN8c18P7Rd3+B/91TW8EqGZ28xmZUxkSqvsaiGrQu7qL78N
qhrwWNn3LDlfn4GF9EPz7QFs9SFKC1SKtgL90v6A9e6DbZkElTgR9JuKuOjCV+ph
ht4KUNIDUZm7pvHBhJmE8ki+uYPGCvpvpI3SBAC1Uy4kEmOyl6jQNNRpYWk8DoEa
75MWUEKYhrkqMjV4We5m95QbCe7buT2d5IcG9pqVGTFbG+EozW+alSeLRqZSe7wZ
y7ZFtuNsAcSDbgC6ns3yfYwva1sZo2kuWviVxHwd/K30ZeMN8aXm5RiYJuSznsMR
U+zwW0BkrDBSZ9hEkyu5AmO5Z+8VqBQSqnVe6WIJUQeOmFer2uF7Sk3Cs9aFZZ0B
+nx/CaPEOWLiwI2KEK6YlN9bO+kFCLwFmLbjFMoRUp0zF3qg+YDU/wYVZNkwzbJO
flcdELJkYJwEi2AMeXjwoeBWb94ZHAT0lAMddyaqXlAhzI1GgLOeyjXDiXh90szs
AaAUfR7kdxlCSrgyPTBTyFGKgNscJ/sqm7LugvNNQDnZ41Xh7Qv1WzzBFX2e7J1g
5xFE4ybYHWuOpd3iF3avyv5sDpV5lLVD5LdXq7YF6HJt0WPmM6Twq4/5L4EXVhW/
8yAQmh4N5nnGjHqalO/SCfs8U2gM1s1WK2XaQ2I7VfojiNa9hRs180O4Ln4tMllL
Cqmc4aXXNy1sw606TXj9esuupUEHlvVeopdTIyMEDQLBAmI76nab0QzTst4pNsR+
aMqhWEsaeDzLLV+ib7gnpXV6Wx0J3qdZi9iuPYlFAuvjBQblxlzDxsqHN9QLuekj
Ajm6bACG/BVkhCMq+XGwvqWHNFiOu9znmsJdxe/hoo77S4yleOkRk4jKi8SEhYd9
PqKFlkQhSGu3uGLzpUrZNuTfFSzPqdFWCR4joEShavmjQQYLAG+IToWcwZnO8OeN
PZLRH0AZ3mUsCSr2eie0P6G+ULPEkjUBzOLi4A5CLQ3SYyPFuuixuPqYyE/rxJ4F
khKVuJhZeSlv1hxJ2u7DuyIEQUTHvidpL3POYB4U/mF/41c1BRjraFCQ4vdiaVcU
ebC61GVfXajauQSZwY6+fv1aZTbGmWXl+M+ReuQuQmemBfgCv0rf2rFGTd3JsExZ
Lb9ZFDPfumRdizYY4Zk1Wwp94Q9ZYXOyxd+snLh2U5m7Nc+WRB9/gO3MWVekJOzp
J2PSUwUzQJ9rFqvQKmSPQFa9dGyCB/pt/7UIKR2/Wpi3l8nyS/hL1bUcfU2fH+bM
zDsezkQIn7O2ic9fEsl+wMWa2FmqWXM3Y/r9Cd4fdS1B6tvF+0eJU037eZWaKv/Q
RLYC9ee2ndI85pQ2s8rrrALFKEmI/oPzCThgxsSvUVQnVQ7EgLjYNdwSfKKFDgx2
qzITGDJfSmAgCK0kDcbnMXHY4fAaN6shv8M8DdComykm0tUMgyAgGKTemgL5oSpF
t6ATMgQCRQqJGJwN6/pPa6rI2lDsr+DuC/43zyAQ3HnJ9epbscQN+/UzNRYTPiRq
YHpt2ug9PvJhzrzyvFDjIH6PVGW1F8bVgmh+67qXRc1d/eY8695lit1GBNfS24Jw
OoW35XqvwVta4DmBAfonFTyCdxfHYs18jOjcigN/evCextZEx4lM6hp9zStBhgKq
817Q6pmMLE/Z8wXI8LXW6RR6zH4tFicv1ytknn/Zthy1MTQ90T0wy1gFChzxCbE3
arYkcAovp4dho1PdfbD77tKEZHkmzUTdjnor/YuelaZ1l6EnT+PVUsr+KJ6zgrm3
fz8AcGhcDyKYrMDNigX6mov9tTu4+4vsq7MRqFJ6DJDwhJPpUHT0OVXsEwMbpEYt
Z1JHAHdaq+TvOWQXVSHGb3rjk5Fle3QUODCL6U2YZR481MfmHoyM+MGYYZmzbVUv
TLbZIcm3GMqfw12FNyb81TDS8AzzIkChPVkmvPCOuL2dl3D5+RMG7f12rcI2TO3Y
D2Nx84k/GWtzE85B2Yp/8q5v2WUGQv0kGGf6t2MWGwjqu1JA2mku8ox8I39OMaDi
F4ijFCc341pGPgmSbtr5WZneoYrd++jF4B+0PH9y4PA+pah7FUqfhuoCa8yAA89R
6j4SdvaOVDVUhAhGRH/n6i4hn0UNzSg4Yv5Qk2K2yDm6XWaNBEgB5xwAe/m3voVc
nAK5yx3eknUcqLZr2Kus7Djf2RmY10qCZIpAv+wbWxDNk9IUQT6LODpn0VthsdB5
mRz7jTvp9Z6Vyp2Z0/6YJalLtPMlEsWR8jPA6Q6JdUVJZ8vVS7+042oN3rpIIQrH
2r38vBLoFqbHsm66AvIvkazpnewD36Vew4IY6AvEQAOgIbkJcMNKVWcH6gBW70zs
Fdh1GeKx27oPBthWagqGcdj6kAUsy/Fjq1QR98p8atCODShio8ueZNwAlMvV9qAA
UwQVvzTbXgkAUxgfic0Er6AdmbhYoNMHijshc9S5uJyRqeNxpRA1vsQuLx+YrNeH
W4unDsa51KDJcAyh/vmJk1j1PO8tTHbggXDvwy+MoOrYuzn4s94P0ZUTuKcJCP3n
oDxeV97TrhBvfpDzk6Nvp0oqiW9oJOWr/kPkhkwbtCevlzloS9pKdcpxwPp30rvN
8VZS6QoCLFfha4CMhTdm2hEQTg2ExxgCGseAlVP7yccWBgGE+dIgAUzB5MUMpFIN
uaO03EQ02FYGbRuzup6CqXEOdfG/1VLnr+58N9V5BtXMbjDmNqrY1SwR9hC/ighl
XC67muoPLyNqUcYaCZ6M2WaukFCmfRZ3MgwX1befKOgpWXh1ur9ZDNPdVHJcL0Tb
PcDNZPVgkntnVzIy86RWB/NZ5q5C7pl6pGyCim9Zm2r9PIi0gKBUamFjGo6/gOcz
LV/UjnZbY9wH6NRMZ0gghpVPCmja7+6TW6brJa6gcM8OibV8YhjTsvVyObt+1wEf
7PC8Lj2egETv0j3ujvSeJpsroXEedOOef5uTqG8pJO+8a1iUvXXXuSdAeySYC6DX
qGs+pY2GstMYmXy7Kasu6J+014CeAGKd8xZ/EtZBYzf9KUw7xLMtqwCjc/c358Tn
n5jcXPxbIxoyREigUI3yUii9r7wLsOBilaG6+l6tMt7kkC35BVAZC7lQHVKmOJfM
FpqUmMYGTIbB0waoOmIqn/yt/IKDXMSOPL3k1ubjQXtV+QZmBIaCap6q+4gzYb6o
LVF4mhC+oV7hbkjdfMufIHbqFR8kZ+rtdOldoxypU+3Twcjig1snWjzQEAo+iGQ1
VJhfxLNyjyHF4ZU0LrQPQiEwanY3YH5QVPW8ojHEA1vBJVh7enI/Rx7+6py8BOV/
e2FeLlHDDkwyP/IZVraWAI6iJ6NeKdJCWbGbKuYxd+idGqfocmm+Z0lzPJD+llB3
BLPiCSDGq2wl122TaiiMQSKMrQF6vK41pfx08ryUvhhcafJxN1xaVYjLbCUd25Rs
h5XvyyLLc3IndQdGYAGDwVoHKFTBP66dAVFkywi1nrLhKwAquYyNBG0XXc0h9f5B
yUvlyXOuWPEx4WlKvBDayg+4cXVifRMb35E+rQdq96GgZsU1G4Fp2Tak5kscukcs
2/WFBUhxEg/GTInhWjhIMIAvQhXzXntHmWoBUk5PmsnjDGA5bxDSMPO2d87G+s46
hYELKTWIpvX79XBlCARewuiBM011vR29L3MiZp2BqFD9drOWAVb0O9of+72XvEqV
ZB1HMCfHUScTRXZbuCcRgXsoe0S6pW8Q5fyIQcUyqPTBqLBvD5PomaXhkkEPA7zL
p4GPqCwH53H6xQ2Bn7YGVmsmODosp6zXjrWdXeLDRzzTf9gO+HZ0kb43CLZcU8eM
CeFDB37QbxzWm3SQ1efRYHHrPPjt6ZVLgUqTo4YeiMBwhQCR0SbTrX0pD24+g6IZ
/0OErYmYRMkSwLBO+eUj0GE04CJwR1c9RG6ZwEW9ZqlAmS6DDJ+0MfpMtOSo2kyT
7oAPhP/CEPl8eKF/WWeR7RbIrkSy3JYtuFp8mZBmZdqC2BnnoA4Y5AF81oJfc3Jl
W2LbwDAKkvpDAXLLXKCXSNxvtfG275YlPxGs35HyEAhgfoKScdUFyiQ2MDE+wD10
WF7SrHex8MrJYachdbrJ5f4v5tFLIA/An2H1prdb9swzh0/96CKwCNbV+YVKQ/qk
RJFDKf7m5aORZ/v+m7ijRzVINzcNqPk0iygVXat9bpIGdNaxyYBUgEwzkDh5VmFU
JWD+M9fasWdFCR98SuWOF6Tj5gA/R5Tws1l0/A3mlkpYEWFiF2B+ENksC70qOhdE
NBCEYqpA6haaEf5bmL6Ps0mJInuY0FKaAf3UJWBwGlr4Keo//NTAEnQoIrBVQTxd
2MLGarwkMYu5m1kL+PyfeajpiQQhElH7pQryRV3U/kHXuNIAiPNKCxsX+/ceJesL
orZGwOV43WwWs8V1qHfCTFY3ZyVFDVrsoQB8g9r5P25IbOa2yG2dIWABUK5IiS1v
khFHtYCSJ8OQoVhgPMkuhsL3LKEUc5/5kC/E9HAuFHAlxNp+NtEo0LYtWM0ZKrVO
rqQk7gstXPBrtlXK4+hBIXRlTJKq+A20CJF5N9xh4XCB89zaady5bTp2m6SGaqTs
BkyivkYUrAsNOQesmzYWkKafmNuW8KaAwIAw1RCuSw5dR6NeTR7pGiOFRk4woexK
LzUqMvHLI0H5rL9oxkhcE8/0G6BEgF2oQU6S4TOfAIznmLpIJOXDp6SihIK39ZpL
tEb8X/2RPjukyBSfmIO7Xqab7LnSCcmQtorNBmR8YE4LxmP/6+fF0RB134CmBdT+
cwRNcANgOQvTJn0uGH2ZzVa9ouEx/Z/ko2gnfQFdF9LJgvyQ+1/g2awdIdjBMN+5
jnQd9EVFSr/L7MX1ncVxe5bCn2Fa0Ba72yK3gKnU9KfMThuY7iMIuBchqVKhXZpG
Tth5vsbXf6yEzhEt76VSSOQZqecfUsrJbcyp7T/UHqU1SBzpzDOlkGpHJpiE31mr
l9xEJbEpZwhtUhPBSifkbMpVOEctNubxSrWM2u3krT2F8bWZlUkXgZY+gCxD+SGt
7e+DRfwRwbGy0+++jCoHpRGoDV/wfsB2BB0e2xHq3HbTsWFabfSQvVREFL1KLBoB
aUAiArvopwwKR0PQ3+vyXPmZGFeNjxg0ZT81OFISY7B6pW/BuXD9qhQGs7jH2IW5
mnE2EzLjlSIVEzQsCuT8/5E1fFMsPrhN7AtBmW8UtOKluIJVREpCZeJIQoH5AZWI
wPbctm28HSwhpGv2zHZ26Do4yJi7jYn9Ps7vQFqxHCjLCOuPzpdO2xX2MisxZ4aO
JqADkwhxUXywfy9U4pFDx2NvHPih1NbP2cbL9dRbHFm6LuxUsyU5x5/FPPWndZjX
ajZ7jFbh4NHga7XLVULdaHm2dQ/cG4wdVgzqG9ohFXo3n2VHprWkqZEyT8WXCqss
FePJZbPM6GUYMWhEw7UQsQooaau4+vVgBDaSIPi5xZC/sR0OTkusWlPon/eXvYQR
vJqhKowEbtLSdTLRBSzvCk0nJ+QQ5ZG+vPYYRKgQNsDhEJOjb5rUiYjSlzuDZ6VE
1C+1SWYauPP4eiRxYTKpAhnDmOYsrYgIimtKwLSWITwDcIB+NUif4OO16EODgZeW
eKsnvM4LUWreTdGqGl2aESJMCvKkptJPFW8YduTX6k110uOrt+3e6onNPgyYM+sJ
tu61J9HNjguW//Z5G2fe0EL6PLsdcGcj212VEs08HcJeYvZjSvfi+gwpBPs/kp8o
oZMYt0q7fqAfw7PQYk+nrsZa45Sznv2bjT5gtbw4HARrmdhFdsLxbn7dq+xAo5ps
eZRAJsKJainsN47jfDXxb7onrOtqjR+p4TRDaxZwQX+EKIQQ+lZt9i3M5vdS/Xyu
qoj507jxmKYbETqA6MVYoIAPPL8P0BXhGLHBG6M4dfuIC1SrWPDNn+upwisF7QUH
ayGVhkx0TwomvbV4L6UalI/SRog8hB87pAYhVP+nQdWE71RiD/b8iQoxSEuTxc2A
P6sfsYzy2jbRmquxdL6nL0A6Ax+K71yVEiAvEz7jGRFj7AoSfYSO6zxOvnZ0gM/C
YTfJ47J6YXBHoqmPJV9N29zrxh3LULm9egRKZdUIzRYPPwt4BAK9zh70RdvvNAs6
eNpPy8kFXTua/MvK7ETnLongVueKx4UC/gHtYQ1db8ckOXJFh01Q/ooP1PC+syXH
9LuheEcjaHZ5d1yYDCYh64S7RpazExmSm8q9abdrh2PRhBL//UUKQTiJxp3lpGob
6LpvwOK17JqZTJb/iHs5rThorK/qClGs4w6ehO5SjwsZHNciIR0dXugpubO0WW7c
b18B18XHW7ScDjk5GBWHJBoXCNFqjwKOrwTM8fC9WefEFV3ZPM7RsztZ5ZBp6oT4
Ymfj056YYA38ZW2+s/MbwHitAIPymZ7i4rwM6NXOCiTwhEEPPanIe2gTegynlMm+
pBzXqdKNCsO28ekfVtcG0bNf8I6IZf1zjyOIniKs0JBhpLq8I5LcRte0WBOb+b1W
i1VjwFT7IbWjseGv14WwkR/d40JbQAu+KqHnNI75oxqw9S3pzfLj8Bc8A+RzczEd
7SVtCM7p0wCp1xaTzzFUMx2jcCVjiACksCmHQfIapjFboTmbmYVYTOE1FowWlIwQ
H7rWlarxq6SCE7fwoe9+d7wVOIWrME2D9w/th3Nr7QKdnhWsLV3HavuseWDykeHQ
NOEdi2EEcdMqWdJR7V+eEZ0tW4vXbvAtPmHc0awZCxsKuFfqfYRX1/V2Z8a62UHh
1yaFatnbGcFP2dm/tuAtFw2FNSsKe4hWvOiBQVoejb6adVQt4oaFxsOVbpv1FGao
3PofitPuzHCLG/ad0B3sLt4jZx9D1evdwncX47Yq4vB1X5EV8rcUgectwqtmdVmC
9Smu48B1A76Rhww7pls5u68hoUjVROM57fQcv0l/Kn3z6B5+UrgVX3kqI/UZgzW4
Z00cI9Qyotk7w37hsxbeADvsjNfVWszGP1PIKN+xChB8gvt8dn0DDm/aluT7rvz/
fYRiGb/9irc7kz8TXWknQrR/AKDTGDG7PDw4BfL//T16UA85VuCM3+XBpR2XyTMZ
Futk1kweg2oggVc9vmjRZVMmdLsqxT02rhhh0JoFwt8DxQmyjf3zTBTpgUbdPZ7x
jna8yCDku8w61tYcN76AAMEfH8zKfOQm3jkfkzHx+6om2GcyZSr06Io1XpZ6ERwB
9cSHBm7F5Slnx2gQPIh+WpvVJAoDokAXRDp007oCCPZ8iqTaEaWBH9UBb7EUOiQs
MugHb1FTNIRz3xQUpGji2wI5ZeyL9ReTFsEMnSGUQL+dJs7mCQjyXGEUxi+toLiG
RVns9UfggTnriz+Aif3LIIUKdlWfonZFx8A6gJMVnA/8NQzTLb8kQg8r6y3opYB9
PygroBY4w3q9Xb4s020snSQc1SqW61wGjtjJDJD1TYjGVj4Ju4PqMB1NrkCrw4C9
4xXB3KZ25BoNL47ndF2GP6BQA7yuaXvGiQ4ZxUaOvBYHxnzc0lxrS7uvU75iusOc
cEXk4257JDjfquxTOSMXbw==
`pragma protect end_protected
