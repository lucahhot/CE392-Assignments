��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{j�X.;߅ţ3n��Z�l.Lp.(d�0�:'i�x�6��dx�N
�z����y��0p=ԲD�l�A�Y~�c$x�tͱY ��!Y$Mˣ����ݪ*]�0h��^�����b�osH>�~G���o�,�,O��:g���s�D���w+g6� � 1��G�� �ߋ*��ȅ5*�=F�i��RVl��Q璐R'�BIz}��/��O54ud�A�{p �`9S#A0�kS���г��v���c�}qJ��*{!�H�Pr������z�M�2�'u(�i�ЁD�S_.d���TP����h�ˑ�̔	)���X�{�<�iQ�����.W�z��������j&�ע�݆�����F�<I^���#.��W�چ͢���8�Rڰ����fW�?� y�d�Un�z �4��vVHt�^#t<��%[�fz�����R�H4^�[�1	�i�Μ_�X�2E�����c�k7���Fw�i�&��W�e�׹���5ħ�`�M���ם�7 >D�����$��;����\�|�~r���J�&}H����2&��m�%��QہLDHF�T�c�����S��5ҳvg���Fl�{IE��:��b<��3��.�u�"� �՗B-tV�p��<>�v$)�̬g�հ�|�m�]�+'����(
u���ҚyY^=z�Ҁ�K�:А2���~ ��0]�A�(�q��^	I�5���9�T�͝�G2�{4����7J��P�K����X4v���Ɓ-0��2�!zݙ�Ni��yI�^Y�5�ۅM�$ĺ��F���m�:���^(�)H��) �X~鼒�\޻�KnH0�C8�w���ջr�17VN��h����:��|��C��~��i\�k���K��g�|�Ɗ�6>�f�j���e������˨@���C�85��`Bn��6>�A�r`�4�!�ذ�tf�ό^fLzni���a��7�@�b���q�
q�Q�2���}�P�X�xڳ_t�ܷ��(@MsIh�`ë+�o͟5e�_�R�y��9Z�B���k��)?8ʽ��2U*��CZN�H�Tx�tp[��㣔&�4mQd/_�T<r�*u����B�O�� ��~r(7�Q��PO�_g���9�"�S j�k�ekA���I�}.$���C�P $�ዐ��4XF�قǜ^C��g&������u����i�q|��I;R��>����Զ���]3r��^�zi�,15���梈Ϥ�Y�C�尯�7C���y�i�����~��S�vt98��fv��&0$O5�:ͼ�/��WbY�_�����m�^�y�d�p-��p�L���+��D� }[n�Z��y1ҫc�Ēա ���C<B��k(�g\<�Tr���{=dC5W}`!:{Kcŵ���yo��@��F�F$d���q�.��?�5?*:~�	_t��-�3�Lq��gW�R�YH�R�S�"I=��o)޷<_B�eZ_��{�0��O�妶 r$>�E�JF0e�R�6"4�6�2�?�p��zds�
�p�h�?R�*�l�4���Po��p�PHi�1	�h�X�Կyu���]�.7�6�[���YV_	��5Gq�C�֌<�#X���-2��Puʈ�tv����̮�fj���w^�&���`Q  [~@X��}�@L�p�G ���;jN�����X���#�\	��'�_�QҡAM#~�b /55��U^�Iu�|�j��d`u�Yu(��	6�-J���*�<yB$�,�+�#	�1>m *�D��]����|J(�4��f7Y���l��;�� F��-ʽ�7�:`v����q=��9�h���	���A@�3���۬������6�ή�
#�j.W��\�&C���eo�̟������_m�����3�+�qP�Vq\q]�w�`]=��@�7N�-�1���:(d��~�ڼ(��iQx��{���<_NPD��O0�q}���O����bZ�#�٠{=�K�)�0o���̰V½��p���rE����H�_g*�������0fB&<�g]3.[�.i~�z��pR�k�s��jz�>�6b��)��@�qlΕYK�nOْ���y-qf[�0r��^����:���Z�r��u�*r�+p�Z�|w��0�a�t6�}�&�A�<�����F�ъ����ĿŒ@n�����1Ro9��f�W�䴑��7�D�&e�-�����^��'$��Yp��m�+΅Y���\^��!�^�~g������m���~ٛ�k(�4\��e2��X��Gq��u\�����vl��#B	'�S�*b���������q�6�'?f@���O 	'�ǥO��RW��[�1�p�Zz�N��L�N.���|:7�ż��w��+��l��-���Z݀��9��y��
Q%�Un�dt�Vʳ�/�Z�M���A����l+bVVm�{C�O��8;{��}`|��ey�؍#�//b>[�!!�=Z��}'���{/���]M��l)�g{ղY�Jʠ�H��r�k��V[`g����R}�����{i�=Y\�ʾN�#ϒѕ[(�2-C;J��"n=�;��6������J�1�-��^2|��M즀�!����&y�N��O�)�M-��]MS(Q�n�>��Tsc�Ξm��qYv����#�E�N�l(8��@(%�3��V���P�{`>s���Hbj3>1�D^��
����6g�Z2���I��GQm���PԖ�/y<a��m������%���Jo��w	Q�$�ϑYd�ώB3�k� o-����*�-9�2��<��
�y��4�YF��P7�D�F������I�;�<CA��x-�I���g���w47��L��Nr�g�نP��ړ�3D�0>C��fҀ�`�D1�>R�ն�aNH.�\ϐ���r?�,Rd��������x�9H�����yn��Q��G�g;ɧMxn����U$Ef�I�Z=\��j��3���H9�S�&s�l�eE���P��!ߨژ��W����M\7d��d�ʭ����-0��3d?�V�"T�H�80�T��?�υ�lJ�&j��#=����eBܷkI^�V����\*�GP���,���'�$�vo�@�I�s�Y��גŭW�*�8{�L���sY�W(�w,(�dc�	����Z-98꼭`�@,�O,��Z_�|��݅x��I��#Z��A!��;���獬(s\7؋�]Bj�hSI��y\�<,�J۽2
��.����Մ�q��vDt&N�R�>$t������Ԫ֣�L�+�+7 s(�J!��=L!4{V"��%�ft��J��PiW=���sGi�L~ L����H�e��� 	�`{��D��9
�r+�p���x���a�5:~Q�ƪ��V#�Ta��]�v/�0�}�i�bw5ػ��fN�u��=1�I`�K<m4���2�������ɧ
��8}�� �h���E�!1�{=��i�o��ڋp�VH'�j�<GL��U�d`�����
�23�}G�1��y��44D����IƏICc棧,���|
�$��q��0FԿ�·�T^���Q�Q�L-����M�}�����a�}�d�.��NUB�%�%]p0�]	�L��K.�M_�P�\�7�Le
:�	ˇD�s߰���<L-��P��gO���N�Y���]P�0��h��C���A�.�㬺�x�v�H�;�f
�.���G�O��*�?���0�%ew\fa�F��ٽM��%L���i�@o�[%�i�i*-X>6{X�q#�E#�����S7��Xd��7�{�w�s��m�PI�*E��U���j |�H_������]��x[?�M���s)`\颌�Q�'��Sȭm�e�����>Z��� !��_S�6xI�?%���9��	f$+^{�	�)��ݰF�%��\��{���L�:oϠ \�v�^���|�+��}�o隠��:!�449�Xcޤ�t��0��
��¢)%x�^/�����~�2���GC�5�Y(��w�����B�'�_Lª<��v<��!Ny4�T7[A��B�;l/=ۗ�z*M�@��ރ�#���71�����ًḫ�M��g�u��2�0���x�v��3��ce��&�� ���WM G����F�V[�"�<�w�Dd��ָ}CD���y�qx�Ӝ�p\�6���wi�Q����Mt35Fz����$Ki<_�*`�"�� gڿ�h�H��7��S���NN9��(47T�Q�HX
$|�/a@�EZ�&P����x�^��!�A��z���_ZxG&������0��+� dO^�Z�a�"3����!�����L���e׭�dͮ��K�>%�l�9�ٖ��i�����Jc15��O�2�*�)-$�ԕF�'Ź�_����Hmv��x���}�;%:���!���,�����k�����a<���ƃ7.\p�y��w��2�+d�Z��6�/)>E���_��d�x�(�Zw~��ٴѯ�/M��IT���j'.���丠 O�<�y�c(0��<��o��s����<U$U?�ϜB�XʛBG����m�.q��ݭ,���Y�mkDx�%�~u������(eM��\��%���!�%*��$�G�a���1���#I31ա{�[J�y�9���a� Y=	=��Dfe��	�e��U�ָ��>"@�N0�?��;׷vr�nGUt��^X�k��L��lN*i��\yӀS�"�6�4�r�$X�JN�2���,�8_~���!'��8�G�prӺp���C3�2QK
���ДoT������ۭ��|'��}����u}3���ME���ʎ�w��y�����~�g���S�y�'�Pw���)mx�o��l��6�Ѐ�x���"(5F󂦹e�2(��3d��#(#���.טXeėTi�ӔBn����h٘v�~`%A�(%)�� ��g5�Hu�fO���Ga�ގ�a?�`�t�~��֠/,�@"0����#�H*�r_?�gM�r��;�Ǡ?��F���c�++�lY��g3a�l�\����c��8�GL��*+�S��zYW!��.�!�Ї�Xx�!��Љ6�t��g2ށ��C5.{��#������hn�!� ��7�I��+�=�B7CtU�L7z�4�j�RZ�Hd��oLr��B~,�n!<�J��@�ɣ��t��f�N;�\��[�w�x}�����RA�����|�/U<&&�?�|���khg�n���s,d(� �f�;�9{(sI����4\)�~��q1]K��F�O?�w6t����3�����&��/�#�8�i�,�Y�5����'��W
�,Q@'��O�M�k�9�[�E)^Q�ߧS;G�]����g!o�\�pq������#@$��@i
,���N��*G����¹7�.��⌞���F�P^����������8Iw �V̚+)��5�����	Nuu��;����j�f�d�<��'���ē�b'@�ϡ։0,ӿ�GxD��V�I쩉}�a_8��Y'V�-��M TT�M��9t������# ns�t��d�Ȫw�P�-X{�6���o�G���;6��8"ѣ�^	>�Z|g3�@��jEڿ�KX�- �)��c��X�_D��!ʆC��j�<UA)̭��9О�uy�&�~���y���D<z�ٍD(�M$Wx�>�Z5l�6��ÃZ=���y��HA��Ra��e�f��I����Z�Fk70��M5[����4͜,d΁������R:�a����A�-'s_���A?Fy�FGJ�?,��歠F5�6]��/��ö�Y�=�T�l䑯��j���x?n^3��b�\6)�2��Η9mޭ��̋D�*5��$D.��.�٪����O3*$�]h��b���n��xҐ��+�|�Z��̮p�M$�y��Y�:��r��F�_T~Bè�iRBC:�������Үc$ ?HH�CC}���N�!�!KYb�����J��5.�Kc90�T�mT?O��Q�{�Y'g,,��:�q�}k	�~���m�e� �g���S��A"�t��<#P��\��O�f�:�R�?�s����M�G�R�I�с��JbW��(����Wg���<�}����I	�߉ܹ�q��\��5A�U	��+]\�+W>9}��N�F�u1@�a�2سUETj��u�'�������PuPa�A	Ȟ�gꋐ:^D�� �}��(V����w��E@]�պ?�b3:��-�����X ZR�0W����_(�Y�7����vg�A|�V�Y�zX�^��KM��e>���fVe�Ө=`����M�ehdu,�*bW���!N������Ḍ��-/��;\#F�/Wp蔟�L�i�9�;WKW�K?_=�S+�e����K?N��Z���8��A��R�G���e�㳪�.��h_�m�g{O$a���ie��}��˱S)~�<z��1;��#R��1�h4��ϑ2Y0Hߊkcb��h��lɩ ���E�o�)9��i�d�ሠ,zz���(��+/�LX�D[Y[�g|�J����������",򑻍�ְ�`)��7Ԧ��� ҏ�a-%l�9R��T\���5��0>ZѶ�tc�B7�N#`�C��x
�w��P��l\ѷ����xR�3�-2��!�heN�Ʃ�����Z]�?h�l\V.����	a�fjr(�tGx�ƟZ�P��(���㒦�N�B �V^�D�I�^�%-�
 ��� ����ﴄ��=e:���,�i�s<�!{)��π%k����a��� P���_35�P���<�@�~x+/����e�>+�d�j>���rڍkN�6x��[���S�	�h7u=�l���ߧ��D�Dj�#��K8�q������9��@ܑYy!r�����ZtĂqPM�m���y��X�t��Zk�����R�P�q������0sz�U&�]ři���|�$��9]�R�<�+bW����D�q-/��<�.G�^Hl�@;%.��M��z�g1̛n/�s��U�8=O��s ��G[�ª��Y`��J�Ҁ����y6�%�;��ve��5��fX����!G��h�=��Z����P�Cȇf�~�W��'m��4p,#��'lM�:�p�fC�̿�s���D�G�_N�?JZ�PʦA��t����m����MдU����^�Е���Z�Y��2I۔��!Ji�\	�G�0��HFp9@�*q��R&N�4��3�n����0b�ɤ,cᠴ$�k#�p�{�o�[�#�5�q��nd+>1o�����^�th[5�/�Y���oN,����SbK�1C�����H�Y7���5�OO�F1`:
�wA�d͒�ː(U6�-'Ѧ�	nG%�du
Z��oGc��3���D�6��h���+opQ_?Sͪ|G�J�{uC�d�;}���©����M���m��j��@>N��+ή1�TN�e����O�K��K[l���?�B�QVgv�A@7���/ :ŘҌ�[��sG���ݍ�'�T��⸧�\5��.�:�3*�������Օ��͓�Pn^��+:���h>�'YW���ʙ	\L3!%p�������_lC�נz:L�
'�}L�Y�p���Yg�U���X�B6~M�d�#��xob�`�eB��"WU��e᠙��Lh텞�=��
�{����ea֤~7��H��C���fn��-������%xm�ڽ��?�����o۵��dm�W�$�WB`������1M��x(�E �||��@u�d��i8�_I0G�ŗ�x,�#f]G���W7H?Y��*ӹ�,b�փ��#?ot}�-zhuĺ���d�އ��G�l�|[L�����cj楥: G#�-7�����+�_繗D��a=�8��H_��a���=����yy�*����e�0P�T��3�?�l�Y�]�Xo�z����*����9�<5
���@�0G]Z��2�ԭ�
vj���u�O���b���[�]=��g����v�4�-E�����mS�a����U��M ��@��[��J ~���_E���t�%����#�lޢ^d�������ކ�h�����>@����Oٙ�>��Sd#�����X`�9��!Z������r?��]��k�(/����F��E�VA>zޱB،ˋ�K�t^� ��~���!�[5��DG���6'��^i��=<�cPC�es�������{�`�Y��� ���x���d��ٹW�4���7�:�o�5�~�u�h>�|`�T8�M�+)��Fb��5^!��ҭ\�D���j��;���s*�.kL�GzίK��TP"��ux�Ք��(���n�ޠ�o㡷��I!H\>2�5@qvڌ�bL��د~��y�<+<�)s��4 ��D� ?.�_��z�.9�s�A5�ʧ���t�o�\�Ĩ����dh��]͝���
�hbE�S���TS&:\��������UJ�p�A`��C�S�!�#�fH7-���C}^"�=�}��z��8\�װ�R�]�9���G��c�]�����gK��f�:�����N������H�* bl��D0��78�6��צ�^n)�䫇md��%���]����>���X����V�@�r<5woY���$�6-P< 싛8���Ú F���s��w��]�p�Q�<�p�+9.�p�lU�m�*����馮�9���3�X1I��|��s�:.���$���kԁuR��/η,�tw�Ī��aMք�}%������1ڐ(a[�)��@^}[�C�f���J{��D�D�H޼���#Y�&`�3�����9������0��>ԣ/�ۦq-U��s��'�>�:Vl)�k��Z�h��7���xT�1����5�^�� ����Ϊ���4�jy�r�#�04��z����%�|ƤRn�$d[2q�+aHl*9��(X�*��q�:�@�%���׻��#9]J�:�<E�M{b�n>���)�
>�ʁ[6����r�+7��;�ֳ��Q��[L�01�Rw���.�:'�ʡDb��D���-mߕ|�!s��UX"�a�f��+�_�iÏA�7�`o _YW|��|�#�B��:6����X\q��o�y$���:p
�J����F#�Ŗ��x�H+	^��|i�QTN�3 �
סE�]�	"������c(��`)���h#��
4Kz㼻���xz0�H��`���}��?zf���N)��g)�_�B�b�=S��i������(ahn���Fԫ�������Z�'qS�L��P(4|��ȣ�e��G+�H�b��^|��=ͳ��y��v��͆��S�;!G���ҟ��o1���쏘8Ӊ�c����!����嬇N{0xHHĝ���r%}�1ջqش��&H�#�1�ᝊ-y������QI&qy�(���Q� ��qD�J΀{�-�U^�u&�����nx���E0��s\f�v���ѕ�N������_�7�'�i�s��w��5zm>��,����?���[;C:�z̟�{�X1��Qe��(jɲ�Ќ�D�
���(�nСj��F��o;�	�<{�	hG�%�����@ݪ�˿\w3���wd
�,e>�h��PIk�y�mIqx�ǁ�?���]�X0&-m1����gl�dKNh<I"0����R�f�={5�_)9ઈU��̹�H�-�)Yn�\O~五�����5A�ѱ��,��~�iX��Kl��SHƪ�|@UX'�+���a��(�£���f!0T����7On�|Y��{���S�F>2՜�kr�
�~SQ�,���\�� FҐPq4���=g���j�oD:y���D+�9ӆ*"�nA�}3E�
q2�:����/�/��56׮6�/ˆ�<pϲ�����z�~R3=DbF=�Gm��Y����5���P7��Ҋ0 �1X��]��]���\�?8c(�3͹J$0Ŷ���j�Ӧ1,���-�n�1i�אq����*��Ϋ���ƽH�Fȇ/We�$�q�B�_��Q��:�X8z���8yI�G"�+�L�I��m�E�7��7��'4ݜ1��+Fӗ�8-��C�~��0mMp�~�J�Ns�׍'i�ֵ&J��"v��1[}G�y4�b�_2�2.Jk��i��X(�
�a?�"ǝY��Z{'�I��|���(��&��EV�!�$M�9�Dg+ 1LJ/�/M3����v�0��x���栙Ǐ�J��L�Jh��N��q����W��[A9�bN
Ãϵ��|;F�� �EE�/��P�� ���;��5���܇�rU��� ��fP�
�V��>Xt^������Cbz��-.�U�'a	�Ɯ�H���yUL l�>i_mP7E|f����W���@2惍��
.U�p�%���Q�1�Ѩ�2$�N��� RY�����!�cF8�Z;�6\��Ϡw���&�\��o�/�im�e��G�(�s�����������/V8����=w;Y�G8�'2KCt�F$ĭu+n�ϤP`�@���@�a�5M�F[T��hqK$;G���A΂ܹ`8Գ��)x����-�=�I����?Z�]".ԓ�hA���BgkpA[�vS�{�&XN:O�D��k?yxF�����V:�_� ���O3�!+�IR3��l���=��r3���#��M',m�֢��uơ཯�c�L}��#ր]��V�> �ݲS?�Ʊt8���s�
����x����r��gi�8΂�=�k"	�v�C,�r�:6�0�)a�(5 =������g8z{�A���E��-��ܒ+�,A<�����'}���z齪�aM��:�y������`Y����)&�z.X@���"%�
(�����r����~R��3�Z!���BW{옏������_k/�B�Wɛ�ﭡMi�t����~m��6�U��X�Zщ�f�V5)�─�_?��6����2<����#�B��*��{�Ph7���B�r���������;�;�`Ѻ����S�վ",��_
qm�V�̩�S�e�[HS1ܝ��_�:���(2�S��2�Aˌ�GO��F������ͭ����"�������k/ߌ����r���Sq��?Z"=;�pZ��s���bBe	���]�t���.��|=bg�lM%�N�۔sQ���2�-�s�{���JJ�[�!Nk�H�Ÿ�Ĩ5&�=	�&�a�%����F�����#�O�����Ⱦ�c-��QׁVX��5���z�i�� ��Wef�s�m�-��0��J�z-�,��\֛NU����-%Lϗ/,�H��j�͡�_M����B�8Sl�%NW��nK�<wf��QU�>M����#�ۄM�:c�qVW��K���=����]<#�7fO��c�D��[�:j�f2�[ ��#_�@��c��qy*}���nW��6������:d��#v���>?�9r�C��sdF����z�)�����Y�굍;���a��l�4xi(���^����[�K%{뜏���m�=3���I�ר*M�[bT�e$&Q���F������zJ|d�%�H-�7��1��)Ǡ*�a�Z�V0Z���i��?􅸣�N��2u�_���^��j��n��x�;����\շ�/���������(��U�D��� �n?�D���z9X��FZ';pl'����3f| �"�HȀ�k��)� ]��xf�0��bu�(����K"�D�")�V�,�,4�r�n����X�7�ŮP��gk;A1�\S$�9Z���8>X�e������f�W�ݚ0�h���2�s��C���wz���g#O\�x��b��v8���9}2�^�Y�L��]��
{*t,�OFږ�#�U���W��z��3�۔�v�'����ϡ�C�s���B��@�A�ӯ��CB�!nX[OΦ�T5vh�M�Xa��n`�1�=����i�A��M�:"�(�\��� l;y���i_fh5$�a:�I����>o��9u���;~uf1�5Ys�_ظ���_���ث����Y)�{04K�Ծ\���3~Ѧ�G({�g��2}<�3�s���2@�0��o�Z���V!�&���!��&2����Z �5�uDe_k���~&ǈ2�7�=%�Mr  ��C�Yt�-j��b���|���,�4+w}8+���,}�� /��� �q�>E
��9Y�u;S�{}3�Y�����cnvK1�f��W�-��|zS�ӽ���h�S�P2�N~c�'�gq	IcyV'E`� �g�eɎ�P���ݴ��K7=� cv�B�#��
���a�s�ƍf�OSuv�ҕ����>�U4��RсRȚ>��Z�����	��)5U)���	��(�v�8W�<7�Np�M�������m�L~�	�i���R:�7S��W�j�����LĽ�?�jf_i����6(F� Px?����h�A��֖�3�F����O��\]�$�|�qߎ�q�_�ج�>8�n7�P&.�R�"����#�V+��d���I1:#ળ<��W��I��mWEcr�L����k���=ߜ�h��l���SH{��%d��{
���LH�]��^�1��=��J2���)ƭc�6~�t�����"꫽��磎�p<9�t�����d�=��+�%�J;��ht�5�����ķ
.����&�R`��s�ϒP2A���O��y��&�C-d�ہyu�(�U?�ieGm�eW�W3ͼ3�p����q���'l)����2Hd�Sl0I�T�Z̯�eM�c�4�ۖg�ĭ� \=WM�r�J�(�*_�e`fװ����,�r0����e�_j�qޜ�tDt)>�7��P�;�9n�7��QI���)9�%�X��b����UV�!��܋uϨ�9�<N����E����}U0�[� &� A:3�0�Ň�*��M��f�uS�J']��[���� �:5 ��q�b`�w(Ȕ���/�(�n�N��^�y�U_���}�S�0m.�����;�9� w��߻�a��~�r��b��dqixL?�ڣ3��}N���������z
V�'�6r����}!�G�L3 �!���';-B�lY��l�����{�Uto��P�Kq����2K8LT�܊L&ˍ�q!4�������0J�龞X�*L(5O2��/v�@v��J"�vB�NH{E89L�$a�(� u��%���7M�����&5Yt� OUd]�;�H̫_Eo+�*��TO�
���
�z����	��g��A�m߀�\�»���`�J�����WoI�o�OO��Z/�˯��Sw��'2� �gG�Dܦ��;�feXT�Ԍc\�I�A���*��RqAm��1�C=s�ێ^�o����ښՁ/�s+q2<��,�3�������u*��i��W���O���)�	s�T��q���b:�6#Kꑵ�I������0��5��<�M ��H�VҐ��'�Oǈp�$iվL�bZWe�ɔ���'��p�n�S��黚pk�AA�W�E��l�uR����РES��V�e|��L(���N���7��019f�(��vB�8�R�:7�!X؇���xo2X���"��������:��i�@q��[��ち�0����	�Ue�<�ߊ�\}9I�ӵ�%��t�Y��d����T	��V�*^;Y�ǀ[M�A距Pv8F5���Б?GUE�j�h�\���B�N[��z�%�ԁ��@�'�}��I(nN[�R����5�w�g�����}J���#��5Ѻ+�A��OG�x���N�K�3��P��W�Os`�+r��IɁkfE@w�:y�5�w��t��8��-��q~�p�a�O���?��qfQ��8ݮ`�Y�EZ��ʪK�{�˳��xM�-C���m@����CK��PIt(��e�4"֊�W��<�?�Aa/�$�-a1)`t=�Uw�i���x��I\� � ��d_�b��v�IT M�eR['�@֟4�@���]��Ԏ�����@��hU��7��������"������׏��V`n0 �r�a����]�M<��
�}>��J?o�{�n+��T��+�7�O��i6���io�I`�XR��'�O\�����WIM���b=�V:�l�����cg�a��vP�		]n�������4x���֊�����
��QW2s�t�3�:ql���h�I�7�v�;�x|D������M�F3F��Q^���je\m���ӈ���W���h��6U�=<�"w~�-�-"0�R��N}�;BȚ�����ս3C�`S��b?	���q/����e!t��@ꝿ��E�
N��Fs�����������ja[YAø�C��1��Rf�4���)��V�	��r0���=k�&(�Ye��w�d���	��yH�*+�{�l:2h��ڤ�hU;ߺc/7��`2w���k�UE���mn����E���2�DG��9�q�$��bs���^c�겏�R-W '�1�X&��0 ���Kbv�D���Be����Mlt7�zT	3NR�_ncA����y[�����y&�ʚ�Ɍ>���
h]-��<����u��%��xRu���#?��A�	@M��وy'z��-ڧ�4����x�am��!�M���6?|>+Oo���`�����]���GyaFB����Nm����2�~Y���� Ϸ d�z<�#���f�F�jvi�knN��o@��R�jˠ'JX>��K-�o`����<Ge,�
��V��7����θ�f|�q��yf/�O����9��ټ�GW���w�B�?���b6l� �[�I}�$��r�7A��FDf��ҫ�na����+۲��}=]&�W�ޣ�t��u��%�wF�jƬR*@��;���".�֡*�M
�����~�봞ʰi����g(�3�AŜ	���+�Λm��	�]�e4јy���цЬ��ηEu<�����y��p_~M_E�c��l��Fn��2���)b����#���|������Lټ*��n�S>=�;�S�����)�� �I��m�!�49�5�`�Q��q�2�rߑ0�P^;�R=_.�(c�)DU�^{ao4�Z.œfZ��S.��E	
An��8n���^��w��8�m�\qO�e�CH�eV��������1�;���Ƶ�ԥ\bi��#!Cq������_%��p���mF"��z`�˲WԶ�Sq���-/���#I�%�h��˗�/���|�Nglr�qky�0��l����,�Bj���|�[�-I���y=˰́����CnX�Ib�%.��Gg�Ӥ��$󶕄m6�?�(�l"vq���$��'�hJ!S	i|�M�%�a��J@�-�zǱ3uK�b�����/K�X��vͶF���*�Ť��Lj�s���Pu�"�q��|���(ŸL�b�R8�zw"P-����ea��`*�U�eq4ս��D�8�9�fc>�#ebԮ��1�����  �),)�g9w����j�R�/��A��!1�� �SZDǳ,o)2xQ�`�7B�h�$����N��b����Ԭɜ��������YB�يͧ��)݈>�t�-�L��y=���1���e�U�5�:�2������#m��':�H��9y�/�|�"�I���q�X����v�:�T
<���h*\L��!�\�qՌ_�*���	���y[T;���$�����y���%=�?�]�4���(f-���m��qV2Y����YF���H�&g�vx"̀��O1$D) ����@ٕW��+[�����N���U����Pu��t]�͋��S��{����v��X���S����I�"��v�A��aW+�}?В:���glx�8&��.D��
s)�#��+��+� ��nR���t���7S��'��cg"��Xl!���v�A�=?�l��̻�*�I�7�/ik��i��9K>D��%�{�b5W��7hH��mWF�`�`�X�T�)�#�[_Ʋ�����[��s7����ln����"���qN�$�c3tru7��-���DǪ4���47d��Ѣ?<��Re=���Q%��� ���K���ͨfD�n(S�w�,H=�bB��zhx�W����)&� � ���Ҡ���_���� v��'����ډ�E�s:l��^f�S�@�ʸQ�2ޒ`��J���F��Zr�}�Q� �0%�ևB#8���a�S@}[~��Y3Uz����f�U�r|�s���1������[���<]ƫ�~�#+�fߋJ0|���-���_��QTK�(TK>m����!W��)���1�<O��3$�-�Ǌǧ�WO�8/)֙5�v��'-|�I+r[b����Ǻf	�óX��v�g0����XR����#:ZO/P��F�����~ ;��w�&��T�}�#�QYr�v{|+rph���$����Eހ�lo	���@Nx�4kFZ�ox�Y]�������w�������B�U�,R�"�#����hl��KqH�/0�pEa��-\�Q(<g�ɼ�ȒO;�����O��s��?U���Ƿ�Ad����+qE�`UU*I8��6s�4�M���:���U�?��C�	��t渾8�ox�Ic�a�NOD��OP��v6B������A�X֙��a>QM,�w"��� ��܉c�E.�7��}?�d�_eA=|�c�����;Y����)�::a�̲�8�q$��qv��Q�h+�Ql��Hu����Ӎl�q� �8�R3[N�[�o1:JOqfl��υt�Zm&�]̘gv.'��M��U\ )v�~>Z����4���/��##�[Iu��N$nh���~����z+R��+�4HA�+�l ��x#�����9�-4BP)���Ү��S��5�"%5��<�U���Ɯ��ym׉��F�DM'3݇�+2 ����=�ָa�.�"CXJ�w�l�-��!�D�+�e�X�+���dn�>�0ߙș�nT1��7������\ЭF;v^@��	�i��S1�,�-8��].���t�7yp������s��;�/����hi� �vphCt��9���>�D����T)B:�dXn�A��c����:��Y��=&�t���Iw�cG'B�u��9���!�wHg�6�)e�D��p���zp��zQ��6���H\k&L���N���ɛʡ���L�_�$�y�^�U����#�Y�]��ޘ;YiT�A�&Y2��b�v�d�<�!$�Ԗ5�I��I]0�%��牲����&�&?c��� �Qj��Z']�If�;b���i0S�y��Edk��e��H9��F[@��wq�7Tm%6��-4Q%��!���uI�#����;>V���T��Y:��l���NA��fjo����h^o�w�o��k<8�@\�l�҆�x���K�n��;�nݏ��D�`�1l��!�|�z<<�|�ݑ>��w�r��)u�w+u�h��W���D(Wq��3�P���`��bO* Skx�l_/��7�b��N���^���u�UNQ�H�P�5o�T���kS��B��6�d�>�!��Y���7q�ZX��VM���K����G-ٟe�[��C�	���� k�ː�2x\�FxEC:4������13�+z3R�w�2��VIb|���ۯ ��d
m4 ������[���>x���7���
p�גE���k4	C�.��=i������g��ak2�w��^�����i���]45��s�"ms�2$b� �N������v���}1�YV���G�+�b&7��v�6.�O\�;*��ْ�F�1|�_�i�~>��aUT�����{6g�F��e��y������5W��Y����T�*�z���I�+O�C��K6�ͽ6�:8[�U�OJ<�S|�����O�o�HP�Ъ5�Hh�\���$�
Fg҇ұ?��`=Q��W*fP�뀸��;���Ң�ka�1y��~�����1��Y�G��T�!�i�+��1#}�� XOo"o��J<�9�H�N�w�gAq`�uLc��}w�D߃�Tٴ�F��	�]|��~P��(�h�7��_��,�_�0��G�7M���|sd�X�&��t��O����q{�6Vc�ǩ	@i�Φ���A�ψ�)��IӸ3Ū�|��<����1Y5����+�j�o�+E�T�"_�������ك��S��C�k�D��(S��e�,+�Y���Ҷ<�ߓ���}��{��'�󚎑�A.�*�d�B����0ҝ���+��l�٠��ɇ�c/d�_�w��Q�8��hx���7	m CCM���a���x�F݀�(uS6M{hne7��W��#��I�
.��9�|
���}2�dLݔ�?���3��RiR�����)���w�v�*E����LH��8�R�LlkiE����ug��G����2R����%��
�P��F/���ҟ��vd�t;5v��﬩Az��+���hx�s�h0��~�f`�`_��}I��	t��v|sy7�i�_���t��s��Oh���a�A��"�$���s��y��.C�.)	Q��-��8t��6�B^�ZjŰ_<�%�m��V���:�j���p�,t�g^w)Ӽq��"qfi�ڻ���ӎ.�՚AR��p^髰��Dյ�k�e/���)J���=6q'ob�X]pɎBP^"֎LН��q1�(��QPd�a ����I�s�-����gG0�&��4��h\�9���T�ȉ~����%"��%��a$a���ə�JsoI�h�PB]��t6��Gp�����K&[u���!L�YYˡuӽ��Y�-�����"f�X������o�6r��j�r��G�/�Z����,��22������C0k�e�4_��(ܞ��`]�@i�����I�Sb�(Hst*d�k��U�7��U�hI"�A��ޫ�U��t�7��?pGC`ƾ�Q"t�g�FPdP���3j�ה"E�"Rl�A�v�M�My�_E���Xz�����/N�E�.��cC#�-�m��������mG?/�{)��Ec����}e�����5`�T�� �s@��~�=�2�8\3q'��>�Mϥ�oz�j$�r�gdH\Y��|�/�gc	l�)ݞ���vH���s�����n!�.�R�v��2��*[s;(�*�� &����p�ks�{�b��֒��S�>N�m}u��+�2��vy�%�$R�;�8[8z�;�7�ꮌEE ��=�=Y�n_�5���\2�ϾY�%S7r�t�~�:�-�;�*'Ҏ$�pi#��x�����D(Q#���[o�@��+{g����i�����b�q[��X��E7p��}'Y���;����kHU��RY�*;XH�b�(?`O�Jb�恣��
ω8>��]���o~��S��L��!tS�r�b�ҩ?���~���vR��gF����gQ߰_$�*������M +�OsM���@�Y1�(Y�w��!0Jx=�H�0��J[�t,�C��Y<Q|��V�h9$��Q�	��X�����xĐ�K�� 2��=�|���c��M��	�����q�b0��˾=^8�� `E��x3l�4��-&ڕԤ���m�U��I��\I�|�Mv��E����	L����fk�x�;w7��\
��L�S�1k[�)�YQ��-C�B~B������|T��ܗ6pTd:����H049��˜�ֹf���;wm�ܒ��I��`T�g�6�Hhc��#0����n�i�QM�O�0-���E���b�D��6�vd������0�I��� �bYg��R��he�i$��;���)pG��������n��6ٿS��~z��Χ��fn�f��j�)7>tz�t��Mdq6 �pR���H��&��f�����&��q��ҼL�L뛾��:Ln����/�����6̧���`�B0��[g�j���~�L��JM�2��;��\�z���8��ۋ9]��V�5����{��9�Ūx����Ud�l�]`�BԈq 2��
�F5R\�(��&(ڷ6�ua������t�	��9�NiO}q�1��M�W�3��κ-뽶\r�������+�򑌠L�={��w� �5Yê�:��K��Su��.٬��8���7��̋� ���d@+��c����k�/8�����OEU]������yd��7�^��̛�����bn��o{C���d��a�8)�F���^�'�ՂF���4�P�V^cO����'���4/�6�u�d¹�B�D�0���4��Y��ć�r�T��#��5��@ٚb��ѶK���A�G't�� ����p}�X��+��gO�1�1'l�x�RDb��;���6�$^�����\{�邕n�|z�BxnḔ�uhuQz�|�t�J?��5� ����+��~�����w�h�(S�V��9V��?�0�G��q���i��U򆳢������y��Et��"�pR�7�z�+�Z젳!�c������#ˤ�Rj���YT�n����9'rc�[	xޢ������	���y�7t�h�wV�l�D������Ab�rx)����!���sxʖ(��e����8���M��*��+h"��2�аW��b�g�5��L
�ȿ$<��Ɵ_�~�F�[��W���g���e�<�c��)�}�`$����Ů
{����)o��!�Mg��ժ�����#��@{���z���}P��t�.X5U�2��=qq)#�׈���5�l��wuk�icZ]��u���e�<bk�٨������i�P�Bm�V]HM6���t��-Tp+���%i��"8v�4Y�8��q�Z%�q�����i���85�9�L�?�e8��
���t��	I�|:�f��8�a�	�CrD�5�=2�ь���w�vl�$����^:�f^{z(�|�I��q>~�_*0�/���`<�N.|���-�c��s*�oK4p(���.�>�ERk:���SK��߯�u�Y��W��X�
i/�i�oS�b�=��}?�v���D��}�Z�DЦz�b�T7�3�D.6���7�j7�ѳ�UhF#S���pP�&��@�+�R���	���wD�n+��C�<hK�w�zRF�z�g�@fu�Cdc�[,�����(8�e������hm��J�p����|o�FL�!ry<�;��{U��C�\�f["�){�r.S�m�RW����9=#�$�@|7 �YkE��F�ښ�k�:����ҹ���u�äN�T'�P��s�H2�v�kow���9���}�Y(���yi��~�æ����#r|6���eQpc� ��7�Y�kS�c����M�r�4]�i��gRY� �m��Kf�) &*����M�"ѕw�T����^������*	�о�,-�]�%4�/���բ_��뗫&�< d�)�PJFLp�@_t��&��.y�oИ�G��N��W��Hܠ����g�v���u#ޙV� ��)0S1���;l�KТ}��Qiw�*4���d�r�&�&�i#0x����.߆o�{�4�AW��|{=䘋�17�G~i�,7��4�P+����|��3�4a���n m//y�+>Ah�᫉�W��NX@7V���-n3�ь������kN�rf��S�_s'�|��WW;��0��ޓnv7�*Tb���#�.X'���&���ϋdE���X����\�#N�aۏ[�I0jQaV��������}C�P��c
��Ls[�5���`uI�V������h�����Z+@�3��I�cf���	NW�!�Q�m�̈́�3�?���k���dR���sܴ��}�/�s�!y�B%� �y:
`D,H0ޙ�h)�OWx��sR~v�F	��))��+?�:{'�^0�-��̯�F>HU�]]@�{�i蹜�uyT=~NoP�: 1�&����M�k�$a����+'׋X[�܍h�4���2S�^I����\)sC@^�b���]Ӱ;E�dsƍo�{�7"�omR�w
8E|�
݇�ŕ�ߧ�Q���Iet��k-}��?�V��=�48kz�_�=F�A} *�ԼX��{5���x I�Z�.�n!�p���R6���9�y"a#S����F��&.�4[d��#���N;|\8*Pmn�|��6��p ����"�خI�b�ƃ�_��a+�x�r���� � ���0C�4n=��7+����D���	J" �.޴��ǁ�Ɗ�LG	r[�_s�$��?To��"��$�![�R��-E^|v��Q{jV� 8�r����zX��{��M"hG+<�w1�S�}��U�e�Z��� �rߪ�F��Ն"~]�5,
`k/] TnSb'hե�c�J=��^��t坨��̬@����/��F�5陋}��6M!�Ehd^���p���w`EJ�D�m�d����〈~�o��!�"����[�?�?:�<SWu���~��^.���(�
r���{����ꖭn��2z��}��K�:��Ǆ%� ��1�� �a6 X�|� ;�7Oqr[�s@��$b	ꃂ�6}�����9���twZ�O��& �qƮ>���|#��y�|��48�	Ӄ�^�B�W�0Q~54�	�B/s���
�y^_X5�{Z^��X�'I��R�j����#2}�����ҟu�j~��R�IL��ʑr����ҽ���D�+��P�Z�D�*Φĥ�5K�,�uՄ@N�c�W��O�������
��������2h��;����kKA�j�\��nf�/�kZ��2�:&;�Tᜰk��z5��t�	M�����;��J[Y�z����_��E�fu�{[����*)�65�}�ب��YJ�b�y�y��w�UZm�k��̒�G`Q|�I�d�󅴮���J��t�Ӑ��<���yo����A\i������e+�J|��#�L����+�M^��$��_��[��4@j\�+��%�'|�hԭ���׻��i`\����� �_�@�U��u'���t˾���B<!�^��:b�u�@���^����r�_Ř���؇�"9c�l�RB"K����/��FJ��lW�(�1z��|'�8C���d�J8d{shR��������.�ܚ)y�)sz�ک���N���U�ό�	����c�ȟ�Q5'�R�+�E:P�n0���0�J?�h���j<Ur76B�����'K��H�js
g4��iG?�F8�I ao&�DS�*��O�a�d썜�Y��Jq(�k凿7_;��d�%�١��0�qКY�ĉ^k!����@���}�����u{�z�J˳���=�qWB�&�q�j��H��$99*WJ��&Ų�lE�%���.8��.�!�*�������B@�2DBq:�0F�3<!�⚕H	��ʀkt`OM�+�2Fc��5�y����|���g޳P��]_�a��2V�+Y�߿��������TA�x��G��ͯ�̆2L��6⍏+G���yn�������1�OП��g�׷4��L�|m�Y�AjE����ttXt>�ɏ���l�qM9��MJ?��:_O�x��s�K�ؤ^�<�Ij�}����?��a�T��!>vy��b���Y��Bȇ# u�V��!o�@A2ՙ
h?�#�d�T���N#��N���o�2��"�Bk^"E^��{�a57H�[�t�O�&|>���Z�]�+|1Q��~�6�J�0;����gSed��jM���	Τ��a㔼�m�=�d_^�����L�h��7l�h,�f���^.�XM�؀��y�c^�C�gN��N�R�y
w�J?���.F�H���c�8L7�b8��()A sZ+e���"*^(�T����7�o�i�A�e`/ݴv�G��:s��&xv��`�3�~�N�����5¬J�rq>\,�d�l�Z2��B�:�;�_�W�#�_ke�{-�?H���T�|sp�h:%��%=�G��Ŵl�������О��d�k�ᬷo�Qf��O�-3�n�u�.!�lt��qJ���	�arv�`����&<�7��;���`�ʗG����L�菤��V'��J��Q$.+���9��8�mo|B&.^=_4?���g���}�'_|���>�����'0�����N[���]'�Q	M��u[X��I������w�JA{�Y��/�qȒF�4�~���F����,Tf�<o?��V�-D��;c�j ����d3�!�m�aq��5�ܗY����6a	qV��i��VBLǖ�5��Y#铴Н� ��ǝ�W�Oѽa��^���(�˜�7TA�F̯�zZX��鮅{�?�Y��=��4�(��0J��۷fFa��h�U����ӊk&�uX!lb���G[˧.5��H�7!�x�[�a��6�(�w��� ��,j�C E��L̙�jI��'�yN��׊��#�i�Ƽ��L�GѴs4�(�Y3G�`z�B���{PT((������ė���$P��D�Ÿ��Os{���s8Kɻ�������|MA�_��2�k���ʱ P�9����k�g�~�C��i#֐��n�m����V��o�+"_��� ��q�7�:�C�3�6�n���ntI P$�q �$Nv���F0�M�T���z���6��\��/t�L�4p�|:�; K��*��洶����X���P����ɑYFǱ 9LF7����UZ��;�{q~��c^lP���l(�̹����.\�`р�y���ڗ� �@
�"�q�V[�#���f_#<�����8
�G^T,VD�{�-E!^R�3���!��4��ci������>�D��{�P-�r#=�(�w�5��ϔ?9�r:�Md��s2D�L��Rp~��α�9t��
Y�428C���\��ؐ�g��f�x��b���r����N�O����7��I)�/�E޳E1>n=�0�7�WK�<���)zt�w�� ?�X��H9��v�W�2Fv��J���H@"Z��P�li���J��˞oBN�V�n���=��]���z��wt!�P)��Bh���(0�"{9�1Ώw�'&�<c�SQn���9�`�&[��ŇT���f�����)Q��dR���Se��!�<��)�ӽ��Z���R���@����	�XkY'���3%�I�7�6��/O�i g-,�f�7�NwN�X͑���8�������	��
U�8A-	@�SD�B���X��j1J����SDV;��~��y�@>���5r kS�q�
�>�rL�d�cB�l^�=)����m�yj\ݣU�8�5�LQ@��jdm�fx@�Kj): 8�z#@���+\rHZغ�-!�T����"qM ��v�/��TW`���G�N_���������n�Zר�Cb#&���vM�}?S�D뎽���2s����Rfyf�=��V�e����@�4 ��E�J��7Z��D��,����,	%ǰ���c�\:[t����A�� \����=�{���-X.wrx���p�(�59s�N,����$D�*Xvx
A�n)��
(��z�-�	�3�S�qR*ӆ�Bhw�E��QX�yL(�h3����S��wp�=е\���m�[?����Go�J��J��uT��[��Mt=��7m�kjH�	�cXpܒ{Yp?�>N=K�o,��/(�y��4����F,*��>��*����X#����&:FLw�l�S!��_,�y���5Ɋ5C?����sA��qhD�ӌ�ح�Ɲ��2Dց*L��y����+!���WWu_[`�W�6�
���Z�)P����v٣[�B�R;ؘ;�c�Ԉ(�'���D2�z��L�)1�����4�[�Ke+�嵨���~��FT����X�M��22q�{�`0��� ��N����4#��Wr|�b��R
���wq4���)�=-l�v�{ˤ�6��OY�T��k:����V��
��]V�葮�@N����Af�iV�I�hz{�i��b��8�O��I^��W���6j!�h�Y����Ӏ���QB���-x�YsH�I!jm��T�/���b���/{���ۇ%�g������є"��g0>�ϡ����� ��g�(bV�@I2��`]�G]�4}d$�"����-Ꜽl�0&Ko刣�Q�$���#�]$�w�kTSOخ����X�:��W����ĀE��k@�j��͕�~^?2����L�dKM�P��0pD�fP�����Wt�h7{��UՄ�HM_�������$ B���mj5�!�册5gX�Q�}
C�I�~���С��T�-�M���mr� �7�d�
	��!��������`��7K��CC��m�l^�5�����z�Alq�
�gb�yq��p�F�L�L��2��YP�,Co$���y��=��*���n�s���a�Ja��}��"х���S�T� �
l���T( �������e���Rۧ67L�4eS��M��Ն���`��^R�VE`X�'�#��j=�Ҙ4I%Q~y�O�b������=m d�;��<74Ȥ\cGq��Kt<���8��H,���ɡ��'����k�������vVɞ[�sB�[�W����Z�J��)����9�Ɇ=��Y�kc��"��R��zA3	�A)')���%������g
�.��>�2�~FE����녳��]���M\����e�Lb�8C���qP9;;D�Bl�0��(��d�h����p[�vO�x���	��^�lc�<�X�3Q�A}�n������\��eA~�piqH��]%׌Wh�O�$Wұ_��{[f�B�8V�@�d�����ɭlv�7'+��vU�ׯ�er ��A+\_Eʨ�/jHf��SCC�ѣ������}�" &��4�~ (y���iB+���j�� 7�a;�� $�P����da4�,�Ɨ�&��=Nf���k��)޸�c�r�����?¤�^�µe��^�f��ΰ�(�Y�H�<*"��i.r�3�<������� ���c[҄�}�_ռ�׵�;#;9/6J��r�%M٬�U[�"��}Rڣ<���=OH.�9��b��}f�$9I0Խ��}�$v���J'��0�Dz|�D���y��q����Q�3C���w��9k��]C^'��i Dΰ�B��i���b7'	y��h���~oMW#a�� ���K� ��ǚ��F����{�+�U4*d���R%�:�]�3c��l!�Y^8��R��y;��cl-n�����?/���/�9sQ�QNQ�3go���(�&� " yvf���� ��3oj� 6s�f�Z�x�mP�	H�;�g�2U�RX��z����a���Z]�L��>��u3���N'�"!���up"m
�~�s,~��ֈ XcB�7��f��q^��D�R�k��G�5��+��d�U���9q]#QQ0��1=���_Lk�yvו!<x4j�7e�L!��V_ݹ�b�qE�����a��y!��` ��𤖿"���G%�I��v��q	��`�Y�n=�r
�E�}�'�H��I�:98}d��N�;�3@��܏�D�ޑ�;���c�t�4�cT&)�>F	v��X������;�Kw=�5' J�
��Jn��M:4Y&�s�a��]��Kg1p�]��ƙ��f�:�0���Z�)`�-�l�Vkyݦ'\�7�ж0��@�~�/����g��Hc3M$�w�r���e�1�J�����>�@�,!,L�6�D	��~�"���Z��D]pq-A��������&us1yf�-c���a~�:%��v�d�2j�D/	<��T�y�Xo���b)�O)_Og��_�&��\G��c�}FJ��ę�}������:�GU�U���^�$9��Y�K�����}�8܄y����^j���㧠���u���$*pD�f^�?5��
?H�C�y.t����N�ʢ�M�y+^*A-�ry428�ܐ[e�#?�2.����=&�8?s_3y��G��癅%X5�y֊9���k����<�����[�T��(���Q�7��·�J��0nN~�v��ø��~ۇuujb�`f���6�:<�>����������d���E��3�S��S:�D]
˰�&�������M���(h����[4�Y_/�(�4-����_��'�&�u����P��H<2A���:��¤�+����L�\�,�Z�_+fq��sc��������y�ҡ�L+#QX-%���~K&w��U��و��X[b,X9�ik�� *�kɕ���] Yc�'�W��`$�I{&R��X��㩸@W�0��c���O���t�뮐������^��~ň�kό��4�s���ʗ��h� `#�Ķ�ˤe�\�/���$��_I����jU�GCꜴ���v��@U�t�lg��K(EY�7\_X9/�ķn�y*~j��:�.�F��^s�<q�p�r�Ӡ���y�]�/�<?�9�v�B�^�`�ٕ�f?)c��:Kb)���Z��QGuK��&��ֲ���f`�����l�P<=�4�.�L�2p4�d�wBT@��m��jd6k�ʦ�L\��1N%��{�#���U&��&y�XW3��gM�6���%�p����( J�x� %Sa�r��'�w�E��T �_�v#�6kn!����ɟE1W���h8�
a��Z�Jg��Ve���B�6�z�=���bj����u���3��AVX��	�����qP�j����!k���J��nڳƅv9��p�/x�$�����-��x?=&r?�;}�wh/�bY�oL%�x*._yb�T�"�s2�9bx��Ʋ�9���.P��Y�%g�xM|��넏��I�8k�M���G�����ƙ��W�b�غ��"�.���j���y���CV[��e�4�X��V���s�U4~��(����1�k$��;�4om����Q��T�̔��%�Fm��@)��X�������X�B����+����qKD�K	W��Q�j��#?�1�%/�:ǇPM3��`���]GCŜ-	����߁\���m��5�K�==Bs��϶+�?̖;o�l�cRb�gY�6IC6]&����>��IZ�1G�{k1`��-�f�c'�.2������n�6`��a�H3�F�:j�X����?�ӆZt��zvJ����Y��?�b�J�X�����Dg��ޟ�V�2��|��D�ȿ�c{����v�f�VĬ�fڊ�Sk,VA�F<gF�D`KFH.[4��MO{@V��oܔ(R󳩝7�݉$��f�b>��ޒ�h�k���p�$��U�xmR�3��_7
m�kd?����>��xʟ=�d�#q�XfL?���y
9�6*��C63�4j~3�c�Ν��yOL�� �����	 �_~��d�0�P#�.ǰ3ŞLRu���E�
/K)!4��Bm��E��n:E�J���'�}f_|Os�n��m��q���}34���e]��e���b����^�$��
t�
�t���y��$��	���h���H�tBaF�ͤ�_c1T�}��8�nT
j緦��$�/@Ƃ�)�Q�.�Ӻ���q�/�[��1g�C�U���_������>Λ�r�#a����s�e{p*��!�eLۑ�`�uDb�qFW<�co�\թ�Nm{D�oT��-����bt��c-HY�a�?�㞔��6L��u��2�d�|�ɻ�X��7�R����|��(eC�9��c�_�zc]Z�K����E<�񔮵4�?g����2�\��-�>�#��W�T�U��>���=�0��g��8��?��%��%$H|�Ս�j�u���(�v��ěT��QUZ�ӑ�g�z8(�'�I��WJdCΝ�}�W%R���o�ET������K�Da�kb��G�V� P�Nu�b{�En�ˌ�O�O�|��I���E�`�#W�i5.u��n�'��X���UU��~�ر`�.�2ed���v>	��PEI������a��X8 T���ET���R��n�[�q[a�c�9�ZL=n(�M�J���D��n��仇��	�*��R�H��E��'c�MK�����r��8�+���k�$��M�w}�l(�Z����~c�G�l������.���
�F��X¨'V$�-�>����7H,W�EnT��n���M-�� �����&U��р��xw�����@����A�{���%�\��"eF��O祳����2����Vvfw�ۜ$�����K���lQ��!�<D���g_���j�o}�y���@9�ﺲ�Hz4��|�?I�XG����;$�/bW�vۼ��K��1T�? �u+�C��v��(���w�$�H�h���Ѯ5�h���(�4o��I�M�۪ͮq��L�&G�SI[_�g����v)(e���4Rʊ��Ƙ(�j�1��b���ku�5�AQ��K�t���N���ꮳBT W���=,?�f��~���+1�;�4��\�<��mu�{/��4�x-Ex���#�Z��B|�u}iC��<"�ˌ�S'�P�1ڏ�m���f�}���,�$?�8_�*PH�i��I�C=��f����={�����aͲn��
��E�	���ԭ�oDd�[���x^NS���b��F��V(Uх���w�������V�|M]O�1UH`-��;�W��t�]n\��p�5!9��0��obix��1~t�D�fΛ<B�f`��a�$ݶ+K�cB���9y���H>�i��"g��@��"K"5XՏ#�,��IFK�H��]C8�yȑF�����|���#F��Ka�k�+�ѽQ�����^�����9��{ߔ܂T^�����J^Yj1E��V`^���K�r��w�z�.���;?�	��9*�oY�2[{�?�j�_8J���0_�#��ҘH��t;�S�ԐT܎Ɉ��Ax��Z���lهT+�k�
E�eq�LUT���xY`�)���8,�J�XU$�~hQ����f�\.��U��=��"#	�q��XA{f��7�,Խ<� u���!gZ��Yt���<��;8�{U(�q0+���規�k3�S5��%m�C��.[��������F��Ț�6;�.��[]�	�$A��}��i�)�d�`bDq`%B��*�D���
7��ІŤ\'��(�l8��*��b�������|���/���X�Ȧ�hc��_5I��x8�6P���1���m��#��ɳ
���؛kX��0W���}ȭ����Y��1>�*"s^�s�|IH��_k�o�V�P,Ӽ N�|=`w�����T�����6}o��92A!f�\�й��T3(� ?)ٷĎv��B,�u^dБTv�3C]Q5L��s�L
N����=�M$����E/����<�m���t#Sw�Kui~�����>3��"1�4��zD �yd�A�W<6�Bک?�k~��ew��Ԥ���QI�]OQI ��%x��3M[*�d����^��dqt>�`��`����ķ�(�Y7�_�L>̧�9��:,23Ȣ�͍�7�ɖe�i�uv�J:�F� +��X|T�#g��<�rG�C��r�N�woC�!�#{]�Pd��3��"�����{�H��s�K!�!��0�壧�wirt�f���RLY��Ht-�3X���`F.H0b�}��ĐVD��/���Q6������J�%-���b&����Ψ�Xto�+)��D�"�*|b�Lr��[:�5s%�K9:�;�������}ء�ӳQ����X�����{-Fҩ��-���(7��ڽME�5�)yn3%K�JXE>l�r9O�D�3�t�{2��ŘhܜY?&
���\����G� /5[�|�r�W	���3DooW';�ԭw����JCڧ�@��#|}�-�$�i�}�Uc����8,0��;�ە�=N4feOQx�'`\��l�v]OrN ��q>S��;�榌D(z�=�����rQy>]x?(�r�������s�T%a�;�g�2jZ���"E&z�u��)?G��K����h�G/��%F4�N�N�ǔh����{���g��Z4;��$p��������S��!��{�k"G�?��'�ڈ��t�r����EV�Y�RL?RH�#o���X��6��%B(�T���=q�e�t���?���p+y����+� 
�&����>i��qz�沜�qvwo�G�T�����07f��,]<�q}���#����Xu�ND��@��D�%$���Ր*�`�����4���Vg�vxaĭ��/zS�S�Jh�W��2��ݵ���"�����]�A
�����(>yT����i�Az}��+��8(��i���c��gKy��)0M8�� W�,�s�Bǣ�S����e��,��|�
\�.v�k�ـ����W��������0':|�Gx��7���F |-ߣT������tU�������bQ'$�ʃ�����<���ᚭx�~W�w��7�G��y�������[eOLMn(�0�O�q�g��t�_Т�)��/���LfȆl�2!<a&@��H��R_������Ӊ�l���c����J؎��Sx��xb���Z��L4B�Z�a�xy�_��N7/}/�w�u���}���l~�;�4�u|�NLXdH(��|��߬ސ��B�I'��3���s�25��8�̿�(��f)Ic�~�f��9��XgY`	�+��lۏ��=�A:�=h\�[�MŹoGC���I��h<��I��� ��(Mϕp'ʎ��|u3�_@^̥�����b*�G����uBo���ߝw���2=��j���;ǜq�>�4c��w;5�cҘM���%M,��6l�Q��Hp����&��t�4�Iӣ�'�WYTB(�I�eN��q?���E
���7�R�:(h">]$���}!U�4LW���ˌyl�_cd�X+R�\�W��Zc�\�phf�����eҪr2���(�C+YA'P�Z+�^�KmeT�8����~F�� /�)5r��������=ב�PqQjX�Ⴡ��y��DW;1#�?��]�����F����TfԤ^��((�ԢĴ�W88�����g(%���MG�^�0��LC��_�	�Φ�3h)��q�>Q���	I] �'��S(�-�Y�X����IS�>H��W��ߢ��-Atx�F�a@�U$�wno@65�8(.��G�F-�F���'�Y9<�Hq޽ϳ;(�0ċ�Ϣ��u-��� L�׶� ğ�>�Ӟm^�t]낽>k�q)y�'ejw_��e�8ș2���RD.s��\��i�9����uo/���Z�h�M�����R�4��@����(Ã��,���2Qc�1^�9H�i@�v�?w�4�/�~:Qc(�#�3ZčG�ʑ���g\��B��t��V<�Np�1=���\�佟�{�ʦ-FԆ��5T/�2�'FJ��;z������W�ޟ�_��N�0cr%̯�[&��l�'
��GXa5)`c������$�8��\P�LA�O\�p:��}ri����'�h�����J�\Ɲ�M+�N ��4�e�,�G��٢���6�7���wBP�N:�66|$T��?�L*)(�FZG�OJ�)$S�����H���!�I���H+�H=�T[�t�����zYz�%�9���4���A>à�$����r����'^�d���I�u{�$ {B�V���}�=��e���F�xnS�?���7�Q�\+�tX�ʅ��a�@��60O��?�Y��fk��X�;d���0 �� J��u�v�T�/<����r�
+a��L�#1:ʋ��|'ݠ��DA�$�l��_e��8F�Ak�Xj�Ëz�%1���$����k]�	$��[�)�+�&|f��H}LkXT��>������ݐ�)�*<����F���9T�^a_d�?gxw�-��*ZL�8P�vp��D�P��Һ�Hȹ��)��Y�7d��6ry/mQ��]{sϡ��d��J2�O�y]N�m*��s뗨Ǽ�n3̪:%��rڭ�㰾��L���?�5YF��4���o	�o�ľ��4�UV���6)KM2M\pM�~�|B�{g��`�L�ҙ1+f7����/��6fIA�j� ��]���|��5��|�sj|�˓�y��m2Z�c���,��W�Lt���I�>{����ŀ�Ym�z��O���A�^,�l�ú��랱W�x��Ƣ�*���y�~��+�Y�}���M:q�����Nl�(�(��?�^�γ+U�/O��\)��W'�m2n &:��(L�L�;��.n�����n%ε@ζv/��M����f�"+Û��Sԏ��m��@f�h�yƫ���ϋ����Zk���ܮ��Mb�P4;�v�	ȢYq��0��QJГ�
x���EJ"! lTij>�4^!��ed�E��c��v���}�K�Bqp�9���^�om���&Wً+rރ^1<K��0��^!=���г~�$h�0�[]m��`V
��r��w9*)Ky[
J��Z]P�K��_0��*�H���3�umo*�:�=ge��e��I�)����l�*�'��i$�x�����B*���{��PB�K��j[Ȯ�Q��:#*�ņQ�9�x���su�6?e? �V������Y��I���e���w�I�=3-N�asc=T�+�O��a(���Bܳ}~W��x|O��'}m*)� $�Dc��B��m�p8����+�n.N���#��mQg���ۚ���#�n�ڝ��+�L+z�ߘ�Ŭ���L\}����ʌ�Xrb���I��/_V�N�Ã��4�����p9�J�|7"�E��})/�dh6�� ����^����\Y�p����`���?��e`D��\�*�e�+=�Һ� �tl��qµ�C����q֯��/G�/o�usg,�F���aR
zm�G˼�`�Æ���ͫS�Ҩ��t��?���x�#�dN�	eqJk�s��A�� ۶[�ml�:s#:�X'e��Ӽ~h!	�ۚԾl��å?H��8Cf��&ۀ�����,<=+"�*Y�e�A�I�������.��(��s%±��e����GK��<E����4"��E$u�yf�a�Q�AV���e��I�y'��f���Y�<c��|��\�p��?BЦ�ˉ�}EˎgN���y���I5��!x��H�-�~�d�+�J<ΚH M	x�ɓ�G.A�����ɾ!���A�R��*|�s��)��v�Gq=,թM���A����8�{p:d���𪾝�h�������q6��I�9V�S����r���16�c�
�bj(��N���i{B}�
��#>!��1�.��y}\��HQ��~u/V\BHT�Ƀ����塦�d܉4p�������ʚ��$]�8�I�=�W��J����R��.L�ݨ}Oh�F2���t΄�)bY4���B^U��R�� pe% Re��F���m.�AH�ΐ"��xݖq���g	��.^^� l�J�^�M}�^Q���|�Iʐ��"OS�Q�+��QD�<rEƄ�(��sT
0�J9�	��~m�U-w��[�|U	�/xFZ�Ɖ�l�]�}��!=>~�k�b��=4��ዖ���m�on2\�s���AO�<tJ��zi©mMT��O���� ���eR%y�0#�o�
��O�ÿ����m��#&#�E� {�q� �l,;��-T[W)�f�ƍ�����==q����XK�V�WǕ���bd��`<Ԋ[��22�;�jj:�9�$���e%��Z��{�^#���coނ��^��Z�����:D�7����a�ֿ��G�>[B8z�}5���Q�Z�{�y�}�&��NY�������R� $'ꀌFn'�I�!��:�@?!G 1o��?��c����r!/�B�<1�1����q/��� (÷`<	�[�݉n��s+�X/��
ԯ㯟�7�H�uk&��K�%jÆ˨�F�<��C?�m�B�=M�KR�Qh�`����q&����O͂�w#i!��ݣ����}W������'�a�If��� f�Z�.�����)�4%V�#FB�Ka�Z\zq�a��f5̌�٢Z�\�� ��Ov��a$�Cv�>i��5 �<%��| �l�	&�"Fe�����)D��6i/�X��zB�W�<��"E��~e��M[�o��A��}7��x�W=��g�0l�lZZ^j�-���~;���iծ8H���goS�e�B&��X�T(ڤ΢7���!2�Hw\�>>ó_}Y5G�(c�UQo0`3�Ö��UnD�(��S�o=�'���Kå�x_���C18�4����r���;VwX;q�li;s�'�B�Sq�~���-V�G��jrb��y�9��]���g H�RMtG�,*����T�TO��t���?y��)����lZ����t�OM���Ė��h�����\}���2��zi��0�<ڬ/Y+�]GCq[����j���N�f��Be�/����@f>\^H� E�w��F�g�W��kQ�4�'�$�|���UPY2cڧ�<���'d�s��^��D��D4�U���������J��(=��� ���܁w���g�_�d���Ff]�
P3M:>r��`Z}�� ך�~(;jC~S���΁���e��9�<2����kW�)%JKQ�w�ow�����A&���VTמDXrfO��� #ܗO6��ԟV�f3U笧7Ɋ!����H ��C��9tb�mRnRʣ8a�r�k{���fs�H;Zǒ�5%%�Hto�?uG�8~X'Ze���k����cͪ�0�H����'}�o�`r��^�~ЪR򤢝���\Ƈ<�����y)j��>���2��q�j�u��B8�=9`�7_2!�R��jG��^F�ޯ[\���3�ǗL�f,J���' �H��*�c�T��ń���4����&M=N)�.HSP�p��ݺ#[fe��N:�0Ieϗ�kͱ����@E��#�&�᳨�b�R��&<*��������p�6\7nst����M���s��h_E� ��=xK�j�>�l���-��H=���N���I{�qFr������82+'�ݽbz<�z����S�$���
ǧe�g��T�IB���l�o��C���
Z@W.�n8y@�Q��m��fud5PF`�i�mjؓ�E�Vx�"���iv��� �. ��J �a��ğ<n�N��W�q��(��ƣ���v�]R�6ɄoR�]���y������εD̉��(�WǏ#��8�����ʧ���v^g��� p�Iw� Nb��(�{|�0����(�C��⡁���7��{�nP	>N�2UJ�j��̸Zl�)��N�&z�G'��3��I<�g������8�<�+��Ƿ����XG���3g�E�Ø#)��j�>;��79g��j^��츍P�2��>Ћ�4��v<& �ck|4���E�p�yB�+cSٯ��G�ܿJ����$�6����t��6��T�5+Q�_M��[쀰��dC��L���n�Mr�鰂����a�E'�*>;��&��33ɄR�T�߸�:P����e�P�^?�f>�q�B�ʨt��P)���GU
�Q`�i���7�Џ�S �dV ��t����!��m�ur���;�`��ǻ��!�z؄T�2!���}�|w�ʾ��@�Se@����un�Y��-�Er/�z���^���'O��<h(޺��RTw���3UI�VAҽ�������㯶�5i����
��� �"rAt]�Ϩ�ls	�l��R0>��@�o�б9�5t���Cxn_���
v��)1��h˨�� N�6M���PPF��CϦ��T��
�YLX���k����1O�0�V���t��ڗ~I�A�a���s+���SZ���yo'�B���Qo�h�U��˼zڝ
�s� >���^��q�F@��
�ٝ3�1Y�;���7���qp)v��Z��^'M��'I��c��N �^O>ϛp�-_ˈ΀�:��Me�qE�f7�lO��Pv�����xE{�z1j��6~�,vV�$�FZ1[u�Zm��Jq�sl�2���n$�ԧ��v+n�l����U��vڗB�O�4]�����֑}��a���G�w���@��e��A�7��f[q���b��O�����> ��~)��:\�BCҁ�B@�&����-�����6е��e���dr~��ɦE�7���LO&�	�ֶs�����/�lSW��d bA>k�Mn�A�lVk���"U��zV�=~�$�öX՟����l�ܮYFy��6���)y���-�et��E�_II�72��R�?Rw��G�˚�x��Ɠ���$����>M)�p�,�δ�9FW�s8����M'X�u܋���]~!6��U�Be�n�!���������2K�H%�9�O~��tM�}Ͷ����|�ƍ�r5��E�+{�#�u����6WN�k�&�@Y�Ga
��s!I��˟2a'i�2���t�ڐ:�%�P>�̹��f�x�X a��2���c����E����1���"�m�q:�fDN���T������Vb(���B#Nuȸ+�m�7�Ehe�i���=HW���P�bu���r��U1;U�ə9�9V�:��9�4n�_%�
��P�F�ߙp![��}��U����ɜ���v�nAq��sϪ>z��{N�g���\}��Hk�'0�N}f�~��ہ{MNK۴j���e�?� ��Eʀ��� �<�A�i�O�)���{��=ˀB����9�*;��:#�^�\���r�пyWp��7� }��Ċ5|MS�K���u�M0��ʾiV;�I�y�s �\D�,k�u�u��&�?翘��?}1๜��O$	L�y���4J��3ؓ!���P�6�2Bwvذ�ћ���%=-�0Q�N�
�o�vn��RD�-��Hj~fFN�W�Z4#{��Gm�r1���)�r���R~C޳5������학�[�D��:�Rz��i�ܨ�ns܀��^ѱ֥�#�h_���aO������{؛{�d3o"r:������X�ֆ���̳�#�ݚ�[<D �饞<'�h�S%�u���AE� �ĐB=����?0��y���D�����~&�{��1���h.�q�4P��+�q����7<�bz`��o�ҩ�b��1z.������t2"�`}f�C�=hvP?|ʖKGt����m��j,�{z9�b�}�_��J�{\E�cx�
�P�.���6�,�C`�^�#���`����l+�1;�b��CZ4�<�8�-
�?����Q�Y�M��O��B�x&#L�h��U3	$�~�)|MI`����5�!����
.e�=Wm�&ݲ�H�|�Yf�!Q�'$P�:y�����P��ǁ8L���v�n�����4ɃRߺ؝?����Obތ����E�x�H.�P�>�1���.+�l)�"�˳��S��U��|��]=�M�!��C�X���1�Ք��ѳ�Βr(������hrb�B�S�R���� /�2W���Rmp�KG�m"ΐI�u	c?� ����d��V{�����X ��J�ͥn��?����jB��q6���[RK/�t$��u]������Pŭg��#�N��(�8���.o��n��v�J��cU�)�z@9kY�-��R���گO�n��i?f���S�w��U�84"������C��˝�6֝]�^ -���9m����D�,G��j߹�3�x\c��w�ߕ�,*6W�����:/����󨒫����OÚɘ[}�Z��iL�b!�]yWV�����,��3j,�R��юJ�&��<�4�$���D��F���|�)�X�ٽ�Wm�&7L=e{֭��q���0{�B����2��A{ߥ�|ŎS�	�q\���#�`�W��m=�gm=�h_�nÍ�H^�۰u����H�կ+d�ɒVm]�Os+~�+ sLI�W9Yx�ￊ�E����Ҹ��
mՖ�:9��N^g�pe4�d�fj����[Te�U>���P(u���l٦��.�EG�&�������2�m��C��4u�s� ĭ��!�l���ǆ&>@;���E���,o���X�t��$;Wt2h,�`�5X�wv�Ϣ,���φz?F���^�B�nm�����C�����Ԡz'��3p��[�>4�q0��6�GE�^���/��1GP�Ъ��Q}C|�"�^8 �e�Δ���j��Y��� �7m\a�9�5	����d;�ă]:�Ȟ���J�
Z����Q�l�����e�S��-p� �B�(�b{�aK���x�C���J���N�� D��w�
�V�u�I��\N�e�tB�/=��I8J�X�7�.�/@a�Ra���k�崿������l=�W����o�t���'�Rg����2y�|�K�*������co�kT�_�����ɽi���
P����>�*����p�0��Z	�2�5����A���������)q�i�J����	��@+(�@�;����a��	*�ෲ��bQ9 �i�y1H���*~�2�С���l�-��������J����(�q��)&�]|Q����8z$�Ê-�.�i¹k�"��Y~}�6�GDi�.T8�����y�띬�s����p�V�O z"5;7n�E%�簫�_o����	��ϡ5Q_�1vm��̳S�'���cy��6�Y�#�y�BZd�g �.*k���Ǆ����������K��C�3�?�r�K�d咃�1�T#m��bW��T�͠xm+�l'6�܎��k��bx�D����zGF���o���E��7]G��wX�o�˗�^IP<��=ip$"�����z��\�I'��^.M��
$��>M6-�ہEM�5Ч�DB�n�qhc9ɞZ�'8�!�S[� �z!�<oǽ�vOt���𜬏�� ,t]�d��S9:�D;O�UXdFz�1�a���0{l���6����Q��rFH���x�5���<2K��W��)s��3��8Dk����2� ������0�J���o����Q�H�K�=�k<f��B	��8害X���_��t��K�foW���"P�GLް0��Lע����a���!�Y�䵆EMp2h�w�=����Rx�.���O���i[lt�'�����ʋ��}';�ϒo_iw!��q�^��r)-�0O��X����9�$�UV�) �ǂ8tZ
G�Ql\Dv�`0Y1��f�D��VE SC�.0����_MEF�Rf��]d����T��QmZ�.�ݝ�%�J(��MLoz�U��D=W�[F����M�š�v��y�R��\ �o�p��&f	��V؇{W�z�v�A�xd���ډDc���c��1﹑돹�儴�[���Nc��{�x�'���kC��-�ߺ}��������g^�+��; <**�����̟uu�{SI	8��@YJ�.�#�7X{�~�����{Kd�. O��7��m-˾�0x���L�f����})����|�<0��f'��In��J�$�u��F|�E�m���,����}3Da^��fp&�~u��'Tlm��/��h{�Y:o<P`�Q��1e����+��rkW&&G��/�Ւs|U��M�6���@7}2�L^����4J,@��͏|���V��į�BH�R���'
�dj�����o��,xbwӥ�)��xC?B� R���o�M�cn�w%RU\�}�5h�n�4����(8o�/eǖ%m��~.Y[��}f���py�/�,[P=�~��{x��U�.�)_x�Ã����7V�O�.H��62�����ϓ��K/s�<�=|5!����$2�wȀ�t�`ʨB��=N�R���n!�Z��
Aw�Y �D���׾m��/WnK�i*�^>H���3'ܔ�JО�n�l�TkJ�B�#h%��C��=�۠k�����uy{�Xt]��@Y�ޣZ�Iu:{j�,$j܋�z�wv�	ǜ�{��KyS\������x��#��#�wSu@���f#c9������I�R����}R�j�k��X�&�����D^�)]��ޫ���D�d
���K׸+Aw��ƴR�_���쯩~�ŵ�2����ô��:�(NL0*�h�À?Z����	QDv=��Ð��P��`�:�h-���šu��۝Ɖf��`�y8/m�(dn9c��-�Bk�t�5��f�v���h'�������;�B����*Jش�Q��4e�W<X?��ĝ���P�ܻ����N�ӱ-�:�V�r��膵҉QNi���E@!�m,��bx��=�{�Ŝ�dN��|�	N��y-�H�]G���a���l�F ���C������r��fsN�y�0�+���[���yA4�+��A�R����d��f̠�8�86�ׂx��:G\�m�w��#d�S��F�.�>8�u��:�����qH&ŻY��0�M�� q8NoND��G�=x��gT��z���ݰ�T�e�}���	,�M���l=������h�4Ps��D���0}D�$	m�tƘ�*�xԓ�;r���v��ı��
��R)��Q9L�cec$��D]��ԆE��2wo�X7� �k�����FbSr��G^�H�W�#~r3�����_�?<������|�0����U@�j�q0C8��M�/oH��Ȍ4Nt7�~~�~��o�n��
�n�+�w �����L�{NƦ���,\ua�v�'����x�̸�� ��7�o}<C[��i�=p�na��#�)X�QB3܄��g�*�{����%F*�㱽��n3���ԓ�-��$ D��s�����n������0��/�b�����3����ۈ�� ��@���tu���)��u��.�����8P�]}�-ԙ�%�`��8ػ��/lm�L�l���ȵ8*�!~Xф�l^�/��_�\�'�
�hx�>��Pg>��ݻk��
C��`�V(aReq�7㮞QJ���D��m���T�ʳ|��:� t���a�8�Y�'�X
v'�@/�	a�g���D.~�2
�i$�_bX��d�����HF4[t�M�P8V�o��k�&B?��\�׀Tw�.����@C[Cj�΋L���;,|q#�Ro1�9ա���=�I�K�z#�,�>˨%8�T��w��'����<�zR*�<U��#���%�>o���(_=��80{�iS�1�{�9E�lri?����k�I�}���}�BA�'�b�媼�o�8e.i���m �x^�e&J�]t�j\KDu�(�N^7u�CS�\�7b�±�7�m�EB�y,�!���ۅ�"���?L5��?��G�_�;�PI�5f��(B�ٴ�cw$���M�H�K����O��Lԗ����e��u�� ��f��3i���m\?5.8!�H�`���Gw�������	��(�L�`�w�8ƅ8N����0"Z;���3���p|�'���œ��*״��x�X���I�]"��l6�%#�����ʠ�3��糔�g?a$�t��bť���-��Y��!����a�\5Y!���q+�. �\8���˩r�c���x�唵�g�&��� _�����A仇|��Bs�@r�����ΰ<sN��nY��Լm �m�1J�������$��_���Wf$b5���Œ ����g��M� H;Ȍ-D#&����[��[�q��d��� /q[�S3)��2��=�� vM6AJc#DAc'�6�\k��ø���Vغ�u#h`�9V�����e�i�{��>�;�^��葏��թ��8��x.]�R�c0 B�����>�7���<�B�u�l^ڙ��GH�yyz��/?�j����pn�Xn�1@3
a� � H��+%�EUqt�@� _�i{�LoD�
���*�B�)�G85�g'���x�9)�]q�8��)ua��>������
���ȌP�lH����w�~�Y-y�=�d�����o�/��g�j��q����ꏙ����7��)��5-1��a jh�N 1���t���� �	u�z�j�U����fN���w6�(��,ɐ�"J6G4�8��IM�I��)���qqo׼�A���9��3U��I)��&��?`$�L��3�A嘭���A��7m��L�B��k�WW�b�CsX�����@��Ҡ��L�*AJ�/�M�]�Wk���;_!��X쏕�����L�Vg��0�g:��R)�h��	$n݇~�eڵ�o:?78Q	���Ϋ��� Ʋ&S0�W��Ȅσ��� �]p*�^��X�bR��1-E#�?¯����|�*4۷�0÷n@,�aA�~�*�_�6��
��@��5�6��O���^
�e�+�m{����Nm��������L���W
)V��;����fGhY����N�S� �n����Ef�?ν�#%E725��#�"a}ja�Ge޲+:/��j�Eh��%����7�P�_n���A[.�Ť^��n᪗�ߡ����q���/��Rz/��G��{ę,a�ˏA��{1�#b �BP�L黕O�2F*w��P�-b�^��7a�'+Ԇ��

���]����O���������&����z=#dV ������e���4��+gC鼶V�i��v�G�f=�\���apb�����wc7�k�����Soz��1�e`Q�MW[kZb��N���k,��0��zD�՗�	A�ǪN�����XS�ɬB��?-�r�r��lO��*������1��hm��W� O�O���:8��8�-���� q��(җ�P�T	�Ť *e��u]u�S�E+���F��c��i����� �۔�׬	��G$����0 ��Af��5���~�����.��(��L�Y�p��jԵ=��b�(�eS{�8�!���:#U�}i�lQ����x��#6�	��J"5?�x���D�}���2l���<%��[f��Ia�疿�
� ?�~�2-{ ?�K�Dokz����������$��>Ɲ�2�e�	̛6��ś\fَ��ˁ!��>&g-�����`� y��G���ŀ���s���.
���~�6]�T7��Ǔ;Sk�����Ή������*� ���9�$FB��ۅ{����xH����s�b�����Yi1���R����1t��O�D�5�Q����fD�ϐN�Mf��R�I������n#"Ky������n1�K�(	�,����?t!��,[*���;�5�Y^O� ����v�ɾ�o$|��Y������Dz���Ƞt��):0�h��aQn��֬���Q~ʛ�;,,B����Y,Nk��͢.b�#�`����fZ�Q"w�9�+���U�V���l�C���ۅٳ���w����K�L����ԯ�^�u��f���\Z��������`�A����P��qq�l`e����ȳOj����G�Y33"��|�]���8��	a�-Q�<���2�ĎB8{�䡚v�����i0�_݇�˻��P78��dM3��'=Bl��Ve�߬?�Y�����vX6XV�9k�k�*�ֽ�R�n�|xF�$D��0��*]�ыj�:|wA�Ƿ��4���n�t�Z�D���^��ݢ����`��_'�y��̌nfk���sO�"��z����������������'��t��$6�g��!�8aѴt�$�M�|Х��P߆��J(ѫ���.�W8Z��B��l�
ŌM�~�oD������P�wJ�p!���)e�iէ��(�|[O���%B��ڎ8�f1���GQ��\e����sw�V(εM�C���sa
���ȳ��&���x�QȍeaË�e�>�'٪��1���q��nֿ�rnjdyT��.�/u�B��W	i�F]ڰ�î=�Z�m����?1pr|�f��GJ")��8ɬ@hz`mz��VA�;x�£h�\d�1�՞j\��æ�9���02=��*)\B�X�V�h,X�w�g�u��ʶ�NsxKz)�-��B&����3(���%�wB�e���;�m�h�WK��H?Ӹ��*�P���o�g��+�?���{��Q�U�T0��lk���+�yM!���bd8Bˁ��S�#�6���c0��|cE��m���(���U��w/W�����߿�����Ǉj�+L�|ГԱ��u�B0Z)�A|nߛ;���&��S��֠>zmԘ<�Q�._���׸�n�B&�Ԣ��\�=bҦ�v��2�&��,�9�C��������{�_�ǖ�SV�f��h�؝�� �*��Vl �X���w�v�N�;܃�\�{׼:�h7�U��'ʄ �0����T?�/{��x����|�8+ ���f2%@��
��@���I�����"D��\�� 0]�3�E��N�G���&���[�о����������qE����0u��*>�f���甘q ���бo�A*9V��Y��A8'�;��0%��?���T�t��R���@�D�tZ�k�U�mg���ݬ�=���{%r�IiPS����f�o��s��I��,n�w)J��JT�
�
��[`/�:zd�#?i��6�,�h>M�_��Y�lG5A;��p�<W�UE�ʆ���l�#����%o�Ol�k�����R���-�Nb��Y3ڝ��K����F#u���B�z3;e��ƣ�mOpY�:,I��iG�4aj���O>.\��O�����h}!��<�H����⣝��ˬ-�֑3�~z��GӼ**�׳-�lxSE�2cѽ nd07)'O�����2$}e���c@�� �im:��:�ej�m\�� �# �)8QW/�u|c�8����ΏAY�O1�:��h�NM���P����������[��C�j ~:zO p��\�1e�j���}�Q�ǳ�d*�)�+5t�'�/��!�z�Eˈ�L�LSݸ�ϫ+VN�4Ǜy�o�.�9ƌ�-��q$"���x��.q���;g`�H`��9�4�\I�G�HV��N8�h��>%{��w �?��g�|]R��ȗψw�F������+UUC���A�\6��[2����ŌR��o�P0�J!���;�� �Vq�ɫ��qE�et	p��=�%l���7�u|J��N�H�K89R
ɥ��G�=Ii�r=��S�^Ӳ#�pn)�h�(�d���ɏ�ƏTq���� )ff)���?Gk�ÀɆ�y%��N �@��ӎRy1Io�P�!_�d��秲X��Wf`7,�:E��&]��l�����x/-�g�h�*��m�>�O܏��H��G+�<�"a����`��K������>~�f@�1/b*�(�2��`i*��O�)����d/v=q�0"���O�Ȫ�;IP���+����5♃�֋e���Z�Pm�|��48lb#�rH[P�����P�(�֞�;�"�<V�%5A�!��Bl~A�3��_��(�������Q'�t�����M��8;[zF��)I8�Ds�:�ţy�U�^��
c+ɷ�U�A(��U�=�L��w�����6ᒠr1B��,i?��?��Kz��{��S�,$�O*X�j��355ŕ�G>%J�r�}T�;���'\���=�,��{�SN�sDj��p�Q��ǀ����J�:/N9��U���򴱽�GJ����� QǦY��	�Oo��#y7�h)�?�@�&:ɑ��w���%���
G!�XF�1�-���&�[�����(��'Zz�^zw����ZX��f8Ż�CՈ"H�'is�<>G�#C��	�P,sg�cxe��Uͮ�`�ǋ9G�2�o����C�	��r�:oğmH��*�IfM2�oЌ��
o���J*��J��6Ӂ�*��)DA����
j�al:k��r��R�Q%X�J��	?���F��n�J���ӹ���_�u�`�����q�*�6��aa��

Z{y��{琻+*S�K�����ackLμO�K�&<��H= ����LymIu�2RF�������a>+�����a��������3��,���s6�7H> N����^�H�<�0�wʒ
�Q�{߬݂.3rY����ޑi��܌�S"N��m����"��왪�J�,~=�VT���5�OwR�� B�1PX1��k��x�'�������9�rԯ1���Rǘpu�j�Y4�1&q$��R��xz���WK\�u�������U�k�,,XG���T&-�l����`���)�$���a�ڐ]|Xi�t@P�}^�Uqs�����4�i�l��)�����vw�j�1���WWDV���*��p^|�@���F�F�^C�'Pz��ze�-#��&���R e途?�y�l��GH�ğ�2�i�h�p�e���cH?r�IA�A�5�$BU/)(rg���ǒQ��Hâ��R�<D�BW��⦘n��7��,9��0��y�u6������L;T&�l�|����kώ��W�����x��k������Q�@������j�Eݼڛ���zI���T拟8L��7FW�_���$A���Ɨ|�L�n-`n��[t�D�_�'1�?�c���=��9��m������CN�K&*�M66�sX�*ʴЎ`RGƅ=X�o�����N�ٮS�T0*���+Tn���
��L�M
>��j���8B�Y�x�����*'��^�24�W�D�Q��\kC+:��_q[��F�xF1�u���ψ
I5��/>w loXgX	bL$�w1�0�F� �r�j��~ך��k%��^@��:(��фoeʪ����誃F|��FBD��d��w�U����e���v ��1��{�������:��h"��c����H\_�>�B{�rf Ǳv���VdQ�O.	L	��z�ւ�Nw�"�K���k	P����(?�?��fz�(�(շ:��U�If�Dh�u5�d�Q�|����I!��AX��?��C	��A��=}^��z����2�����_��o���0n��������3�`Q{��zt�`j/�p|��6�X:��zx1�[E9����F雧Sk�E�_� ����Ҷ�]~`L�;5C�ނ>��
N��d�hu��|Ui�Z����h�n�L)BPA�G�@{|"������vژ���$�k����x��n��PoPQO�Yظ�5���c�������*�]B��QC6���V�
�y� �S=ŁP���2buZ{z�b�mU���p���gՈIJ`�ف�����q�f��lj~�,�����-�F���L J���C�u`��t]�E�IR�K�w��V�����:�P����'u��l�F��l	4}�]�vj��j��Ň�7�n^�U��}��
�$n�f��TV�����pw���ѵ�􏅯>�g�V�N%�I>��Q�q���G����G=�:ױ��q�����8�A2��мkRg��c%ô����nV�x��imۣ�?T�6fy,�}J��{�U�J��g~?n�T�1H12�IF��	~x�� ��� H�K@+�:�IN��3<;�5��b!�=^<�ԑ���G�_XIpUc�w��է�0�n=��/RJ���O���X��jQ�"����Z�vֽX\8E^�?�q��cV�֡���X�D�٠KΚ�b��=欕���U�q��|qz`��Q���6�"�X��u�~d�5l�h��NmH����L?��:����)��5���}*����9)��*QM�H��g��ޱMs2T�Ϳ�L�Y"&��#cYC��cyM/�J�D=ޘ	� /���A^�S����$�
�R_Z w<e�_Y�����Z�U������d�x����0�x��S;S�m��pi��,T��d1��v�|F�%u�90!�Z�0�c���u7�hK�����+� �a�ēH��)��V��pLzXd��i�ߗ8�V�L��qNf�P���G"��9!�����f�u�Y! �K6�q'���jS��ẋ�.�n��	�c�'?��M�@Z-��� ��4��㐶I@�B;Ȅu���F���fY�z���E1������e�N����l6��E��b��;n��i��َ��Z[8y�T-i"�D����e`N*'㛑�R F�,��S[���j�	���w�n[�n����uM�`]P�=�TI(?�(�`4��]r�퀐�N�/F?l�_P�L7��j�$P�@m^+�O�8�m	�!I�����4b�	��c�q��VI>O����K�%�d�s����e���e$�?o�ܙ����z
PP����R�ck1������L���m�e��{D�%�Ϊ�w�����/�{��{0zd}�2�T�F�Yh��#T��&��/ٹ���6>ܬV��Z�EOJ�����r0���Ц鯊it���M�V��#}�P�oC�DR�h�mo��=��ҍ�6�ܡ*����P:�J��� bD�B7<�NR�tT;"C:`0����1i�t&�/ ]H�8��$��iE([)�B��j��8&L��1q3Y`�Ns����ۏ6�7����z̖/1ѼH� �6��7����k��� ���'0�K^�}=�СB~
[�]m�oU��2n��"�F�ѧ� ���+�����p�9}������T��?Q�6��!�7�HHZ���x�z�j�}Y�:M�v�Y9��$�n}3&EDP�ʥ�M��Wةy��2ä�fu7�XDR��Sa?��J���qy_�,/��/�޵�����>Y����q-ǒ�{�5�Ѕ���p�[ň�A���4l�{�P����mo
�ᣛ��m����C 7߆}Sʦ���qHY��T�3���a��i_�y�Q%"vm]��3�Y��:w:$S��+u
�>�D
.;~��Ize'���Z��#�'U�+�f�4{ԋ3L�U�]+/fB�\q͑�v����Nv��\�7>2�p�{/�Muߖ��B>���7i�­����u#����DhT�ۄ����tk�y#e|�+���{�k�,�&6Сr�VU�(���D��J9F�>u���%�B� } i�|��1�� #udUB�����x׫�4t�5���of��-a BH5`������=� &�b�ي[m��|Wm_r�ϗ�+�~��F� g�.wd1�*��~����������o��sE�̅AɆߣ3�'Qm7�٢����]r���7�(mgM_�?�����0��i>�:���ōE�3���e<�����>��+�����&�ΎZ[OyOO��r�*�@����~��f�c��+.6���k|Gd�Ɉ0BwSR�>���_��R�����O{��8�0�"i�߃��XK��̬�@�����Y����������u� ���*5"�����դ���o��-'�E�C4^��5=�Q2Q���G�� i�$◫��B�ve*��?&�����U��7�N��t�!��l8��L�H��:>f��?nӇ�c�Z9�X���S@��{���kI�Æl�ԈF��_���|�����x��d����:%�GJ�T
>P��*_O�������v�!�0�Ln�\�O���ʂ��yQ7���d��6�w  ��PR�,_�:��[�����t�R�2}�)��O��6p�v���0l��&2�h��θxա��L��=��t�-K�k����Uu��tz9�I�V�1���J�]s��op�R����!?R�˕5�͆�N���tΈ������Q��1o�|8'��HF������7�1E���S~"��*��XK�l����0�@=ec�)�/MP��[��o��m�̞|�
�\:4|b+�A�f ���*2J��Λ�C���"9����oCN9S�>��X�h�P�����^�&(�>k�0c��[����& �뎠�#��/�9���=�Ť�!�(yzҊ����/� E)�b���z�QM�S��<��j_B7�	!����_��	�/���:	�?AA;���C�P O�vͺ'"��o�0�/G!D�P��5MB&(�@�{Y���L�[�+�}��'�䍉''���+?�U���܌P�Y��x=F�^��*b��"�{Pڟ������g�V��I�M��Fg.Vk�43L���O.8��kJ�5f��W&/z����T5G��I����Ϭ7���di��nZ����,:���c��k	��wR�� g'NR�gl�k�-��$~��l�䆦đ�Za"(p�y��r���{�����2�c.g�?��M�t#��r�4�n^�����ȅs��������f*Y�n}*Z�]����2�J��+�Z/>-�oyt�]��~$P��:!��H�zX�{��9�N�)�=�.� ��ͤ��,4��1qH�8�<�w~���̳
W�BU����3���[��=����ab���`&�PA���T:�V�C��mt zj�a�~ ��~E�]"�"�Y�F�r�t�MZ��ĭ�Yٱ�F%�{v��<���x����lm�N�Ҍ��-,Ҩs�w3a�$kM�,�U��<���A��u�(WLhM2�/6b�2,�	~��(��Q�ɨ�-ih�Ӻ����OxȐ�婎�eXu[s��\��8τ�D���)�u�(bb7�t�!�3�<V�DP���3T��k� ����ۀx��E,(g%:֩ �H{������|tO�}�㻲�����,`Q�J%��q�rHN3�V�_���h�Ē�"�n�tR4.��3��V��o=h�t�EysD��  �c�ʳ���o>�}S���+�8!'S<Ղ"@��-h}��F����<��
�T�-?ݲ�8���-c�'�k4���X�׬�i�uT������Dv�Eu�2���ܼ��K\p�"Q."�g�D"�wق�n�	�e̔�L����?%r)��5޽K�҆���ep떥�\�J\�� <K���Ś?��PQK l���vt�K�2���h ���iC<E�vd?<%�ލ"���Ρ����z[�]2��4!������3��f�8��C��;����8�(�W�W:���>���E�����)t��z���!���囪ΓkTvXg������U;p_����r�V�?&qŃP���{��M�9V�i-DKf�>�&�t6V Ai[��Ҧ�1sH�41���R_�JN�*��\,�s�V
�|��O�m�dk���T��>I�o�����
&��ԥ�E���"���n���*Ո8v�&�/���h�UR ��)��&���A�^���rv��&.˹-����ے��]�榦����E`�[���������i��J���~�ͻ7���:�g�Uo�L���۔[}�$�r�
_��8�b�;lʄ(�,�iw��6���*�W��Տ0�JR�jU�C_����C[E%�L���El��ȕ�e1�t�
��M��ɔǬfD�m��7?|'��1|�G���>���tN��_�w?�%Osh���o����ָ� ζ���7\���Ȱ��-s1֕n/ohx�nP�9�_Y�3B���"Y��;�*jJ��!A�e&�YO����-13�h���,��Z�-����Ø�">��q栩���~�M\�o�M����w��]R�/i(`]u��3���y�q����?�/��|�3����2��3X�>B�4@5�U]�ZQS�1-�j3ʞ�S��A��4��������eu0R�U��*$(n��%+qg3HD�N��e�lŭ+ߞ&�)��9/.����G2%��.`{x�_��c�C��ң7���O/���q�c�*!c3O��l�M�}��_����Q�%bsG �$EθHN`����U���ugC
�v�d�[��2!�Ż����tk����+tM�Ûq�Q��s��E���Ip���2k�Bh����M��	��U-wϤ��٭�9�����8o@�ǆ�nYia��O�!f��i��-�{q2Sյ:�@Ł�#��y�K��
�U���?bכp҉����m��̯Rl#��٩ĸQ�?��>F�v�-!�HפV��1��Ё����P���}����0G�:��!���Fk�o -�(`~�x�J�`��:pӱU�X]剾/���0��q;��V�s�%,٬&��Q#̧k�i��Td��(���/n.��iZ��<��8jd��Q����W����w�͋�T��w��;f��r�ͻ��E��;�j����%�_�/<W�o7��ҏƈ�S�i��v<�8�����9��aˆvI�a���:Ie�mYӌ�T�p�rc3�˗�V��5��Y�ʠ�]TK�O�����h�`{����c����Z��N�(k��4���r��bqC���H?�`nEt�IB��S��O-�S�����-^�Q6���6��iᬣ��}Pl���Jל�ϻ��	��ꐟ�'S��\8�m+o@�ue1_���Nqo�#�[?���W�p�Q�l���5�D'�����GH�Y����џ�>��f���ˇ�;���Rw�x�t��!���������E��r��\�㸣�f���J�2e���h��	W��*�� l�H,ب��c{QΗ�lR˹x� #K��G�������v�;�Y%�8P#6P���l.L���W�K���V�^C=�i/�">��B�MTٖ��:�dQף��d_�,Ξo	w���#	��[����֤j�[�Ad8f0�rGv�PJ@�ٓ��&�/E,П	e���ly�(|��f Aet\��`��2��� }M���)��hj�����F�NT�XA]O`[:��_��3̻g�Q��f��c7>^���x�@�6��~��Yo�j�v4�	��~����VǗhDgV��׬toz	kY:x�$a��\B��G��F!�7��:S���@����,�f�y�n7���c^�U;���!�kIO�7�5f�6Լ���7��ۆ"�:��vh"ӊ�YH't�ͫ"�� #W��u����b������>�u�D����"g�q�^��3�[!��\�sǍ�Z["j�A�L�e��M��H|FA�U��:�T��Ʌ�ӀM�^h���/t:Q5䡸T+ <�Vau{�ͭ'DT�4Y,'Xk��>�"	`~إR�����.��81�\���a���"	�z�	�b���x�7�Z�?fm���>)���D�_�d�e1���tm�6_��f�(5͎�3`�ۇ=ӿҮI�Pg߻��>ݖ#Y�u��aEq�9��Z �������3�9�%d�M��`D���KPH�(��q/�.ج����q&���5��د��)��$P�;������tx��D�[C��SW��Ū�ǚ�J�{��U�R�ڽL�^�C�l|֜?B��@�B��� $���c�!�۠�C<�s�Ds��j�Q�SG!z>u�C嚷u��T�6���U��o,�V6`��y���9�1?�!�3��?��z�B�e�?s�zO���t�mzM��t�x�����~�G;��Q��ͳ����M�<�n��~�R%xc��fSg��Q��!gM[�������s=۾�Ň�>b�|Ys�$�t�h�Ii�S�"��^"&z�}VM�,rV@Ǜ	�u,H�G&Eg��~nx��6�A��fth�����̌CǢ<���P/��V� =;Ź�1w����,��*���$��)�p��Pʨ $	����f���u��h�|��T��N=Ws:��Bb����Hfғ�v���~?���]�N�(Su�<�5����F������
�$Y5y���щ���l+��Y�5ʮ�,TΑ���M�8�_�����K�2ڢ�oЫӬbM�_կvs(�:e�s�vT���F�( �D��\�Zo �.�r#S��=�e�;y\g�v�m��Q�[$�?��IEl��)�����k�|}�_U?}B�i_)p�C�ְ�n�	e
Y�Ww�sy=���0G��ÇE�01�\U#Ow�8�*�,t�7�2f�=�ѷ��>9���:���z\96����K:��|?؀�%<v(Z�I@*K�jh�#0 s��A45��:�PXi�T,	𦫍�+_�,��ob�`��qFb�kV��(K0�cv.��
@�K�by��dc��@7�#ϡ��q�%5��E�*��:6�׿O'�z���i����0�Ю:,��ɕ�dL֓
�_��7�"��,���(�wC�k���ʼx,��6L��69xiyt̼|�]�֜��=�wy���cҒ	_�E8���/��������/(�����⾃�>�=�;��[�����K�ι�rY���:�Pxi�ь�5�望�p�1S���c*S!v/�t�wt�`'����5�3����q����0����w�sd%���}b���m�6�7��0H��vgz��p�G 6�|e2��bd�
o�a�H���۾�&#�6�� ~�9�{,����������\I�p;{� -�Y��G�N�� ]� ���3%�.~��d:@X&n��'>�eOpNLe���M1���ܒ���{�ߞԉ��ӱa�	
�l��[�B����=��`!,<��%�o�n2�s
EG����fx�$�8wG�ܙ�]�I��K�Tuco�H��w��B(�	���, *��l,�C���ە���G�z�(�w�V��{Qz��K��&��a��M����ܓ����<=��^�۠@5`���b��o�E�XRƐ䨫94~+<@K[ n�U���)�{pNZ�5<im�a���!>� .�kaگ��<qc6��p)o�$B�Y�
� ��h9��Nya�U/�%��.�5Ѹ�i��C6��'�k��gUc�qmFEd ��^S�'�Y���������ۏkzuD�FȘ𭂪-��q��b��t�����4D�cL^U �?�zH]�`n�>Ĕ_���k�6dYtvkr<Ž��vrbKU�<��Ցo��[Ú��S��LH����_� �;�Љbf���I&����_�\l�`D)]�ĵ�E�XI�y�n�cL}���$�&��9׾Ϗ �.
b6�UuҞ��>%/� %���i)���E�$����A���^-H3�Y<# ]%�㔿0�3U�.n���_+�3�(A~�k��3T�[A��5_�c�r9{�[N��|��[,�P䅂���-B&��t�6,G7�l=�(���b��XV)�\ܥ���[������c��U=�q�6�����G���)�l1)�Aqw��ʰ��Eb�x�b �`'4�DR�y����$���3`���rwIM�>E7{K@|�Ǵ�x�$B���sЗ����L�߂M�I\s�P��sg<�y~�vi_��Hodө.f'�6f�ml��.�ݞ��oݛ���븇���N�ٌB���-�??��2!0��l�2'�"�G�)��+JvA��=&�
�'D>%� _�R��< ������OB�K��>Xi�t]�k?����58&���Հ��+gκU{���������7�r:����8�c׫T(,I�
�͂�1�'2��d q�>�����6�H�J�X�?�/�YB��[SSv������2#�;<���BqVf��湎�^��J��.0/*���-��##3��d����-H��Y'�˘`����ER]~���6C�r9wŪ���`���+ׁx�{���N
ٱ��h��:�w`��9g�\5B���)Սk�j���E��W%��վ���hC_}"?�9x�Szy��n\N�7� P�W�uM����{�'�ӿ�9����*介����y�3h_��.��ۂ��8�Ԩ�6�/�քI���e2p�� Nj��
�6�	U���RǸ�g`�0E%fM�u䏭�;6}�T�Y<���)ô��Q��w��j*)�n5œ�c@��9��K��.� k5j�Ҧ���6|�bG��Q��E�dG"	4̗�ŠX���T��������,�&9��E�g��4^��X���@�e_�'��|VkL�i^�u��{�[Jo�����lz��9lZ#$8��;�"���# [�2]k�EKB��� k���9z���j:�v�'��;����V4g����o}3F�2"�'LX�Ь���צ�_fz�l���O�I�Zڣ��2�z����{�v�lr��D�2.=��0�8��W��}�����γ�i.��@���2J^y��"�+u�F�> ~|6�Tc�&i�-OU�J\�6%��"���n��Q�`��#��QԀ�۵��'N���	��8L�B?H�����_mpz�Q�˚b0^�<XaoN�H�le��?�=���Ŭ�tE� ���A�w�~��l�^m��K�kw����w6��z�T�ߏ�����RrQH�	���W�K�$J��矽q&Et���4d
w��c4~�8�ǔ�q�PhTk�w��Hք~�^~�����͵hU���"�ϣN��!RuNt��a*�ä$լ��L�:�b������4s�y�A�h��!��$�����Z�G� S�]b��A��ڴ�P���A������S�.���u���]���h�����>v�5S6�e�)����!��� �?m��g�ϴs�T��t][P�?O�F����*��h��:h�r�U�> `9e6�|�_�X�Y�M�W��Pq�9|:8�|o��<�Ɓ�]�_SZNޙ�F�������7oD�J<�&N���}]/��$m_-�aM-��	t����я!xg{o�,�KI\m��u� v��Z�ݖK��[E���7�J�mde��+������8�9m���\zs��W�� ��͡�����Wㅉ���h\����?)�i�A�iw�s�-�0�d�B��n��Fy�A�
�Bt��)fB��ު��V�0@=�BRn�T@����D�X����&��ݪ�������!���`A]�K�?/qO�S�ܟ��x��z䲊�0+u�]ӗnТ#����bEI�]�>��ee��X�=\�����
�qݕh��E[�׆�H%2!>$�2�ȳ�V�I��v�i�f�܁�-H�{'Se`�O>�ʨ�oc.EI�ɰ*����RD���"���S� �e�������R_�
��(���D�x����z��EܤU�6n����|vB� {Ds#�ʚ�[��T�"i�N�(*mx[��$>�ڒ�A�h��+��l=�F�I~?�}>�)-a�͵	ؑZ��#�5n�~~��g�F��?����pA J�����n�O��uYxh�r��C$]�2GA;�����y5M�X���4v`^�o� �ScFu]��/_cU��hU?B�����6Y��L�9���d����sH�9�f�l���q�N���*�i�)�H>�p휣w�����AێTE��j۝OQ��1��{Z.8
�h���3_�z�@����o_B*쥻^͌�e��Մ&7P���?H��ҥA ˗�{Wc8ܧZDu��X�պ�� N�υ� z�U$�Z�G����OwL�Na��`�V��O$W8t�Bw,f!�M#X�Z��x�kة	��U�LQ�j�:���N�A�x�e�@��#L�5�ѝ�� *pXCҚK㱑�l����v2����X��9U�
�w��zU��ഏǒ�8	���HT��#8� A>һ���dӠ������2.�6|/�#���e�s���#������O�lw��(S�g���:�ũ�ї;5�a{���Zz��E ��B�:�PDl
0�uT"�V�{�m���z�p_�=�q#������Y�&��o�p֠�yW�43\C�Rє�-� �s����teċ��WVuW�@����ۇ�pd�����i�8�,(&Ĵ^�k�ۺsy=oCދ6w��7<�:Ԉ�
��\�H/����e�����P;��6� ʙ�{��H�i �o�rz�f_��ib�
uО'S\�"ᑾ�C��'��}e�]OFyH�'xh<��mO1v�c>vG�j|�L��vz�:����&ʫ���t�	�,��A٬^�`���GDy�@����ϳ��ؘP�-��c�άp�VF�~���@�-5��<�Ś�E�2�����U7�<����E�Roꨮ�����Z�D��PL���l�y�SEC��%*�ꩇ��ϴ1S�����h�lL;)�Kن� Z���u����îdi�c���Y�h��Z�u|��kDnGz�����a�����|�^��t�,B�dÉQۺ�J�_���H£�<{�.�u��8Z�����y���ִ������.Fٮ�>��W\L��$J�l%|��t�c���0��`����֜<�g���`/g*���5)/�Ixp����J%�Jn*VCOm�桯=Ue}��cLEW����fp�m��C��6������_,�
=
m�[USig�嚢3.2�s�� ͋R�\qV�Ϟ��P�~�c���f@�|���*F�X�E��e��9�iOJf�{54�?���[���u_�8|�(GU�s�������oڷ����K%��=5%���34#���Ǵycc�0��$�g[S)����w:�p�]"�;�vu�0�$-]D���޾Z��=bϢ!� vs�Ќ��PS�4s�U�z�v��kt�+���o3��T�3��׶kc��� ����%�?�+q�	!��J�ᢧ����S�G�V�P���A���%�5���"l�Yy�&�|�b5_UM����\�oZv�
���x��D��vo�0;O�I�g����#��ǰ6Ԯ$�3~Lv%���2�O����[�E�f�%}��;o�
x��'"��˪ �'<��0�t�mv��~�.SG��ҳ��ÖشIx�KDd����D�;�	�wn�ʦ��?.�?�UR$I`���ݖ�{����3���T�����BL5�'�d�����\�v>I��(gm.�r�V�wd'�d������	�i�r�LJ�u�'�}�M�>H1�����7�Y�\*���>*�>�jK��R>RC@
���zΆ��G������)R���5ﲏ*���ڒ��Ew�}��=�LiD���t��s+�٢!Zگ�1��/ZѶ�E��>�Ⱦ�3��S��,J��:�"pv��%��CMȃ�y�g!�~�����쁽�X�*��XM�bx�'��y��<�B�]�cO ��D���UG�g\�Á���tm�*��Q��qj]i���ڭe�Ո%��8�dv�0E��3q"Ρ�8��,o���c�����d47M<2`}��Uh�Z2�>�B� J���*���T@{U�Q��J�Se:|���-�e����LOj��peˁd�?M��A�r����V.���Zl4���k��f��"�� Ύ��F,U}��SoE���i��Tʎ��	]j@�O\ThB}�xb8b�V���	�QF�.Ȧ�!k	�.����X�	��n�0M�f)_~��3p��ĳ�/[�=����H�l��	�u�$��g�Pt��#�[���/r�z���.z�җ[�d8l7�v:(�Ñ-[8��\|�x��k��܀'Mu
~�N_=��Ö��z����X����5����(�["!$������Qɩ��r.]�O+2����Rn�5%�V�$`�9��Y�W �hO�� � {"�ON3;��A����bU�,�7����Ɛ��q�Υ�������~p��dj����|�������|\���;�p�{��Ƭ�O���ë�b=���K���XqE
}V?�Ak<(�U
<�q}@�cX?�x�T�1��M���I=ڿ��ZA��&���9�0�?O�e�� C7��L���]�8Q�<��?�4�&P�P��|�*�	
	ǽ��}�9���7Y*�@�2��ak�{S����M�p������u��3���u��c\�m�d%�UK+��3j�{��*�59ĠY9b"��Ң�y����H�۾A+��g�����?���9AH��#�d;6��$b,�1S>�Osl�/3�����-���t�wE�w�Ե����e����ٳ+q�]�Ē �*6�x	6�&Ѧ,7�9*Τ"�eE"M��5�t��ER�q�
/�5�a���d^YK/e��i+!#W�+N���W�`�G�j|�[�Z"�㍸0�пd�Gg�	�+�r.���u��M�]�D�ʖ��A���{�q�2l=�khkp�N�-s�"�!-��\l|άv����sJ'D�꡴l�����dѱO`��"��W>ǂ?�L�I���1A
�p�d͑x��9֊����'iH�8�R���}L�e0#��s?�n�Ou���A��ġ*E��QP��tw@�g���$���v}(N��=�Q:,�4'��[�G! �����R�ڳ~Yr�٢{�^㇪q�f�{� Q���祴θ�y�C��ós�K��7�-�N�ӂ����Y��:��r�f6�x2��m}o!/Y��(){q�L�q�:,�8�6Wb�E͟�z���^�4�@���a���m|�]��l��L[y��\}I����<�i� y<0X��������jz��ѵ H`~��hBt�P�Tf����_a,m��u!�傪
�ke�A^Y(7�����n��3�R���'g�(�26s{���Dj�L\YNq!)At��J���D\f�2���fd=���A���-�֥��3�K�S���ނ2�h9*�_���ýE�m����R���x�_6��7�K��{}豆T�Z+N3�3����H�>zc�-��(����6%Re\~r�@��9��ytG��\�{��3��v�d�.������Wj 8OX�S���3�<�"#n�7�w/`�EE�w>�Dr��4��ABs���ӝ��w�z�ǆ����<���w�Ib<=�g4�ٳ|��TP}����ꪢ�a.�3�	Ayf^���7�^���x�h%Cw7q�J��_�7S�K$��`��Tܷk��ֲ��2��6�˯1L�(���I����i�KA�}9�f�����ՙ��W4'�R7����A���D��(���/g�hwk4q,��Qwk �Ү�EQ����T薏���5�dķ��e�¢ҞEx�WIN�P�T����y���P7�x�X�}�z��Q�E5L�*����K��*��`�y���hś��B �
C`_G����23l����.CҘ�~��D�����qK6�� �����dG�Y��+JE됸i>�W9!Nz"1Q����>̊�������/�į�����7ET�(��V�q��*�M~��� ����eρ��`�ј�B;y�O�Vx�Q�	)Ϗ�D�}m����R���O��c�^�{�):�oV�:��7�z��6����f"#���{ ���8���/��Z�<���F�V׾.�8 q̢ �'��|$1t�pa�7�o{�q8銵]	�!�]�"1�֮I�)��T`�Q�k^d�Dѥ*&D��x{��)�~Q�N�o>�S\�\���$�W#k�+6�C��J:%z(8�ћd���])�u�3� (� c�X�K���K
�R�%�}U��/�����Jϧ2���
0
%�:;��I���b5P7q��u��֖��$�v��!]�m?�p����`�U���a�"��nF�n����t���4�I2�l��*��x�,���-��LņX W�V�������t���Ȭ9�Q�_�I<�6���DwB!����(s
��7�qh�G@�|~�<!�㬨'�Տ*?�XI� ��#F�v6�.<�s�f��f�ܱ�b�*j�!v7�5��bo�'>]��j1r	�iQ��bĹ]���+�\���\�����!e䫲S���f�9?�km�q�P��H>eΌd���b��4Z^n�#�(P�?��w��s��Ω�E�ega��������>:��WO
��_��������՘6Fn��g�}��w�;0�M���A�}w����sx��_��,-#�uv�>���ʗh��|'m8���u��f��C6N��@/��3�k�p-(��tw���V\�������m�$�5}�U8�(��m�v�T��!���-p�A�w�:v$�eS�8�l�5; 0B�J���Xw�{(�(�[����'�?"�ؖ�#?��_(��0�C��s��W����h��֒��q5�m6��~��fw� �Ϝ�6Fb���R���KO��+	�$�H��H+�f�}�(���]�S2­� �6�C�`�v���팳1��&p�GS�wa� h׮���R�bb`R���ؚj�I�w6ٷR0x��T��m1f�	u^N�/(f��Vn�~y��/t;�S>�I ���r-��]8}�d{l�z��#�L�1܅qI���x����N1�n��|!ϐG�V�E\v�U�,A~8�0�W��-����V��]�]:�wY˫�/����X�!"X-#��J�#3�Ju�X�ϛP�l�hyL��y��i.�O��b�(�j��1�z�6��8͚�,m��ڶ;�m|xu��r�)s0�*x��~���{c
���t��H@�Yc<�dC�U{'�,?��������M���`N�q @=_WSUS�js�����1տX������Hn����)S�B3�(�󿖻r��t�é��e_�,;x�MV�X�=zI,3c�����*�%i���,��>Mْ
�-G���Ȧ8��n�e�X/���=��O�I?��8S�K�ؽ5�I��iyV i�4�6��tDr%�Sl�K��鰓�;�cx5}z"F�ST�YD������3 �����}K)~S���D# �mb��t�{���ҮU�������b2٢H��0[�]A�e@3<�z�?F> �"K`3CI�{���:����5��W������d�8�����S����(hՔ��^��Z��W��;]l ���w�U�E�T苌զ�2�HN��T+��SaC- �++��(T�s#��i/���jS��6k�4:aN�<�+)�&mS�����'y������z�}�_�I�!t�=��u�M���ܒ���V�u���]���F+*W�*PI� �H!��U,��ܶ�ꆣ=�CWTaٙnY��
���O<]�p9�Ъ�]�Z]o����վ6(h6\�
\��h �V����e.���WA�)�Q)4��)%B髉��p�*<(E8�Nv�����zR[��խJP������I�1t5K$�8BKB!����<��)>�%���v#��o4��P2W�|��8r:o�;5�
wȖ���&?+�G֯�����.&�(C ij;��o�*�5]�=�q�4���Η�qF�M;R>����f�� `vc�S�h��� 12���&��w�^n���5y"�jh��*����k[I|�*�a�i?�xm�wq����~�}�@*��U�o�Zx��Y��Q��ބ�G폾�N&Gk�߲�Jl��-9���4K���o?D{�r�7k
�A���q�焤_�k��=B�H��!�o�e�2}����* ��<Ý��.w��tk��uQ?ߪ9N�zO�7s/�إ5��.�&���5���h�%[>c�I�c*	�o^�㟏Ώ��d��'j�����y�e���i�7F���}� � ��7>�3�^������(1�l�}0���T���W�J�� ש�oRX�}Ȝ�OKxz)s��L3-��0��a�=Cd�� g�S��pE�cQ׶tC@d� ��"^e�����1ձ�F�_���8Ǳ�T�ē���y���O!h�V�.��]����)ї��*'���13AD�J�������M��x��&�(���u��B���Vڰͣ֩n:�����|௖�ՎƎ���r�Ͽ���d�I�F�y7*"V�x2-��eK)��ث�\=��E�|dA�o����vKn�T
�4�jxߟ�WKvT)��Q�hg���XϬ���É�̯�<7z]$K�z�TV���&A(C�SC9ޕ��:��p\�>�/ˈ<;���M)}9��Mr?�j@z�s�W�Ј���#����&]礈��}g�f�B^kk2踴���T��܃|��'���WkA��T�k2k�=��3S��l���o��Ʊ��K�r��p�-�&D--t���$t��j�##P���S���"�Ăa�[;�KǼ�;e��6�5��m����y�������5E|�+�iLF�Q����uO�����c:���o��5�SǗ�=��4�sH��v!8)�r�3\��\W�¦{�UY0�>��A��.;�����8����#b߰�k>��� <�`�����4)��yX�G:ܙ@zC�IQ�;fJaNU�Is��g��TG_�N@���eu�:�s��uiu�H��`����F2���o'������ț����t�K�����
�F@M�R���_���B�o7�:��6��!Ϛb��g��%�g����o��(Z�n�6���?��}Y�(�<����~Лu�ዝ�C����r.9�.`Cd�u�Z'�".��)~o]+$�Zl�=�4o(S誌�,��Y��d��<A�����h��b)�RR�k���w��r�A���Ī�Gv���5���D�|^0��%|��o��7�r����rtF�^�T��7� K�|6B�VD�1.�ι�-w
�� @�|L�_a�o�Zd	�	�pS.���`�*~��#7�'.�b[uE�^����
��v�,>m>���ލ
�_���Y���.�����*�P?m��;(�{�"Z:�����`a;o�Gza~,d��A?K���WF��U��	*i� �74T)�ǁD��a��>�o83"/9TI�}��:I��/��ɕm�Z�'��);�<NBu���t����M:wp�j�%�4�e�3���$g�z��ߠ�MBN�(˰ٶ[9A��B��2�x���47���:#ԯ�GA�k�hs�����&��1u�;�O�b�$�q�]�4�+�:��c ��������d��y�	�3��̶���vOc/�w��S�4�=2٧�h�7���!K=�KK�	�H�\��$�y�����]Z�d������[�,#oE�[B$ 5�k�)Y��(J-��;�Ա���p��/�?��Mc!.��+�+efO��:�8����ȉ4g���Mv�Y��ק�f�����J�j� �I
N޶7���
rT�����a��=-�Eޜ&-Wk� �%��fH�ޚ �S����T��Q�}�a��1uc�9�ҕ���'CD�FG֟�����U/�4�0<�#K���l�#�S� ��oy��}��U���A��iU$��fLh;�X̊��Q���x{s�h���s˛�i&b$�l��7�L�T�<T�X��m]8o�݉%E�%�[y�$�L$��S{��u$�&jk��ª\ #�n�n)������T����t="%�	��0z 2�K8�B��ԑN�>����|U�^� He���r�Z"�6N�%(�g�`m�������m��p%�D���ܜ]�싛����4)N-��Q���D3:t� �V_F�.�/��Xy��9�r�X��T�Çz$����P� 萗��i`�Ï� �==�����x�Sm}��&H�q��w,� z&����)�4������і-����+�@�p�dl��յ&F}�yRڒ-��1w�n���U�O[�����4p�����Kt/�� �{3��#�6�N�I{¶r�A`=V�t�9��U�i��:�k?�����V��/:�p�ᩅa�<q�o ����>?!����^���琦v���$"����( 3�[-qe��U������y*������nAa��� j�� ��E>�o�ua!%�[�ڼV�qP�yi���B~�q��嫛m�rvcl�K�I�߻o�\M��Z��ߎ��
B˩g2���e���q�ĭcq�~"%��: �He�L\�C��>�GU�����K�|h��S���л��.@$����O���8�-1������ �,�n������õ���p���Ц�����.C��oI��`��-��L�F)�)s�]�Q��X�=+4J��Rʲ���V������>#4�����ȁ�F�l�a�b�6?��Ń�͐UgBT��Z�.��FKJhGF�VE��m�WBV�q�e4����V���+v�`�C�JĶ%U`X�fA�`����=��'�J�R(g0�k*��]�FD��Dł+�5��f<��[���� �Q��Ƌ��꘺��͕CY��Җ$
��Pkv��
����q�q�:&����]���j��>4G��F�ca�⻍5�k���������SΔI����T�_ B�ƽ�>�y�i;M���FS�F]a��c8���5u����=Z��P�����u�3�5a����zĞ���b)�i]�@�"�q�t��~I�%OC�V���0�c�D�Ģ��ėFM��X�Q��D��#'�fX6%tQF�Yi�|��i��``�[E�v��.nv&�3���7c��Si�b7�0{bdo�df����AD���I��;�Cꥒ���:gMɦ��4�z�U� �^b2�h�0I��.�<�(�7r��{��A�"��F���g��z=v���J x*\yi��R�jbSئ�,.��,�;e3���4��7��p(��I�5�B���O�����L��x�
�|u>թPS/�E"��<Tl߆�����ė��� ����W�)lQ��W�ќ��R���<& ��8�\�������bJl-sP�_�4
�Ug��".�R�����v�Mɤh	��ч}��O��^(���T�����$�y�)��cT������8)�'��I��G/�`�ຈ�僵{r�௦�z�[��.�ccʌ-�fX�5����S�$J�_��Z��Ġ�\��m
�f�3���?w4j�M���F�F/8��4Z�h�(j[4�.0-��Y���r�ozhsg�)N(�:F�D���wG�E.l_�������]��\��5�te�����Kr���|j���#�3�I>�?D�"l|����7�<<w��Y�v�D�fVY�Yʽ�3���5?��$.	l��#A6̮;�@�r� �gV������tU{\���>,�ĶX���#�Z|�;�W��w�"�X�|��n���9��z��bdɿ���C�xX�	a!���_p�i�g�V]^�f�:&XJb��p�4�Q�^7�$"*���K�:Ӥ�^}+YLcճA��G(҂YO��?W_˚�g^bxRh�y�_�\��?�kAX���u�̸|����2�^�4}߉G��f��W�P�������r���x'���zk����n� �~g��Y6B$oV\)R3'd���{f E�������,��	1�<;q:�~DMw,�=��T�3#.R��²;1N QmU�Nt�z�dzU@��%��U&U/ �=��L�.(��_��+%�R�1B�lI�!�#()h�a�X�4�}bu�4���<��Sad��-걵���g�k{� v��������Y+|})ȞM����)�Q��9h��g�G����#��&/җ�<z�������b�',s���PI��y�1 ���-��U��|4��Kne�,A|��>p������=�/���KISrք=k���!�Su8�U�}֛]�#�+�촲�2�������pJ�X����Պu�Ywr�&@v��'Z�x�P��B���\nU|7��あ�a��u8f�ϐ�7=V�V�96�;3a�����+%B���,���8��y_r�6�!���u�U�,���Č,��-K��vK]�\h'��U����GvLNC�<�~N{L����yC&�K�U?t�@������_�� YډW\Ð��ۖi;����>��_q�<�ԃU�,��_�d;��|��UYAh1���*��6��qq��FG�>���f��W{�L��Wk�4p���3O���s�<I��2���C�������x!�t縮��
�co�]rJ�0�Q�2E �x���o��k��M�W��카�<�=����9���]���[�o�+�� �m$��c�Gz	?�qc�D�y�^gqĶ��c`F �_�5S���4س�H��4�n������K���D�,fQJ�8�,#�V���Ce�ǈ�@em�2��������݂�����m	��Kf�[.HD��8~�:!���07���e T�&���uN4�B3g��Q �"ᡒ�{���h�;�{�!�������^�ҩ%�g��xrj+�&[eLk.g�ΩR@�ZA���3�U��<-��>�|�?����	�mw����������
LW�V%�@n�3� ��4�6�S�z�
�!3����\�II��~cp�ZK�bV����'�L9oi1N�uV��l���� �^Z`y��/}�-\ҳ����`ҋ۠p�';���z���g)��ڹ�R:��ܪDg��{[���Ӷ�G�+�� { vs�2[����\���<�&���Z�{z����N��[&����}������,�܅�9_y �����~�v#�Z�N�0P�n+	mv�j�)��ؑ��H��M[-�$��˳��c���71k�
$2c�����{����M���b���/g`Q�&�o���Kx~K���OPI�H8a�r�%>�sC�� #��h���)�4A��~���G�}a��B�H�oKJ[��&���@�V@_#x8A�|����=&�}�]�#��
��YjzWfq�;��@���ZQ��Z�en�F��Tw ݿ
�G�[��Y
+yht�`�!�.r���G��sƴk�X�!=���3�k d�a�R1�rY��U�}��3Twb7u��%D%�6���:Ɂ:%�u�KO
�����Wl�s�˿�q���a�H�Q���SG�W���@9s�]&C/KEGj��.�ԇ�'�k$��y�:>��pd/��ab/_����'�C2���^��������������q|q��� �l�nt'`�e1�4_LnY�T��Ӕ���B�C��m4	�m	K1���W��ˬb1p�6��8S@��1"������B����K]�;�������5_���v
Xb��W}�b���wc����j+�v��������1��\�Q3�\��=�s��,��pe]�I�O�*������\�Aa|������CR�6��������`Y�Tzȹ� ��0��{�n�F��h� �g�R����������������e��������z�ş9�-��8
�l��o���@����hzp.���������g�Qj�n�N}K�(�Y�����{G�]�߭�V��_!�2�?^oG����-���=��⭟g'<��� 7	f43Ο�B&^���Mr����BKv �;ϵI�q�䌵��"���^k� ��v���Px�B.*�K�PW����F�2�Z����fU�HZ[�	�T8ݢ
�K����E��h;�힞�$�g=r�p8��)��Wdk􈈗��y6{��ͩ�b�,k� l�{ʤ��ǵ'{p�q��C�&(^�ABv�[�sq@Vi�N��'kd�����0V�x�c ��ˢ��Rr�JD��t�+5&Ln^���dٕX��I	a�H���L-Xm�ߝ,��^��y4����t��C���� ���w�5��E����o���՝�$
�'{"\'#����x;����
N��j8�Q��*<�1�.�vj~�xc�<K���v+	`���ԡ��~��S���!����4�UC�Q�U�+��M�,Lޟ�o�J�)�d|�jl�B�+��3���+�k�Q��Y��%;�{�>��eu%�0s�S�K�جТ�/<��6@����X
��� G�T�|���)@\�춳���[} �����;�q�:�
���6��PH|t�Q{�2�Q���wd[�#��K�R��Ә�#?9�uC^.�Jƨy��F�i��)��W�=��Ʀ��;����2�0*��i71]��1w�����s-q���ux��J	GmX8�[7��k���^[~	oC��x�ߩۇnq
�+r9?h��B-� �J��v
l��_qMN�&��F��>���?���E?�!��
��9���s���@��:uX�[+f8=��'!ݮ��z������N�j�������-�ǐpI�hţ౫E�s7R�z�T(�" C=ZЕ$�9����ރm� 	V}S�@.��k2�(�8y	kw�0d�m�nu,~�Zx}���+���˟�w��5�<�Դ9� �P�R�c(2��?�|O�.02qfuB���b4�K�N@GiK�h5���35-�V�@� �X�A'�Jc���TId�s���SP�BQ����X����$��_��'�F����̓ۧ=�w�P�w�;�wa�e�O]Y�U�Fýɗ[��e�ih�**����������1�T~�z�o�{d�b衑�3HT�0H���_����z$/��{w塪\h���97���|�[��͜j���FF��Cz!'6W�p���%_,��*-Q�/�����8�!{����ПN�����7Aaݧ5�:�zqP�S&��r����������ߝT�.'�ɋ���Q8��p�%'Rv̭�%n�b�1�6�V����Ȅ~�B~�v|5`�����ˆg���U�ִ$E��F�irx�5��;/�_iG8���:�r�=�9��C2��W��p��t�!?̥�tC�d{���f1ˀ�;�0rR~y����:Q��� �̈��Hc�Zh���b�e+��'-�P�~�#f�T�꽊2-S��M,f�:=�x��Jjx����^�gI{�(ֽ�yf������%����lc��8<��#剤ĐY�3�����އ���!S~qN�m8y���y������O�iNv7�wn\w�.B���R�K��ܖ�ҨEQ�[~�P���ι����4]�x,�}�k���F]�7!A���������^�<H[}%�I�E�Q��	�Q��9$@:ҫ�5K�c_���d��>��~�fe�d!��N��C�������A�����Lm�d�P�Z@<
�����򫸝��&���Y���@����ʪ��F�M����!�|�Y3�/�@��0@d,������`�ڧ��1��[L�"O�a�V��Oj*Rl����6'㰍+�.��*|e$��C�+�����<��n-�$��ajf�y��j^�0��0�M��Z��b�9���&�P�U�B���9D���Ʌ��V?^:u�8��-)+	�0�6]%v�c�k�IM$���Ʃ��)� Ǜ>����8�*�*dRUܷ^5:�cI��ȣ5A��~El���T�e⦊�����ؑ����oV��5C������2�/�����fuc�>t~���Gl�Jo?�t�@g�L�Ge���fQo����/��ȇZ�k6RM���ϻs���@BL�e�zU-�*W`T���w�����Z#�D���o@�8��#�N�(=ӊ������	?���E,�݋�th��å�+�@cTH������)��q?U@^�-q�_�}�� e$�sq�U �)H��T��`����+�hަc4k��4�<E�Jy/I��$�Ky;�?0�<K#2���pƳ2Vt���� ��ܪ�뤔&n�U��yW_FU2-��[i۳.v%�J�a0�@g�4�p�>_.! &#�pҴd�jn�R��0�ꈚ�х�/~v�XW���2�#}j��-C�L`�Ĉ�v�^n�@�l�B�}"��g%�<{�p���[B���Uos_�s7��*N;�O{�)˽
,D�Ny�ݻ��i产<n�j��}�4�����)��{�y<
_b����M##�0P(��5nH���E۲#����\YD@YF�K���ڙ�1`����TJ�( ]m�MnQ��5@��>�1����﷖e�`5� IEI�K^in]��98�����c�Cۼ��N=r{=R��X��Q����P��l?�k +�9���m�r��Q�k�4�c���`����l�}���a��
�c�z��� G�p!�����J���O3~�L����[m��Ӣ��˿���Md�N35��]�YkB��@0[s,e�й������8��bp�J'�{j��4u ��E��Pq��U����j�,]��e�bp��VI,'�u[p?3v̈́5���ԋ�f��ͯ�m1�n]����X���2�r]�xi�-�]�)_�̱%*�$]
4��}���,��W�!���H��	΍�ȳsq�^��E��73F^��%%q�Q�Q���0��Z&g�`,��5�fT��^�W��0�(}���������>��d{�KF�3b�%P������s~���J��^�L���JB6��8�iV@u�WO�	��B;y/jh���p����`�{��̞��c�7�"� |XM&�Ûκڔ�si٫� Oj"=>sf쑀A�GO���۞��~�Ҹ�d���L m���jK�T�J�%
�nK�'ZL'y�� ���V��s�^�(�V.�X9��GDG��K�u�o��Qzt���6)���w��~�={<��.+�dp��5=�j5�������+� �/?+щ���!~[��ܶ���SO��g#̧H�#���Q������������u�@9��1�Y#����Ύ��|�j������u[�|-_ �w.�ܳm��U���hd�!�<��s�\)�3���nϰ��D|)�	� b.�at�_g��zHZ��}b����OX�M#_f�)��&J��-Ld��Z�i�E��I�yS8�T�u��d�g�T3v�ĵ���̑��L>���Qdo���u�	�ZSr�5����\�%��Ց��=��=$I�1�Q�0��K��,���e�����.%��I�)l���#�kg��-b��kwR���9�
��>K_2���l�"WU��ﻝ�`��Es�;S��61S�3����l��tlj��S�:w�^���f��x�!�b�H�ɲ"�"�١W���a���\��� 1�AS��L�Y����!e_z7*B~2�׬�C�dB��9�j��50�}!�Fp&0�D2��"E�*�F�=v����JX޿ڲ�z��&��Фm��*��#^j����8�8�֫!�nr��UvB$���.�vg�a5ԏn�XdP��w��E3��+ܙ��v}�$�:�!�9t��f�.` ����%�������=���	�����so
ko����l�N~U����/8�@��>�Q�k�����V�Y�||�����R7�&O��K�"�����}���Bx<�����_��O#	b���X*"��򺫬/[��{&b�4�ˎ=�2*�'A�]��F��$sCc�<��$?��*e�#��
���
���eR&��uG�fC;��Up 	��o�5�/z������q�щ�����{��Y�����?�X�t��+U�_U�N���+h�8e�/�ˢ��!{�\�G��X�Đn�nu��1crT����� ׍}�A"\Ƿ�8՜���V�֋��\d�2����a䨥 >���U�0*���|Z�M:�14�J�^�~�I�b2��C��o�rF�ް��R�����_6w���G��6�3>\+�C+���U�9�t����� U&ӈ�h�}�*�󁜷>q{�_h�>�FMI�MC���Ԏ�����M^����je��ۊ�۝���+� �	��G�^6Ug��k�$^H��Y��~(����`K��_�ulk-����f�rb�/�Μ���?,fтg�g�"�ԳJ����ZD�f�Y�P5�)n�����w�S�E�?:���Ɉ�9�	����3lҪba�Cz�����S@�!�� �(���ʌ3S ���Oo$ʅ�6�,7:�\���I$���^d�<ՠM�~���pI�+Ĥ�]��2L�' �Z/(�o�)J�kn�s�-��X]� |���e���C����:m�K�p�!��v��o�����%8{x�]��K�����~W��~��ǂ[�\+�g�c��8�NWp��n'ո{֪���\|�#�ʫ�i�R5��{�;h8O�+�{�A�x��Ay /@�Ѕ�qb=W�E�O�7������Ns��x�L��-§�ν��hQ�pFQlb�\�&R�Ξ�`��پIu����`�2���j�p�YWM~wf�7pM���p5:�יvA\����a�_��q~G�g���GG�!HFa#EZջ`$�ʗ�"�):�9��/��\���a6����Ӛ#�q�Y���Gv�jtd��̡ЗO����Q@N�哄�h��3��u���i�>H��ʩY9�f��˓S�ne�o���h�����;6��|:�S�`FDp�2��T�p}c��$2�\�Zi��r�e/�_��%'�H��=��K��p��"�񞀼/���a!��b?��)�qxq'�S�C�����c�<�'��l�����B�)�*�|+H��KҤw��ĳ��c3�d�Pe��c-�&qh��(��%�5�(`��w?;e�.n�V��Ԟӱ��D�?�ė~����xe�$$"ƞ�0퓄Ρơ5˥��>eLw�n��-WW�l��R���nGŨ�h���MP#%���Wy|���B>�����	:�������;��2_ȱ.{w�����꟩����A��v�b�/,fIK��V��l'���&m3&p���1ʋ��p!�� }�@�m�fo.������sh�)��s����և
�����a��� ��M�VA�'8���0a���jR��NGw���1�T�M�� �	���5Ȏ_��p<�T*��(���2,��(�>�1 �J�
��~�+�#I�y� �w;�ŀt��{�Ê6���r�$��}]�H"�Y<��'�h��[@ ĝ0QN��g;�n!�>r��(��'6����È��+r&�3GQ���rG��h8i�z��\k ��ӁGk�*��^����9X�I5^D"�i�OVb�a����eGշC.��=��Ӈ�N,�J�cy@��>c"rt�2�A��Q�3j�A���`�����t���'
.���T�`8�Jwt"�e
����&0M�
�@6�f.�k��OidF��J]/[B1�XZc�oL[�=C3�Ĵ�$��f� Ё���38�ޝ�>"g<8pbx7Vr��Cn73Kz�W ��ˤM����]��w��!����^�����w���yK����t�N;_Ҏ��~?��4ث��;�5S��ˬ�j㞲v�Ɋ����j3�W}�2�׍��3v�m�%�(���4�=�huNr(�A�x�5TN��k_g*��Zw�.�R����Py�q���E��]3T�Q�H�e�>�g�yz�-�������eV��y"�jf _&��YL/��g�Iy��ɲ���%�/�X]���(>u����u�{DK+�mT�*.�՚���/ۃ\� �Z�2�Dk�*
Aa�(���kq���u� �A��W0%�)۞\`���-����#��L�I'���vƍ.[<�z��K.��q���A��F9Z������(2�
m����U�mR��::2�Q�+��|rFV����v{����UNea[�lA�t C���2��?>d��)���:-(U���¼�a�͐񈓒���T�1ŵ9����"����W�����Q��e��π��-y.��rѕ�d�Rh�ᶱ�=��i�ۣ�n�����qwV��\�r7�HP�f����I%�B��ޟ`\�!���Ћ~�)P��Z�����9��y���
�)�g��-�=�1K&JTKţ'_��a*ш"!��U��F�4W�3*̬�i����w���jj�ZejBҠ�/��a0�Nr�Ͷ�"U�]˪���t-؏�`')�"-w�KX!unQ�LgؒX��Z���@c�FZ:��U+��2t�?�De?��%��4�P���p����k�2Bwm=�u�i��zu��
�-Kg!�0ę�Tt%l����-9����a�Ma�
�5�I����)���L���`=czoF\�k���ﮐc�9�Tp�x��~�:V���>�0�e�i!�B\[��xԵܶ��U��b	���d�=v���k���za8�����,���q�#-�j��73������=]{p�5F�'�m1k��``S|b��΅[�y��R��PI[��������m���T\�������4t4�8�8w��f�ٗ��/^�ɔC.�\���?������/m���7���o��&����#n)<@���w5�b֊ek"�w�_��s���[�+�U	{.�]��0hxI���(��L'(��,�k�닔4(�g�#��d��a5��bzǱ^d���G�6KLXO�WkX�C��c(p�� ų��x����X�Dg� �5!ݼ�8Br�"�=E�{��@�&g�
&��Ǻ}ѵ[��a}<�L�T��#����q3K|ګJؾ��}��H�h�3��CC��Dɖ{3����U�,}�����wI�.�������2����޵'����ݤ�Ԛ��k�[�Fr�@���Ǆ�^Ƥ�J$��>5q�?�<s ^�߮ӳ����K
�ʚ�vf�X�q^���Ih��o�弲�e$�.�&15�~��� �XLXF%�2����� �Z�NLM�SJ ��q�]�f/��/���%&�_��>R����2M��A,g�(� �	�c�ˈr���T�G��ݜ���$�o"*�>�Ёp{b8��R���wS�m���&��gN��
�a�Uu������,s�|��&-��l�Gv
S�6��ӗ��>r��e�n��U��>��(��J���1��$�����l��W�Q������KCq�� D���ۚ��r���ҟ�$�#Y`y�O��ҟͿa�	���X�]���)O�Рa��+k/2�Ւ��4.kAw�R�L���+���6d���o��*J����F\H�,.�����:-�ۤ]���ʬ�%��������h��ՕYJ�Ʀ��n:nel�+��C<74���^=��{�������S`�v�[X�%���帕�\1_/T�ɆhO6�!�7���O�yn"�&gW�P�+���!��nCx����R��f��my��C���&=��%T��{b�`w���?�As�*Gc�yu,έ��A��0�a}��zw\]+����2���_h���>�ˁ��o5�gZ%�(Uc��0P����<s݌=]��戈:{��fY	n2���
����*H�>G�4��5_4\��'Y�с��pՄؗU_�9�����%�-�g�@0��
�wG:c���7-��`ˮs�䚃����-v��,1�7��ԏ��jg�S\��1��wޫm�I�v��a��ԑ��ݥ���P��G�03�2��N�ĳJ�x��vO�bj=6 �mcg�@�*��8͢� ��w���OPP�^�!ujE�q]��J8�*.�3;��o� �Г���:,�{�ǇG�z�6���k�(n��;?����i.r�7粥��D+��+�|N�pٻ��Z���+�(S�(�_
��,�|��g�`�y^��djw����3��9
>���A�ݨL.��K=�&�(�\�kn8��)�b]5���oꁏ�<0G����W�P�8�Lu%�&\�V��d�@�n�@k�9�ث.{wM�k7��٠�p^!B�����9�W!�����:M��+���`Vq��j�w���@O0�AxtSOF�Ay�N�~_S�x^]F�vP*�TZ�:�KBvX�(xp��z�j@`j)h�\��mj���.�"M����qW٬4l������M�H	��R]���8T����v�/���DO&`H�vL�Uj\�\���pD�:le��IH�a7�����Pt��w��ߺ��>!E�
�I$�(rh��Z�*�x$e�L���I�YzJ���hqֳPD��c�H��]�ĥ�l\*J�w�~�3�у�M�#M��Y�С��_�����ѻ��y�U "-f���աJ��b;��7oPN�=(�7h����-�EK�شq/'$,_�?�arF]!��{6zo���W�≞C�&��8�����!�^�V��m�*$ڱe'yc2og�/.���D}�%�i�a�v��GqQ��q�n��Uq���m�� �bs_0k�i	�7���Y�7��<��\z�������y��4t��/|/hA|��mZ�"�\�-yq����q�C鉌�B�ZX�����S���
^_hx�=]�펿&�c\�1�^:�=���n*�C&�*t;�t��NUv�y��C�y���$�}ҿ��^���e ��*4��7�AQy}��'��eYT����YS�	���e!˫%O�It�$�3��%Y��ؙ�g�g��7�k�[�����,�G	���H�þ���G`V�TXv�\�kԒ��ȯ��'�-��e���w��.���+"Wh۸t��L�*f��OM*���췕��Vwwt��\'��F�w$Y����$��-��n���6~��@:B���9_�z4��1~�`q�s19Ǟ7Ս�tJ8T|��	|A�Y��"(�v�O�)���7���=��A���@��qn_0�%p�Wڧ�����4J�S���y@�qP���f�+d+���^#��٧��(i>|;�qNͿ{gt�ž�E�'�{�g����G\3�3$3](��C��P1_���W��=�&v8�1O����d��+�f���o룗�x��	ah�+f��C���7��Ff��]5@FБ���S.�&��?b�wcnZk�6�A �	�4>��L%Å���)�����_l#��]	�Y][�ӬLT��� �a�������)�����+�YI����i1��hM�䲯����b����̃B�¤�e�����6��<s�z�^'ب/$xW��e�5YYٛ^v*��sh��#�b'�Q��ti���t��U��1k �	f]5��=�wa�Sǲ&�hs�O��o����� u��e��L� ���%{ �t�b?��T��}ʖ���q��׏7���cy_#h��O��}��8VMfԇI��rM��=@��Q'"�{�~/w��þ!��u��N�\��0���昪߬?GxA������!�#��W?By�H�J���C���b=Uֲ�>ʲ��Ɲ~��3t;q�9��H[(�]䌝g|+7^�z����gI�a&����\�re�,f��X�w���/XL�5y�)9�e�~�	Y�} Z�Xb�چ�@3�f!8�湒�g������H��u0ѕ���2�.gӸ��7s=��D7�M���ֲ�WF����j�HJ i��)� C�䒋!*��f�Z.µ��!�Ӥݾe�K|�Ȳ5U���/���x��r�n͋|�*���忡YyGX�'�\����غ����xsK�x�[��,\�с�c$r��%U]> Vr>>�Ul�H����Ƅ-r8^;x�4��m�q�.��B�(ٲm�gJx���u��d�}�"4���銝��$�rk�+��E�EM�5�@X����+�M�;X������j K�zws�;��'-33Lf8i-=���p\�tne��6b���(�� �t�5�IA���68�r�8�;	�І@�D,�0�C�`��nk�xD�߲h8>�u��yͪ`y~F�2��2t��D�8�����\�"K&�7]r^��x�u��=��Ȫ���$����v��: ���-k}�t}n�f�'������x�b��~;�NJ7�?\�jF�ٸ�Ѩ��p�ͼ�WN�-Ԉ�ah����ꤸ��a��:�5G�[�*�A:&��q��80�ɞ�$�è����)G�ʹg�0�rg&���9�,̔Oj�_�t��E`�/S���bIZ TӬ�c�y����H�<O�s����@�CT@F�Y�	�OO��y���Ҋ���g�켽�#S����,Wm���"����Zl�@�k�i+�(�G��|,�/E͹e�y����Nv��"�8�����;hq���{_\�����f⢽�B�����6r��Dȭx �H�����	|��}ٔm��Zc�'&q�~�b��Oq��[]��Qx��s�`&�o��ݺ(nM�x���o�-+t`���-ҁ��«[�%:΁���wT�ըͫJ�v�v�C���\�l��S��m�*U4i8��X>�VzҪO���Me��^���w	���g���$���6��P�j��<�7������605��ŮuҎ�FMp��?9�P?��A�~�`uMg�n5�U<Z�ܫ\�Т`ʹ�4����O*�"W�i=U����Rw2�/~��R�.g.�䆡P�u'r��D��7Q���ҬSܙ��R޼�LvBJ��3�=Ѳ�<�p�B(�=�"�AW�SG��I�c��&�����
Ȋ\�S�r��Hy����Y��(��#$I�����w��`������Z�a���|���4�H����� HP�w���w��K_����C��j��O�DT�&��Ħ��Х�����+Ϩ���[NT�3��1}�s)��q���8�mP��\ޱ ��r��"C�u�<�9�ڤj�3!@a��.(�[t���|��i�F��>P�3�r!ly�P�9��Q�N0݊�J���&��#�۷�U W)��M��f�V%P��$� �'S��LvG��h1;5�)%����/Z�n�[b�]�0�f���#��Մ� 5Fp�e�ى�*�����ZP���^7�_�)H�J]��譵ujd���m̬�wp��#��O�Z.�S�΍�Q.1K���&GOJ��p�m��L�)����x�Ě���qI�H�$��s��"�y�1�K�<��("Ƌ��aG�sGg"�>
���h�d!Ěn@���)>�,����^��2+�r�I��K���"P���i�gS54��>�f* ۫Ưb��q�N�k�����K�I$���ݰ�g�.H����&�'���V(�z!��?���e8(@
J� ;�e���UN�h���im�S��F�6�1Rc �^�6K�;9�H��8re��@�nB��.4��Ρ��JeT}�����)`�-KE��+e%dL��.(ӳ��UUF�v�1w�/�T��4T�Sz�
L�n�m��̣��\��=��H��]Vr�aZ�ԓ�ٔ"�;��*�T�MuzN�$��Z��T�?�!<�I,�:Vս��:��X��F����BÕ63�!����i���gx!^d0�,�-�vѴt���v���N�Y��������bX�	}��q��Ü�.�|ǈ;t0c*!�G|&�O�6e����v����e�`����6���U
���0-1)Ζ�\�jݪ>�OpW� �UЃ�8�ho�����-�y/uB�-�7G��K�q�X ������)�;T��שpw]�^xǤ ��qE4��k�M�$�8i�d�zI|?f�pwv�����9��k�L7�p�c�Jo� 
����E�gg��� ڽ�ŋ�șƲ���5IN|CTU{k1��W,���s�,&(�j�:��N���n�̘��ޒK�����_�>��)�m:��_���k����_Ϥʆ$��F���	W������p_g9��'dS!�"kC�F�B2�C$^?����"�g�1��x�}XR�t��\�<"�6���$Υr�3��A��=dNC�,>� ���J��I���o�u�X�J�Y�Td{Ĝ�*7��ǆͯ*�g�=}��"��)�e?�*3g�����ҀJ:��t���H������dfY!V�G�gc����ڧ7�]g�H{����M�*�� �t-̈Q����L���.�:w~�Y���+$��v��Ύ���q��֩|j�^��Hs��=2+�����h�5����]@��'�a���2C���ڣv�	��˧b��R�>�wD���^���Y�Y#-����$�'/33K���W����"YÃR!����sh\J� p���o-�k��X}y��d&hQP�����n�ߔ}N1����X��h��2ϔ�hOBG",���P��]�9Bx\�l��+�n2G]XoF8�,��ʷ��x �XɄ�$������h;��5	�����A���%�|�9S|�"Vte�)1vh(U��9\�x��W6v]�[^,e�I�3�J��-��b��ؓȽ��)�M\Rp�5q`�g�؎�R�Ԓ���&~�OG���s���H��`�C&}j,]���8%+�����(k���W�Ȋ!�dG�3�dm��X��e�X9Pc��4��Ύ�zS$7�V2�aq3X�.q�F�6ė������2;�֜�\�����((�׍�"��:��x����ixՄ2��&?ҬDۮ�=G���2υi��TټMz
*=�u���	8 �G�p�r�l
�	`�)��K�ۃ���6VL5O;�BE���j�ۅ�8q�I�|������n��-���ĝ���@ymJ9�:�q�A���MX���O�Vg��{CCe[�ԣ�i�W?���u}cڎ�dim=FY�U���hY_������$��|�i��6�kZ�I�R�u�{�Y���x~N}��A��OlVh�< ���9J�T���ɳ�5��gj���b�o��.�����
	��]��T���P����}Zl�7N������]����[o�^ ��N*�;��
�%B��y%��#��S����8�_m\��� ���CD�� L�A�H9�F�I�L	�w���y[�Z~�6�X�U\]�}7������P�ܺ���7B��.\p�C!L�"�鵹����5i�M��a��_���_?-�٭۬��OF;|�]�rf�,���V��z�s\���{ao8�� �&�R��;�7,C3�@K|������7��b�!L�%��u���@H���(N0��w�&5���z�Fe�9tN��:�ɛs��"�'����l���n؀�\nZ;d�R���ev0"c8w1�,��;���-����ho	M.io,�7\f�8�̶�^����Æ��^3��K��r�P�+���Zw�Ǎ�=a�*O����O�J�U�rq����c
KW�<�M���z��&�B��QS��Ot��9Y=$*�����bNV��X�|�o�gnY��{��I�D�&p�}Fէ�d�{އ��C%����sP��@ڀ�+4�d7j�g�-�bd��w��F:.��"+�B$	|���Nb%��&����w5!�O����o=��^~�b2����c��4��^C����<�`+辺�B^����F���sF�4��B�^J�rX#�ъ��������2[�.����{�] �ـ�ζ�������lw�S��dC
:h*�09A�p�e�ߧ���p.5�?�s$Һ�p��}��DW{1�j%:�􃫴�k��
P��:C�e_�oP�Ӟ{�ut�A �2;�4]L)v��p�: 0h��#���DU�]��nш�u��|���x��L�E�r
t}>�[�u\��K�i�J���r�9.�� #'��T�q��T	|���Dњ6&���҇+�|���d�_b
��;��s�z=O�}�m��.�s�ȴU����j=i�JhW������,���`s@�3#�k&^?�Kx_�45>@�$�\&��܋0�� ��Q�[�����?��@3�5�eKƠMA�L��EgɚO�Y�5a��F=���0��%..�K���<�'⁇,��|����� <%�����]���^�-B�0YQV~ݷ;cUyO&GO���k�R���E{�J�q�١3
��"+%�v�BuU�W*�/�T���J<O�5��ɱ����|۬���>-���N?��d$��:A�m�5%p0�
z�S��X�ţ����"���[m�d_�@�-=yYmn9��T�W_Yl��]�p�&��{ɐ��I��B.K�*ɗ��/��7넹ma�V��\�J*F9�#E{Ӏ��r�|���1`'`X�_LCz�67�%��(�q�B�0�W�wX��l�F+����#-7e �Ty�Ve�p����rK��� ʄ�p��`�;����P�}\^�ִ�)��s������w�e=N�W��TQ��*)��aX@�?rz��}�6q�E)��d-����]��2�8�0��g�Ap��Ԯ`vAe"�q� �0L8N[	nϩ1��$Ɂ@�]���sZ/��.4>��c���mvZ(<�T8��sn� Oy��h��(��&�j���_��#a4�M�G?C�t>|��;�s(��w=�FX�l�oi�A�z^�y�@:�v\S�P��5�ϳ'rD���j����e�n����:��x��#g3�R�.j�64�}�h�����j~��>yP�2.��(����R����Um�A��S�Z����R�0�\o[�������Q���X���,�D�`���� �ڿ=dIM?5%�zG� ����όDas��T�Ǘ�ǁή��MD�J���̈́�8]^��l[=Y
�%5�d�-��^�r#5w�5z���� �60\�������̫���gH����2Xc��+�_���aH�%uv�IBGfD�>J?����x}���C/@���9�S�'�[�Ҋ��" �}r���L��D_�Jm��F.��9��EP�d=����Z~7
�������)穏�~*�*}j�nV3N Fc���W(�Vv��T��UXְDB��v~�����g����b�S�+��C|<�N�r������Ɩ4���4���覴c:;?/��\���ee�M�ME1MM�4�`a���u��y�V�NJ��F��,텆�ي=�J^(,� c�nu�Kv��{
��3No���<��e_I�I�$�?�b���	T��30����[�i�=�	��\�L�r��+��x'����V�/���]��L�z�P3a���D�����6�5��BC$% pO(�gn�_o��8�\��HR���>N�zt�)�%F��Cj��>���v��yڝu����D���� kK�I����A���CE��
��]���4Da�^ x%�A(n?J3��vi�XO���ȅ�%VzK�� �����A9(�U��a��1��x��HR�d��Om�/����U0�``�t%��n��eд%EҽqO��Tg|�u�:s��a@>3��lg16��c� �f"Y�b:��o���"�r�e���LviQ.bu��6�[)و-w�u
_�����&�Ԣ�:v'��6R�.9�#TE��ހ�']�$u��e
��}%)������\��3����M�d&�3W�ȊD��N���ی�,]/�t.������6�撝u^7�f␄b��^��-�6���;��4��~V�Ebз�1]�xHE�sa��>�U\P�-��F��HNM���w�S��M�\�ʱ��I���[I�b��H��<0�I�+��C?#�-�+zGAG�*�͋�{Nh��_(},:50�v�@�[�@��+X�y5�ܻ���?�3޶�Qt�R�=����aBQP.���֮y��=�C.L!�9aټ�yX9�1�k;�y?�&h
�������Ћ7��K�3�b���,8V�]:�O�9Y1�q��6�e1J�:��Y��a�SB:��M��X	�	=�_�0~Rh���Β�	���~��Gз\��Թ�	zu�����~��T�*���B�k�Ȑa4N�/S��Vq�+�$	ÍF<��zyK7����aL�$0P��8K�R��pϻD(嘋���(�oٵ�vj� 	R�(��D�T����\>=YDY�e�]�a����א��W��Ǵ������k�-���2�/kLsYWK� ���ۉ�?�h�5�B�A�$�����!�Ҹ��q��a��^M�\'�FQ�Zn0\�	�H_(��M)�k�Xj�X����pJ3���W�C�&�?ES�� ��#-�]da�F����Ȟ����Ec+vQO2�!N�A�~����VX��� d�i��;���˾���b�s9�p3㹠�9�-v(
����f;��Y�����<|����̪S�}o�~��<a��pc� �N�Iدs��MB?^�7�������x����Mk��L��of�!���Ɔ�$�_/f8a�I�
vOP	��ˠx�޸��BÀ��hȟ{�VD���SC�����Q@�s��G�c�d,��[K�*Gp[� zF�� ����B�]S�dK�̦HK�M.��H�;#�����f�L���Fq.������}n�T�I���"U�:�C��2t�Z���7d�T���(�
$�����#�"5��bX��?C4�{C�U�G���7Z%-�w���G-0�g�Ӡ� ��s������[']:&22�Q�'�ac�wf�\v>���\�׆l�}�%�3�ȰoS����w�)�-���eŖxx��P�{���^�e��X����p|5�{)�IF�Ie�����ak\<��"�@�>�d��wh~d�y���[ �X-q�2�C�^ \���E�J ��Z���+�V�������x'Zpv�o_ib��#�猁�?�cA��3���	�Ȝ�ǜ�-��JM��j��v1��L̍qe:��E{ߋ--xZ"��֏�?��⻶�j-m^�I��-zzu�ex)x�Q�A0��8����@�A��k��q��H�|��I��Q�V�vvc5�x�����ݤ6�]�nC0c7�Zi���c��O25������H��>Yf���'/9�n�ZcI��		�a�wՇ�Ѭ�C]U�J�zA}�Y����_��Tj)�qM����w��V�<�Q܍x�*�KB��T��MT�3�p{3���т��
��`J�g
|GG.��H�>P/<�������;N/�KD
Ҝ�"�C1��S��a���dH���qN�wl�0�P�`|�>p�ȭ�	/�K7����z���"Diۥ�/�Mݑ--�8~��o�bKj���Rh
�m5�r�'O*}�v{l�����k´=�!ʫˌ��İ��4�Āq|�=�lC���yO�����Ǥ�$�^Yz�y=�}@TRv�.E�0�}�gk|������ck|2#���E�b{�<"��/�v~�0Z��Aͦ��yy���E�2\,�NM�b����v/�д�6��9ǒ�&��P6��Y.r��$��i�;����g�W�ut����*c�?MV ��<�	�`�a����P�V����4��F3)BLIu���$�y��!�����~��b`��s�H���₏�S��Y�GWG6"��#�����E'��#=�8f-�	p�@>�#	�d��}1J�[g�[E��iV�oi����8�6�i��]?N�n 1�P	��ɦ߲���,f̻]d]���'H����!�My1�I�,��k��OL��x˯����J��4ɭ