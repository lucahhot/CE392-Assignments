// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
7hqk+5fhpfi2VYdzvSwgwZmSVgU2YB9TnsuQYpXzzeOd1m3//Q8X/gLuCqAqNNy+
iCumvN1rCx4Bq/huLPEL2dBSRhhiTQsNIx9nFzOZLnQncW5rQNe6HMUFRPV4JxmF
iP5cAxOKrarMsd1UEZYAhZz7N2ky2TZwd8f4BolZ25jkCBRrHw1FSQ==
//pragma protect end_key_block
//pragma protect digest_block
9F/++SBhh4G4OQGRWLkk14ubz1M=
//pragma protect end_digest_block
//pragma protect data_block
ymSo2WrccL7fPgFSs0dZKEvFLuiUCIaWt34InfH5U0Oikzv5u8A6wi7nkvzRLy59
ocJAMwP/nX1sol4KafBMtuCYh1UFJA3h19cyt+U2Q/2xpOlgk3yhI1ZdEQBDDCuY
LEbDQ2VChR4P0WLr1tPE9OmUisfcAojc6vEM/aWQZuHyjeq1Ap3rRc7W/JubmNbZ
sGLsPCDQxk/tnm43UAn62E3dJCdqxdflYfURfwbUsKernoqFLnfxhHjmG2VxoL/2
4YQ2NbHImQe3bsDaFQk/LHC58lQA2+6024PmcDkHVDj9iEBHjESGZ+ScCkdkiovi
uKXogFHqSc9v5hcFRv2mErqyJ7YZoVW9PFuaQv671D2GViX4lHrCqoUPE0+f2fBV
0s0FU7XWRQowXP0JCjABlusJcv5Mt93dRdaA+RHiPFx1Dve5kVFnYTG+Bb0d/tnX
DPJCUlOHuzh48T0MERzAcdGDh+K2nTHPZ6tpBhgsDBipxdnCAFHj8JdoJeYHeDJ4
bb5XS+OB7Nxk54rlmrr14G4AHxam/tgHT53j9rI8PddLQQN9Iq5s/uwspEeMSVLJ
3Z8iPkc+EylmXB3yw7IKu0wR7WF5+5vFROk7QaQKgfpRgkvbOIdx3opk6iPToKtn
V8Q3ChC5EjHCRuz2aSUWnnxT/sYjHZBUFCLueJKMopjljizBY6n3HThoWi2IXgq8
MVs220wvAQJWTgztIhniKsIpn9UVy111H9xRXloqcubKc13LbT9cb5OWEEKka/DT
/9oQlFwkamlvskqEpFSsNL1+f/EIUMiqgBuXEOXaNGiB/tupRXAa6LL5FJw8QST1
AiE+QPzUcv8yWZ7C8Qzl7oQDmEnHkkLyA9+7ZpbR0UybKydRBE95nyVK4kRle0E2
VxJTl3nYyQyLu/ltFKhwe1yFelFKSJvyfqcWvuerW8MMyWYGnncyODOzPYJgMFyo
/QjHLef7ZmfBgQAVidSPO3CEkSkChDVWb7hfRn+TmOl77CWOINjTb4pZDihj9W3c
qq3v+nrF0+9o0iiSjjMA9Z0Doj4w4d8Tw78KvbGSmPL7aoj437YO5KMZyauDC9ZH
PPIoFlcWrDUY0v64n39GV30CACaYyFID2hG0ShdpMJNiV8MqeUt5JIwOq7UdTW5b
a4IkowRzZKlf2dx2h+LtTmVnEdcr2p/rpvGFsE27zRhPi4Ph6YTU6HNkrcr8ApMa
nv+sAqRIrYxk7y/WbdOyau2MHcGv0f9Qf0G7aLBqceGrlNZ8rYet5FsIimjTc4kW
ib4/OpmEJdtkdukZlrKCdwgmAwyi+c54nJfFcIiXt3kZheyMJMcb0F5WZ+NF8V9b
t17HNPk+K2T9DBspmAJi+w2xqjQQXb0gPs3Asbm3rUeRZB2DemWJhnJSOgkJdg1a
91WFX6RKowngVB9Ra1nziqRtonw8M0SdBzL9CfScjubaxIvkg1gbG0+8wawFz1QG
adFQ2cbw7R8qb8c3w6LB7v9xWGzxprMEcPk/zF3dmF8VmN4kijKGieDwNOEnzVZq
4K+bwwqSshAzSjCx304wr79gQ+kAnmwq7CU3UosJU1lrglP+uD8z8Pz4DnGBLKKC
624f4eKZG4oVJYnA/QA5FEfu5sw1QBu9QrFpy/jYPkS7OSOCUV3/U1em9sNQpUTq
nXviv7mEN9ZuBehAIWbsJXbLlPVvKZvMY7asMZAF6IRD8S+F7IRJnQG7sLgTbmik
9VDhUuQK8MvK/lvqZF3/zl5jza5fU/XKyxnl4okV34tnoJ45aq3QAwM+KuKS7k/w
gxA378PLmCNnpRq3JYqFLOXeZ2HPPxTs5Jv1/OsgFqewrFqRgapYiTNDss3A9Uqu
rL8ge0Tu7TNMGkozTo47Q4PF/vl2mTVgobqs3QGiOE7DtVfK5aRHT4GqTrtj18uX
Q+0sNBNQb6+ppC8PqRfCTbImNoUUuyoqB2Lbe4DT6Gbfs/JJd1lqYWyReHlStSfp
FHq8zNnLStYtqP6z5ooP43LF4zNon7clqB+4qZkhgDbLlFiulb939PQypx+EYBY1
UpXTx3ZRYC/IfoFdJVtqU/tgWTFC4DDLZs5KVIH0zZER0bETrVuPNi1AueR1aMh4
+V1y1wLT2rcxbakp+0nkYDzb9DgvlreRxniSHw/P6foT7Bry3qHvV7zNe6SYiQ2E
hDvqF8U874rS1XzCBS/dhXB3RoSBYP250kW9heFFGqDG2ecK0uTdXQiXMO8bgR32
2lhPnLG7QZkPcJhirJw72yyDX3IQVWbCG4WVrvsYbn94wS2oUOxi1M6HuS3yih2Z
8MPL5ohtggLJH8mC171W8sXxA5Sx6NMTTt/tij9j9NlQNfJGFhI5C7Ton9VQNiWK
5zL3g29SMXJdVE/rgzVuDceB0c8DP/nXbXU0JdIX8nEXzlEG9Ps99+A958p6D+Fe
A0FVaryY/c2+irJuBV7qBZ5SL+qllObTqHInR2ZOExAjCHZq0dVKQy9mMyIGVG0O
L0U0fu2LouHShsNsVpBeUqSUq0LzHPMP6gVkL3ZSx0dLMua3BzM7w4umFmJ6FVgC
nTqr8OjH8Z6uG2K3XRLlM71pn/d1cBKnSx2ewMUgxR0dwZ4wvoUmE42Q7c/2L0Dd
+31cWPINTFvrMdpJhDlr3FFDaht41Hs7yrMy/HnJ38XwrkB5wb5dI0nMEZuQ2i3+
qGS8b0US+XXFZkDemRYvz1oVmkhninVIyfBSLkXzZJFJtSdvlbJ2t55hEqdAL7uT
SZAdgvAr2UbTfd3IHk4lfXofFltradpVunjtYZU3z+VU4gMT2tnDmYBPK5H1KEx8
qASjDBTmQmRGMXdHol6XaKm3Wy4aLufP/qjp2aLru56TgVv8p7Q8sjHSH1VjoLay
o6QWkhuYnIQXXHZqrLGvpGyCq6lFRXkFHpV/1iD+2XOQdC3rJYMwm5hcoxtzFON+
l2bSCu5j1yfm2Hop+knSrBO7+NBLOsXq59cn0EkpWKImwLvzMJ8Et2hnXO30KZEC
onWenIhJ0Xs4ydhRvjRuLWiQQv+ma9qhoJqng9WoVuwWrHoRXAM190LkGtRQ9uX7
UGXNNOhjwZWXW3DxnDSMcaMkOcEvkTAEVvslDRArm4azqr6pse42LcAdCuu3pC52
lDv2732hN1xSVQPs4nhJpG342NHdBosqEbrgnf7S5oKz8MxdpL5C3MKWXZGzmo5l
H1Mxi6IvmzGYAS48SpUIj80fHVAbYF4PIe0EyzIf3zE/tJ2qRsZ6nLIUYiNMcQ7b
Ifew1gM9TpQLJJAnsdAzBeIFs9HMShrjkx2jC0usTozH663PdD+ohuk1vIZ8dfR/
jLRaTzlLv1Obs96hgu0O2tg+r6n+lmYN5gtRJe9bnQzTqs8d1a1RPY7SCr/7zeVM
eKgJdzM4jjdsVCMEPBR+Ud57yq4HnZqDce3pOIn1eGocojAUTJwuytcaFBJOWvuX
+QlbSXliAajn++5am/dtf3iPSmuZGJGIxd1Ay8VX6at2eBD428fTD0UVoRWvYnHH
IY8q4kAAtixJ6ckwdhqQpCzP55RDQlsOgQ0yXzH2fRZw7rJVAZaPAH8ptg7TGyNA
1xslA9ycd1mhLC2sC6u/Ll1d8C43svkI4noZqLGlcFnxtmt9Tr/BwIW+uNxriq9M
05GnLBoos7T3UUSMVva7UGcQ/1QIIzyyXuDZVsas2x3TPP70+PYvviepVR08gjnB
DJtDUyhM2EewkhGTcndsPrE0ITRLBQhdQOnWng4uQf8TEzTWeC2iQsodgEFRoBeu
b1Sauhz18BsloOBz0QviOwGwvd/MPt7Xgah2qrO4z3dctrAaTOFfP4EbW9ndVsVF
kqvK6smDVfiUH1qPEYeU48vwJYn91q8nCO+/q8ag38ZmMrlm+fPZ2BDcbWBLvm32
ZPQd6sXPnGjPXXHSPnlgn4CnVkzMELEPIYvtFSLICtZircNMkxbWMZ0IuDTJthT2
gsa3+hRpBBBzOesM2LYu7+s5hR8MLzCSxvf/WxmiZ4843QnPrjSFMcrJxRmE2zOx
Cxn5Qa3jVS01PPu5dguOkE7vDwUIWh3BeXmSbj3nPi/v+xWXsqvh9bc/JQVK1kTg
+3OvVTj7bYWUiyUmlmxjC/js+sFCa+Xz25KQDcubWY61fqiXIziM3tv947x74kca
xSqqa5+uf4LbPyzy+a91nSzu1pM0p04yPTxllSZwQkBk7UHmbX4MckeZqpoZ1RxF
DQdImDBP4pvEvV+fbHvyVvnrSQOn4stP3k+FkeOkOCpG0XeqYjxkubCJ87dFQvHi
sGHEzcgLcrV6RiX31PAAG6bUbQdHbynjnffNLjtNpCRKZohNktlXsNPj5OzQam83
YfkYr38egiJQ+ZuIS1jH3OsEXkRKUApcGkQ6jUTPFjTVzN59B/0xMTt6J5Ww1A7D
0dAsraekf1brf4Yyymfpklw/8dG/PB7ogZXKd0DbaSzc8CEPVEonJtRl0zDl2TIM
AvTxspF9qZIeg3swK0DJOSEzIkJ9ccZ+aHUUb3SbW8r5fByy7sr5R++mOgC1oLGR
YcsUov89bd0vbraVhqOzEqIo2jt0/ri3K1MQkBQNuxZG4Ocb9tsw4c5oIGQzse/9
LoeW3zH/Qpt/sM2yEza4dU0TIOSpAwRkk2UrQGoIdzfaMxb5qhnxXRoAkx7ltUKC
S5gYYtfdhD1GOv/E/dlpho6wyVtCrwr+TnLF6BtccJIdiUn73s40Q2pyO3i3djP5
/2C2NIrDnqGCiBpiTOzTJ6CEdV0zjFneFfBH4ByTnhwIlNvh7uVIu7Uu0jEadOqQ
dH8EXZgVqBJsCKfwrDL6bVkBrhvqVZem96HYvKGbt7hYJPk+u0Ly6F2cY0H/seGH
2O3pykMKIZO907maVt6krFDp9RZcjkJFa5Upln7YcCKKmXOeft2eBeDWK6qpwky7
I71Law4L6RnlWVhE7YuS5ZmhrJ4wVJIKVwjY6K2zeTaPpOlobmR7yOWUG2SEQvwM
7sDIF+H6AfiUHLZe8+nuTrOC+vvkPJdvzb1nBzIasUYGfd7jK0CdnotKFH+LzMb6
fGGtCflXA/Wy47Zt9SrIIaXgYM7idcOug6tV9R2ZaYixtkE4lUFAs646oG4faeS6
Evr4wEMdlamTKfHd6SzfQncwuyeUF20R+JED00mQdotxIgXvWZfUz5ezDwP7BQ1D
VSqWtSMzZBi7AJ0BubKv6Y5q2PZ0RP1ftFCasW/vAeETlK9qLvVcUWGgwJ0U8yG6
eS64syOFT3nT0+aiYXtv7SKuR4Vxg9kvlwAA6RvLFmc6NVHVq93SfhRvY0cYquHb
ZVt4TfeLV3ZUmr1fqWTUkcDkLGRFcSOqw9Q6SXDj1Xsj6nXUbkWFqPJe/qRAsEBC
yNwNdWPHxOurTDUAwb58Ijf878FbwYWiD956fzmOH9U1MLRjBPGsaJzMqhiH7Ewa
i1GjpmXk7q0hd954BOnb2U20iejNo0+Y0dC4y2YnpYuz8d90Tkjc3zokPSD5uLgn
jufY3cFpcca4ZS0KQ4hlpFARCa0TvGNWim5z63L7yg9zE7sdqZAtHKlXhLwzK3VJ
hwBolS1JRV7J9GxhZEuC1PgId/7RwULsyM19pMnXA4m+8MB4bcLrxu2J/OWgOqHh
uem1q56AtkSc8QhEJxc3uIMMl0p70gOcUYFiF49WTNObHTlcpwsd3l0uzoWU0xyi
lcqour+QEe6cti3KqTDmaZdYv0fuHdeERNOsy6ZY5qlXRSMf3itUP2XBmO9+r5Wu
bWw30jpTq0wLitQ0Hvb4GgSCJaWQRNbPiNc7/xVFrDaBCzhsJkp8+8/suq2/Ak6M
q9YO+XFe6HWVt7qnM58pQ0nybP9st23i9PCwzLoc8RXxJsf2qvj7Lew0L1eKGvUi
LEOdIHSOnCdQF+inzJo0lvf9+ES8afkmpKaqaunuSs3F/uXJhy0HzXnabDxrd/xb
V0J54I1xpASwIHxQr//wAiv+c4QK1yZcCNq0orgqC0XmE9F1ogrLMcegBmN9mYWx
Y6K6cR8DwOcxGy4EdPXSlZ1Che2FMEPmgosA4xDAcYLjetNeDngVKK/YAKsfJHUs
Y0Cig8tXo9wcYrevuyxfCVXT+M1iozIVTmBRwytWAZfGZuQRMwYwIG7hKbCaxPqF
+QpSgLu15PHSpFiaJTkBQps9httDXOIH2x8gCU8ZnlI4f4MY2nXSFqIhzyY4j2rc
s9MVc3rytaPjhwPk50sS1sWuQ98zdqkfC5NDUUgXLwwo7wJcYAfuYb0YsJIk80MX
DhUjI3EpXu6PiifSOwBON91nbtIi1T8zXLJpW3tqW+8bQAVsCUZBquHAavGguDmS
M/07xZ8k/8IiWQB9U7DD3K1glE5p6GoDfnoAPd4WSMevnZ1VxwanO12KZ8RudCJ/
pTObC8Q2CkeUS4k0LjQsbVTO8jgqwzgNvdA0GWgu/pCCjws+NSFkGnDuKjO1yLfW
wBAzAUJpsaFYCs/STG8ZvwOAoRI2Cpc9dr7tLS72yDwpxJKvdbbJEhX8gWupQzvp
lyCeaN+4KYGg3DWADaSyLCr8issSXkn9Wfb1Sfsl+r1ik8wL5zNoJUtCZfS6ivXp
B9F2TnpOHeaoDoLLyHp49VKufxRxViKQSeU1nBhVHuv27G+Pwz9D1RuvI2zlT+xN
eRCvUrwKEZrMQE6xBZk9l7dvQpG6bYnp5Db03Z8XN5HPtP4qwYv1Ji2Wansbx76S
c/U91HgIqe5kNBjxHMeRBsNGZ0x4X/hw54SBQpqH3cLGwDjpkhUxOYfmQLSPfjgW
iKjd8TSvaZ0ll7140HOEF5Dd4gqWnvPczWZHnnGP2bs54Po/mE10rMqDdWISbS66
3PRt3tB0vJb4i2hOJacGnwtbxpb0aI31lxbzAGnBE57unC3TcH+NkbpxmfFxh2xA
Ng3rp/S186LlgQkhR8kjGGqeaLPV9yRwUmhDODX6p3scCOc3/gX1FoceDdwSH8b6
bu5A+zX6TiCHpkbsgx3UOjOQ/p+C0uK8v9Lij9IlQo8WSjCU6RKF8RxJDAZxQ2Ss
c67HA1JNhV8yN2KYt1mjhjcjLYfS/Cg5x8b/kNbdCLzB2MJ4B+L/ug9Ni7tQhMU4
zhD0yZzi1dXZyFbTX8uGKKzms1OBFCtHlHqGANicGJaCueSXGjoVAGCqHRX4QBL6
GvSUkoBXzFx6DwtzbiwMIfyTR6XZV1lwshuOvov6LvecavpmjjIUABtGDic33lj4
7il0OklUc0mhzN/2JQ1QxFMHw0s6cc1Ny1E+FIQ7+x5wj3XD0o656/vHto4vx8RK
L0RYytoqgE9afPtKNDFuNlroWEUMs/NPibkecYk/diZQO2HytA04gGFf4GZ9iEbf
/d58PYPWm6wS7qWNMZl6eV+kV+EDMOBx92+O3Py+fxaKIJiUahHKZ/SGBSA5kZYx
jReMe5R/CWYSaxPYqmYwQa7tz+taG/HQzUGmMtHSvmU2PXWeZPuiNFNAy3fU0nur
7OVK5cy+9Rmqn+H2cVcswevTbphUGqH5utgzCUs+BuU9ECCMm8oLmhE6sz2vQxJC
GMxEQf+yxKam6VVdW910d1CWef4IY56TlSbj/5EaDwZ3LJdJorf8IBK+XiUzGxW0
PlPXohr+hlgRqyArhfUMQVhw2ltX4PYY9IFsZFKucdqCbjQlwvdr8Y2Z67EmFySv
TGQ5PVjU9m9/iMkFJmPk6dDvC/15rOZ9mmuRNjW4twEqk46yrSuZ0wEM+3NsSUbS
8/zfDchp+OfqFRKsjgWhFAmwp6sFWpUXhWrxCx8kZyo4vE7ytCUTi9xnSWpErj06
Mjtv6SR1Rs1mIY4FfY1l3URCmtLut2H2u9E/ap15HbJF9iB3BEQm2glw1yKZ9JZc
7OgcJTgGswbg3f3JZgqJHOX2TLtbszOyHB7aEFDqli0SFE0e06dhVd6WwCCzWnMk
qnWTJjrX3/eLW84CV5eTY4uBiuNyPWtcGc+QrNkGa7qcsvnH2oYLwNZ4gbE0Toe8
wYQAAA/NJedncgmtOhO1WTLiG5i3WQGUJWWc8NNKDkStUDDwjAu1XEbHxXcD57qA
xF3dR+ohg/uyedo/K2zYs4ITtPGmxFUo116LNWb5gzlwpqSmA7bkJI7oh+195bKt
GhNtBnPqeuPemmWrFP13L+5Egswg7hTNkmH/fw7NK1aGcJP/uvftQEhN1Lj3guBX
gwdR6CNMx57t87zANYshGvdvA/II/2SjKHwYwLCGahLBKtKRocDMSG6eh0qFkN5h
lm27vAFSzy5WzA4ERv4jH3zY7jKbveM847vKKWy4hxLdB6/Qdnvet++wZ8Tl2FrW
gQPBNcrvTWvNwKF0uRejyQPvSyF4Y4UZoUxZh/S2UmRBubP2HULLAEhU34if0vBf
BwvBkHzE4JXRfMirTOS0GMKKOb14di9HHHcAlkf3i+RIMGDMdGhvnUUaNkVoFPaH
pGiHQ0M6iuE8QWjbfVHYsW534W13CzT6I4gNTS6kWW+roPdn4BcI46lBMBWb7Aho
ZRHQmZNzFvAQ0+K++WQpHlRNeJjimP5fcsW1SsZPAMPPKcsAawYxrA2Iim71HV1w
2FhcgGaPPIeuI6M3XWgU53NjR8h1wBFdCwm0/n0MT18XsPvlTK79KQqB8reVbRnX
HVTDZjvZ2S9URIQ6COPr2UoRla3YrYWefy1sVaVShKF7IKvmf0iXAmL2xPDwDdhx
wvoriLn2oPEWIUsNLPiKd581DonkfojCLPEx0fLFFSCdpImKGFcEmk2MdiWrmMQR
DG+6MtmVREQkY3uE49jYN05qPwwil14ec8GMffsRO16n+JFIDrdN5ZPWmQOod+ff
k7Ji4Jb26ZdZYqZJy2Go8jh/LCp/DVzD56qxABsklY5iJ1rZ03IAdPG8Kx4Z39Fp
OmQEWccqQSqYwPhQh1UCMScIIuHZb0W6caAs7r6otlY/OJ2iXi8/ligJeSgwspD3
LktFgeemdZULZwFbCLX65cZao/ar5S0R4fI2n3X2f07MM45uV712GMVKl/NgixOj
H92sMb8hQKm3PEdd9xVpWFaHFYkhqJ1arr5yREJga5egNUSSt0/xe5w2kX8sVGnk
14vWoE6O/e0l4APRZw84GFMgbwUmOcQeyfnAQ9YniEJPCqAYdLgSapsRJmFAayBh
aBB7t+2FerKcOu8+J0K3i4fvxtPU/yFa4m/us4ujUYNQdRCaVvTt9fd6+nfot5HL
LmKWC3oe07xnx0LwO60SaGy9rYZPo9awk9m2y2alrIGOYNVqXbECnYWnn2cTuXOE
BAH/MyZkd9EpeD2wdg690+jrFPR3h0caPNLBmTzjXTOHLvNvrkNNSucfTsEkee2S
oEOdHd7VOaqKDrUWt1/Sq7MNqTt+qZv1qaGpzMxcnlqW8DtFt2wkGqohT7h6SWA/
0bhoxajTee1HN8gkjkOV4Tz2TKnMRHh7RItA2AuHwTjn/cKaDreyaCKh0CnGkag9
3DwKWoLla6aPWU+aDS6rK1Bb/J/+USlAqXv846hz0WO9nCVx7QYvWN7V1pO5GzTC
cPOVRfs6snHfkOPeXLZ4VCtSrJ8BE56ADYBNt9115x7G+bc+GbsTg5XberhNaadn
xNEnd4E1KT+kx7E7VM7oSKOQIGA1q8Vq/9gE42Hi1pwe6D78gvn/iO+biPdnxNDq
Ukw+X1tCHk9bTwW/nHj3voYXo3WLMOFvV2ANxUyPHKj4Yjj89qNIrEkmHZ6vHbx7
g26zwYapwngpAzvela5Nzpk8dc84ST51H4tWFD1TiLtzZlSsRpmku02puDXUmwNV
8dV+ExzG77yY2kdzmAcD6sTy1kDMw6gPjZC9Kwt7HRGsZUr/OXdRreEX/ubZOlIg
hKHLN0eA5/zfNuDFPQ/KiAcP1TxFb7xFNsi/QGu6Ym02WxCQIoJ2PNbOYt4QyyrA
rjSaITy1VW4H1+yO+L9nigcyz9pP6gB/pn/WIWkFp5R4+pcqZlMFqTEvqHDzI/DV
EWGTVCTsGCyKKdiJPSa7COzYOIC5QQmy5FA5jtABNFRRGLd2KupVymC6z91DTBfZ
hOyLlnevTmxMS4YiNBlaENqJ8VLII3DR50DImtEoy65kjbV3y9tsLYCnOE6wc8UD
fMc7lvXifyO3wiW0AUCI9BcsTfnrqtTwkqnOhjA19M9ziLFKhteFmuiCUSw3JiL2
qMx+fZfhMcZ8QtHHxqkvqlcaAdTnC9QFmXiIFQJJWbhqGLnGKg0k2pKEBi3g0STs
+KzHglWJDNMGrgFwc8k6RqdOIG/2Hx7vcLlQe6UfGqH3bGtWUTeCDGEYQ+DwW/It
G2x2CLyXdXtlRiGqiFgrWSrZEQRwIMcV/U8VRv6GjAAqInjEQxezBJpvOBU2R7rM
FsEVsMYyA0c0bhEAZ/2qrpl/KUY09CKc2ABb8JZ8LzIcrPTKQg0Wh14B6ZMuStGr
/cAs3aLfAo9pjjZg1KAmAQDSY3xpVNwS7awA+Ncm/QK1c3B1jU9og3YMtp8xIBKg
LbILwnstHMpuZgsbYH8j8lVJc0e4W40sVYijdZ4Q2rocR8ZM79SPRU6nZiO0g3Uo
wkvBAQRA3MW6KwcwDK37W1Gap1t/cdWAuuCPBCJPofR/dklUvPlHWjPj9D39sO1j
EPhDHC67i/LWlg3lGYBcBH6OZIZpTO8zStLbKYOoeW4QT1KoLdOr3I/qZBkbHq1F
xltTkORlilN0d60bMgmMYnPwWUDKiQi7Gv6CnwCXxDiOHvC/zh+2l38L4eZjbpGs
9J+HqahDdJqIu7LYoF1YsEaKXTL26J+XEvtjpgKSESEqiDnwP4unewOfG33otIlT
Rso185ttol37zkF6y/2V6wPyKOLLzHtha/tbyeHAC27H+jYkyDoimC1VXUNntvWy
2GZfJSTLjYwqb6O8C/iGua1xnr7eD/UOspbxQu0jlx4Rq4bFBbrRCKNWalu+/Fj/
U9WFoW+u4SQt6kWvmpS6IphQswi5fhl3Cr8G/KBnMwMhh2TLrgPx+dbICUGtCiRY
fH6YrYFFhyowdMOdV8iccu9EPqfoT2gaWVBqXepm3gMXHTkHDtIQWStvCxoahdkx
JNL28nxiPLNHtGKJ4R+XUuFC7mATAYdTB9WFW3hkAmOJMyEmeOamcn0tEicg8e4M
n59QKZEvKVy3nZs4RhXcXn/4LmUVpvBqeTYUwYd//zKQ8YnIcwPZjXJuzBTvMhWQ
zSjh2PV64vhTGrx7hP38LsfvxNK1YAIoCgX/zKAM5djAy9iaIdCEZE4gb/rTs4kH
xSGLdObtlsITQZE2LWB091Mhzl4xF0HiGeMUyvsBCjgupwFx9iP5n22F3pcyS3W+
BXKFXLvbQLMqVJ6L4FnZOSFxJjdLBtObzCWS/fVEPGxZhYjmgkQNGPj9p5WeZK5Y
S5HovAtGnSEaLwv7MRVpweHEp5FgZ1Fiw7+21ES0M9NXDw4c4EDHN7JMKOh/G7yj
38IBYM/akSOap56ekNW8uGwakOVHOYuFdQ4ZuXUNi+j3uSrojHAIDOyz4l53VpED
xDPxBjCOP66NcskAfvrBPFcPM2N39Q2AIua5KpToz4USzu1X1WkzXPYbnKA5Bd9o
x6VPJDKoSh0H9d65wp3Y6KZmkznOH9N3Elo/6D2pYpX12P7xGYsbsZtEv/tVuVHI
hj6hQKOgVEyY+vR04cmkK39GMsDLbp+d52fBvYxTmCNdzHVOzuS5J496H/fT+QIO
f0aRIHLD0YVEuIrykb1vOgvknsKQD3/nS/hozK1VkOqceKQq60Fsrj+G/3ygIJoy
lhouycdItaYrngSfHzOEKjNoxn7OfyKxvOMzNyk8fdG81xPMKKCpB0d9zYYsptXT
kFXyksEJfKtMJ6EUl9huGsZToaRUY95i19E9vlswaAdMHTvrPI9lyVgamjvl3e4o
OIyjoSgXIeZp6RH01fKxz6I9OCtmR9GMr5g2mqKgP+uEjnCEQ2DAulKZoQlxn3Vr
s6QHu6sOuDghcolacPhe8YUONehrAXBEGwFTaPLbTuwSYnHo2WRYEC1kAIrGMZQw
yfnnP/FMVyth81IfArg45gex/XMFu2yIsWW7DQbIFW7vCAJt1m4qE9LvqsDKvqmJ
vc/C4tIAQ1UKFAHLosN7vaorcI87cIMcrN5PZ3bbonduPFaru6ooGz3GMpqcP0wE
Myzyx1BAK1iBX2DHzsvON8iFO/hqnA+AqxC5kd1aZ7wJk/UI9xmB5VamGOv7Vh9+
aSZ2Lh3Y3t3LmpZTR6MwC4Qq9GAH1zByFP9UL6ppB9gCwHvnZVE/JhcWsukSB8Rd
5gEKLw8f5uprmIQjjitX1i3e8RW7erKjYLtaAcvwSXIf6BjM5tOHd9slEz+lLe2h
m2reG4IKvVHiR7Hcb3QeF6Kxk02BuiKIkvMa7wVnknZBafTKgaWs+slepYkb5Mpw
xu48xCx2D/z7GovtbwYLiTxkndD3CaJ1he1DvNQxijc6Xd6Y63qNJ/EqxKY6kba/
JkCwyMU+EcknZLsu0Ac/yxm7dss+qZU7cWQcBl/X9SWNNdbzR7PAivRIrHyCLQW1
l2TFgQbrt3v03Y7vSTjN7PmPrsa6nyYNSK6YsoYnhibE8RifsBJ3cclb6xEX2ow0
7RtntmvF99IUppIwfuDnFDRkxGOogMv4s2kL9hh8nnNSEFd2N9dnknk+3y2aNGhU
4JQKA8TW7AtFssnXWhus9dWa6DCYRkMF6eIKOT3JXGXvTx6VoC7mJStYDgzJyqbb
MIICcieHn+5J/E3OErmZlHYaCsqUn4lpKZLkNC8gviE/pMLshO4oCCOzGaWei6D0
wYyCE1iZYH5GoFuQGDSXcT+1tGixwiEgeaFRUeVjdiKPtNOsOdx/mK9tn5OAn2pS
kgjh22KJ2U4NabcfvB4STiGEw3EMWgrdWuaMpMudSgYVqCwCTIyguu6HgZuQlBBb
PJrzdtIEyCDEYMiTa2Ix3qAvtF/NPNfEvPSVIEEocfmIGgWSynsTfx5yWnyquBUo
7KG2u05DJ7oY+TJOW6oZXTBLlGo2nmjezxZ00WTj8QOIKL9gQZ8yaysrBck5G7jN
BAkAso3bgKHI56dPR3jT2woWyKgg4br+JbQZzvoGNeTvEqz41RE3EFUDSTH1dbcx
5/SafjTtaehjqFrms0QJ52GmVlxhHAphm1VOOLqkzGBlCaDkchAIJNR/imK0+0xt
l0bJn6vqF7pRZcXCtt8ye+MCrOXwZ6O6E8TA86Z2eE7Zn0fKVz0TwI5vuFlwbC2v
p3rubjnuNJme+RC7KXtoNqXXns49WT+C7+JjVHXUeURZdcfFsS7xAL7q+GsZENu2
vA9qLlLt0xXdgxyu9hcJpjEkFsP0SvN3wJYos9OIkj0zqKbtS9peRdM0kh4K4qnh
yfrOZgohoNQYY9GAG+f64qXg53kQ0y0Rqb/8OSQ5gw25JcYMvmaFqVK4SNFhtI6y
BMInYrQXTfl6SbjPPReFFjC+txnF1OpiSdMpwX1+bYRAuvkVutPqoeFUEnct5X4b
nQiTNysn/f/96J5XAZIvKczk6dHLkEK0dzvRxDTHTi6/k4cXWG5jeAKDYgUHTvUl
UHt4F65pXdfTIQMxACUeK+bPfygv+2dlxXw6ZlAFIsehP0de8dslrW3FsAeeNKYJ
LVRDxS3dsCmOMdK/QeSoMhOSfj9CuwYyuBNPhnFtJ3s4fhO+X5otbedg6oeL78Uj
EpjlcgbIVJsFwxIW+7gnQCiyy64UDI+dp49x9Zvjthe/LEzbFxfcRuLUuKS1zgrx
0DEIw43WOFUb502vQTjToJFhwjzu7nd1P1R1NaTW5WhhpKrgfzxWoh9PtRmr7zlL
6TL6Gad5H1XyASQ2xEW7M+0PcrN0cJ42PvAGZSlzu9zNk7ER0hB51sqF6dM/SWwi
XKPWmRuZRcs7KUc5YJO/Z2SheO2lghFu4qJkcQDpba1oIiukAsz6NBXbf8eu96Jd
mqWqvQpV5uzdPblRvVLNGyEOJZd1pohvAsH4hxKJZeB5qmXKXsfuU1f0USLdHEhB
Ik/Zgp6ibJyYkpdm3FA8++5HU0xkrWcOvch4aMUlt28B1jkDAWRoFj6rtQu1ecyr
g3M9OrttZ7ufXrJxa16dSdFB3Co8FBX/8jUrV66qDk1LcJ0YL2yA8xAijFzop0yV
lFR42BYfPxrUa5/ZAxiu2ubJqIyk5QGvAA6X9CAIgS/Mw2Q3FUJsu2P58T9wFbsB
9kE61FtwKznO7nc7InRXg37UUdyKULFOT/oYWUeYfI/5AbNOPl6tqDpYmVldNEYU
s4R0a+9ix0PvAVPuGIyR7ORHo1xqEFP+zYW+aHFdbYBhyEP60wLgdpOhn+JVczsG
zcT2ImPJ3TKB1ZlM3hSn9/zSaLhYCaQbCNjtNMQ9DH7nNvbIBLU4qPW+0s0up1FH
OY8dtoT6F9UGa8H81jkJg6MqsPb9Y/ReCmtgC5NERsSGtlR8GrAiAsH4jxw/0RgJ
PFH+AWwiOiw1xV/cu7p2mTtgJp/MGxU6TUkDtr9JpoTF7l9+bhrDYJKAgPD1Oqen
bIgPaoXwMZMXBqVgsy1kVLBiRUeVjSX0WBRB98Ub210a3IZCuWKUoi2cdmNgm9kW
bTXNxkFxg2WRNmOEztqXWLRNhu2VCcUf1tE8YltkDds4/mYPhHuaciqBru8//8KD
W2K+nwFdIoDkCRE99pXWgBcYtp/7UKyEK0nqWB/lARthkabd5UC+gZ+8EshTHXHM
Eog+imqOqSeCy8LwZgrPIdLpl61igrldlRYffgufMpRQ0jMe4QP/dPU4XxqpmDPa
91ksr5RQEu0eF37nY5jYUnW/l30xQ6yAPhk/ZVsTlgpVPK3rmYCDyNOkzCaUHn3c
1gUb3JWIh2KVLFj/pzmhSxKPBkgY/VJXPwa8Qk5jynpYW1mHp3NSds4eB8b9zRLA
SELD1rH8mYdCcleoWTddz0yyN/JDcPVP++Vrw8/jv/xsGN323GOgxRk1NaT25bxD
Q6N9g64T7V9TcqgV76iqRUc/2xwWt/j+9GjwfrcpODpFgdLp+zsK1oJ3wE+Sjj6G
0E7PL+I8nJtw52vA3T+wIBJDhd+/gvx8gZ/Kjotv43996M9hBGJ106RVXR8CFpmy
iO9fWJAn1eWYnPe0Q1WsFtC09+swbWUX5CD+VJY3JV7wlDjPY4JqACNVm2tN/Ez5
YdxVJj29+eSwJ1cnxOj57X2Qy+fL8xfKwSKJveMbsdoKhT8K7fdI10LFXpprRE2S
/uurP6FhNgZodTH68dx6zW204IUrK2ltPHTVTg7bY1Pj+/bllrEOtlzXmBygX4Qe
m0tPRiAwb1lnpGyHDFVNo+2M/zaiMrlAgeX/jHUAvP8HxeK9g81VVVXVviA2sMAq
ND/wt8GBFN1vOUssDLnj/7ynWEnU18FlrWxB//ajOsMCp5eR2fYaT3tXU6rDxY5b
mKZ5MzwwZbgl2MQ0oylTXJ2bOqPUrFWEHFRwVV/Uh3qUAdmceYxgQ8NI0gNUXANA
bRC7TICeGXSz2On6NeRJa7fzVC6sSc/g1t0hsG/nThuVPa7xZyjevKxbXn5BO1L5
PRZegMAcZwjCWufJhDEW6hMNBIb79pqzj0Dw5Rb1D63Uy8g93roj+0R+ZQCdKx7b
43yIDbbFXtR1scxQRiJlUqhetZQHT3RmI91cVaVNnNjwX8pR+hjGiDetzDhRhc8z
vmhWWleL1kL6Lf3CqAbqcD6bHxz8q1ATHvxrLHDrSK7DNviVrfGw9WfJBCyQ7sOA
qSeF5LluL7LT9U/qZk1jWWD9I+ENRjrO1BSTSWRVdmwLOeGRajPVeeiLkBmNLJsG
qi2tx16wZNWrAw1Jey2mERV2QTH1oN2RKQZcDHFMB4kqnHA3HoboCGKKBvl8Y+6b
uUjV16/X/2YXdfec/c26t7paB7q43htvbYOYGVagDJ8bebWFoAoisdzRDlnxBTzN
WzU03R2YHqI9Er0vC1qqjdKVL+3VVl/78Lr1Jk+IBLjouh0CJYw6wkIklUBtWiAd
QNWlKtzXZmcujYZXbeE8QYq2WozpWE/TgHfSqnunuFZgh/CKHV1znYtEf5IqhfYA
NBRH8E81bekgo+Zc5TEH7hm4yNO+5fp2qGgEEpX8f+8WmX14yhuIFCCeqQnVoQS0
pbtUtyLOtB8NTWIxrLZIrLhg7SsEIw3UZEjSftBkD0PIAbBdXeBzPJ9SRWKNBy+Z
DW3K5VFdJzDI43Id3Eyez7FanBh/7gHdHN6qajxMXPUfSTCYKn47N+/ubDbXB5x8
ieV8XzgbSOGts2Ao1dBi4+qbkL042DhnU9XVZbd9H4z8JQqaG7PBIdT68DBzpbFo
vCsXfCvZ7Xqz4/40UIBGeAFDBd7jaRDgQGmu4FquH5KwGksZsjXGwMseAc8IRE8W
rlCyHej3JUFRdyfyR9hcc7WNXBBjXmYDVPwFYPwG/npjiomT6zRlfE8b9Kpu5XfU
MSF4igQTzGZyFuOxhlKblkPTsRXF/D6OCeCyCWEVaxBdxPwyWj+AYCIjQqGNcHvQ
OKDp46qA0UhY3sN2QxN336KjEeQJLhymokrogt0SKw5cVSGzIVN5JkYe7k2bAW7F
sOvK04v/A/FptDLuHqEZb/4mXkHwmsHEM+Un3HYRhRtRkLvsHA6M6SopkzHNNQS4
yY94MMIaxl16LOPRGUQjs4bbVMoghJE9Zfg1/+JCoKmNUAIcTW1QnRDstmPHFAfE
ru4XHFL/EbT9NODBoadLWlUg5bXKRXXw1UjJDQImxb+OzlC0GtorklzTlb1UN/zu
VkEkJTTRoRkShNTAT3Yj8iEJiVac0FWUXRYsYusOhz+jciUPs+iBt5tpfpP4ydAM
xYkcG6/wZ6nf87I24w0V/vAw3bo3m9Akwt+KnGUPUeRz0Fo6KwRc/RkougNnm9wZ
ej5CkYK+ITI9C5RFAhIHyfij903MfQ1PWvLd/bGuTaMZBbpkdHoOl2F/3RXGi3Ou
nE4pDUqBN8qDwiiuJ9T4NVmnlJOackr9mHIuUlygFOzX+dof29Mf4fG3x0khLU2G
yxOPFe4Q70Ve/EpGpR2X7sl9yI5/9nYbbCfqjfjLz1EzOuDszlOnn3vZRY2qqccH
b3a3AjrATD9ltRmBRPGP8/F/5nG0Tnp7R6QNtrWvkaP1SlqNaXJBQDe5uIgwYteT
1QBBMzonC1WUYxA1GyW+fR5Iurpfgv7+wvmiecw5qRYmqHGPJYMD39HXrEKajHsn
t+C4/VyzIXLQp0NTdbVfmUEv0nTpI9UPpRG5bGLFBoxt7f3nYidMyM3JPcoP0YRP
+k9obXrIHKjfSGevbqVmi+R3f5LQC37VxxJAb8YI3DUww17Q0thuRb7LSKsTZ1TX
i4TQtPG3n2UhzEmvsG0O4eipc9qxALWQJsZMKWI49xfcQRvJjbRtSMBUhxdziEES
u+GzRqVWErvOM5ZJbMfisWqaPGjzlIPiBXf6ON+s7zBnn+Gg9Z5LyZi/wZfErArX
Zw9weT5dnxbxrACnckVL7Yh06DbsEb5y7rcIwM6jL0M21Tb1y6U3ujgSoXUvFKX7
7Eeg3hTHp+5FQgmYjIDGzk7LeX1TlOH0LAktPOKKddL3l23UKGx1Xxu2ZRKcf44I
5MCByB6Gey+xWa/9GhbQozUyvLyTzQgAFa35dEXmeTOOfbY9dd/4EuomzHFbXU6D
HW/WDcjBsMczoqZAipXDXBBwKae07xGqNZGO8++bmw3ZEAd7iCbl/rOJub6x5Wdh
4lIjN/bTIrgQatS++X/0pWpkgWAVLiEgDastFTu8rezt+VjmQTTdpR9XHHONEsCQ
HeuTxU/2h+UtM8JMWEe+Oa6B1JzBPbXtZwnKXhCOo+TG0+fTgQ+r/CqnuY+TN93S
fRwEojVWhkXYpuhiS3u0g85zW9gTzVkZjlZWFvtPs5fj9kPkjAOUycUOjBff4aTX
7p0xDIDYS6SSzpK3cZLXeDTEoP7kNDMh81A7gsMTW172Fjy4xJaPW7RKuqa8xy4W
Fq35hI3ypoUj9M8NpDdgBEZgWqL2HfpEFSGdRQgVENkm0bSeaH1PBYAjYjEeUDYs
/9S6k6/Zk8ZrCTyVQYBSdyi/i7wVN7m7CiYbvQPXTiGl/5wItqXeSeMAPGotf/Fg
dlenUtuvrkIp92yvA3D4SbQnJJKY/7J11GSB4NwkOWeW5gNZiGqaQN1ByEnaF37A
sZuhOscwCGrtzBQuBPoKyRLrmvs1pxwEutaNjTDbL+ww2i57LonYic7mvLrlEvBd
CMMB50WveeuvvNOKKA0oKfU7NX0VokiWnkBN1TEFlqRjTR7HoTRIC6wvLIBJeDpt
ROEn+dsD5+jMQ8qlxdiptGXtGITs+tgTAp13H3viCA4XsOCT64KmRarYDDXg0p8F
+zjlDBMSfnyNRBNs4UIN6jpGu49jFCFRDFRwppJ8HDYS9uYyZUPNblxEFofmIBdl
PXPe3enKqsghtisxa50vfxSCzHgQLe18iM/H3tgtBVpP+IS6O44qyiXr1KVGm/Wh
1VTORR496LMTB0O2hrFeWXtIu17xH3ApqLc7A6pKxskirJkGlB0wUIfFGhL0mSta
9aNqbJQ5Xda5gWOxITR4CL+qHyks1Ye/n/iOqezexBszsnKrAl89KEvQqxkVNjNA
B3JcbeD8oNIZRpKPUpeTRUJQhHry/cPtG9qRJYy2oCcACzIis4+ZoRjD92zrz1xJ
bXH5zO1LJKl3HgFVo6WPjOBVjtYAaI44CR1dsUcWnVZhhtuMzzTjjLrGOnxpq/TL
TJw8DgXgdSMzXhU8/4tXXpKUKDgrsuvkcickEL1p3sUZa5+YrycaCAAzQXnvd87H
ctl4eKI1B/wKnGEpqjfhJX6DjmcBUUuf/DfHy2TZODV4u6s/h+oh9CTvwK2wNBS0
fg/WJf5PWun0wWJ0DJKw6JSVm+6Pml0KPnN0cYuAPJMCk6h5LEXBk8lYpyKBy2L9
a1+hcj6ottY7+wTJdLeDX51WQS4ravn8TglIc+i6AHqGKbuiIZaF5p6uu6JOooKI
5c2G05Z8oLFFeTDgh7fEBVt+uaFHOh/4UVRpt+2KfPdCb8h/t44JSNwXlwY8zyAZ
qNfUGEaH77hTERZfzrgIRdhfkZLTVNktXrvpQBgqMVPiFhrcaWvEhKsY1aZgEKIt
i4tUV04Uc4LBwWu+gjJZC6jeYrpL6HKXT0n9I9yXAJkbnuSSYacbB5U11Rn/WkBh
lbTBSZcvXu+FM/LSldMMQbC0FC+/4hfxUaUS8wNDS3K8y6upiXE9A1c7hRVwk1Vv
BuotYJBhQ2ZBsE7Cu1uglZbjM6LMAsK8PCCzPhTNn22I/PPFwd1JQQ7I3r6aKz8y
HMvCDV7nCbhYTrwLOK0wU5/MuEEdNDQczQMh+7yD6/Xw/swZgPcaK+3kLxKrzI6R
s6jFXN24B9MSyOQyPVZZRSqzBJHFB+GneeSR170VqZPOtvl2bXtuL976F0OJWvO0
xkdT1znpMiqL2Xbf3PyHu3rk3yMZ9ypAfZmRuXOdw4FbnuRR21GvZbvIpkfUwrEi
fFbOi4AThtLe9kx5FZMOvp/ma3G+K4CVg7CI+QZrkS7YG+wCvjZqqZSBxSNBJqkC
C/ySAMfFgF2Vmw4n/xV/YCyDL6FQAWknLCoAHZCh3efuWUWSlZzrKw+iaqRjPao9
BG9UPDQ1BZE0DZakY54ifMmik/n9qaIBp7j4m6rNHKmMbK7hG4+mTywYLpLiWvY1
bDi6CNAmlKwXcJF96pGdvX8Lv+Yn6AemthQ/rN0GatCr93g3KRvtQ7iTagSnL8Ix
XXP/4Tr9fI48Bx6hCDhG9FE7AMUgbFdzHUs/+sAF38nOChc+S6uAWrkQfC1AyuIG
c3amsHnqNcZ8lT7QkGnEKluQ3ZJg83RqV6srLudB5t6NGNajhVuJKuF9dGRA8w51
EoCk5JwlrbGorQLIBQNG/f1IQfXA4Ys+Xwr706nW12l/SIcBrskv8mH6GKBC8e+e
KejcZfjAlwDu8pLJK/FHn3gIIj0vxALfPlEVw3BIdLIvH0Lf+MO5rlk575kSdVJN
uKvsdgN0psbxJmPITzjS0g7aGI6Ex2MHUDTd9tSwru+DA7na47oskthC8X+lWIfx
nouLTmj3QMFo3GRgfYj6iAsFEeF/vU7SXzTRQLiIgFDTFs1nX6nVH+aPkoB0jOzW
GZv4Hfh6HpgFywrTKIy5fvHGJNX1+j0NOQNJG66AyTUp37d5Sfcamn7F5nl25ooJ
gj9tmQPfPI2vFcMBdvPM30YB9E0MKU8FoCBo3QGnEnO5kmDkTpKo88XYHWNBJH0A
NRlTLBawcUj3+JuwlCUL0U7NTx1WTLivHkNcfwVwPy7vGSy3SoJLqMw4nQjFrVxs
TQ591qFPKogPROZ8DmN54pA3/eRatg19QauolMXnjYjssS2/2epQYNS9etefTHh5
9RHDDeLBlngSgfThXgrsmZLtsmzIFvEkOWnSHNra4vCPfj1BAi2KZd1NNfSgqEJE
KTqPimdv0C98teAwGysulC77xfvS+6Px4Fn0tdcpaZz5GK+lc8VnJMvt9B7G8dj/
G0Vp7mLIJ95Hx4dCW9EBGkDHnZbQxk/46kbBd9vzR/2C+m1OtTfVGmRwNXFOOxnb
4dyQRBfCZTFAToBJmNoKKaxwCJl6UcQPPllc/u4zK2+ks+kjqnqS03UVhMdbKftU
iE73jZ4XJfSkDm16WgQRQj23f+9l6276oh/v6WEXLCSFQJTSWJDfs3cd7b8Isej3
6FJoxXJcinAbqu0/qc+foXYUdewLjmM94oPGMNkPJOuwx19wzoF4sKQJbMcPGaMY
4IxI+ID5u0d0anHlsxdyiXRVFjVrY8ZhLug3/Ig9ogp9JBQqJDo+tw93juzoQq2z
LuscCqrVwHqNOqWdG8WyNwsB2eM0kKiMHgNtY/4vhXsa+cJkmIgcZSVDIPa23vSe
zIW3Sbc0XjJdNhlwPkhLBbgbdHDm5r5Fq/4coJko3caAFBsCG3zGSE3JD+RVY1cF
ZC/ywvbpJW3uvMtHfW1cVW4KJHwjcqcid0Cmm5OtMeaqCYgiwRjqZLiqAQ5VyyW6
QwU6d1veGzzSRdH21KiAqCwlBCZzo/qXNWsUs9vtM0BFHhzrcyeps8XWtEvDuuFs
6vznmViwB4sWAyzf3MWl++foqaY8vzkbQ9Saf15QCWOahJCk7UXiu4eSsynDWkKI
0q7V5SF8iM/khESUmrRj1UaUJMG9V9v98OhNhBF4xn5TY3juGEerEb2URO3i+hog
kxO2Zzd4a60cBj2ICzXv4yEcqWQDn7e3NJ6gvlLB+LAzq23g7J2JD15EAaSU5dFy
bxvvZ02xVnzE0DYiwbs314YmYNn3vRtFbTCogqnAXr0qHWGTww0MnHrj4FjUntmj
4VIt7xhURrRQXW9PKpToi3dQiz+fVoS8pqGHG2oJcPcsEprl01cAdOfjxRIgYLyq
nmJ1BvjRMPGp8EPki1Q+1dgkN635iClD3k293Xk0W++bwI/iSl2Gzjz5rEuFqcdk
4OwU7o+JHIb3fSx7s7m0lqVnThqZNRx99NCKicvZfNh6M3Gna9g2doDP9ct9iwas
zB0rdKpG8JfWTSgazWGb3CpnoCrM+v8Q5B4k0A43Eq1FxM7D4AolERkLUJqfBmE2
cO4JPKedqBK37qJ6Y+Yeb72PPxhHGtflQjPkDuaNCtebUCZwKL9451cT6JwxVje2
aqaJjnA41Fhk2mHLM+yeLH29FeUSzQuGt7M09BmfpnC7De+WzmrC+ctJ+N0t9Rwn
+3a9OTSrLBcGVXfAoFauoPTaS3OVTp2b/Fc3irkt647bjAfkYXaKFE6BqlctTuTW
+ok4N/iBiYai11Zwkv+gpscrCjhWWPPBYjoMCmdXm6R5TQ1NEUYVjKhnHPfVxnsX
L5bLxB3SQQ5BoQVDq+HUIqjj3+r1hr9tf24Dc9QENLSgkhQA2FBn/fOjSwP1ROP3
454IOk3NER8IvU9i97b/0sKvnWQ+mXhWVv13Hfcqki2LXX3Nd/wOzIeD+NuYDIpQ
95Ws8SpnT0wxEmvPwTwezVh+ngYsmjYkiAcF8WWO5OXHKqgoFApCYEWP0PXoMr5g
DSK1n8sp0Vd5nFTXd/ECh/iSebxJdG5Ojj0ecL7LK95K13CDASy2aW/HuW/1dPXV
YbRBUzd5KFB4iYb0baselntnTDjpoRPEKejCV3pursGMJ9l9uyzSwe7GGjkWmXeF
cykMyJonjbk8eKERr5xQboPwMMvkirnpryJb2XlnTNoVj4GwhkP583MuJ+sVQJqj
QmTl/962fYeMP02xbZ+A7I04rnFCSWlgOwxC5tUXyo5/NoObzvw4+lJK5z4J/NCw
qlC6IngP66FgnkR0FxjgW8WmAAghci1o2u5UxsqXFzpip2xUUYVit4MqcpaaL0yu
P+wia/OFW6T9cGzgHklnzUkWQZjH+RexB7mpgOSt4BG3o30Tqii7cbq2ucKAmr5u
S1BAe769s6c7zH/6bXZR5dpeyYT3m31L5iMiGHT48VI9wae4F3CWIjpWVoDgGYM4
jZ6K8KrxuAcwmr7yRy37y1//rDrFZWIh8Yhs8ig9Zhhzi6HaD5O1/NWsjBqI7ESx
jNxQzOfBU7oMo82bIL527IHxsSQp23eWRHCuUb6DKl4SnuOMSQxKK+RkyK+Kq467
837CqnJtnUGRE4hLSBpmwRihO4UKQ/dqrokiFW9HUPcs90YbxHiREhRcPTV4oeM1
Bnqze08G/EApdWIsBG/3MBJqjFLRt/UVM0Pko3i6HE5wWTFvAwxOoZ4nA9F8gNtH
ElE1zP7/Th+VD1ggiBrxb6eBccpt8GbkzrpMokhL9l0jXoABE31hKi92Xr2vLU22
cXUlzVDSQoeFMuOiG49+JZojs1R57L2/HgPaMIZbwWlx+As1ojw+Ecr6EwdkUNVp
SqIgKQk8f+abkQfIcXm7xSGgdi8hLOUTAfZMXT11wA3h3In8IkhBwfeWhwOR0JHw
iPeYAD3Abj1gbnNbifEofSBgXV+/MD6qjpndsH65PHRwifgvXQy29BDWOWMj3AU9
1RC1jyNBVvMWMdCTRHooVCw2474BA4imqMAdn9fHwWnh6xPehSlCv9bE0SIF4I0+
ayKarmAdCRtSx1WLkRFVURJAOzrCb/pnvs8eK5bbDxPmlZcrkSBaJtGHAPjpv/bx
rPvw7YNAIGnLlGK7IACgsCud4i7F0H12ekEGYxe+iS8wZ7k6hhTBwqRw2dhfc3oG
Aerh2HNXZCCBUi1wuisfUsA989oPJSgU67rR5EK0wmDaLudRqssFR1AB6XROU4CH
F99guEHaRWR5M1w172KbdmW4dlbAfzHuoa67ELjNnQJED2UYgz2zkBaXdPXS0sMs
qSF8E+LwCEog8LflD/Xxczke0oLT6tHwNdZLRKwNWcd8/i7wNp49HgX0XwBKF7qV
B5LfkXjuHw30Acq5INzzlGMKiDUCg1hAgOojRXYGb0x5oIaaZjK3gd+tqjRLOtgW
/kEzqb0JWWYjyRl3kHNg6MISlytyjtqFVXomp5Z7fPCf7yE/wkCSaQoOCyOEiXvq
xYJnZjl+MQZRN6mdGbSBazhNPSxx6DfhPJ3MRqjpYuJ1mVg06YuD0Nx5Yslx4P3v
wCCyg6HlO50D2JxSy7iO+lrw6Vz21lMoYLE8qz1jAmP08OLUPogMH4LnZYiVmJ6p
qUuE3idzn133CppC8YNGVBo/5D1Oce0QeCH6zpJJeEY=
//pragma protect end_data_block
//pragma protect digest_block
DSr+pSlOCVdZRIoLGJSK77Yc4RI=
//pragma protect end_digest_block
//pragma protect end_protected
