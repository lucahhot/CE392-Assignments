`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PBLVtdNY1CBHasnysRHiFM5gXfu9jPbfJgCiBVnZ2yprymcAhloglDt4dpeRyTJE
igg0eJ32yzW4iPu9jaNDvnE3S4xM6wzfLSHdm90qMbAjNO7tekXg2iVDxNxvNiyH
kBMGFLHhWUlVdi+xMLYBv/QmFjx9DtNPWk+fBQhXNko=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 108224)
dXbsoprMQtMnkPvYwCHBPncyRu99/0Y9Y2P46oNUYQ6nW78ngZCjnZLLcxMSVNfX
wQ5DGWc9LM4PulhtMtwv2WI7z19Q07P/SX9QVKRnNRq0x2QwiytUio4HSyTb9x1s
DmudzGKneMIwWbVqCE3YeeUmIjlwKKiLwTplDtyGeDQvYEhmvpJsHkUfzs5JIzfc
iLhb+EpybDDgFMlaxYBfTlBKd1p4KUxD4pA6az18M+lRL/d41fgbg9ssPK4sROQT
77lBGSU3JYvwnl5TdRfhR9doBBOdUMO0a3kk8kro+dCrF9Ds0z2VPJ6XDRTRJo6k
CmhkcJGJveCCw1aQwy+T4pnBQleSlkfi2vkKxoU5yTemw+PFovM+L4lPyouEX16S
XjX6WXPhz0fsIHZggwGhd3N7SAGA2zBWMqdp52MbhMrHK422EIN9tEOlBiZ1Naky
EKuQf+deu6ZAL1mXZTpPy45o3KpsvOwlHfhzRltChiTPIKu3/ANsR4mZZ+e0I8WT
dXgLeOJcuBoHY8Z6bhblpn+z7dTqEYLNj3lWE8JprvbegKeC5rRut0u/caEdk/5C
ATEnyR0yGVvkA9eTEpsTcTJNWFq3ITXqzzah8MmzKv1+cbT4qNdS+sATdXHl71Fs
/4WBSVfqHXmLq2y1ehO2FlqYSh1yGA7HPd3Q0hMOMQhAIy9lH5oD1StX3KcYk2dw
zwqstiqL6TD+iqWlTOgxXCsO1CzbYzvUuv/fRIw32WiOpfuetKlzRe62xQVGHuco
BbM2uMG4531m5+phWSrNwOSftga/NX5KwLiLBI4AQgrGs1fgyLtz+abNjZIfagU0
KiwgNcDSh2sCf8Fap+ll2i47homff5VyBtikKwpkY/tuLNJ18/otNDTg9dfpz+RN
SRbBQzTnZRQe6QxCg39eNspqxEn4MMNpiPjz+71GliHz7AqX71Nq2qI42jGI6oKu
hHPC8VCzQNCRJHHAAkQjnHPQAwUl/JCbnAINMOCdylXEFvC9qcJpKbPugOpnYQ9c
mYQqgS1ptWWNV86PdIP3BMNcVAB/eBvnMh+NNYSGtgyBf8afPsnklDgUCKWkxvmK
M/o0ncY1NtOMRfQk1ph/L6cVrcrSAmVYuntsM82ENYJUWHCCmwEDTVYxwqXx8arR
fwaw6yMDRPJio8aoHFxx8TL6a7CLkSfwOgJFhBvWmAd8eGnWIcp5kpOb45gIcglM
LJBYOb+9E9s8fhXvutEIVxIYVgh/JGQPEWSXAMNXhwJgN2CR5nuaiI/79ny5mVQj
cy2zxhE1J2+2hl5xjxruxuqBxm2wkvQyygPADyNC/fR0E/h9zIGDa1D48fg9aH/G
8T9APcC7XagWrexHUpjOniR6Wj2ErCbysW5s+DaOKktK2tfdRJyaBT7HVGj9UiP4
1xM9G5q5kb8Fq5/3u4widYcoE+C0pnZt+72RG80Kit7svR7kdsdgBrW9W85Y116S
kZpLZ1xx16rbZrpKufDrXN3Z7wgFp+wbXrXTYplgH8gJtjeOhCjVYlFaRxGvv1OE
6YNM/T9Ny1FKj+zd2lT5SseCvS/aQVDb98cWtSCv1gTZaLxbn6p/5oAFS/H4ozYl
nJN7rKdQkzJqzcEBfKSmszIVxhc30FmJuwG8t0KCrcmiwtlMmM1v+P3FkBLQkt9w
SPBLzIrR1dU3FHO55M+IpVDhxzx25F4bC+PqaeXex6WbKfnLezQgY9Z7Gh2B7+Eg
WB5CYilARdAYGfd0xhgDEj+cux8yBptWgfbhXlVEcbshwy0Olh2Hvz2gljXXeZoW
4Ls5iRH+xd/3Nl5dCx+7EwWHNSUOzXtqAH6Mm28chBaOr/ywe2cETgRwqjWvyevw
hLLP71hxZltiyEw9PD+YQlS5vawAub5RfouYdDrSKSEVDjsoj6QXC/7yAr8y4M70
vWCHbsQfHiGz+73FH+DMVv3mz1gB+vpajxO8vzq0tP9Q6Imsg+hYJTj+WkRMqe8i
1CUFkr9otFskcKIXt77zU5kJIN89+jVQwmdSrsv1oewuj8wTsuh14I4ZTfj8/k/4
Ih2EegDN7xYoYUYb7G4mYGzAxCItnb4J6QKu626CwCknBw0YyQv12jE0ECPFAz5x
ki1BzW/W8mY2zGOt5HWcBZt2svCWaZ3jweYU1slqWv7VgexxMVuIwSKhJGar9n+W
NtIuy3aGPBkw5VdnNBnzLDTFzHtKyxPhJV4sCNhwlW1+rrtzzjUxlSiHRmvypQ/W
cBbdP3euruvYtRxuNWZfH6c/vQOufubQCWghtDsPNF2Pjr/y2MUQn5AfSY/gN3kZ
du9ncJ1zTGl1UnKCxdcpzM/Ij5PAt5VcRUNcDhwFfBXCcemufYyU4ZmASWyNEI9S
1jJYgjTJfZXe2/lqRB1sJXS8uos5h7h4Xeall9uMigmRIK0zBACfva1UOqft/ZN5
wH+3IhobLmiPx8IPHHWcXoSQ2CZmmWW7TD0OaJwYrB+AEreSEeCiaVHRJQZ35mjY
bW7/gitlwVQ+wCnQ+hMZkV7w6zGWcfHclvwUrv5kvXcx9zLN4tVGY5VRLZRgqX1d
9g/JhB6YzUytXTz8LmAipk4yXGLT9d032wlg9BaVSxXu6+GKa93mNcKuMfGRhB55
kOjNwgGW6iZJiK/m5m1IiouehnyQfJ1QI/UvZTOSCQYz/Ueogo/Feqj0uiUPyVpx
51A0+IUnUWdjPHTSd+x5R1LKvEpjvEvbvbhhkeP4/D0UMwyfO+bE/aafCkiTAQf9
DioG1HVro1W9JyvEMyRIumSDxxNY4eyEONTNn402ZbfD4UdtCQAOdIXGzeFpQsv1
/LsDS9q66zG5oIQNCt9PrR0HNrD5/YN93rt+65P1oWPH7Vk3r8WQyT1KbkDlLL5g
OkR5nK0PIXkVpISXU3E0+qWB2fV4RqWh6T1T67ivaD3sWJVBFAAtSImJlccMeJXM
XQBOAoyAYRgZ06bRlv2cdOxzndgZD00u6VthqoGcNDBeVbu8PmyMbdzmPHXNDxhX
vbcSHgTgzPw0/eapQlStWxzXlCAcArN93bWrUzzWplbzwo7qFLk5MZr02h5tiafA
edoWeVI+tHz+vJeNl0yruZ3NzNBFEE0Lw7rpX/WxwxVB4Pqm1RSap6Z/bytY7IFg
6NSrUK7kAEjA0p1NTqTx5XkBcsXyLC5JunX9/LB9OtxDQoXWPpD8j0tOy+evrBpH
psocoV9NGqCgyd1DI/kX2kyECgR011b8T7mCjYDHUTUH6ibfXJDdZWoqC9XJYkma
T4nNtg2noQ77JgIua6Qxf613SGO1OjtiA7nXqQoDBIvLCcB+FXEs9R8J3DBXHAoz
f9HHgcTndPSVy2UXNBa/+b9f62bwdpJ0B5HGW/1FpU8iyVQWM1gAgFDphjJQE/0/
ZxDxuT26bXpy0g6NXlkdbWWPksCOrDB6QmfjCURfLa9SOx+eYkTLp7OdVPwh9quQ
aAv1BusGE5/xraMETA97n6xeNA8f4v+PcvFqKZTdTk1W9i9d/hCHud1TfnvPG/KV
nEnenx80zF8MtGba/iu7AqLoMkLX6Tvz1bGqT6DM/HtGovkJeVuknoZnULiHmWJL
2TfU+jw4BErP4+ilXdDwnqWtd9y/U2T0FW1M/oPKmEuDb5e1IiWqto83z4P8lH3/
WFDCG8V5BB91Lf0EBUR0VRB34CSpGk1vdFdwWqrqG7y0QoVvElwKPFHCVp/HTpNS
ko/GHj6DBlAXj1YPHzj8RjReB2uSFL5hKylVqaNifZJxlCOWtSWHAlqjxtmypQfW
LRzAavXQK9V8vKgQB5wUHKmYWx/3jciLirxpjC9QhtemdLJD3RLMrHfseUHQxBXG
8qul6/CwRP2KpiWsvWpmZxijyw/GtKePMgepLeNSODFV2H8PseN5zIbluL25/rgO
3iyOpaw9TyLdCebw88n6YLfTzFpzsr65FBYEGDGclrZvAKHa8LptcLQ4E3aB8jIY
6aOGQTMToEhQ9J/S2Xx4gA6sksWxRevxKhBENPCq716YAo2uza85j88U6GAcTRCa
trXxA44x8lRFGjWBgxD7lb+m82aErLojKb4Y2HjQ5gwDsv0Vwpnu15/TyP9m6CSg
2GqOD5e0hPTJJGemK69fr8PHE05qSvd7qRA61Rv8AWFEFWF1E4WnVAX/ryZa3YS4
eHO6pErapKJcy09sIrSwyKGJ7zhLzAz/WxEcHzgbrq0rgvxtxBG+ekmtuqYOhVCH
9F4X9vcTdpoWeBPVEp2gf4Bb3HnBSZIkwV4uPxhjNnR9vil+YvB8+XFqUIl1X2fp
vWye3KVuobPGePOwmw4CTUMVuKRw/yxc5F3Cn3suWsAqgWKru6TBPjkldFwLdo54
sLMbJJMS+fujCO2jjY9wqpHpY+zC7p3osZseQauG6+nAV8akWVwLvO9cZXsMeF1t
gskDrJpxYg1x26NWp/EvrF1FjOE+h2ChRFqL8WkUF92btIrxEM9reQ0ZqCNZELHf
oQeid3uRW/9u7XHNLMyqrb1OEtxz3hzO19ZGsMhf6IaQMLB0KwQOEqy1Eslxk2sF
+NTzfVHa9Fe4GWT9bUKu81i5gOXOLWUw5M4kGhV9FgosGQ0WK+GFv71BPdzgtxp5
shsimvqfu54zCRaR/bRKmu3HL45LzxGkxNjJMVc+4MX0PMUTU81FpwMKES+A5gA0
dSH62ypb/Mc+P70ppCKiTtWgp9m8XH1NfE+h+PtNpvlbTtz/NFVIRsM96iHMDoS+
bZCc773gdg3cX1pzv1FlRBXm98k0YVGw1NZhXWBORsdXAdZBx64QL02Muh7tzg7R
sb2370fVJ2B34WSDZHf41REjEZ2rlRLwILNq/Jx51BSEzaaxq1AxyUOG436aM3b4
Jm3Cav8MQnd438HNf+zop/9Kc5l7HzI5/jDbIcPRpeYdIQzvDSgat3NI2w+hffp+
LWRtSNVAVHWh0JfbcCGlIMIXencSYPffU97bimom5HlMApqBivkXFEUouS5zMTrV
MeL+ZN1QAtsZUz6fUclCQFZzpdMDUkNGYKiHCEAjAHHpBQ+w/W4ok2/BU5JUJa82
Hear4XTX6+lVrK2A81PymotZqhzq5EwbChXFa7vYp+gkMVwZ4WReuLd+1NvkwOmk
5DVQnbL8wnaneqgtFFVG5CzCXd1FGB6hEDXy5Ova7lS+8k6fdrRGIplANHZ3VmOw
l3zOQhdwpr0rneHMI9zEtdO8cQYAbi+mCHn+N7O0VhQrgYZHD0cn/p9yPC823JeX
0RGevyW8p97Tk0VYAk5Fe+ZdPUm2eEpHxOpToJuMiLA+BUhEKIF6Rr0Fbccust80
OYTrVok6dqk8DKtov3dyZNYbfxnMx8pZbRdDvv56ic+DpFc3m4bc6Kgqb08B6RKJ
MDTIU+AEOR/lLYr9nGmTwq20eNwO/vZVflnokNXdx74aLo1CYp8YsOPYB0QhQhFF
47vReaAPa3aLZMaVt6ynRJ5B2nJ1+u/yAGdtjWzAKIULl9I7+Qyfym7+Iqdij/8a
fNJsRnP2g+oEnfqZ67bh/WgMA5FDc6aPezgT7IRmPFplGTpa2WCsdjvarur+259u
Aeqm1FNK7woh7EwxCA6SAwWKxy74PhXhisIGnwqQzAy42/hHKZnm0+9M3wO2pEbl
bqFy9p00God+GT6nB6VL1hRBqEOhm8FlYt2WCoVp7+7Q8sAKMCj/hVn934tw4uLY
1dPrwxXDRrlJ+kaDjYuCdvJcdQHEK4o3avj3Hu6GKd3eIbutTuazktNen3wJeXLs
xhfZpItBbtxMhJF9Gf5hyCuQ7I8bQBZ2fBhm85I9Y1B4UZu5ld4eXfdvKL2NERSD
Ral6tIfxNKrMWJZZKH22QvUTimJmybfiwR+uT8nZxouRexFukc2ZJKqNPqwoGOgd
nL6tcV9e87zVQfYsiB+v9WW2+4uo9URHXVKMaJBu8VVYII/of2Bs6g6VOQwUEqYi
9OHKcll3trQde2RBr0lmnB+WPaBifbvdr0FZo5rDLZ6BAulQVjqLKUSpVflrhYoa
HhDwzI52T6DTATwjHk8g+n1q1S+PFCmv0RsoFmrEsdQ7p8MuYl1PUf6tOCYgVzmv
YKzul3dFViuU21dagAd9fRyEpAd+GwCKv6gvGDXFtlwDterIb7BZV/uawmjpLpDl
LNya5cV+7l4odxK7PEzF8vFC2EHDdbAFtrYmgKlRc9hga1SFIvP1CUyg0slFD1ee
fcqQzWkjIa3waJZ9Z+d3DoQNpySW06GeQMcX2fqhfAFJH0PpNzNhShvm167bL7hQ
+Z7vDHvPUPbOB94NiAjJXzgKAudqv784jYs0qstnDWhXgYb9sKp+lRanB2yMENBH
9M6HjynxZlyQqD/Ky4LECKu9TbJWgdlomWJjrSkNtp53gl165yzzrYJtt8jGFdUY
1JOSIBlnr2n3T9ErFuPurcz5GW3pIYnr5hvkXL34Oemt/ObZ2Go2EcEYEUf0DSb3
FucydJPA6Aj6LuWX4DyV1z48v4TX1AkIrSGgRe3Jl67rdsjl7/86HPG2ki0kQX7J
D+vMFNtDXlmBfFiXcUvHpj018/MQ3tdl0sDujmFHBbGqVdtrPBnZV1sD1EeR+Xn+
UUlud7Y3161qjHX6Awk/HtA6jQAx6BO/mFQ8ion60n3hi81kDM6csWPV54AuJiPG
UrV3lcaU+1qzd/dhfgiqWebX6QjBYOuZTrFO0ZJpVRSRseo2XpWiBWf55nZ02sTc
2+cGRZILebRJ0EeLzRx4tef/LdEeKRcsm54yWktGrk/mPuNV+Z3T87/ekKNsVemg
ajESbfrEkmzIxbUBTgwvUG7qLbiplxM9hVLoCFYEKAYE7IuyqHO8L8QDJUmP9sT4
RvDszADfKS2k7d8q1rrS0Y/orX+DwYfoEGzntrQDe7jIn5XhwpykEvlG5BQB6ys6
GrviIuhcjCT0RwsoA9FZIkGS5IjEouwtpJDJBTp+T0ZDcIMnqR71Py05WUGeBk+D
Kgk6AHjzFYsDsVQC9a9Z6M4xLC6/YrJaGaeE6DCuO+rr+P20O2sxrSyPBC0P4tSg
2addMvnetAb+6RxaAVfEGP31yCCa9AO1RWE3148EyFlIxFkXR9EPLie3Ot9GnRjE
7I2ivOX/GxKZh0Lk8b7Z6iGTBZous3t7YMJpdqNqDJ+pjky7qcDFOrdtv9Q+FosE
NZTdqPK4ABGfbZaNaGXU6Ae3BwCfEkJDMga8k8YXtJ/QWFRVRzKigqxYDgbPxMVq
pxIfJt4UFlgURBbQePf7ko3c7NHQ2MFXq5rehBZHwpJnlsX/06P//wS+KvtqCKQE
67XAOkKL6Cw0iDlXBKXJKjvjH8jZzqdC6v2T8AjPiW32NeMAMSpgQp46/MTQ4giE
0L5P3/G+MTnmZScCoga9mOamd0PIAIZdTYjxOJYZS2JkHxM0/v5KF+EtRc70OlSI
guO4HJUe6pmT8evsB3njekwWuudRqdPQgtidcRwab4diMDgMOtaRvrWilLBDcRgy
BjQYzSkX7Ov+HQSN8XPfruwL1T6mstztUxPqjcRKmv11JAkLxM9Ivz5dKohKFXzV
1dEay+lzaAXPLA6+KTAARNcsmOw+OTDTAZ7iICXlDBNX53AsRDNXf2w4rniuy2Fh
ko4ZzQ61bGcSIqo5ARtFrAHGgTKo6LMc6KAUZ3zOASgWJtMM7drnmt/HjWVDd9Kq
Egu+xdBMeiTxdyVxqZFOy2IGdTTD2czpbD4vH5s/Gb7+Aww2Smf+eVwdUc/eXB4B
u1Yd4ImLtdJDB3JKndYaQUqa1xajQ0rp3tWFKsYE7mgjPKf/ii9voip7s1OlUtqO
N3JVxlzzlolRiQr0ycNa8mU/H1oBUTdADvPz31LhQGgE6S7O4SzNoo0omK2a7Hi1
EYPcDlOAj/4VLeIS1/QFFJZa891I2b+wzCbJdQtL+3UTwOUlfomQ39NSaQ4FmC1C
WcE0CcI++B9zOvjl0qFk6cixk26hAZo5xAJvHIhA3FVlRVwZH+roXRkXepMw55ha
voS/TeRC2La/fAHMdihwr4pU0vElxv+hMF1/+7ObBXUiC9tDt6d5uVksd92F76PV
81TK0xZLz11IvMxg9Nz8R2/diVIuQuAX6VLkllnO7cY2WLhFkrJDn6B7Wo4CelbI
rsI5QIvKwP7s81ZYSphidz9ZYpRQ+dyW9UNunzO73PzFSStkka9EAiUvZ//kBwsG
irsGNqC4fhh93KPv9CyX3ZXZCN1xXgOrh3KZUQ92kGNAwiilyk43lbnmm93BhgDC
EtVWYbZrreHpuSp/wntsFrMNJrral0o4fndCpSS2YRxpD/grEfYcOpHfQNk4yjJc
gbLyI8mebW1/cg9/CgH/EDTsydWKA/YZtcJE456tYib8Qnk/SC1TeYYWCaYcRtCV
+uWjQrCGlzyIyT/F/BJxZvWjvxvHTa6jKGwnJnWjO2evETiRhB1HDHSw+sKRwi3B
kfH0DqJlFSfbd8+ocPQrznbTOPOrlJJah/EMXXEwy7uAgmS8OgzIAc/hNBygMydr
U/eaKZQR6OMsSJUC8VFLPwh1Cf6EfRj/qEt3+bPBkFr/xVEd512jfFlVv1blHyyR
/RdlK0JJCi1B6tCRRUdkYmtWyci3w57d+D7Pi8JmQQLYkQsAYr7TUL79u9qEgrge
Gx9aI6+Biz7OJinOEodSTUTLqwWN3W369kIcr1CCrWFNElLKlRxIMQbtoao+Cq+7
ihOoFlNLzDFjdIIrlPpTCiMcgr6lJkMlG1DeiXDdGVPwSYnZXqFq3XVIqsScVRtM
uybAr8fRrKw/ipN8LWKoIO+EmR8oAENAGnhinzsmHwFVud/NIMwmw0zgjy+cxuKh
89jj1e1yyIQ+PkVEHnOj/bdsxiEqUVJmVZkZYbq+cNBGhZg9bo5eUOr/MHKI72rP
Az9LJjvuguYL0HkCnkNpPmGIc7ysW3dCwzxP3xy1D5J5yzU8m2UpP7Fbx9UvBfkE
EVfTm2t8wxxn+nWIQLuNAZc0YstFScXneRtqv44/sTn+gJJ3D6pV27nOrmioLQUE
qPGalOIBuWLw4oEv7hhw8v4TC01w4U8cZbqNP8jNbhc1wBotIzPmj30PSAOcEZPE
xLD4tynNU4HCMW4rKp30fZsn+NPN58weHE0V1LAXO1vb4xp1R5ojmzqmoZQ7a1AW
AXA4yxfU6kJ8DTqnqr5r5njyaqhH/SrLARScy2EACMHuSY6N7U1z2HZwNC25qOrD
M4VVpiV1T1DYt3JOyWXiD74LGK1f8pNF3OkKPYqrTKlIcD+llyc20osK1klXjWHf
HokyX0T33Nec/pgYTpafcR18eqx37bUdF1heb5rUc4RBjlH2qEw+ECecig4FSHxI
15NZtPbrb4qpX7VTvcK6xHLDAJ4+zGghQMIyoPfY/pZNWQgMpeZRCkmfGE+HXT4i
L1DmNWeN6K9q+pMfBTF06P6XAEcD+ZiJ3ydTVGSsaBQk2OtqvHLLOmr2gKyn7DGA
FRZpwna970vyC2bso8UufNXQ6j9YVfglHlSWTMpBOalpLmBIPF00qGXfmmnQf1Bw
a0ZTMSiv5Efrs2h9usRPggueJhkMKW0ob+4Vq9Qzj55Ny6DCn538R4T0kSoCin25
SrM6kN6VlOl6HCAgKiJYx3zybhP9sNSH1qwlrEXfpz6+9dDakYn5T+7kKS6Q3LD5
Txu8np6vyF4R6UaLRTMHqcmtuULm409ajHGhy0tGWmsHFH2ATmn03heFBj8vSffb
6jYhjkhPmNOsQQL5M/dVutB0KWanAoXucFu6xuT/vMYoBpnfm5rSAwH2En2MPBF+
ESDzSqG/cQl10rJK4sC4hV2McU6tdCPaVCVeZ16IuDSzf+asXm5i3Kj0do1XsAKS
TNMNhJXJNadp651o9Tyc2GGZwQz42R1Mp143/p1Rmz31cIHj8mR0d/H/76994rQ4
VZJESuUUVNkmTgGNmwQhJoE0Yc7w/56IzDT6XRCDmhnQ4Z2JB4V3uZkFdGE/CjoH
17Lib4YkDXOPzesL5EsK62dssuUO3gD2AilblrqirWLjREpVraPUdy/k6V6nwiva
wXczOnaWwKXQubbD8IiZVadCrUDmDWAfAvSKfj/6mGiAsfc1MrAVx72l/hEY9OIm
JK3DNAiDFZ8NdsRY4NM4HMHuQ5GYkPnaESWIsg5psaHoRlStyDg+4bf7neufNI5b
oHKIKwzkVZXpDzmenbfUJD4f45j7pKrS5PBTEBj+WOZXF9NJJBI17GGm6h1gPVi1
iW4icvgmbGO+Hrl3U/BazZkCkD7+vJlOu+6e2KcH749koJ3BbeASW9zvSSOAhlv+
YfqXRLzGKfC319g4Qvgq2YDbPzwNsKKK/JtGURExHl0RwmatSy5nHAjtB063BXtG
HNw+jH6ZosNsF14syveV/Yy4Om511alRM4+VfzGgsPzoU/3cnPVXOkXtgLVNgqBr
VXgAKP6R/rx7jScYMPXbVz9AsSXUBvVX0dZA7qIGKNyAVop2pct32bML+mNwcsio
mf9Ni8paBCW1qSQ+vEvDUac1mclE0uboUvS/PiRVA3ynwek1URB+miMZqbkwbAr0
cuMdp2PBCkYvDpEUOsbq/cz1W0GWzJ+LeOg1+3Em3Oxe0G0JQqh74nEIS52gQINH
hhoAazaD0L7AHgcHd5fqMOPPhPZG7YFrZzlWf9TjTyGhUoFMUZBQy+a41dzRkpZu
T99PBfEAW70NsjWZvpjh0J4uXfXZq+OvS8+KA1qEe0wzTdfDoNjDQBr3f/UnDxQL
t4stBQykpQFa86DIhUDRMzmZsX3djlQWd+B3Co2QfLoIQ7O37cACskHgbX5SL85v
c+RJzhuiEx6B6Co6/PhdxSNaKVw9+3/cmRkx3MTxqmasoHd6t6YR95ssAe28iTGp
M48JU2RCDP0ojexZt+WCxtjtIQxaLEJPDyAKJ85HKfA1gX18iTxobQjNuHEvQgUk
kXogZHG+5XHQO9xAmFxUKB0CbiY4Dg6wkQRPZ+I5SF3vcK7d15sPwTBcwzwtJcne
j25f0t/LxYBxqxxEbZW+ra2nbM6xzY5fHz3/r2nuNpvVTjq2uGmYmtGNsRfABJHH
MnmVBYQZL2r2KAP2njKR78cWpOlJ3FgiJ8UuLm2sEgwaMIQcG/ShiG6hXeX9vwhL
YNAEaedVNJB4VRasT71XvSz7m8LDZ8w3wOIhlKWAB4tRAytpHcGgz7KyOYJBzhEU
Q7kWecbTI9d65wPkraow5c9XBrPetBokFCkSEl3KeK2n0m8a/GZ3Q2YfA38k2JIW
PDn7J3Pxdil5GmQYIy+CIICV27+Ls4UG8l3a2mTEE+VD3Oqk7M+9pymU2gQ7YnAl
9+0OMqcGHd68aRUpU0Lr+k0nlOq5fz3fXiBZdXz8x+pBYDkjR2y9JFjil7zDUuG9
0IIUKdMO3F5AHf/aVfMFjo6H4HbLBEUIm7ISheX2au+e2o1dnqY+AAHaCHg+Qz3m
Bwci7ltazS9aKYuHAE6FeROChpmGxjXV4DVI6AwrTx39/i4PTYF9mubCwWmIckPu
yp9z2qWxvusR+hXZXSbLY94byuKNLVJ/NZR4AHEN0q+5a+WvS0/WotyeJTSXaFR4
STt4BejxtdFW4rH8Dp7a2B+IELCIx/XVLoC1Al3FIMxCrXADJa8B80xEtL2O4AXV
FQOFN/Op3J13CYJJ0/N2g2+eQ/83sNwEGVWLDetBkKydt+hpDvMs3yjL1SB5L/vi
cyePKC8V7906oDJdVSfNjF246M/P7DS7vGnU+esG3LsfwPE0R5g/zv2Y1hORo28W
B3HmBhHn6KGeYBXE4IiygTfW7hZviwwgkX3A4+B65RLhGMUx/13OAuOtinl/IdUU
BdqkOsSKe8aHLfubXQjc3sH+l76I4D2Fy9/AaOoUmw3s+SVu7B0VUal4fI8AsBhQ
yKHL6EWIB8RDcaI/fqimCcajRuZeIJhpDyQeCvN3sRib7KaXxXyfokvFINT/LbvQ
zenUx1aP+f8GRMBoOkqILqwyTgK1aMQUoUpTpEsqBijBafoJ+UqhiwNipNDZ2FmD
pT/qlZMb+MC+f35BJsr+XHuBv4Rm/18dZQz3Qadu/bZ4TSHHhGJd3+Un3a1dMDt4
uOxhXQ8S3oGv2SOTRQFiKwXS7lm0hM883FY32WnxtkqN4MejDliGmcCGpXifv2kc
lURvtP5zDtJyOoN2WgiZy8HeEE4aDBR0rhqJtQP3moJ6B7CyvHM1NWEwMf6iN5A+
roj1MM1+WgEVxfbEEIATzg6RrenCo3Vv+w0CnfFAeA+Py84VgBBCtLhE65jeaWtC
QuVKTcsFHnV2WMivvj9rI77WaKfrxlBVPATx0KQD2RBiZ/MCZ3bqAcnwlIdTISAV
bOSJaJ9j70mlSCFi92Hiar7vQDs2r0mt/DDatI7Yeps6aZtx9pjfG7YudnIsSXzo
zvPJ3DBuUPnr5jZTwAyfKcpuLnTZPGY0MDgtLS2LSoy/AqRKKyhzuKTuHILIfcJS
SBkJsr8VHQ0vSMWpQ1MNtD/wpMOuRp82aWDxbcTArT7FE/zgxRtgPj4usJvJE7XX
MOFnwCv3WPXGRPZzxIfGK74dS084z36ES2kmV6brbNuJU6lVmkvlaJsH/hEx+mRA
6qegK+IMD/4h652tyCC723f36e5qMxG8yXFQamYRL9azxlxguBsRVDabPKxIniaT
DfJeY00DKfyp9NbQtTh7Mqr6iHN8dT69xPOsoiUrGmCLIzI7aLBn7yYUG6gA/nsZ
KENtAzOUajWl0u/KRGC9nSUdEh3kuCOGpVqjzdJlzoBV3scYxJV6PcO6e82rumZU
4saaH/2sR1OyyjGO/Vk59xhSwWzjwRe0dOUFNpsQnbdktr7LMBOs1K1D5Phx1lQK
7dPYqRn7UWLTreybQuU/CKDrr7fBj9i8gdjhSharZslwYOEBlqVTwQfjv6l3Tunu
Ib4xs0aPtVLO5fGqihO6e/7qxMOrpgbHkcDOKoxJnqjXArYWLq471o1sNImrRpMg
nzGEiOj5a0bhH/c2xWXhnYbAsUHu8DBOKb9P28txZWivwE1OYjRD9YtM23YNDaUo
FIv+LQwoEAbRyMpnszHsrusrDN94QVCgiaPpzR13ZSlOAIQ0dPu/6Bq3faunoL6c
9cQbRz7bntySAzOJ2VmsFLFvFVb/w+x04XyNLRHRFogZWew8YV7aynszEs9FO1sq
a+jWfUONKR39RTecgKbZUGK9Gdf4M1x4F7TkMa32hgJqC4zGUtpT9HczQUXfhJox
1aINiNvYiF8SOpr70ZRry8+/PmVVZophzalYWjFzWdMSp1xHPGldHPONoTuK3qYY
xnqiV9DavQl2XIb+G0j/ibSoKH40JwYXhtku9wzEtwZ3Ty0Wzpfkq3vKOZLo53T9
oQELU0rqKsEKRGJKt90xg9NB6t15E8eXPw343pNrDCRTQH0z98vbqkoIrgnCUOOg
p0PkqT0nzP23KtDghUNUIp7yxFI+WFkJxdrkFzgARv9HDTz7apmBj+2mn0gsg5Ne
BWwCTmKZ+xjyIQDbtJjhHAU+9a1iM6jbelamLPOH7M7z9JZSEsIBs8OSnYNURWB/
0FoAOhbEXWnrHbO1UH36kOYUw3t53HYyzdktzMPYEcWTxUtuq/vLZqKQQtcQizqv
Mi+E4RB2Wga0j9Jmsw27tplpy+1NBM9dfMLayacr+8VPTbNeUT2qdz4J3iPRSQLb
4zLqJdhi5IZcKBwroeByRHSyB82P7dY/8Wz0ercq1effICuSR5J0vOLmG5qbpaXf
WeZKQPwH9QDsHccjV49G5o8rA7QEMP4APGUfoQ3/Htn2HcBw16F5yjUAt7LHqdIU
slmk6i1taWLeTV1oArBAe97GEIyeS0UOwXmz2xv/8w3gbYF4MtMqxpVMc+CErTuK
yHF970oQSMQm2CzzaGW+EBX9AdUzyHFN05o9sXHcOobip5msjh4zgrbIH/2u4nwi
CWsmnyR6o5capnDiOnp5ByDlhbJzzsYrub8jtd93XWPY8n8UiG6Eogvp6eN1fYPN
owHHfASmpDeplQh680C2WbKBb0QGwwjA02fxCn4EqSqu2ZPgkTUMbaIrFN7th79E
6EKfpEHiXN8Rq5n0QmFePTnTCO0csXmvGEtgytLiAod3wOmDU5Kpsoy4NnbuIex/
VHxJP6Z8fZ4K+VvrxLV/VB8j+PNOG0GK20iZcIYrYt6Ra7tqbKO+4nHN2rzOd9LM
k1IOfe+AvzBxl5JZFoT0R+OEJYnsZFvJ9mT2GAGm7XpLqmCH0nQeIc1iHR5u6/2z
6moDCBTq5qbai84mqvTaUfRGQb3FFuSTyNmapXisCFQuZwAGFwcxqveDnXrkxME2
vtLuqNcW6SzEaVdsWcOzO9tuK9BiTeZYjIkDfjZk83uSpFV/R1CzM88T6ByaU4hy
4flTmzBtkY5tinUzijkECQk8e63M2g8lzRIveo8TGxzvhncRl84XK6KmOtjN1JUT
5sXqkDNfOmm97MtDGyJ6bnrtJX4+TCky63bU5xtCczlX1Dv8viohitoIx5uoYJTv
aMeCNogXyOdjuq4CBEGFhkqvJTOC3t9Na4UedNjVZWhk60GrSCQD5mfyl+5qtSjn
fW9ZN1D6EwaZp467qpy06N3dA9vMMCecT6+0A6k0rKfQfoAfMkq16IZvjVZTvpdC
99jFUpucXVUI9kt7QLbqlBI7FcPlOrXjkovGKgmIrLX2YNJWQgYHrgm2z83A2DJD
5Ra/dXIl4POGTqts91ellCibdUKdQCHEukPY8FV09/jArHqKBEUOeEDEJ+VvGMZI
N2OZ720iPV0wEx2DUfQmdC1JEJ4qb6A2EnmM09nb/3zoNEJ73CCsUTn8qMXAM+3D
rNqfdun7+7d0XoFzT41oQlRzX1kHTfTn4J1T1TbTRXrvDnO6vZJqbZ3cVE6rD07C
+0FPz0N1kewfKg4LoOmXiuIW1eD0MiqLmu9BuwQvwEJU/UDUCC9o+hHBwCPOpAHw
/l/Oidqzpcx8rsRK/gydbsVGi9HsAV+FJ9Gm3pjUYThfLh38OARWPOsK9UK1OO5+
H8fKrjb9Kr4ZenykjexKx+TPgUoAvOCTP/4um+jOsFG+Ui32p6DQoAhYlvqYCTbI
5bik0SFDxCu3mfezwlzyeNsD8n22f2wmbSEBG1jvsn4Fc2puXDq7gct6TGXI++zy
0yRwTW5aalOWzEZM0lHsnsbxLmOnh1MR0CMnHzKW7rpCsoXdYRzBr+BdoZGfKjaE
F3liwmkmnZrG1K4x6xFmS9PuCjbM+95+BmgneCbQYgd/L5Xf3LN67rOyFgVoMxcw
c+wWqkLv9Br1DwoTmb70T6wlEIDCNet5OvP1KOiWn7N/6ezAX+a1DN0Ni/NmOZkH
VVjRGhCS0NNhab1fsSlIh/7Ye9hprfx/Y+x8ad1blT32WCUudNDA+AfpplZJmoxs
9EmOhdx/+sjMhZF2uH8hbxthcF5EsJFR26NIJTosePiuboVgSvsMN2dwO+CYuBNP
mgyNNX8LLO8fyp4RVlY+uRYJ3YUaJGMOh2hBnf8jKN5EoZmjVCrHB5uFrc+UmdzM
Sofzq+GILaoOEbNdDhS1/JFMnkLutFjxAJWPRTNOTuz0yalZCkHEFYaZ/d4Jr582
vHb67M1IzZlmjSwhA4lW0J2/L4JzQekmuMzeT0OuSvgNYRPDVrYGTJ3tzab8a/hv
YfK8qlY8+BqCwja5bWs+pSqYd3kLWOp2BVYerzR52+YxtkVxz7AT7MY1i8fBoDW/
TRiqdFZzV7MzOG1uC59nxfZKwYRFj9SqicnluR58zn2KmuiLj13HgXhEPwLFwQgp
iKdUyrbJ5XEEBgK8ELDhGTgMj4/dWN2jK7K9hL4ep//Ah9eU4tC/itaJr+XRGFq0
ZcG1dqAsPsYmaYFFmY1vZ49oWxlep2m6vJuHkkf2sRId1NUuhmKukqfHmmgOjUzZ
8AurScOngWOaowA3k3mfMxscFSGC7L9qxQWIKQ5FOjSI0tNw0Wp0jBnbyVStlO9w
zbc5LQy6uNguGIwnJHxj1JLkvxozJsq8y/NJ30G45DbD1ZzLHhQcm9PFyw+lqjgu
H4yZBaHShqOOYP/utOD4oE2SRnk1/muHCPUwTjqbYi/WTygNUb3Q7d7HiJA+fZVk
63HDHQqxqnu1B9I6REn2aXaFU4iYWrBHiWBJUFmMS0RDG/lfqveBSPl1IXtZw8G7
9WhUZLZCDaxlGi4wz4/B4xhhXndrwYTf7BBFnL5u5TpF/pQZtZ1UVwUwUrlyRskq
nsYr0i0PmqVDP682Tp1tGJp08qH8ZtDcEmQNZCHNYK/YU6cPH61v14nsCjRrcWcw
iVIKKOwwa+By9yqwXbpiCvimZOSJGILJTQLrDKpr25LS53sRNdVpauDrN6h036ob
Ww9uvSg2E54scTLnhM0dpZDTPVfTONy9ssOjGOHASxv77QyhVWYNCXAqcIHW7cTS
jV1yvXjwrKN2rbdBP0g1YsjkFTWwlrddWoVb1Z14cympLQhrGs+gXMrxgYshvmYy
mZz6ecKikcX9u0wwzWjqBDLQ6+VPipuLo6KrQkrwxWdUozo/uE0Ym84t2M32jL+J
Hyesq0SE6Tdcl+XF5VsiQWgqDxPCy2JZz5TQkKhde4fUi8tecQjunqYln28Sip4n
pAUmDJDzhVC1owbU2l/eYloWOeAMODL47fNm8gOiNMIeoGXxECm3Ku/Hm95zVSGW
W4hCBFGcFPkdbBO2cgur40SpFu8ps2QvRUuqsWrMUamlDOyFmIMgjYIyaLOsbhaM
Zu4DHHpnEOj00OH5lzX8bguSzLwO9TnHh+ZeMJ+cR/IdCjh1VNQT/l60d4mME4XI
IViCXR0o5+Ek5WkNUywNsAhdgevgnfahmnixfgixUCCjDtpw0j1/Mnnt8dR2zlWF
UH/js1cF3bseU6jLBEnxPUTLlpfU9YddG3EvC1/St6EOxyFIdCvStFF/51sGuAtW
r2XfQN3Q0mxsI0XWEQ6PG8tyICs7+4wCo9lX6dim8PnucJd6pW+J2p2pVJQd2yVi
EN9Wq9Akhaf/knC5a5RRDYwDTm68jxpp+Y+Z0w/7U97NTqIQSU3zr5qvzzoC0vwA
DXpvF+YOGUsXKmOPHi1XVB7uzTEZNsGB+r2N92ADcH6mJAY1tR6uVAlcSMygXF/D
OYU9uVZNjtGJjf01F9xsmJT9eH3DxyMNP0KER1xeN5JGCQdjkRAOhY93cfxqUj/j
eA6JoD5f4CUo6yjFvz68vl7PzfVZ2IIrykWv6O7TwpbLt9t1ZI6aFjLsBBiUw9Gy
BeU1r2ButO++I1sPqIobv0B/0RxqwJwUlrKlmVKv61xWyW8xbW1ucUMLT8xeb/Q2
JP85rZyyp60X0HTL8QEJoDdPXl8eVPK1c2tkNlaUbvXhvgzKyVrG6UVNaQQBGG9v
TRwgkB1oPgjnn4mw+KgdTyqJNPR0PJukBkTY0TD4SxkNN56+YaN66YQZLBiMUDft
PBafziUI23qyEpLYqajfLjhjYApeQEHxUSLYdHwKO3eM1jg5v61ZPoxhjwrITYa1
sRJLPeN2p4ue4yTSAUl2uGgqGT4uv5BdNtwc18mXrxczgc3XomvwQ+sBpLsIc6Kv
RNQUGwJTLdNJ3WitlHgFXnV8DA3mxr3KW9PexPwohagJoZIKn3DnZBZXPQ1OdTiS
4xNar8JmNGJBS2Yk0fJTtDnZWQjaMV6hxC8xSfdtm1Ef0nwF59LprpD2q5GG3Yci
7GIIjGVT2TbIuYqaagZ4n/GPGFgzsz6T9Ld21X6797mZ4frUxlE5Z0B0e6J5ScPV
1+MgbjoiDidS9FhVy+PjCWtDjPaUfaCCOdChHNLDRuNdg3SMqb15e/2F2kG35jM5
lMesqUjPeNY6lfGXuF8Msnrq0NpMPKozAG+tIbLo3GhY0+u6lmxrxlpDg6IwsAYm
6k/BKTpvoCeARKSfWzO2GvH/wdZTO2g6fAinX2vX91ne3Wrv4BzVhLCaonXe7eCI
zR6zBIcVWUN1FFPQCq5hIrBgv36DvMeeBpvZXu0w5PrScykuSKM9kOoa31XQVbGQ
DpsyZtR5sB3S8ATQPKvk6/kxcbedGYf7tVDZEYyPqFvlLmMbR00SJREn633807bt
yHGcDndOImAymhNLg2IaFfNVBNJa96GAx5+jpmpVJ4zFyLZ0TgZEmSQ/t6DPJdUA
guzA1gtA+vvOkr+eOz7L9FfT7qweqsQkQGfZPjVohFaemwT+Gua6YSO34EEZEwRq
GzidRNnC8+VqPa3SMDSz3+4ceLx5CEg69dhWuJSt7yEiYsGiW8FsSROgMNDaLptL
vFa3ehnU0kXlDL7wL107wMG87pyFbmtqO/x70PkNjU958Q4NOKYxpL0JCWeEPYZW
AbG1P+jNxWNvidO8b3t81bJ7cTIIHszuCnLDZJF9QTnvjlKFCFCajFuOfywmGKmM
6pmB82rY/8q/UEhTe56Z4Iun/FPluqlJg8q83pIDLtKWvuByVRdhMpxp99WxmpAw
m/GseZCovu2FJ/jsOejSXUnKrAExZv6NERpUjTQCeNr0eZoFZmA99Wiex8gK1ERW
RGR2P+FiOJHDpln/wUOaq4N+qEolQ08Y9uQpstc86ruu7KGJODpEHjoYHZvHlTJT
5/HiHu0e5kjRdVLDqQL+4xXXP3Fy9Gdu9hSTzZn2JEyyKbGU+0UX+Zj2HMXfh5Dw
DOUoEGIXWW2Zo7YU5fVdX80jw6+0MO/QD52ZgRcLSnTifBjnUmlUhzQhCXLjxx8d
EIo5hSb0d1vGfQHbK+5YXAzn2iKaFE0Ykz3bwlIrmbqL36YT52JOdX7EHLEBc3wd
LPH8eonPNbZj3zljRJcPf3d4zL6ELQm7DNOEHmblUEk9PrQGHmFBKP2Nbw+7epyv
eLZF0FfVNO+QjU2wEf/vjodrqL9Kbb5Zd0HFjn8eOYi9EsuSEwf31RPgcjc5goja
Pid9MAI2g8I8Xp6dCHDxSiKYbOEWkM/NjfR7mRKOk8OruNH2mwYd5NUD04TOw3Iv
aXSA3Wr+CGkR80Vxk5dN+6XZU+aFtl2bdMrS4lV52U/RKexBOSS0nbjbjO+qJO83
XOw33446eVFXEfDGhmjaRxJNqq6lo8lw5MCrIqJElG9emwBHFp3oR9LYFNc8jv5k
ni/KQlh6YnsYyHy1xnOKpepa9t3/r2rT0NiJ+UV5cGeHWjlFu2UhA0Yrsnp4vnPq
WUqj0nlzBMow50gvIEW3mP3i14Q+1k473uroqzowaLqvZFBRsLqEghrR3lOxE3kU
jppp0kZjtlJhm1SBHbbtQi9hy8V5YL4D5ENWo2Evyte3/OJ+Q6QcRcwMZLVgYylG
WxKs4MhzoeJlxd6NFwd+DC1tcS7U4JU4rUjK+uVilEvMcfvXhRsWCb5l6INesScM
QYbNGZpeOMSklkQjd9yjgyZwVZXnoeO3M+2Ca7JSmferuqt/1aVtFDa0wj0zs+SK
OVj5vf9VAg4xlP3IOl3KalCLpYgPULZqfcF8bChQHbsW1AKymxGGLBd4tZmphodS
UHulKOd41bTtUJsD2Xo0V44m+tFUgLl7VBCz0sO2hK8y3O6FHi9qY5v1I642phQT
bKbL09ij6fyhw+3nZeB21sYqE0LXYIfp1atmzjmAz/rcK4EwzDRg4VLKVNVtaoZ8
4i+kyEe51hBig75TxhmJ73FaQx9BppEnj3jBmwAklBJJI+QLnqNFs/nsGRfGzWYP
g445v9YvgXMT6JsHur9qPYE9rn9WOcVLapRdkVVyTmABGh4GLRSRc7t/zomEryew
f/8nIBE7c/GZUoOYKssOD73rDlLbgqCciei6wLDK4UBM2SXUSXwTDEympa52HmZq
eU2JB7xfwiTyPIw0O6Jw8sKV8GcNpHfWj5fk8li0KzkbfiaI4Ct4LIK16fBjvxHk
H+HxptVC6/Tj0rOBKdS9HHupcNBuGFaZqQW/ADO+Iu1R3aFlLMAYfg6JZNZ8DyBz
S5kONo4Xz06wdy5bGXe7khlMUQ98EGf+sGiz6tdz8cLoGb786A6u8H0lLkA4r9iG
rYzW9Wv3LsUPcdPbYwL/m4ZYedqivsaDXG2ZVj2m4hxjkEdZPR9CDwLXIfSH4ZOk
cIwtLD/5tY8ObE3P7GpP+MVbkhIPE9l/0U8Ko2xP/Bikf7NgkzTJUqOkMOfhlkUz
HdzuqFCPTCyuIM9bAGZgBoc4+R5CWRDzAqfa+G4vZmui0puS2SuhRB6+uiXSNDfE
95qrHnF4FHlXN5s+6btxHMF82+fYsbHvc9htM5T6x2OqXyCDxE2KlljN3voai9pG
qUkIDP6r0M5ZhWnEV+geMpgaG3xgs6dzNcc9Opcqsb9kz/lVzqSWs7Hkpb9SGtsX
k/Y3CzJopm089TZBiKbp08Ow+CtW1NpKd00wSHIJ21mjysVP48iOyQFaxc2gkjZJ
flpE7oA87J2LRrD6VXPyCsvglo0ruWzL6XlKojzs9WPEFJJn8TMqDYQ6VpuU5F7T
XBPrRU1KpW0cnXgfe1ERrj9PPpgpd7S0VXm7Ym8x25bufFO8Y5/jFlUrKXSvzoor
bgOywiV5JlKATDs2EBgseNBkAItOYTIB6/sIUOetysjUC8EJkClOQ3zp/uDcFHZ3
OrP1wdTGl9pD/uMr5v3Nk3X5B7JgnA6JPeNiOCoHGOBL8Fx/L87iZuOScnYtR9bH
JinGCyD3FVM/BesbHMhRH32NFWLLDMQ0SlrzNKzE6piyyUdHPyq1fi23TSF2ZZtQ
N1uckXTPsPtByLfdauDD1uhM6CUCCxMbtOW5zKpKiQZhjvBjYPPFweXoZpgcLDiu
o5rKXrvSHEfX7dr4k83PUapoqVokDP7f03EnmRvr9BZ0ucv+TrZunyHaah0TT2A2
iMy2eCZDVcoqi1bxYKBXRW2rEj7N2oOqq06TvszQ2FBTmXUHgou1uknwj1z1q8e7
js7dhHv623McG/YuXQe8FTeyECqd2I5V4HkueDIjdRIqwJbhrlI2mdc5jzY2wUyW
ilA4n7+EztwkjZt7BLq15VUSrez8e8P5vMeJzTeKNpO0XY9lVSH7PAtOVdadWf8x
wpwmGeCYgZFQfz6EApeMa1RzW86U5BnfkbBbBa1UemNZuqdihbcv2HHrlzTkWJTB
/zV6KZooDFIyfmhvdwcW6zivPTftAMnoYtZJ6I/KHO5qy6hK9FLTua+C+OCDHgCC
uysQ6koGo6XbYws9ZWcl4cxROfzkTunVRLeMzS3Fbzc8sdmyy4l3mloKL+NWOoO5
R0uZi0nw/Zz9gwopER90x9BDOKSWSaJvnwOMYzLYWqiTCzcsg+nQGWM2vp4H1DNn
VyzL+E1cHmjf7wC3GnKMhG5YCzlBbAXbMD2sHBCSD7iLJYevgy0qpLyaxVo5aZjC
nAOz1fYJYPUGfqaaieNfquInc+WWf6IL+ljE3Xr5RqqPk3A1WFcVn6xSovz8tDml
PZLisoFapsSrIDBhYG1nHNkeuJhTTe3/+b7kKH6fvChH/PYsy5sX5E5OYNeiS9oL
Q2Q4I0mY5Q2b+P4JrxeCLayexylX9x01uEQyQ8xM13LHkkSTm7WWvLhovbv9i2Wy
hmzHRy9vyM+It2+DDq8n2jzUfDf07gRE3kTXf3F1qoXZuPNAuQQwf8MsWgC2Q2Y/
wqXTIzXJiiUfDpp+0PhDEhjVVdREf5fs/7o0BSEwTD5L0LZxb4yzsJ1XTHN11Sxd
rnBoTWeEV3dwwWN+CBCvog5t/QbBaqV5Gc162XpJEKdwbQxIRQte6ptsOKoBAtHb
lEm5wWkwpNsgp+vj2mPtVNbZJofO5POPoi8DtuM+OhtDWo5fEtHtoLgJu2EGWfFI
lnghrmay+98/irtPftBdSR3t+XXc7xzUTT39UXK1LSUrSAN1NLe5+ofXNBm+7Joa
DbFCRbAN6HEKHKjdOSPKIHZua1+SIuSBwrNNQTm7XgPgfr11upDyo21/eBCqNu7l
TFHnTXcHanl1ZfP2Ag1rYi3ZJtlAfGmkfWr5av+Nkc5JabpmM3Ygq9MbreydIv9g
pjDu2yiAqhdqBSEgqivHUJMha96tJ3s65b60LkFBQVMGJdWCst8OPD1ycYnuztcK
7Nz2eLmm0W/l9eHfBKtKzWX5HZv+FsHXCLqUi0IJ7Lg5iN6ezUIecFKyKBcaZwj/
amRIhppc7PRXWzxgbiWMeXF9beafSp9AJ0hWjkDXnj/xScD2ARpjTJOqixor722k
cv4al/DrGTmIwFVtThcoXer1kznbGbOL+SiV1dBhq1wjzDEuFmZJEbwOdB8n/A5a
9X8o/FCP6OdzVn78LG1NlVqcKQaB00iHzXdCa1X+ZLFQHco41b/854PYEFXufxOf
lNHBMzkcX5mNYYkZkwLu7tALnbk2wvRrCNLDZUetJzBm8uiHfguPZQzegEmiAYBM
tWZBmkw30HLlnhGR1qxsc1hj0zCv8K2/T2wWoRZmNFe+1XuyxTTs1hfjUOjhy9n/
cNW4BI9D/cU+jK1VjTnRXeXwdF7Abk1c/O3aESoDJRwKMOvc2sZNkDC0JzIDwEoT
LP+dQrDPMDtI8w3e81CqGHr/rS3SmMFaMU3Efjt9x6iR3cblRqVCoibdnEVkfya6
XxN5MqRXHLq8asC5wDqaAjl2RtFx4P1XfYsSb8nhyEx/Q+oecEnJ8Nu3HL0yV4HL
c1tGf7mzHtxtkBniTAG533MbHDD13qB0ZFOcBRNkUnw831h4XQaqOIO0kFLvh+XG
uzOyJ0GmgP1fpvzKnE21Dfv6M6hh+SSWpaNhfQy49BhkwnYzozHzVlw/vNsikewf
NSYEWJqyHmxyWCgr+/AnWCqGFxE47K737/t6RUGRkDttRdArPbzzMUELJaHjT1jX
7pMC7Ch53f/IUYfcwa1LXYtRKXCxSs2ZiAD9/9bHJgeZwU7hAjA2egFEn+GGMbHY
DjAL8iwlCcyT0RDqa/6+d+P0EYL9uE1gXrMOulFeA1cs2KMFQQXXQaQ2MjIo8gKz
PjhnQQKKrros8xzgi/ufYCpO81HewxVi773l7oVQe0AeI54KRp8ikg2kKdbiCAiZ
tde6CHN42hd2zKXso14CAeA+DfBwu96MO5R9sJn73TzColNN2OUqZM1+YlNnwUe5
3rtETHA7sLdsjB3Czn+iODjz0MD1s2nCJkbOmKgV3qwel4ien5s2Vpkl+RvYW9Oh
408Lf9y733b45eIMypVDkFYwGTshDPZpjt5jikvaX/+s/K4RA4kKtEkfiPt152zT
fyy4K1/bVoZzPCPMGjJArg/2lp0hF9K0879mPUYLU8B75NtJ4uBXDRFuHKKNYEil
7te4Rd9fH5n7Dc8Df7fyAaQgu0UFHnbDotljreOrFfvhWn+QDlMMenFc1vNj7FDC
keV43Yvk6dXIclIXQGG2SqtJOwNPbpjAfWUR8MaCcxm0v+YEQ6lCG9n2vL/BNMIj
oBY3Dk1haJ1v1clAdS2b1qWG1SwpNKe0CqCh3F0bM29DaML1fQbQTG1bnY05w8bR
fc6d0tJZc2M6u2APXAWu2n/tEskEU+vFK8ImeCPxvhvA9EKqnS153DAYLBooysTU
O+LvsDPTXUf+yg503gUhud4SwiKygvxHsu+4zMk5OqTry2GtZCbPHMrc0dWdoqIB
JRvUzF5V8dxqrj3+Up4pfC4qM7M8kaoOU5lsvsQRg9YgOoF2qBAvGLke+7pebspk
ccfyJsWNSO6c87ANXB2EucX33yG9BUuBt3NMe9ra7GutCNpOUHF6O6cRmgTmnWE3
IGuWtY/WWxpU77y6Ye5HyGREGSykNMIX9UDpLSMxLYFLvvWBmQ54IReA6jNPokk7
0KW7Qp1s/3jowWzU7knuoYptANAxz9BDlCDCirAp6hP6dZz/4ENh2VL5LtnrGXQm
QLcx6GJL2GBeF9qq3M4Y5bZAV9IF7M320ivo0hm7MqdRvW8eV9Fg2s5+QFNN5vtV
jnLvl/gXr0H06BpSZfvSLHjyC7NholxIg7Qi/YL6U71BNEpd7R8zAf2PNb0pjoS3
o+yAaOQ2DdI+Z7kFmkbT/3v5YQC6eXCBDJOrDf8g31l99GAWnjLYKY+DGnIM8I2t
Z+UC84J/9wu6mvto3KZuFcetIkIh5z39HVto45t5UqgLw++6xAT/uULX6VF70qyt
lR9q1FOdnH2ZkmIts9+l4N806+Ws0l7g7Yqks8siOYdHwWIdQZQBiTdEV6GmH2f9
Gj04Ci5sN3bpXG+pxvET3RUT1oV6vWk+qLUVUIvQoZugTqzUL2xsYtlDrJX+pgY4
A59eH8P3UMEu5EErw2vRPn+ajgsQfSGv2doLi9N0cb77+/hx6ov8G6gfHgoP5XRS
sxjGx42wuht5U88V1gzyx6b6Azlzo0hQdtkpZjqUD12n+8Uo3x3rzFedDyr146IX
7QaxLpDCIxsGIDqi6DWFxE8uBOomWRNxAFqoBC/AciW+Nxsi/+ZY5nIVssXUuXWM
vxOdnykuhgMf7YRhBN8fMp0aZu1Kh5peIcEB//lxHjUXTeQWFcZDw1F/eo5gYQ58
zpF+pH/+xO47EaIDDxAW/8fRDqBNmI7EEldq70dsSXeIagR0sf+9VfbBADkBxZgT
tmWYssg08cCRS7+GagM3b0mREEbSeRlW5uTRM8dzLRJhDtZkmK/9OOE/fky61GbD
BEnV5XGij3wBBv9AcyGBIa7SCmz+ewhnt7K0Tv6t6PJv3ZPfxNlA5DlIT2v8QSkb
7WGDwoGFDIBHXKWa9GHuXnClhbotx+81Zxc/QTr7mulcTOdn92sBnDF+9y1MFFvl
Lun9qdDZ8UI5Co1VSrYx4IH9zlCN10fQm2rsVk1EGDS5q6KHoPH0DkoamuWDTXGi
z9fLggr/HfCwH1+1D8IVZ1UcosCv4M8cBwV4LfsFBJtkVmKf+IRHfig6en4FKCmI
4QooQAfols8aLU24bPMXk01wx++VkM/b7QmjNlO+yJibZ6bGKAij20NIv7pzIa9o
99zJhBda5n0XgseTfLerzy/jpu/FLJMnhXJMCUvaTByLm+x+n5dNBZp2KiJMuKQm
lPZNDqLH4h1hCBHs3A4aqZ7laruvOJvHFr/MPHqUg0oo55oPm3pm+NHIiMqMAQ/e
GFqTUDBArt8P7+1yNBQe0HE3V0a8CoZcCTURknL8li5za7/ea8CjQUOBBJsn6kOy
QcGcvOpHUxNCOp/tWGzVOhCDS6M63y47pfGRhGh3BFF//P1+lKuZneK1BPf0uqwM
h8c6lUPkKMH8K/vJsJGpuii76FTn+eNEZmGhC4wWuRQHxOgwHSYQTED06ZytkQi7
RosXfDWiOpD8GykGBz+pApg6wpl995k4cv05KMFtJwOUYQ6xDhCxmYVjmb/2Dld0
ua3SR3bvMapagJYOggr7DecoFwwFBZ4IlW05rVYDIZSrU3fyDcioEfSfgwsiNuDC
H0kdXxQooA2inJzlpcdvXLOVeO4YsWut8RTSpSXQEz2xk2X0/oSw7eAv+vLlErEf
pECvtmTh4sKsE09BV2chEnLlwUa11I9X/szpZowMgEf7F/vucI1fu1OxDyNTnBGq
i03dltgoqA4+lsKk2cBi/Xf85e4YX+4YS4QMBkbYv16x5gocWV964XB/ndSrHhAT
auSXZ7jKifS8swdkklT3HbdcOAy1m/6iHzTbZNajxx60TgtitHsvz3ASidP0vgEk
rVj9DT2QVuLf9rzizPjhg5JEJ17M47xu05ZiCMCSkqIrSQHLmeHhtlyGk0HtdblR
nMP/dpxRMsnO/UEG+G8JBRuf4S2vwu0DMI3U85nWQmY1OSc+qqBQIHABg//FHgeT
I7cBKV9arPWU6JZmVrLHhKZdQzvDOdZYD7rNnxYr9NLB5Zdh1lYjMnseNqVK5hS2
zOJAeXbcl4iKOVKZbUxy6HCVc0Y927iS20gOylFqxATjIcod/BpPiY1GBDDGDokg
grPRyXHTmPxSBAmszGdp6VRIQsVJFP3XoVuTQQcN9pgFvnxt+4CI1VxToM661Wdg
4BZq3OweQERZ/m3DXeoGDTMDkYLnro7VABd5TrJdlsE1LdD2octY1LkkUh1OaU9S
WmdMKafKFkEvuPZ5pMd0lqPXnm5lRrzHR3I+KNn3tt9jIrpZZpJDbrQPbBk+Rg35
jvMv/MIQRGKKySI5Sc/4CvwrBcJpG1H5Ls2LHtL37cKCe0Js4hkbksjyN45J6bCe
jmzepS1kJIojWFD6b0rWTP0CHa3ay/KWVcabFuKqjQP11ppigJ1Ym8SJNr53/ex8
84D89Ytubzu443INFEDiyXHZJ5qQag0u5Ha55Mpwymek3qKVmkbvbQES4BTnkcdX
AC4/3vKCoqk2NQkq7zT9oGft7I7Ivm3dXKWLgvaPXGbz1dQ4tm3fH3nVczincKWZ
ygATNd/Wn8wE4RMLaZ25mdKBzB8KsbnP0q99wa/Jtks6Zm/X8UQEPWzbpaTHGlSU
WHUfzZlvGEXziqjplGrGGk982Un1kkXBZoOcbh9wX2zQsnsAW2vYEI2s8cjc0r0r
BtGFiwC1qVlKhCkY6sxOweLeQPeWRsqakn4WP+JvSFLSzi9/dJMow7RilAFnWBC0
fYqZWoSz+ykT350ypDtP4Y5GzbUK2ygOGWYH1PkOxG1Lng54irPuOvrIRhpCrl7J
DajDcWWxX4UplVB4Ng0pjyLKfrVkYWX6JSoropvW3oWAymwhLcmkTVEnxQUVucmX
g7ffHc/JFJfTz8ltrEhR8iO4p2834pV9fOqC4N5Oq4Jd2tWjiGQ7PXT8iPNFaDzv
eAVkq0FgNgXJk7b5U6idHUxF/khHX/OB1GCxZL6wIjPPNI9Ay7GmDHzV6yFQG3Rh
E4SlDdc2zkHY6L0MqSgN09MNzoyiPrOQUZvBB2ibDu+zS8LUJvW9XWxPRf7dOj49
MD+gR5k3a2glmvzNH8YDIJxPNDFaUTXY/ItrLdDxy/NcZ2T+aVGj4gWdodeSxZRT
mpzTFYSta2c/gHNs24l/lj1WpEF+OCaC4PnJmFa1k4rgHnksBlxvN5L19hnLp5xt
3IBJirtJDNoJMWoZVl4HlpbXHFJDJqOq251PCf32HYPvwTepjwDuB6HwYNDS2ASX
mVIOkTfUjCHSMuY7CCtpkjnp7nq50N+wmvQGTp3QLGhr/f3Z72getVQaIsFZJ5SJ
wCDDRfyIE857MJVM2ekBknVhgBn6ipbq7047v2toC0NzKuHuIZfukCSLiSnP0Ysn
hDvIX0rwOngrxl41UCok5TRAZUJDwTJp+PtjyuSIA5MgGS19+3tj88NSysnSritq
oJ45i2WWz81e1dOrhx+XcynWC/ZjqUlkiPsmlC3JBZYP1hOkwhPDXgGNYPge2POY
V87+Kubbgtw388616b8uLwkbLEhVKVHIGe6vzJ/JpC3qepjf88s7PYABZBOTbeGR
afI6o7gBJPYSZGhiXZxWg9BNOvcatMAb5AST7QkomtKOhu9K8QhbvYodE2dq99SV
6KWfKAs9S4PCKpDOCRrxuUtxSogCfFt+QvyPWe6EmMvkeKOsgmn3bgBtCrF9T205
hmvZF58h3hks8IbXylqse7nSUSnGrUwnh+IISY50f929VUiGqoq19r22nHFNUxdl
fMyluyaNNPC1KVwpeKxKV38rraxgrP5K0y/jTim8MtORSkN4HPntZyEmZVcofMzW
nPXVOpJM6E6p3LHk4Ch+iH2U5tVaO7mVyxo3KKsiRciNVsC1jnwruIh+iDrOmotn
qi0nz9ZtwLwouRuX4rVfjeAVKwVYga3C0CBQgpUHpG7M1hecS+UrFaCsw8GwpPv+
Z1PFe/AkIAKU2SGdfSL8Q7FstOEwDLWtsTJ/hYF8HYn5KmhevKwEtpTQUemAOlsr
swr1DJkULTzk9i77DHRVlUyUdEumOv26NrEck6tjnsRq/Fzv7Lu3pMZkaucEPlxH
B0TBalsEzwZ89aBRbPdm7rkjm8HJgHYl1lGDkpQnJhObUo4ctzpDaqstSBiAZlXT
zJzCCQQE9fdiLxLgJtaqkD3Kcg55KoB8PoQOJn/nrpiyYbvERd0GUqJBuEvEf7KF
Mq/ipTjVrJ12RAjVqYojhCjlKzMbl0dniRzYJyLCiNU26YmqTGKRFFRKVRXiCEZi
GkHQi7VYc45RWxrow62gHQoRC19Wk8ECJMelYO2xhv/5yG9/bKA1Aa/LCvCVKsJw
D24bhBL7O/sxKmH16vAr6N2w2ZXZrYsn6gWRvAkUD+a1AjbvNxFjJGaxdE+lwwFj
RFlAhf+si9Tn572mnV8duwwhqGOmK8DiAJyCDGttvbLDbxhWYRPDi96iknextPCM
jcyUJnzDexjmwXQqcUnYMB+swUJcgKxyCpNY/W5pIiiind0ZId1zeTljdgi+9gZq
MD6EUya7u7qGEUjZOncVMt6PxRegaKei5T/rF4QUs9e3xeCNGNszsaXbvvdoO7FP
kW5u/YeIVdC9pM84yrhm2+t5pwEvBGYwrEr9VChFSx5xT62QWvqbDYLm75sAdeA3
EU6L/S2Tozw44fuZ7poMhYjIH22g5O5xC4TYU00/m9Y17Enx6ZnCX0UXCUPVrDd7
ottLD6nTddWvE/GO5iW0MQm2IP5lndaG1AH+xM820BnB4VkbLYodvH07G9vx/h4Z
bumSai6wXhOKsqjBOdO8xjDMknwHgFp300+qduSfJATjDPsit0qFUp20jWydDp3e
zjCUo+t0Lnumu5heieyfJjQikxiQSSdbENoEHSqJuNQGop0/Cjae0xQ2roOngIsX
U3rtL6EqdGddHT1SG+DfL1pyFgDt6YouHE6RDS3fOJ7tZwZV2TQckZ7d7O94UyYW
+/K5zohHlUOIqe45zYQojzlpkzKXaAEzaP0em3gHjpqQMO+6MCbvbk6yLzw+B077
UBTLxsBqIJfeoDi5OvUcrMjcpykCPwchrIHwunB2v81O9EGt6oUhJoZ6LJRmmK8s
4wbiTZmi7GFl4fcvsJXUG7GMqNnT3Z3lw2zplzdgxIVaHAwkrV7Z87r0fIh4129N
Y7gXW3+skxMMnZq7OZbaVy04n1S6HzgCNw2I9aURDWKlWyXdacj7aeLflkBG0dUU
nubGu/vRE/pO5TAUlC9k+1XQvQBFmkE2KJZ2qhmJAfomrNaZCwKnuBy7hpxiKk2z
E42OerHaJlw8SR1oa9FONA1pBckQJxVbo9JLWKS0bfZJXEvDAGQwzg2k/Q6DT6SV
5vtZCQ3TyKaAW6qTfZeCaT+sJajFV6Y1XgtHIN2HqA1JSFYLmlr2j4NedWjEzf6U
c7KkAPdCFKsAcFXHk4RG+283yPEe2B9KRtSH7MCXeou1Sa4dkLCQBeN8O17S2pQx
qLyCu6hmX3WeBeQ0OcbTtdzjrbcQpCffRyB+vz5za24k2Bijt1ThObIR4E2osV0E
uZviUoBwglkKXGu1K+cirYlw6oLnQvI2mXBejNc+6lNjkHPCikWyLv1gCVWE/ya4
r0ffiTWIOjXNGxGIMnhFroAyfeysSN+ZBViRpN+prOtpXByLLRkSAPMyIOuOhw27
+9Dl91G3rRNaSuTNNHjpb6fB7xUu3XI7p0csa64Tcb2YYMQg6fBZtNUpaeZ8jP8M
XGMfJEk16U3Oos6O1whJjr228p1DO1lpgckVkyRmxNE4lhXI2WQh8xNqo18JOWRy
qWdPlHfSbYGaowrKzVscMZLHD9t9ib4NQtEv8roDV9foz/io0SglCEgordV+/vNI
nq2fP2ju7gTnNIoxWgi9oxoRI31nJzGwBWUDm3PPZiVDF8eY7c6RDxubI/a4Rz0b
o/nyrBf+hNW/qfZ5JLnV/BgY2Av2V45FkCf1Ff640m/qQE9owBx9UlTQ1DsJjzZO
xCcvGV8QVSRcPclH390s8P4ueFZ3gG92AzqxGKNFG1rgPhtNEemUt5mH5zHFbG5p
XgdFllmAPiavblg1phiqccbbl2PeBBztyLi4OL2V445PviGiABitP0MpUkqKrrtv
LkSCFlikuUiNNktHy1DiNzMv7kx/DpXGlTyiIo1u4p9MGMZ1+Mlew+t/SZfjRziG
VNzK4GXCS6Cl056kAOkR03wjJYJFKJWxxE/pU4cpMfVV1l+YhC3N/qeHo6Iqt7Al
yRU/15QQl5gRSBYnZcTX9aob64qdGof6MGHj+9oI4NSzVb4k5cXy/0fI93Bi5+BZ
Y1X7XMLRF1ictrr234Bng+771eFmLnRZQkKhQjOJ28F6rbU1ovpPQAxY7NPX6zHT
ufwXLT7CF0F/FCH/s8UTMvzL1jHs4YKtdxnBKYBaVrPitDjkHR8QWou0hSaQt3CC
oZ+6EN4hiG7rjmxv1yDcqiCeAJdGh/pVmy6jQVgEPslCCIawZCAGtER//QgPyy/b
JMA9vmJTXSc3v8r3TSn53KBrAVe0QuBUsoJmKfUpGeQz6Id3tP3iPIOr0gPeMK5x
ZNdoHHItLZBY7cc+kkSDR9jPyY1roOZHwP3MbRevInnCf4U8xMtpC/HGDjH5a4kB
Wi1LjdyK8Xb1IU1dG50Q9Qs4qqkiDq2UJN/VKeENblZfU3xaU8RweNPwq2qIaevC
9EWbfxgjoTe6Fuuppdgc4zR1Fkje/5ZYv28qeRYor1s8qIWMvc3Ej77ypJ2W2lKH
2OGKSQgNKjEJv6DBWG/MAPntnXrMRbfnrg3zugdbrPr1rc/FNibDmRJ6X90DFChf
RPoEYHy6MjvDTJQiCRlLq+JONn7hDMYxNBvxtv3MiHft6R5UnoQsJ0n/PquAn7jv
es4Aojrr7WsX/sP1btQf0xqLW0UaZRGDt49IIS3gYKENP6jWD1h/mEh8eQCLWd49
VgeGivOIz8qLWw6XxpwOJdK6tvTVjE0WGvJLdZ7EdYQVfOxXn2z70Q+f78zAAIqQ
Es+vI9W4EPvaMgHIeQZ2anqLeMcjeGoycT3JoKpUwLWsNjz4bWh4NJjpIVKoEIk+
FkIg+o2mFAd22vywahwn/J8VqBugjLVwgcR48WyAs+MwlCKIwa+ggfPqwJOFiU4q
HngByS35rcxYxOsA6sk8mWtridR4DT49GDYGrswFYnJXKgngeJN73cUGhASVdwe0
ULLnOU+MhwJPvXTtXZPXD5PWBRrQbr6gM0bCFQ9AqF5qsjt2R7oYy41Ugd9Wwbrz
ENv+G3G6QHP8hJvMRgIlb2zOHGKd6GX2MobCXk60MCPvj9HxJ4WRSGs4DN4jmpYh
InpvFqVoQ+T+iqnszF+32897qOYUYkhPnjwVSHzy2p06AtPZkoxiald3uiTrKMyq
g33aPHLkNLzViVXHAxAykvI355ifoN2K/fLjFhbKTmwSri/jQHfM0EyW3Wd1Cg5B
PKR19x+3Gms0drD3ZgE6cdvvdiHbL9q8ToOJSWqsZ/rfV2E+7B3Y4AdOHv4NAq9T
LYEUrorjfHQ9gaLcPhyCvDtmmmoQu/mMgKdVHdwtzmLRTBKY90A6/b7AZfbSYniQ
AyFXPVOV5Xhr6GeVpDnLUFJQJRQ5NfqKFu0/oOdlP4cZAdmzjNdmvdrdzFDfoKp4
+fY1UNnLkWQQKkMH8YriAktmTyBV4dU6hvTlbKDUfBFBvAQKqU8QlRD5biLxKUcg
B2G8NUusE6h/QN+YRSxFKMVJMbFboP9/AQ3pl5JqAtJAM0xdSbE+KRBzPpzVHcem
A4SlEh7zg8LNk15mMi8LnRgkuNceueYfIj4wPjGbAEuOswJfRHFuvyHWkPrur2C1
tGMUgHpVRqqhoyNmpPaOYpn5Ahpst4ni5nZ+UNnPzBlclT5ne+7STH8XHr0+kiIL
WAzo0a+GPAuadb7hun1TfkB5smHjlkkrnRrqs44GDMhX8CABvdzpGWSil2oX6BrZ
5iADDUBJESjCoyEUtvLgW5+nojQYiH1M4LK1DWGbscfRZnp26u9JafEqt5SVuLv0
Pf/xf/m2Hl921j2WOkhd3qtuRzPTqHsaadoJ6VkPZ75SM2+R4EL+qy7hPSeGJcry
MDF6dUv4SIYJc+AONAx3FWQJrDIJT5jpbHYtOwKT4VTb60FcxeT6BGoUi23Pz3CJ
IjrHHre/TBB9LmCWgqZG6MVZc3AWF79ksGlV6YSZiYVz2y5OsdsnjSAc8E1SfK7I
2wrDdXuqFGtjVlyZzdUWXLFZlnE35Hg/S+CGjtz5P40HEbrJ+KpEKFDmkQerpBnF
nUiOXZlGCQRBxxANqaiY7K6m7wQ8NQrawRmJLaKJ7IKQMESCj5RDUwAICsgvrXKu
BqchznJO8WgGooNG1NA71kzzR/hylH+DSYm78OxCYd/Vq8BeqDU0Sn2B04zDw41Q
JBhrt1LIJODEKnhyiLjOvwpaURSWB9jbc08QDfUJisemHQRceMwqcKB4iRv0Db4X
QXQM3G2buj78jdAwfemXxd5HoF5trWvjv+d4FDE/oXiq6oATx7SoO63r28oRVUG6
QHSq2ZokBHh3f6EkfPxTqyaEg348XPnN/W0qDBPuz9TjZbEpp8coSHQNLTMcng3t
pPDwf04vYsZtYQm1n2ih7JHx/vNq2jxSmLwcGFeDL0Lgfz3jNBQpvlZ/T23SxylV
tVxC452np95OerAzZv6UkeBczZtNUnLFJBT97cuJo35g2Zx6WRuIJFvmYQM5Ypr3
2VeQbCrD/RBdiw2px+YAGEGn26tWJfl+K9Lp+3ScTx/YgPArT+5zqf8csROzg8E5
/TwLaXTyPMaBXVUeoXKR07y8mDFgtpP+vsBsuM4UfAU+lo4j24Cas0Enz9h80ygE
Ho1B5Ep4mfxeREfWuMXRpbxwo4TQ5YfZLaBxX4RT3gIrjRBLH9TPi1SmHofwFsI2
DRFiHfYN9qQ7oqhVLvmNHo7oTp8hN9leJnDUm95sce5SzcPvV8COssVRLbUbuZGh
kFzwbSMEGkXFB9t7BClX2D374z1zLpIq0Bga3TjZMBzaY1//deVx+EfVzZXgMARm
LxrJL0oJosA8yk1sFXE+vKcskruoLKT2HKI0S7iNV65ZXgQtHqfwtnPdPjgTMU7z
3zxeHyvL69YlNujdzuouFn/jVzEXs0yAHQA5QwDsfOmQM7LFVgLSHlaVhEBPEd2V
BcLlfYY4rTdx+oVn/iaR4tF5Mo6GWKoy5I7w92e9Ppvla17mtQQ3zQPbDqlhuPym
gES6lMFTE+HFiwmbEOTznzi3Tp/Fnl9dHSi2ymeLvxTjkhql641l/aeqb5mzaBwo
43+CpyEWqxd0HB8dk/pjUwLzfLLB+DiPibuRPSK385/PvCJaBsLufJOmzMDbC0h3
g6px0qMh8hXq+V6FsIcItBirO4sxZIRidEGQRGoaUS14L32DQjFocCX+SozDVnYy
GRlk0922reLItIoPxFMBkgdKzhIUT8oYHtaf4kCrfINhqpQxPT862rcttiudV3Sv
wPwIGWK1DcU3+0xYxW/dupUNMCdu0ZCaxNZsJPa4A73r2WzskldM6cr1u+H/cg5d
W1rROx7hLdDMuSLiH5NHINJLCMBTYsLwFS1j4u7jbftN21q9ESSB2KwDTdkUHJTO
5JaU5uMxfXMtlHs7Bz6GmiP8XDYYtpNcXSkam3AxY4gt0zjGl2OyzAop0UqFskx1
7iOvSCWq4gIHBN9yYGHpUIKdV058JyQl2MSozWCIGyFxj4ME5r8zn1rHP7ufOxQv
/6YgcOclegcfni+XTRElqtP6GFPMC8u6UhXdVo8QpP0Z1XtOYu+cT8JfAFYRaKoI
5mkJfVS/syfghQ9d3t2ICNTIAIXjGdO049jf8k3hHwZhC3ww8Ww8Du9/AGvSfxau
DsWXKsqw8WkG9k4XbScMsVbV1/xmWan/83zJKm9W9M6eL1w5O4nePy91H0s4FMEN
PTpKYf9n+uBUoI3nwwTNKpjltdweelsCeZx/i4vfQBqVe3fSI4jwP8ke8NCK9i7C
GmB1sqsdpXgUBmGPLaowJpohHsxm0qAsC5A/QVwZ+aYdDtAqXxfQeTcOwhsdnqQP
RLKb45cpx2e3kPRCKpCuDIU/sbBSXf5UswC0fBkdZaKDoucaaLPA9+VQXJpey75p
XMSU11EG7QFV51VVLPwDIwOKQYSmT/lsnyI20DxJZLO6gxJaXpJA14Zwy6YYL3t1
0u5PvFQBfLbnN8wJaOdfqZsdDqpnlzBic0gnfgsqytEBQ8CEG4BUT0/9arhf8Pqj
SQJWe0jFCiwilyDVNhzK5CbnGNYEPunHbCQ88bfc9WigBGBxuvyd772G9vxsdU5X
oWBXJzuwiddKA1o7bbi2Km0AtbKab7LXvi8/f5IrYq8pioZcVehQk3RCmjSrZee3
HPHwnaQJU8qnI+6K1PXpeNKxlVJjqsTcmLUv6nb1PHlGceY2UdB8ueZJTgdId7gV
KvuCWTCw4zqdx97nourNHDvVpCsbDPm9kYUzbjyKzgIYDhoGt6O2qosIfw3qcdHJ
cjo30JYAO2Cvxgo+dl7n1cCGYXyq07J4CFlcwIbNyJPw5rZ7+Rr64t4IlWjMcR/L
6xvSJZI1Wr0NgEzv9k0ZtzO83zQO47gE6jM/YSZDBCgmOf3wJ2pqy0FyT263V2hK
HphO6UUj56Gk9Ql/gW6OdDF2koM+EMHEU7ATGicZi+naA6iTd1zAFj51p3MMM+sM
IQcj3oyPZ+zpKESACHhloOrgL6v5pwrszBGFZ1lFK9ntrTs1aRqqkbG11rU2jpNI
j2csozlR+0ARATxxUR3QIvZEhMU8yU+3xeupPzeWYSefVRkAlgiXjLZpu1rwKR47
cyKDIYM2MmF/6aySq/hNYcxVGh8gn0nKa1oWpJnylxXubMDNuqI4bVRHro9DeqnM
OIJJBVu1PXgbGYqTrt/GJ/b3YcM0VLeYP/fITBSwrqOnBkdfFjrvz7SdRpuHOkvd
dZsG1lUyi35DOF2R2Wt5OQdWhtI54DpcxClG70I+dV+GDDfaXFiuMYMful+mrE9W
ZIAD9dDLWVyHu6B4HcE6pDPE2WrR89XfQPM4VIXDttwyEZ6h8Hor7b2UJRjTCLvQ
+lIfCzsuCOzW/kWMaOBGq1BsXD7RWile6Ou8jVHwps1Js8PjUiFcW1PB/+P6Sf7R
HYe7GRFT2O7kI+TldqAKUgF2mNgycEsHQbnQckrgv7EIN5/DVUMAsxYdjPMq1Z98
2Zlrb11gwqBRuzWJ3hyA3B6yHP79yzeBZKo+sWw1OXW0ZRoGEDA5HSm8hmWmch25
RmEi9yzBF7gwu9B/7XDfgTtw8sR+qNnqehV89fVDxndqj+8vfSVl12SRlvKWpVHC
D9tOZ6lyKDaWRgP8s0i7p3FVTx5Zg4HbKRlcBzDHb1FZEcukOEdnrYEiQ5V7iTD+
n8BgNdmEcvsLoSlGzvz+FSaQmn1LeU9vhOTcBQDe3Vd/1e4jykbrj2vsub756idg
P7SFGes42kpZe86YriAV4+nMLpmzUq8IveUuyRRLnUWydnKP5kg/Q5lnbPXNSLK5
75pucdBuaXXZ9ZDF/7/5DRJzeV8vfPY+YDlAVuKoeeLl9hLt1+fEIAHkPfhTXh9F
kces/fcOqMf43TVun2EHKaXX0qblYsc/PUTXLaEeIp60JUC69TKn1gHQ3WIPTgNB
d02Pdb5OZZMWZsZQBByUqi15ix/N+uIhuyxHXg9NI3Kk2EWPf+UKvA7Ot/GGWdmK
3vf/ilK0SwtgQlbNHUMFofw0yzb8RQItovaAit9ARiQxSvb3zzPdgQjqCdlI8mn/
W1B4MdHZ6bln/EGY5EpaqiBCdeGRT38Va42pALMOptzc7VgJhviu9lEDfZgO/jEM
jkUQOkmlLf0wIp9gbjoylVuOd/SlpSOoA4WrTH8orpXDxWyP3NAT+HdMUWT/WrTu
OfcRMDI3VIg/E4yELTxyEkz2WvKzzdI7nI3eu7pUY7QehkwMx6KNMEoM95ztqYXb
tHJW+6F5OUaNWVy+HPYWL0YzKir8hmtUX4xjuiW5cSAxxbo6cALBtAxTAygWV5Ve
NiXob1kAy6bTfYNCINGlFKJDl+zPPxNalFlz3cBbPK4a91z8+fqqiTl9yb7JEVUb
k8ei9aV+vSLwnb0y69bQN7lUeYC8Wpf2AwdGgufteWsIHapkSvC8o1SivueLdGgD
6cP+9z46Yn1mXwH/FkD0GyCTo2WJW2fwO6va5LXbgY5l7EnITOjvslYVmetWmJsR
W6g5unYHVW9kNOWh0i3cHcp/4KpLmgdlbZgs9tjqY3vnf4iW8tW9ObxTMJRUhbW7
jwz5zGW1wc2Jx9Hnp/on5RqDUVN3734XR0yuWvm0fM2/lfjg4Weh5Tx8OPEcyTcQ
3/bQioGM/h57QOhun2mbPeTy4lbEIbvjIbwyDXWrUMRURRjOnJ/i4rn7ahPIPUKS
L41DIid/T5wR4XgbqdwvnMHB29Faaz8Fmv/tBjM8kKnqd/u5qdWtJ/+3vYQm/xEN
OBj3EKsR3LnFpIgN0U3hjP0DVbVGgfk7hDv4wS4d5qx1Jo1ypI1TSIAoJCJv0oqR
EjSe2GjlLEp4aNrkP879tLDODEyV79A3LpJ/thjInIPPqtbfgZ7Z8X4dLq7PWUv0
BlMvplfJtT7HZW4rX4+bWDOKIU2PEvFM/P1fqSRE/+IyBQ771B3Z3Ny0NISb8lQY
4/fY70BExB5/R9gphOPyXRMKt5Cz6vzjSBoAlKHUeH+TZvUCpkaE6Zc6OubZ6Xyh
UK4qwcwpqLD6BCn1LxtbItrci23+Hl5lZoa33tPHKq8tBmrOTqU0q2GRqdKkIjfC
SC/P+AT6p9zYE7ZAm4m+fArmOUwaJOyUrb7sfJHAD+LX8qqzIxJ/ggLO1oTQoeev
eY0ZDYYS6/hWOGC8yXjhoNK7kVMgYOBI804+YyEuZn9wvtgpykgE3z3U7iRXPDuW
fZWfnZavoAAPo0deQWuzW3K7FgZf7A3isB4IVLi1qr09m0aKyXTrfPCnJrYefksm
bIf+7OyFQo7i68eEAhkbbhfoQ+3QriNAc0rCTpf7C7RWuveiTDIkp8tvFtKHg4gl
xabBhMooRzhxFAPTg/maJL3eBg5YVaOdYG97NMfVjggQ20ok/UsEihCwuQjKno+e
Y9UvVPBuhaQvXrtf/9w7D7fz9Ens3wOABugmAhlTTS1pvtDAher8GlPrWZ7hm9Yr
FGswu1j4gY/N57S5PhL5477s4GkMHhg/266oKV3OsZFiiAp1mGxKkjkYOm98vQHY
3bmZWLI0Bf5M+wdmD9aWWw7jqCezOFcVc7hqjql8EfyPYQtz7+fWxuD7c4DEkuya
GDctGPyQ+YlndimLn4skY7YP3B17xVSnZqw91R73/4ZKvDqPsnXC5zMmtKrIPDFR
xiNrY/4j+tY2aJVHN7GNkPVOtnbX/4FDNwQ4OjLXDv5p7KA4NX+M7RFOL3E4Mgwc
2o/RTuHnBV4aiPtCipKw8Rv2wM66tK9Bzob0JkJ5TWrEpwppkuLsvGyk7DUWsuwV
WU3B+VLpFEoe8nrqNZ0Pp9Jl6DeeVZC2V1UH7j7d5wKJN4dUidTJrak2OaPxTP9M
elyjymIvpIesbl+kOxgEB/KRBKy/Pd0iX7Ectjaix/yLV5plE0CQNu5z1hJJzCZW
Vz5B0Xr+QwQ78kwvDx86OoWJl+HhisOdRFEIB80t62nWvhbZOIyzi+xv/WsZ9KcB
izSHOOrWSZOGXQDZMCGyKMzb7rXYClJYFzSzI/LyijvxUY9wGPB5Or1QpCPUGHba
6t3h7GSQOQr71VEZocUWzC9hbECoddU6dwLX4V8oarm/j20gxvIJ3AQLCEw2ytmT
WFkyp+pSMbiEjJ9BWX10eOvTvz6NSuZ6a1ezYCfFd/tf7sWYyBU+opWh6uxyc43u
EtetZzSt9/SzkztW9kSd5ntT3JZfJxxL0yVQw1NozYzlk7RYD1lC4y7M6Lga2bLi
2CsR7UYXSBZSG3e1GxKDuXtxCZOX+86AqPORRqu8d7iJWzQyDHzmM2jXT72sA08K
Lij+C7CmTFqapIw8nDsGIe2Vrv/IprEdD2gIUH1HL/VEZc0y4Fb/GNz0rXtLLPdj
22dQMnxve9tQpvTIshFTaV4Jsrv5oSAQYUzgyyAVvbFj2OVW89/kIpXYVE/gbOsy
3fXp6iyQdza/61hLGlX+kpcU/LJ4vEHDgb5v4Cd+XmqG2L6oP2Xg7SmZqc/hd6pN
NFrTDJuePB61PEKXqt0et87Nyc+r0v+istz+xx3VVtKezG5rdspEnK3dkEGRW4WV
2X0Mk+uQR7SxfDxRrbSOS7Ww0WfobIF3KUnRwz8syZYgp/93WbvW0CwbVf4BXMKd
rEjlQOo9OoHjc9EeZsemn5zONSiay/NqeF8GVw+tbO8wLCoVEFR7ta5+kPmYhHlz
5xx2OS4TBvf8xd+d4W4xGqcQ5Ntfdyml5TxS8E1wbv3iNYB2Nbxr2CobfUsVBISy
/xRTnLZOlXPVt3h9JkoFUKeMjy3If6d+YCia30+48QYwQQQO8iyLC60YhOfLPPC1
eQWzhycWN+4f7PdK1lVK/wnVGTa77f4jxNiIE/dbYCNuzau+NhHi1bV7UwJFKjJR
Q8m6lv3RTJdHwD08MTGhXBAN0Aa48qSxe9A3ZT6ZdhFu4Ib57aBsfYkT9gA0d9Lw
KCtDio83f5vGII/+3SG5JowDHxKBjrwbEuFBendpDAUL/naSwrrC/gtEWLvl0ZWb
oRt4NF3EnX2fHA/EDWRmzC/ehbmrP1BBt+VCYkjfZ6ldPjr3oSXtx9bgt98t1wXO
Nj+iIlkCmAjpVcyo5+cGi+FQjcxIM3UKcYKenQmPGtw6UslQVJyHQMvZkCyC5UAl
YWrspMq0sdWjPpO021KJll5ySp/Ycj2WEasI+SDVcKBhnWHJ4mlAf8RYB8iJGHWY
AJ/0R6MT1d9/DYMrnXspgF4VR1ZpHAWD2kOw5TwGwFkEFsMRpgECyRXhkl1Ro6GW
TUkbXxJQCGJpGaF9cK/Ip5IkbNw8O5DWYWo7AfcuhkgrTeIz9+ByvqjYNnNIbgXg
TRGaGLv8v9aTKOrUN2XICApAeEvf9rfRebipFZwI/M2mOt7YaSXFeb1qx9sJ0/za
CIX05MKhCgJjP0ZoNzWdCZ0ah0TGPUTI4UBcwahqg05aTA2EHZNhXWR3v09/CyoT
A2cLRyVdA6dPgpjUrlcr5mnMh+TcEsUKOxm2ihrd1KA0WBr/zT2BhRwk7tfboanz
gSZFW8i4yf6vqlKwS5cD7/sABysyiyHyHURI1DVCFnDIWjrfvM+KU5tND9CF2LVw
YDXrcpx1gcOF3EX2LrgVRRVyNh7XTxi4xGa8WI7xX2jkwRXBcYUpDK546tAMGANC
OevJG4FzMAMeSEKuNCsz90sdqF1zK/9Xq8QVMjYEFqq7rDxql5rsnzIKQIOOJHOn
XiIEMJjKNn0azkjKJavkLuqnXtM++uV9MxI53FJfVXA27j86F9z4QvNzVprdswhc
LeiQPKzzFH3JUd18OOCxcOuHsYQAfZkmlIG/QXubLsNea6jApO10Rc0nIsWcON3L
xUx8ZR66RFWXz6hgIpi8Fvg2p6aERjSDXwpaJVkuY0SGdBLo1fggy0r2ykppyTRR
8/neLCBxPLPlE0AT0RLyfcpzfNZZqmToCkZW/WIajvObKW0Cka3VjBqfzludf9HT
MNLTxSSzUZbEwpnpiTOesojeMWl+GQCxxPaOSNTwCv2oUYBrX+DB/kbTj0GcLbda
cFcBp9tyo5u/hnzAe5OJ8YS9FsHUJ/+a+CyWyTqdgiShlUe0SSQMV5Mkocl5+Hhu
a4iymGFMkWbYVNFiNeTT0lohyPNt9b+lYeRW1wzy5+gCg4ZOgo0u2CLMEIImzP/s
NWMJ9JsD5UIwYlDFftx93/AKuXKj727TPD3009CKYKP/Rk2dq98+gqHI5X8wLBpd
7+jbxl2dd3zPC/kLpNQMqbbvAuiezkYHk38njFp7GewR9eUv3QWp4tf7m1hCIel9
GBWqFkxF26NPs/Rp9p5R04gNaAJDAysHatbSFg4xwB3Zkdpmc0Blnu+8BoKyrvz6
6aygznxEW6DJzq8py0KeAmYdpLNaP02xNJ0+WprYzTz4V/17zGHHEjl8H9IOXo1h
sJagGEOIq51Zg7tVnp4LCpH3kARVn9n9Z2IH6PkRSTl65/ZIQthW5nXyV38utRy8
ETMcLdO5h4KaFUQsE4P0BUfKr6kKMg+ehGcbyEwJzMobfMqLqITF9VFVR82GB2qI
KN1Dp1Ev7su60wzkIGpxn+rJvXxw2Wubgf2sy2ZjqGdfXfOlAWJQYNwMdAGK+vk3
dZafw2LPRK/hUlkpjBrYm8YjSZMDnKbBgeSj28mq0lXrk3RtY45JwUAO5HRz5/3s
gpmEGDcq/+hRPaBAhXn0l516to4tYkX2J5/1xEC9JNY4BSL4jQXSlp6gYjlMbW4s
zCP+X9BfcCc2VysV4gX9xM2q5YCAc7kW3HDoWuAADpvbA/QnJlfC3fZKXJd6/S9u
MgYwlYDrg5oToN5ZHCNiu31/mH8/JRhenJut58u60XfVsYXiKVf3OoG/1QTPJMTC
zhfH0IOJOOW7tMYnu/WOYR//yTp+t/nbvEm8SNSLTAGrKwcIvviB06sKeWOyLIfH
0DzJAvTF+P+/AvYwVcZlyYGWypH1pFJTZwW91XZr7iBTohLgTc1mgtrcvGDbp5Ni
ofamjxjiZkBgiHRLW0QuOzHQnMWrfbs3VP8riUiG4LG78NOp+wiAGuC/7/fPUY9B
wkluLsTmrcabfzGCDCrKLcGT7xUH8q8oIeVN2RMB25swN5riO98YYjBhs6fkMZ7q
AvvZMrNkY3SozAotd01WLogj5lqWy58A1nJW/BiLZ3MlR+A8/NhBjc5hYwXVt4eA
hPAo6x2wiuDts244KZWzgu9QGxFdfJHqOK4mOUcOV1qfwS2gBHivRLms7JcBhWBF
pLo47CZJI8N+NlZ6Uohuqy3tIQsh5PtcYSgAUDNQXYIWdqP8tfWaKY96Vddn7PAQ
ZZslH2e6JQaapo93A745BcUZJ6pULWPrNLsgb8Bwj6v0xCUk2afs0Ngkclo43Ns/
TtkRfL0k0B5GSNX9+IOVg8WN6URvvLwW4+iKBt9FWz4TbWyucyuPy7SWMOiOgXKP
RlP69R5UHTEDtvaeT28zZUC8XfM3ggbkWP0MhE2uAGi8kXkLMNtxmRXWL6S9E46q
PO1PEj5UC0z0rkhGWlyqYU/nmdsirm4KulyOj6koyu1cSFlz7BMAEfDh1j9aTcOB
SqruRPPlOcHHlgFrjJlatDeeOeeT3gUnS2yATutnImvrEHyfEZAUxjxqhnyL9TjX
6AYgBXRwDYD3tNOLzoDC8nEUXXU0bhZ87pcSdoPGsBLcHPgBYNc5Z5+jxXCn1nWm
VI4UPzHXtD0KPhDipWxi1kAf0tTrXpbaOTvLGZtKBbCsj9guGO3WsW0cis7Em0Ss
hXnF/HH0lxM4M5IwUWeIbUzysO50BYpTN5IbTZNLkpK8CugNFJ54wiUluS0Iw9du
3pnqc6EFRiyH0o8B7ZMdjxF+ck7g6/a3IApw0MNDxZ3So5X5+JGzh2yTtrunraNP
XVztgBNGXCTRoIeOvAHQRQqBSlP8AX6u555MuonDCGHQzannbEmwwM6T+AUQLaMp
5uIohSOctEC0CPiJyfFpgA1txCVGnsKTiB5lqwwbzGZ8QqZqAtaAorvlKLNkcakK
7FN70xBIIwWNH/fBs333CYDENxZzfEZgt6cDXAI39vhibpT6VwziSL1y9ua8/32J
rTOu+JgJ09dbSJIl4UyEoMJq45jq2EoY3L/tA+SQVsR4gNJdlPLpipX/U6NPiXXB
V7MTlSnxqUnnBr85WwxBgYznZjKWQC36YumYMqJWAi/k7D3MfjnLQ+XsG60mfPdF
6ScQwT9qG+5wsG8nzryD8haEi4uLzBpDeR2o7q6rZuMtecJ4wazGUBemnnstuRtz
yNk4EI3c2LGTYJHyvFwe4a9NI0UKAMQX6GfhZRdezsobLYygJI+yDtjaAT1A/bkF
7Bz1Q9xCItq3+R3TB11LiVXOoKfyTN2OXHH1H63sjpJDPskoM9aOGoLHRZus4GZR
GXXVQGlDB7Le/5f1vNAtBaDWZwT2uGWWCReRFWVo6zx5SqXtbita0tPSsX9+80WN
x1XNcXvLfDRURATlXBuJXfBj5sybWCA1aE0kSEv6YGu5ys+EDmhmz9ApddjRyvCo
ir402dvJqtAqT7h4s0s72qld7ISlRJsn4gsSPmG3jo4Dfia5CecMUB6O+AA3B87g
IgeTDxV7o5zxUTwRbq1QSl66qy74ALgavkOOHpD2dpkiuSTyCIPSdDHgg+Oo2kZ1
YnqBD4yOkrHhyXa/NkqGYT5B0acawDT0Ac1pVmkiP42Wue1DGDVpOGDLyoElswVB
cJFqysxQLy8m70rAyv/tntJmpc3G2UbM8E2WLG7E8x2KvXO7e7CjNhBir0eygRWZ
P5Ybq7oxpX0ZFYeLy8Yc16NsVSsGnw954OYqbV0HZmSHtz95YmKyZAPIhYdzwJOB
C6oA42fQfcZ0S5L/yYh14CCY0ZXB7FU43TbH3/yODNVBDG+CYLKUe8F8Yi7dDpna
cViEa37j0gnrIbn8fuTKLIzF/0qvKnw8PRdXt45RzvHExd6S/S0o0DlUj7A6HYxZ
t1Q6vkUzorw6Ed9CMAKzA2HbW573FkarXlpltnhS2rRvSBwFjPIHBfg+IPN6FT8C
DHPYxMN/HOx7Ctx0Ew+ivZL8yIwwVtmml2rmF1pTO3+kjgSyIzGwq10aSlXLplB9
JuNKhGOZHNV7jFNSACfm7PU7oy8z+1DwPeYcs2KH3OYnkV+vsVmgI7TMGOBnNUYg
Lvj1dyutOjYIBYgMRi7S8DsS872FbxSuWbDq9H0HXjXw7kZi6NECtmuLTPwngkfr
RDvm1Qh4lBA7Hb41jOIHxmcrVjcUBA2JqvIfbvMqLgp+jgGlmN7rfVUhnOt3v0qu
waV39Is36lRSYviQnj3abU7c6nbzq/D9BfjjNgAWTX20ovYfOGdMCmsNrfGl9IKm
wZPPLsv91od1lxvUjoDeIlcPLjzIU8h41Et/bD+QiTAryA0Y+wycxvT4eYFVxwYl
R5M8sYxu/5Tq0j+vl08kyffErTKmaVOdn3qsOBTeu3YJUCktx2CktvlFL9Gp+yr2
J22ct9akZ2pq5007Ow47Tvap2hSTDOnNkia6ria5z/KQvokvO/uxD9Z/Y26PHI2N
vb6xdvnBWkqi0aEEghT7kKSqm73QFz9RvNrGjFyGvEo1aNAops9z89s+HUP9pu0V
VUfl9IMqociNH947yYXVBoXsLoN5boalGs2OeE5OrNsUZCE7jYCP4VbXhAq0Lvjm
1yKq1pyMxVANgyE6LzoFqw/ga0a6ebcdQOsb6fraCwIzxV9UCwGD8BEb/o9g+svm
V54hP71XUgD3ICD2EOp5sl3SLOEpuvzSrd0dybjMqJ2nlPSlaugSi7WtL3f67ApD
tVnidXyqGfX9Hyv4xBj7qWoRQCs5pRX+en0581I0YTTmuPEo0gRe+C3lgMYrEdGj
KZTDm8MXiiwDDV8Skrr04icskHOkiCtwcaiR8PQAOdgLaxBjJdkOi+6nv+znM339
A48HSGUOJhscWwgS6wLRClpZcwk7wkErK1XwFg65C6HaViYUnFJtEHiV74uzeFRs
1NrqrAIylEF9fPgdiFc4I5PTGybkLVnJ5CwgdAnfZ5BfNW8ZnFTI0J9CihAyQzrW
CuRfWtd/9SxTFY2SMOVH6r0sP7ku1QT2yHHRplH851yqBqLQEIMuLIX67UAU5eRX
uX2xELoaC9bO2ycPrwJ31E2NTUnX4udGb11O+H7NhOOF62bx6vF79tQa5jZD25Ba
1mW0roXO1/QRONnx4PRIwZnJE7TJgbyXSwDlr5HbdNYHa3LulDot61pXNpc9F5nO
6PD3Q+ZNgz233aZD+WW+W/yVg/1dOeSgkUvNbrsmOSsQoEnMhQ4Ga7Qosqwnn2IA
fJuoAHUyHMtqv3FBcasYHz3gpPMGkJmh5GJ/32HH4wteb3b5JWPrI2DAs198r3dZ
1ySycqfLoDASQ/e9aCGIS189u/KTjrmu5e1Sd7UreOZ1twUB+A0anFimch8lsBs3
0d7SrIv9dWsuc6HRfrKvJF9sdkBmpX4uKMAZDdih9sEQ7LZQgAGplfqOw0XZAlTV
JPRd7r44nfVhpQXJzxc4XsIlSjY2At5X7lWudbhrWR04dd8vWrzdU+RKyrZArbpL
8EJhqun5v1pF++CoTbljMo2x6OTdnss+Rxmd8uC6q81u/yC/WE7KDNPTNyee8OrH
pK6g1RtUbNwDTkAlVLcsUnaiesvr8hd1P020vmJpigIaHS29qBcWdo87WGc5pbba
cGwMbWS+tsvcNGIjageBmzony6u3H+WYE/u1pFcp32kDGONjNdlEi4gBzv0BxWbe
pvGj2lvFY1FDIjr2zJp7d5esodinlLT8BKSFYm4ITIGnSDWtrPC00axMXnGnpWER
KWXaW+tjN04qps6jg39zUyQktNQKdfn6rh/FAcAqHWMWFpLrTljOXFTSLBeiBMS9
DFcCNUPHoys9EdV5Z2nm1Za7BdQcIehyWDG1GblQ5gMu5Vi5BND8KllkdVtwdX67
Pcb9REznTJJ+RCJJuIoA14aLNYdNRdalAefdk3GZXlfocddcaZyTuMv8DXqC2X4R
08nnt1ccRRG/YaMy2m77H3W1GdWto2ufmVKMK3SGtoFMeRumdptowH7uFmMo09B6
kZ26PEqk6COnieFm1u1a/HKuGOG+p8dxonhGloSLuY2TOSgU57Eagi9GAoAB1p0W
WP3dPrSfYPMIHKt0c/lxkscKDRqTUQa1BULkB9iJY69SDMoUym+MFSgk5kXtsGNR
iymJ7X/ESYD0JJ+f29mkhdwnCqIyhdxVQar0Z3iMgWUD+EtO3QOjkUpkdMgBCLsw
5bxyMJnw+MTa3qs/Tj+JHQakIKIVnKyQhbkzmUXDjHEHodgclDxytX3woJDkt55S
tG+jD6RuvwR21K6f0fhEGfxT5ddnOEpSsfZfeXawpY4EBevpgE95raWMiGFLvbyw
kH5Busiw5/jzl/5OZ6ne7RuT4E1GKwJCISDcTfS0aM0JYLGhHI8BIPMXeaGELRje
uZj8Zvs8Ux5e6vo+PbvA5YGVOuyaN0uGtmvQdynq97E5yu3PNzTkyZWM+MFxUBFK
2XnDHktbqFG1RKYk7BOUKM1VsAvI6pmzSUrGGyi7h+K12TRqMSahUNqdRIH9rJIb
BeqZz9kIlMdU+TUdHuBaddrIIJCwGcdy1ai8G9hUDkCo6mtTO6Ik/nFkjp86RdWU
B3yhTHm6JileT+cC81TXe7kGnPZyyjQ8yjDKOEV6JOGy2EXhwANExMoFv51Z93W4
Z/zXErOsy2e6gYx2/AajW1d58reySKcC8KlyW8JLXiiWMUr7EHErDAZJjK/oWajg
VMDI8foLZSUhgcEUSlX/CF5XlzkbC/UwWMDZmr2DmWVrhCsv7A0G5Jbp/U81wCf8
XLFvbxUQ2nCJbmIkv1ym9XVb9mNbSWG2G4Q3/gRIJQFhLTMqs0dGGRS5MWkeSOYu
kiHbauQubz96Rtp0PvrotufJ0X+ReVk6xP9FRba8jJ/LLzEp3P0gBeiNv8G4Z8Ek
1eOP9KE89KSVmlIs1S98w/byy0M30qdiR2ckCbWLONHMlTKwEw2lyHGtz5j+1kn8
RU/wnfLzFE/Qrqvw/456fiRG3yZ8Y/KWjTOuf7ZVNb3x+6/gBdRIFYE46EWRiasy
ApoM3BM22YyaXiD/TjN1zdoWGX2gp8p4H9P07JWlFYX0k6D0VYXyrLMIGnNY0WIA
lEvhtyYWHz1ARpTdLr22cARGWMNJNB9gHYluFz5fQqSz01y0ktyDtKQaFhEI7D+N
6a+QjurPdzPYKyhs+OXbziQFfbe4O4bc+I1cbeWV1UoWecMsXERGvLT/xD876PWb
eWWaq+CbAbHO+Ju/TvroaavgdIp+SuKxWHeikKuqkwAcx7o1LGVrmNj/AAnno0vM
4v0/xTbYhLfD0lryGLo4fK8lhll5nuiTCEjrz8hMbdD0R/dC4Ic02hpoWAZBS4Wl
xWEUeEZOTb78E9kb4NdfvuRg2NtLuqRDuneJmvUGEWcmLaBcYwH8i7hS1PokuTGK
TtMaWeUgZYIm15Iz9h+j3+qZU1Nj1uX8C3LURSeRixSoFZGw+WZZnIlj6XBSCjjF
CifhOBxvZv3NTS1XVfrOChWP/8kILNrPSsvvlzYP6zkh+FqeEkP/bCCibz1iYEVi
VZaxvR0a5sU/RGhhOZqAz7nvqOAy7sgbPTcs4VKvYkgP8dfZXZpFffFMFGWqZ2/V
WP6grwMzmUdYgcAkv5+ctRaMDOyh/eHasb0ei5u5w+Prcw68dBcpHsxKMZ8oCV5+
GmFoAGNQgkHx+GpuXnwSMpNnzAxWXgA5+PvsSVtVo2FX3IqTmMUl4dmT4QLweJSJ
wx2tftOXC28T3h4T4oBSDZGp5XNT+C4ujUgzX4JpF/2k04uWBCfZxScOTfJBPwde
ulp1rLLrpvoumPUtPlWYR3mlgyYoHZB/A6JPwli2TuUjXkRRbX0B2KGmfBD5oNXN
+oO9grovxUCd0N+e1oyKDxYhx+soH0CSLyV5m25dljdgX2VXUNzFnPrw1ova8ni+
FgegcQVs2fy7F0hkkVd+L/B9Xmwzc1AVVFP3NZxfcoE1h9F01KOdpQ+PYImPVXax
AtBZ3raKjRYBAICOqp1wa2Ofmbo6Lg2yMXQzOHhq8OvfpxXkzCK+y4qC55tARkrl
uo0OdVMEnjRIJYYL7Pj5exNV0PU6eASE4rgenQbvIDcOsBHgUBLHHmwxHOxmK31i
3teQbOv3KEGzRy7MutpvoNH9ywIAaWar0hORDMtL/88boBa5GP21SeY54X2zuZhK
2M/alj0sk/L6OBW2NxATqutPKbgTk+NKzYGzJsHzFXT6c4Teb5O116KYGHPkqWVP
SM67mJO/KO1WfNC0/vfqGsrBOGLPcVsz6ct+SBQGcz/Ob5GwkOn2vjvOFcH1Y+An
v+1soKMXcoYB8cc0GqkZigQXl8zIOD10aHA4MaEyEdKGmeGFIepzX2PiFeQAPMZY
U+Z0zXjLtAhKPbZXLOM2btfW3FXIP2tFJ2mEIXR0N5RDvCVif8xGCS4h+UmDh26s
S/mCCofLmIEypn1U1d69RUroQVxL9dJoTW8h6pL70HuVYvWAn3jFhs79wIX4itDk
hjCGQx1Mo53gvESd9F9O3lFtoFO8EvcvGi3G98vRacX2P5+yVJWV3MP5gbVQZZeL
IFRdZswleSnLVu1XtUdAVx0N+7DbYQnM+z+nDOhnO0XYUdW0GJxfz3kLEoSbtIC/
Yvoax6FGd0t9XGRAURFNGq1g+xIUzFvK7QUv16wIJhwJfHg8kyXsQuEtvO/yTZ/s
cLvs39Sba688RWrIAyW6QiiHStVr1GuF1E6gByJu/ubQPUBDH4yhWs5G/AIih+cf
UJXEjeLyyGdeAYV8JW/t8tpM/rFw753ZDZDTF3LuLw+FIpCipHC0nAV1T6CuoRd+
X9FR7FIrfnEtjMcv76hwK2xjNkd0A0a6iW7I0cbN1M+WA6LJwXPR5uAwdO2SgJA/
mWHjUZkTnpTMhynjXpi7SVuXrez2u2kxAKWG0JNmqKRABQas4A+8Nr8SfnfFItgG
F/Y3tiZ9n2Mlw997VBNwQPAO+hFtnAfdGb9BjAdoYF69ztHlEX7d9WFrMmrEHuDk
1CRepLba5i+BuoYd+gGhSEwOZlfNZSIQQTz2WTAVXTlp/wgZjnxGZVqK6QcTgM+P
GqqJQizMsrsWliBk9VSxdHWYDbqfv9lvjBP4iaqjavgiTa5t2noY/HLk9QNhN7pv
zVvEEEu7tv75G1jOEJ/D3XqUebwjHdheUiTwt69oI7u2yI6yVxP61I0QyDhHmN60
bFvVCXKf1fiBdrB31jgeV0MR7NR+qQM0GIHJgtQXapOlrtHoBx2mkNDF3Eu9xosT
8L8433FoF532/4yl2ujIj+Z8m7XSvqkhRMVRjIx2gYUfzqTTrby4+WbR22wYdosU
xlLWbL0gsx3FdFde9WnwPn+wDDzRwDSw44roDcfp47w8TlDe0s1JAwx5U/afNA+X
qEKVbSYuiu8O2HxciYkX+YBmv5DbaWPpCtCWtXngnPG7Wr3KMxhNiMik6WTr9pf0
QaRiRSwW8XSR3Zgdotq2s2AD5anLkKZAZh2EMnszPseX+qFNRCiumqPre33iSFJl
ZFxJjoWmJP9qWsXJPV+vGqeUY/fffkn7mTt+bc0QhvXcrDFCfey4t+OZ7f+hqcxB
jhn4hT4GRRbEDWBqPmlJn8EzXcMiWrrs6IrTj6GkV7xlJrKFm4bblSj2uGrx8401
2xqrjtAN4COKBzpFj/SgRtWZiX+99+Pw0o6qLxVxi2upnzXbR5sIh8hByiU5yZDr
RCoNqyOnsEqF1LLn75aO2nwqIZBHTrULN4Vk0ACbyAdZa97WpBmPsYlPYY1XKmM8
fcLSb0MTsDQysqMKHxo7uj6Tm3kpa/U8/tLFZkUpzUdVZy8djLOZuSmHwD2jhJWn
4Wq7iM2OS6Tace7nooNdIys+XZ52QmmnLPPU326qaSlY8MrKpTziSd4TeEs0FNNo
TPtvme4C8u8L/xdaMe54x6nwujorph3hEQWtQNHjx5zVeUaFKEqKnLxC2xUDHPiM
LaTqFXJSPrpdr5GonF8Vrrgo/cbUsBsyGkBHmd+ClfhM2D/mHx1pMyqeoSC77Qag
cJ010hZbWusU/pPflOOjjEbQvuNCBVYhIEXdVlq8a0/TmjuuJF2OUgYLxPCSg/KQ
r3Qt0wn2SRVd5gE1bld8OQuOW5wcxyjIMDB2hBMVMHmHDhlz889qd2efffk+sG/D
Nl26drLb5uw5PsdI3iuaZ/mrQBwdRNexRepX8yWOb6BBBwKvhCjPZflp54xLMPH0
rQ5o21XaJltMffAR9y1C3HJtyaUkFDdzkwAMBc7akvgwQWtghLcnjR2qiIjfvr8L
yqG5btQM+6lM2HlX2l8L8iLr1pWOwz1rz7TbF38gYQrR1tIY37yGE7iZ1UeBzE3T
ocKPGiO490AnpB/jdLtJUc61QBeNII6XWBUmFi22HgRI46YUf6G8wqpaUH221yu4
RFFVH0GhQ1MYqVekSxtd/hXXkWhu5TCXA5HXEXTzPupv+F76Ks0kt7YmXn6C8+0w
zbzfMuGgHR0io2oTIz9mgCzYqcxAxykdd2ZGXD6PZk7BdvU5AhHssMYHKHHpNpG7
Y52muj5VZE9qyWfPb+YxFI5/lHRiRAD/uGTkh+pwz2EGkkY9S9sCB8FmM7QbIopJ
oOUsLXaDTO8YNJjDCaSHmZE5U/iXTNfoavKxmOF2vI+UVuaDpmgAfVcLhsyUMuTG
UR4Hwwf2YWJXbLJO3K7R6OOOBsnIUbpCMkAgaWHzLQmWkGQ++da/NX1prXCuP4EC
gUpBg09dUDkLtFwKtOekiDzwIYsrBrQoLsYixt9wYZs7wq4usfHiX9ZJ4tIbHcUa
A1xUp2K/sB1gaSRNSlkOpKxCXmlo+q6TedxXtxFskTpLm7dohbHqSaYyui5wX1WT
bV2/fY4q+XJJ32+g+7Va26Yv9638NTDQhMUDx94hsGq6F4VWsVMI7cgCXq/jAyoR
U62FINyGdZmR8zPwWUjHkDbWPX+JKOAIOMwdANuS63bqp8frX8as0+bkqiV1RYFo
IehDzeRo43K9W+kN69AC0v2qRgbjsjtOF4ci/94YwJhhrrM/6sa4FelFXgJs+uPc
eGkS2m84lDHkud+5OD/Jtjmb6iITxNyzUlvcdhhUzpVcmyf4Y8ysW0G0S+zBs+/x
BfPpuTjezsTO0cmNfwH8yzyIdf1x6yUtQHF8mu9IGABHRtD5yEKvehpPnbhzzjTP
/zGnWlRP4IKeU+q93QjPhpueSxLf3kIgs47e/8/7SV4yVhMKd52FY2nGYAVyDbu9
uZIhR3B0xchmqWOzYma40PXbqR8ALXbzuu113kJl0UhaiIL/XeFJdAJDGg/tILhj
YMkQ96fTwNoqk6i6ixk1ZOhbuRcA1OS5SLbbfnyBXl5Y1bEat76+B5VjfyjQYrDC
lwOhfmpLkJ7rj0vm68OKe/1joPlIKC4OB9EeNHLpp7eEUFJH2oXjjMY0EXphDYtb
OXUUESsabveulFNbmHzBpWWOn2TwxRoOSyrMu8h98oePaF/uQFH5TNeqbgtA54FI
IEumDNL7jBwdVUPrfw7/BqpAV1xuINOT16FhfrSocPceF6ZE/8O7f2fNbgWja196
QiP4wczK9eEu1gp0WY/5RqgVfi2gRVgegpCL/7BTdIkxopF9vpXXnz+nDZInfP4L
U8qOwOQJFbrL0unGOVkSG1BHzwHuEJgIli+RVgqXS8q/rAZkmLp367p3/s5ndFzn
HpslN245cm6XINDRYpzPKMaWdCsaaVZ/wZiUogMNKiz7a3m+47Mvr1Gpvm7zeSDB
ljHqSXk5qeKziv4QAF/OO94ynSZ3vVBesEKTkHNx7RE8k0e/9w+6fywfoY9AbDBN
RItI1d/HZzp5tf6GCEgipEUlECv4UN/L0/RtpsZ3A5v2Cm+u5mfkr2uTZJ7lBI9g
Dzz5FKbluXL4K/uJFu0KVxw3X/w1ofOgHeOAxMs7ivTNKb5xgXQhiNl8yRlu1CvW
XRplckS/lAehw0LvVVkq+y0Ph0Rynuq6R8YRya6cbBEqT4UMgdhFn0Ioj+E7a78O
vthbjybFjZfp8Z+5+BCX4yoRyLtQQZT89/pMxX4QAoBRVR1mmKUvjcGQ/CTHncmn
Mtg1v/3JbqNsbau3reXTc2wQi1u5Ai7kKjmIAa33xCbQW2pFlJjHDTc0C8oeO4pD
Ik5UKz4oVWCt0m30l6qeXrTNAnQ9/ZtnYotDrw7qBbdDsc+52vxfzumjPz58/5Lr
/EZH0BRVw7CV3i/6ge/f0TigKx0IJvlH7gimKsKhhunhnSBPPdZOi0G+mcwBbbQu
F/XEKcyt/Y6HLr/z6dcGyUr0QlENal0L3OO11ydTaNA+Ey04QHaiYhsCvIfYoQRg
P0a9LxOdoLAYlmVHE5IlIkBIugYJO0ZzRYQbEzOHW7nZ0n3xvZDZgxJ52BLTGiJ6
JN7uUxnfhGH/KVaYXYIWa4pyq563JoQ8YNWHTQzNXUgrt4rP/nz2movgNaDd+ogE
vuhGs/RxZ9DY+olGsTmIJ6sLsog5Spgmi8F+7EXyXChvWNZ4wFu41T7hvPGu/ROP
eb+P1cqrAkwyUIBW1gayiRshaZlfEmiNP++13GYSR+ybN3vdteyAdiU0gDajhtas
kC7jGH7vq3VhBj1oIYNJIpRRJPq/bT+9CFRjyYnXSEwJnG3HbpAX9aNwtS65XaqT
r3znCj46PR10SNQjO4qmagvkgydNBBq/8tvZcXf/PCo3J/VRSrbpCgevWI2X6SPk
e6pECUeb36vJ+uieFfTg+v8R9YCJtT7BmBGS7XT6sPsUNcoSgi/86l+T8roEyY8r
U/t6B5pt1xurYvrnHsWO/UuqjMPQY7MyUjAbnlJSee58cr7OfaBHR0JEaLWOJIIo
4UlmazPjrBQv6knUIFANE1IVH9IVZyO6QxTZlevQINIZWImH3w/g+iAKtMqgF/RI
YnQ/E7A0e4IRPq3Lvt1c0l/LpfOfoASWcBGDBBNHmVfI7YrbVHuMibtNgtAsj3xH
7RBc7BjPK9TlM+yJerwscjq6vg7d3M8kpbRvOGRah5fe14vyBLXy8rosTKiOWaj/
ohbxisXpwA/+UQzsv7anjUpowQBOkx2TR49InPzzi39VSqqS6adqrRAmvxewITj7
G3tCbOPbmg06EFXO9P9De7GOZcwZ1PHsOZT/iZSr5kOUd5w60wnRkQBkNj3qxCtU
nkxQbA8SEu4MSsdRj/IZok8flyPe5kAlBmS6yEqq5lFYYURinQDrfWGxVCPhzB08
65nRuMFj55Q+LEjKsIUw/oRK/dMN4WsAXdvvoteENMEYw6rvc9o62c7wlp/aIaSr
+ELo7jOw8ueLgSKgp3CePqTzYuDLcK12YEtydz61CcYDWhpsWXVtNbXmLyhkYj0d
wk16ePsOJOMb+mGenCNCcwUE7GGJBBEwwmXnvofmoTJrSvq8eY8WHqMkMgm2kl4T
u0n8MQ7bNCK6BVUjWmJ6Ugh0k1rX7TuZC1di7rkgNcAdRctfrDuQFdRlj/NbP9NW
RdAxfr4z45bNoGSXRxacGg8E7AhGcOFoGOMsXF+AIQ6Fvh344nrBzYNEKfHXOFPV
Wnn1oSli0azUNCuzrmFh2vA3jzxB4/i2KZ2VLi96/MV8XPoU5cv5s1KxNmBvFREW
kr2eaWzckS2TDmpsK9FJiADdyDFyAJBUOniogdEpf54zQERVj5m/Twc/thdvzeRj
qK0X6kfl3StR27N9BT1RhnuG6No5ad+Sij/V+nBwo8lUcS9MVKoh1QAxSvQi5QKv
ZptcuMiJ2LKa1GzRCPiShJzZ5C3hN8ahaNdUruA6CfDrR9t/JOdHsn61c79hIz4L
/hbIadKV1HlNXFHIjCpLPin0oa8Wfdb1Kk34NAdS7Axa2wZf82n9oe4Ulm6EeUAJ
YCfdDYf1gzRQi80uQh4veh2ogm3lNl1jjDfp4+wcWNVgp+jVSDdfqNjPAoGqmVTF
Gh5cpZ3Ss7BvaLz7Hq2U/uG/ljdVeZoebJ3fE3+vS0U2BRgEINk2mF37dIDkT400
WLUDzFPU/O1uObVkXfI8S9SGV5rTfoMiXWUOusy0nIePBRPbO0/snE52M6RHC7u6
f9ajmTSyMvS2T7kRVEupczIQ8h86+fjuLf9upzw6ScU7H3Lhqedv31w/GDwdaa2w
SH9raVcnFwnzjThSK61lUWoL39w8NxqVpNOHnKPGc1ZORQI7YNg+YIeGTALj20Hf
zisXT2CF212MjHgOfMpHS9ByDjGOf56ElSxh7XsWSN/JQNVks8+SYkCtsK7YmvTu
Qw45+rdCfr7nSjNBvYVhBbMDPrgxX9Papo6IoiOTttf+M/zJ23TUUR2PXspDdWbO
UcWavYwgZAo+xTNXE28S0Lge3bZkf4W9b1yiuq9aWSkfQWCjhKeOhYyTTAXzKqwv
ARM7RSdVSuFchxMBC8UbwmLuVr7a/ziCt4cwpbOCnWgZD1Afw4IBXOmZSKyKjuNr
nIuH6WdZuJ5HjcNfIn0wI1ndy7lJ2NvIsebpP5KNz1ZZ1V04A5sU2qcdvsHDc9n/
5/XxnfCuSRzZqLW7KlfzOnaswf32oCQYHsPnFsWTBVMl+6XIklW5XC/McASTxBoi
qH4iep0Ib/fP973bB9UZ7oWmb44u2cnw0EvDFftXRhMP+xMMXcuVJRXmTeVS7Vuw
wm8EYT1x+CZGo0cslIL/SNsigySyOKeFL0bkLaetNiVip9pJoKOYl0lay2Budib5
p60DAteQKDERynuqS6bAmezMvFg7kaObvtNp5iuX+QyUPPWbeWTVj5EM9BwbyM+z
l2pY7RCQ60S7wlgGUpEYEJxjjfjoMocU4wOVyHeA9o/8Qk0K6BLPOnmQ0HYrpSuv
Ad9nvdB+vwBjcLHcw7DdHVq80SrC2kL154UQEO47f8WSmVZ7UPMPjnJbFmYwX6/r
ikrzEhYMw7tan60TN9Vw+PwMiJD2rgQRnyATPkpHzb0ncTmoeNadh3rPau6ewAGV
gnBDkC4nZJCyalcezI9OD0SzaReyrYOoj3lSitR6MhCI8akLJbKzXfccPFRJxmXr
7+zZruZ0Vm5bCy11HDHS5y1A9RsgC3D7snqF32uO6QWmKK0j38HU75VdRLknP35I
BYqvCaQuDxNFEj9SO69tvH+JApQrRykD0dkNr7MZpAI0FaRDgtgDCEkIUn8YJP68
3Yrlo7HXf2QihZoH9/ApVMFos5KexKWQGZeLQQb2jS5XoNTpI06K8X6pwLepxWg2
GehB2A5LaKoukSsD3U7I0ZA0CXbRsBm4GHy6QfRebl4+nHh0Zjc6IwVi7ozt1U4P
amqIpVRpjBLRp4db4KTSrBeHnOI3Ztcgb/30WyBe+gBrXIHm4Ny8BP5iq98j053s
gIYepta9K/D57E0h24Z9IExbnGmhm0H7BaUkPtiGxop5NKgfna6HbaGmoaoXQZK6
e1yiMtD6h89vxzfb8rcBTiFq0smvuCm0vOdlSE4DfnndN5SH/a54vaUZdUuNgD+Y
NZx7vShpx9B6duvp7QQxE8QzRlz0Su8HclCSUEUNzcim4y7rqQJwxxq4eA8W6yVU
nfmcImkTHVUl+kv/dYadsJDg3NDNOtDK1wpybHfwrX1TP9j6x9wNfRN4ko1wOi+V
lrNvyX/JntTADbY1PLpq/8bkUGKuHikk9bDPmRmlq7egmp5fNQLJ+bYz6yBxp3rs
MzvioacoRnPxeSQ9sBQol6zZmq6dGPxxV/aGRYmVvzgv6ztqbm/YQVyvw1v+RPy+
Z6h1jzyMEhjs+Lp9flA6jzxHoSnaOnN/X+Ee/X7gpxgPaCvQ941u1qti7mpPKGYg
Aj5XosCBTvJcVldsYgCJ+SFEeb+Nr0S47ZSHSv2Daw9bC3TUD/LnTNz2PysLS2Ww
IuFYUgobpie+LqjF2VpSsNfP/MvzDKUndzsVu4nd+lL7K9qNMZ+t0AyD1Y7F73CM
7jfn9umFcTcl7nIZehXuD6+StEMXS2S3CaNlRe7mSvhoGSz2GDFI70uziqjQsLka
MXWwmuvtDC4f2xi4x2VjlKh/bkUkm3DrA5wG7eQgrAbLcVU6SVJMzYXOSkDGrqev
CmqyGey8GHZWfWDCDkFXJuCKWhSsOIrqEwZM79FTtEPwQx6h4NBXWweqH2iprEXf
V31qexYxXReuBXEVIGOkwGntnqgjK90MyOfh8zkST6rFc7jLD02OrKXcZl9z88bN
FkoLjyrasRsSv3DeXwnpQXJPVA8E03/t1ioisIEMXQrA+LIJAzhOFLNdH1K6AOX2
rsInZMEHSl/vn+Eqh2PCIrQwfjINz2Ih7iMcKDi6qiU/eHgMQwi2kcf7aG6mdWVH
FJFCGqMsvg0+Sa7G7gdN4HfwR3qFBEnf24v3+UEDqzLgfT7o/J4ZQSd+lRfjeNP3
KxdZzsOp8Ip0pgUBaiF5h73p/VM2dIwddJRzFo7poCv60eOhoGSi+YwmPPENgyt4
TuDEAdUOGmV8uoC5n7Xcc0XtysgkGqkYyFv2ViStSO1DP96hNMPmq5RaI6yxsM0t
ylTWN3NXDkg0J7YJhZaRXM3g6eieqolUM3EevXo9SejXLyMt3rLMpRo3AX32v0JB
+NwG2NwnEn5ukub7eTQ03+vWR1dpMT47GKHaoVkn0ooGwoKpmmFRCz7e/MyVyyll
0ypYrnMZLUbWEsOIExd66rvmXSaULitL0R1YXZ3pjFJ+VL9gdTlBId1vytB386H5
QPeuPsKH6a/HuLUvMtMhUh00y8ZKiAfcxePTHryTEh2PSAIiGNnRDO6tWNAl2/26
riSRcAYIAGW9CfNQTK+BveevJx7YfRR7NgEc2SsOku7YZC5j4uiU4WYfSJBPhL7x
H+KikAVnIO61Fx9aPcW20NRsEScMKWuIC94v5NI59163FABPFO6NZvtLzRQy4b3l
QV1N7J/odCX9COSQ4dvxBzRdhxcYJUP0/fXqBfutllOlF1mMyfK2d1kTAArkTwPk
KVBU9gKNSrw4LgneNAjXoXr0/eRvBpjiL7+sRu8JUoWdEkxZjqjLVBwwTDjW6vWn
b1sSXVaDdS3OCbZot14wMJgrYcCnZOA3wFaHIQNmoCvNNrVTQE6GXwSwzDVuMKQr
dwkdvDStZihQoVzSdY3LrIRBAe0N4iuHXfO5x4xazi30JsTttAODkFUr5XKcZ70J
BmIDFhjtcafUeIwNbbnsPVmwV6Vs6+cGPZchUpeyedNtLskEOXTCigWnVA1hxDcM
3t3PgJs4eEj88bxYujmrIU4+QYWH3L3XGPRniKJH6Pfa4C/P4ur3Lc9GXCl0lGSX
treVxXuEdxc/bw0KdeaJuy5KQmyG3f5hgsisg1S4ZrlmoHCm4GavrV+jRoE4aclk
QH5yWjEzQ1LRDA1G02sxDZvB7Ceo0fTNMjh2ElRmlDFndAeVPGRuxGZ67IYGaOuy
XLwi8Tnne15Jkd1+I3GCt4owCowA6w1Kmz72CcPPKun2hxo2yOSifulLVk8RQ8Rq
t6m2oAhheosjqmAadgWE3nnLuMITF5Don7Sqc7zU7Nsq6FPqpZhk/WUfFFkAqPPA
2ZabtMZFPDKGlgqVEfVYkcbXCzaywGgaN3ql74RhtQCkTCmkQo853CuRBDqLUFwG
CkA+2bSO6l6JB1bFvLvuy6nYo0Vfqw9MsKXMMXg8dAXikK50EvXpqkz2JKTA9Akz
Q38Jml4ctDFZST6TWF8BhckgjZv5OKp7mHJxnOPRtEpKgg1sCZekbwPBZ/P6Kb+1
SuSLn5XvGXlYdg3nQ/V8I9bI1qyuG7/Fr/o5ApcFoWfNSp6M8C0ZizIvvos+Z45T
86lPe04OrKYD27TTe629xj8tSbW75vQOS2Tw6/V03zoLeBVQVwXPgf4Xen9nRR/Y
naCXz0fm1D0dZURKhT65xELBn/nOeQsVfe0pSmU5wiVeD0EeB0A5fWCwbhTLokns
G/P6MFnJz+c5rE3plC+Q0yvu3JuC0XyrZ0BrROaAhQumd64wTUxkEr+flaoAgkNS
Bti+10Rq8AMAr6qk+J53qU8RkG+g5mogfD0GpmtEtYf9+9xK1O8N8RXiysNhC9UV
eE0NFZ0iLCbrk/VMd0rUqWsFoLzBxrnh6ZTqINnngmkAgGwUNNZeg17hpG+I5Ynv
NaADtHLhsZhlrmzf9DWyFU7bOKVvBr/etDz5AQQHvkNWb1wkGAdPEn6JCdF6fuHF
pOH0vAYdtzRY6iwBPljXOllNm79wh2fzMca2c9Ey+ZLV0nKykpvVkXVW+ddI/Tk6
3PN5s9f4VUR5iWOiK/88ZcZdGwNP8Dhmj5jh/Wbyeg64+1Lu7GzxCibO4xJiegKs
RrECsAQihYHgtR+pERq99UCrw7N3KdWADbqqIXiovuupgg9gIWexNcewbpXctEge
Tsirbczabq9S88KTQPPUjdjwDGpZaSlMNZUg7LohtHb23CDprjmO5qCeI2PgVRFN
9secgMGw9RKDPFgCy+3ajIJuUeeef08canFyUVuX3n5Pw0HO7psn2amOgoJfp32j
A8WDookkhc2FcTxECWfsA7vmp3oMdjyCv/IEt5l+KADe8fzh1R3UijPmAaU7JaRZ
w+Nln7zKyspJIDKTrLWX1zxpgjcJrCLvhgpyU6nKlOXF52z57o4SzFJxj6vJn5Ux
Gpb0Cwihtn1KlBcYe6LwiFCm//NtCLeQNDuSUPpM0K4XjgmKaomMiCgRjvjtxEWW
cuYx61NkRolT3kxn9ITkl8CfUTknUK7Rd+uSBswTZ7HWP5H9a0lKz9/TCizxmqrF
qB/qvI4zungBt0qxgZALrj53f3JFZCYIHswglifJxjyu0eLrZxsNUiUIBNjo+q+C
IhVmvMTzRQIkjOvMaOXeVI0VMWxCeo5al3A3wpnAiLHyxQZdZjhNaH7Yjhh3hXmF
FZP0UvMyYBLhh/He7qNsRLa1YQTa0YpGEsbl1EZFn4QAOg4IWX0mQVBAOgQs0Mc8
uMVUo73XeUQhqAsxg4L8EsN9NR0oybGEFYSh35hMjWW3X1JZITCJqLoFKTgLX2sf
QkkUo1ooLhGOw0N+X1IANUh44rYqewOqlEW0V878ku+CLikGpV5U2K+D3jUvjsl8
m5iuotKn3J3kpXULtfVZgY3YJQs93NHwMtqRXJcd3tJQ8kCRiSM3//XTEI4qgCgL
z0mnbMrZkk1w//K/q/ILBsph9qj1Es4UuxgCNXzes3fTfdBMOc50S7lL5faJn2Ef
MASI10Id3BBuvgqQZuAsaKnwqy1cdQCS8ZLKX5u10OQQFh9eSH6TcJPk6A1Nd3En
wGsX+16EYttcEhOKn2dsVqyHrqrzy+tTHnNBe9G3a7xN/1507nIFZe77juLycU67
VfTz6owDJzx//CpEkWpvV3wrXSNj4fBffpx7XZffzd+H6D0dQAwQNMdulem+k8R9
ER8t/3dIicfG8GCeiMfobQRVKTzBQFfspZEzxTX0Xi4pq1qMNiylI7zFsvd4toi9
/laJd5PrjI+Gb3mnL4nz+zBk56rMZ02zIePhcLe8/u1wGcUy0vsPcKrWE0AJrsun
2h1rXP9OM/SB2nJoJSO6ybS7t73fXpLJAlP8e/J0Q7yQ5vFCZ/uFP1UxbKlYe2hc
blvXNavAzgMGM4/Oba59S6Nv0Kxm6x3Y7CVNgzodspWCMKdP67fuY058L9URRIZ3
IYHULNZe3hOHPM9rPvzN6+y6mBRhkGBDDFcblOj75q7OEHFhzuQCzff0zS+2ajD9
50pXX5+ihUDGsXFgOdbHxe1U4AS+Lh29yrIT1sBv3V97DajnYQ5jjmnTDlPBNjwq
Lrh3qHQMrKoXpfigQbRhe5kG7Gm+0Na1UIUTPsgeb5KQdl/Ke1RmDy7o+zFS/t6Z
QNEMOzPzGEoQKWAfaUKZwznTMe6zMnAouTIH/KAyM9O8MHK1XCuc/W2QgNGyMi2W
XvFpWtUdUA/Peah/AyS4IergF5ChlVTOlvWCcxIM0FnHS5ap4IampLJvC63lEtAA
U2J1ZeL8+FDcHG+rzpCUMi6ue3jIyAHc0ZIj/zk42ZSxGU/G6I6/2cmQlTwJMnSf
GY3T1PqQ4+gZnZUum+q6kHryphOtufNYaDARB/zKxk8kHG0qOSTQ+EpJ1PmTbKsR
a6sAp50MIFHqQ4OEXmpR0iOtsgKhjKEiYfVvQstzvKiHi/XtahMqXU5hCbuXvxoU
6lJCpXWoCuLA8PhZO2a7mFHhH0I2CGVGvsnssRN1GlnyHfjloGmkXFhZiEfvlovQ
A+Ie01t+ehdsbzxaZS/EE1j7nknPKFQLNbURR84qeetMZCcciCLFrf9tjczae9Rz
+bbScz9jYqQ/RxtF+o0B8l63pgSIezmhX7+J+WdyoRG3KnqPuwMgQ/fpTw5T8pkg
oX555w93bwESiwPW7gZAUi4RinxNHwbfJMKzLb5+AHxY19S+MQzIoEO4ynuZFRfn
2PV+xmQ2XGGEj9fN0qjD2qNqQU+DQgbq5MxoKUEK7OgiWsfmAeCwy/HheHqh+v+d
piLfnj4JEq3b9GsPgyGGWt9xEdActuWz3/3+PwOe/9xKLddaUpW5xuC5Lix9WAce
KyS99IKYBxYuaY9pwE+YDKJqILhVtRE+tAFZlxMBlGoJqXPS9Y8G5O/ra4Lp/NYE
X2W9nxqCuk75uPtwfuhtqSR1ZGRcMG3dMqtoT9SzOQK8lTPGCeuA5NJgbazJfzvc
pp6rmQgT/cNPzIU7tro8vVVuCaGDaiF/HbPMBjWIWa8ImUiypSu/krlpFFxOBKli
Wb8LhXbibS8ElUMPp0nh6qEdPjfPmN29IKsPh9h7BD6jRAdQYTruUSDvwF/gLJVW
cHFgI74nsVIoSWJiWl7qkV/q7wPjAQdv8id1bEpAsQHGPUMu+ZgPmzN4jirAlMBI
Q45c29tH7w+CdFfI+8T46Z4PUX5F57Qk5uKM7RQ8jtgrqOJvtz6kcK1KT6y/cpS/
k5QdzEJVGCePUnuDggIBrfrP/O3ONjoQxxwYo2C1ptUPDCM07Vc2aIMuy8LljwEI
ceR5dXoaSgFAqRvF1jGpC62ORjCXK6/Gv9q5hg19t+jLMOM2T0T9KZLW+2pAlgKw
Xx14hAr3m/Ktm9MbLBRSuKl6fdeoNCxPzh0hSkZ187G40Q8Nck2xpcZVjonwNbE8
gVeDHCyNfHLnB9t5Le/MI8v7O+KeIF5sy4Pdbku6ansSPHiSmG0labkJe0oeXVGM
IpHeeJajsdYLsNo94Er8+rThD5H69yzBGaiKjZy4pZG4XWmgF8avg8iv1ykF2QFX
HY18q9QjRDgIG/+AI4T3Xur9KEeX3QXwOHsPDHHFEItWpbHdz+24tLjJSiylwBxQ
vPGxNc7AdQIptIVbn4uGJY6u/5k0bHNC6g8uVGlTDnKS1pZZzs5l6dcmH1cmysQf
Y5FM0A5NapxfqbH1QFFkQlGNuZUKz9MaHcj0Er7oi4gMem2gHm2UZJAmpKG/IaSR
Jw46PC8vFjdAK5adyVhkvpGCXqmPH9unKb1JReFvhEJijhjrq6RRCQ5oDF2Nti7A
/nV8lVuecQNe0I43P7GhwCCiPmne2oOmrysq4AC4/ZX5Uz0smxvdQXwmlwvRXIfJ
QrPxodUyeh1qSmJJP2VVe+CP8JaLaPagg9nvIBkJcRAxqxrlRIeTvG28fdJ8Uw+t
2zR054IzMiU5zDsW2teja4ohWvIGM4Edv7LJnmGZ8e8hMAnA17jv9UcSWHs3YIdc
LyN4cdfoQrtvEnsNENs31yvP99hwonCN0Wstbb22ZF6TnUi4DPF+ttdSO3L3O3xh
JY0gl1b7EZjcbmZnhPMCl3XLVqtn+XxNIDy6W00NDcxf06MZ5KReER777fm3w/5D
7E0uRLpNgBh7OctqsRqQgiEhJ9s6LaL3xoEXd22B/ULn9jpqbq+Ba+KSDrZMkfmq
IcNVB10UXzwsvTDeD6Rcbidu1GYWSDInJCW0KfNrcIkLfJq7aRZhPTpKNDlaB3kD
O4ltH+LouZQCTnDjDDqS7RzwLxQvO62f7C1fvAADDzMhhY9r5bYiIRby9pbLQINT
9/tbodx0Xyp3oKy8Ckg4OwyjVye68byOjMG63YURp4t993d5UV0g4hLkTdi8wW4Q
5M7EvBKm9L0cuU4nBd+mu5Ta4csJ5xW2tr2dq4f0wlarWGf7UgIXEl8Qf7dIYdJb
m0uPlsQwfFad/pzV6wtBOn39P7KC1+EIvFO268S3u0svoOmzgh86BPx4CDkboKrB
NkeK5L2k2XQVzDEiOY2XkLKra/QQat+fjYTUWKngLm6Nr5LBWNA5szjPxZyyNb5L
CZDaOCJuqgkBmefwZFcHOBdZ5wHc9O7nI4R+I70acDPzNge8zAI21Kwf76j/4Pn2
P3YuX+E/TbbFSvtKB2SF8SIAU5pCvgLMGEM9BTbU1ZbqTf++G3/4gNjsOHhX25V7
1dpBQ8ydfuPVvxG9itRIVp4RaHVOoAzcyTC/0uB5SGEPwwmC1Sm0bbMsfAGisAnB
wWoI4szk4Ga8B+ORZeeKglS6G0ghEFnY5nJ+84ULSMksvyGJPB0pBVDYKyqelZLA
Euk/E1EqKieLQ03JFeqNPzTnM5kjzPuxAPElUETdNHKXz9fgVkJpJ0pTp7an51fG
mENkKwGUHnae7DkK1OYVdn7XvS+hPIOl/Go0TU2tiobhsp7vVXfgeUkx9/u5v23W
43OtqOe39i7CgjkMGEIFNdSVTh0AQ/6t32+hX/lx6A0rLfWY+FGzfvkMbG5mioa6
PlHPX3tamS6TJxgZOPymh7XU5pW3FPTSr2/7NmwEosYg8xxUAuHzFEEGZ2lSc+0v
8dzfEgxdxGd+uymuezlfByH3bdCU4MUGoPPEIIJoW+6IiuHkUNKjTXi+l5X/WGJ7
EHnANQ+R5kxbx9vjHFh21R7NahundjxPm48iXjS+Yx2yPyFFnxBt7Qkf+x/m+2pC
30EQEfoJ68CYFW6DVSO+ZxvtNJ3ZbNZrpvuT2vXaDK8jkka1EhSp035PTUkvX8zL
PLqOSOs/N7WNs38xqJhtqqIimskqHJVLSl96ld7D+XNHYuBG+o4n2Rnke78Nr0x6
SQYUxUymXc+aMGP0kTDXmtIJSVM5YjTJpcyl3dh7jpe+4SkzLlCn3C7JGHCdDWSk
5Qui22UHOSIMstn5FqpJ9iamMjQtIPXGhua3wayAdpth+/OCTrGGcXA75Ij81B3+
dkbd7pNYuOEDejzSsIlOV1voc2pZLID5mQZaD/seKWDzcel6hgqRRBbFQMP8JflS
tR8hWLD7jgHGaX2mMUtW8ci/8RqviHk44IiK/1nwv23CAHfH3l9GA/UItv2T0Emd
KVaqGA01mqE4zOq1y89Rp3p8yjZm5XDXeJFzSZTnknTiSU/uedOn9g/KK+VeFJPg
NUPIGIXNopCr4JjcWUqP5B0DHcO1QL2nRFkYGLp78lUFfT/l+gCgZVeyxKbjIoBP
Idb3VNFSNwV0lt7yrqGtkGU/nm4LgHDJqSw4GI31wpm770Cnahc74Nvq4QbtwEwC
MED/WTuatohE14s6s7x90jogAy4R4vxUReUQd1byiTsWnFBxgaS3isIB6bgGuMPg
YnoeVIkJzLwkHcwTUJYkmmH0u4VJvSEkAsodRlulEPhY5aZxOYq9AIa8osUgOyLX
mChVGLgH9M6RJu6iRB/lVmruCV0C0Exl7MNX9cMvWoTfM8FxmfCd7zWemiSSqFSB
0jTHnuIv9gNb5Ip+jJTjjF1XpgVcmqVZ4sBdPUPGEcRd+oglM989gOml2lYoyc1W
bJa+S0Qcm3vxl1w2YXyJthq43BC3YxM+ngQEkJYPZaQxt+HzTEZWk7+YEoFdHD8E
RoDHwghCg7VrxLP8aBC4mEcAnb+zs5CkbHmSnLQ5ZK3ume3H0f2rgrOLem/UAy6w
fJJJuEdyDAf0VmuzyTvv2jXYm7ryCKwUGACjzDjlcKF1gcZdxZ3XvdHkPhdBsIy8
vT/Z1uZj7bAyyp74XXDzZd5OT/gJfdbT9kJKjAVDClYmw0kc7SqvnEQPD3LsEUIm
sv3/2PstM2QCg2Ts3l1v/bLq6TYbGkLlN8Rv+cBW4H0wh5XTkP/ceg8CxGxujNMO
eFR1e4VmTp0vB3qW6z6j0ERmB3ndh/QsgKE92ee4WySE+dhCdxDN4rHFgsxcBmuI
BR51mNbZ3sqaf/ZZB5pvnJACG6oXg3xfow9VExnvhCy+9E6oRW7DyOTdDqfaksYn
2UQEqmUVX3My0KtVyFJ+q4CFFH2xLAZe2Rr/8kF9tv7iYQgs9CqnFX2XA62Vn3P9
gCR92MbbDzWLll/5JC4sL7bYIPsPREheL1+fSBX7xoavFFAI1EvIeoFnWQxNsA9E
z6PdQBGrs7AEbp/oSPKaPjm1KtGq/eOPNPAcpjs24+DukIQPjg9ZbnhDJDBAEDS6
nmtrQvztC4JlbuuGC4UUxK5hytUkWu5skkxOLFaIAKiQpy4oguulHHFncGJjIwDf
xMIQaEVroW9vD/XFvGh4xoHV31Fg7Gr6JhUKe5NDckAQAce5FfXUL3+aaxCwDpWj
N8RaQo8bEdTDV1P5C1Z6poioek3R/b7gGgl6AaZ056GQB/k3Ow1uZC5NH8BJdej7
GtMW84CbOxTlSZioCuXMfLp2nc+f5Y1YUtloVsqxg5TsDobSZYaUZAPtOqA7xbAj
7gqqRQEi6MGUkbW9q94c+JqVVjTShhGoeEGuLu6f4vgK99FsyYEW8wZw1Zbzxh4X
qiF05ypYnZxxWx5OMP3JlQTn5i/Xui/EvtJY4fl+qo1lYiHMDinJtCMv9TNJing1
b8cmOfp9XK6Hv/9Ws/d5pMpO7TjohM5bZI7iWMALBMhFoXIqh3mEFGxq3w+mZL/P
Tc4ldDReqeO9SZhVNBsenSPu5zPiddhTPCVAXLEP0FzRPyluEaSEgBGKeKkny5xH
g0KBFBADIIxfUj6+bw364yo+tMwKxKJWgYxkIEibAWusMfBt5kcrH3UNTrVQZzG7
4mYZHPPfb693lPKYqpNVaMAYiaCL9Li/zaTA/URV+vjhWJx2ocJJswArt+/9nxa+
of0/oCdumnqhPqUdnr//xS2sant6QnrcyioqMgg+0NkyJJQ2QQHm/l5LLH+HijIg
bbA/sJKCpO4qaeQ4H66y5YzU5rI+MdaOp01XiWJ1KXShouoW9lZNH5zZgf+YdHvu
qx/20uUmjcdJkciDP6REo0JvXlWnVZueNjylgdqERRrhxoalbeV3Wwd0TxuLSr3g
FeX5fpa76ikrHpj8ExDaIyQ3SZ7DAwK5T+cqK/4iOdChb3WbXkhSm3et0AOd3kEz
6mgiKMt21gJYb1XR8iI4thTRrLhbZjPiLqw0W8mEYvFBTgBhLG18+iBrVrTrXdSq
aZpx76BmeXazHclS2P8zCgYsjKahYOyKC8bZvI5+EbTS6CbAnuZLNnEpdojuBb5f
ZmariuzwoAW2OWdo77nyWjbh5oU4mRTEUKwW7C8x1su3/yQvqngiFihsOY9HYRjp
LYtnC5jtXqlq4LKl16eWRJABGFxKwCHWHXN0tH2w/Hq5MlMk3myiz6VeloUJO+OK
Tjga+Q0ffqew74JDJ5Vy0XCeZ+GvADaNpST6taJ6ZJZJVvmiVEEZC5SMv8qHoM9u
CEScB25FZ9HySHRZTjMyL1bDxT6k/KBFukMnE5/Sj5+nM/U1Vo/RrEJft+IqyI3z
M2hdB4OEhlNk5bRn7v8dB+IbTl9Bh6ZKeLPhY6hDfi9+0dGIo0hh9iVARcs8oeER
ug4ufJ47nIjG5FO4+IcxQ/18fsJUln7va5ZeKe9R5xC0pI+uo5d5oWW5SXh4+CsA
BgVvyHMnLE5a/OONSAIVoCDmQE16cYDHkNZHUjpQxbEGIckr7XTOVkvamwcd6q96
mtFampcc9RwtDaYciec3ZDcc4Bx4k/qCqjITrVEg7OxvZyUFt+tYnQJdkw9eVOCd
tpljZFYzDRy2IkUraFA43euYBehfalKTIInE12+LW+A8gnV5tPLPxTLkhn7cfIhK
MOcXOUftxhXZtydzYwB8HBJhluPClObUdnCJbxGDpVSr1C0wR4mQpITqDal0Dc4/
9h78j1i0hh5MjMwDcDhy1l0oKQhkOT3IW4vQCNvjl6xSEG+T3lc8aXJ+KFinKC+f
49Z6HN016dC3iL6aNc+kzFXXU5YRfEuE+0ke5jkK/Aib2JSNKqjPn11q2qcBhrfu
mTIDDOjiCVA8kvfQZM8Ex0HVuiWy2mHLnicBRqL8KZT7CQ+2TFgVklHBqs0jOC5Q
VmeVB0meqru6do0Orkyi1fhhmGoA5l0Xvb53yPLP6cxoZ4INr996UmTBy6QEW4Pr
EUbn29SB/xuTIUWp9di/EoFbs7pHZ1f0CPVAx77kSPHveVJQ6u+FP07bK09hlAV4
D4yyuufTdKCmMI/VD22Ml0x3nMBcez7kxrlI/UZ9nOkwm7kkDkIy3np9pc+NkY/V
MngRcfl+DRP5oOvBMC34ZFR+sviPWiURmYXDqlhXS1ZmqyuFOMLJyVg2zh1/p8Lz
eJcLRf/jaR6nPjAmduLaf5L5Uo7mkovQR9BF6bJpehLFu/G2Q+umLlHumHsmmukg
crfNkZIle9kyNo2KEf/mMs4mvL0BqhZzlI7uXSDrmH7Y2bxcU49aqbDVY3McuJ6A
yWTCbN08X7YiABKpd1SRA40z52AtBffVa9mUGIE2RQxl8ms+NDvknSavZsKkYMJr
8J0b0684hTXg5YhZA3V5gkdq/bwZlxco+GoYF5PCXVMVgFAT9vt8FSaCyHAQBrzX
XLRPrnvkTcpEyZKBa57ulFSgGpZ7sKVeIlR5QqFnv+IOd/d39kysr2egOBR+zWwu
KlR71fMH/pMFfpN5EYIVRKTVDmWfOr3UpxVDK3Shndhj5lcCdNBVvBooKQTn3aQ7
LF3oPdIBsI3drUIP4GjVVc8GVKvpYsEF/zCwWH1BbfT2UJp1+zvJ46cgY7USmqSl
eISfASkJ1pAvdMFQBkIGSDpPvwf0kukh9NoCJMfM5E27qNLIyIIk3NtNocBnyYXB
CaFMgpvDK5LZToxc7GKSjRUatGpeobu0qIMkyn47MgqklXCe0rjcmZoH7kQLEJdc
4afqcxdTXc1ItoVWK5CgXSAY1+TQvN0k5CyZVaSdsyi82e7C5DtaHsN8uqoMpiko
Glr5f8OT1FTkXJylEjZlbsU3FL4Kn0o7I7MahE8K8VXsonXgVPdCPJO507e+peA0
P2ATTnKikEFfDSJgAJ9N54z+UMqICvfTFOLdEbxvp+2XjFzbn6Rqyh0FiGqh3ypc
LHZe22DP4Hw6H7aZtnpHqQnfFutPkn4zo1G8k2MbsEctH/mDevHPqdNzLY7itUb3
Wp626HV+2oPLwYGkxD9LcJcuSpT3/SScthkTn5wxSfiYOJeCP01dZ0j+DymWJ2Hx
DICI7xjF/5sMbsXO/R+7KgqAf0s8gtFzuY/MLj9axxYxl+gwQfCN5VVKJcfXvct0
gLDiz+0N6oXZhByKARnzvtR6q8+AzNtK6Noh8lTSn39T1Vlk1uFPvReBj68vaLIZ
aexeL+tHLaT991da7ayW1YBqMg5KNTfGyOBqODMASRG505jAXyqywSIccFKHR7/8
+BpcwLzL4D7H6sHmSITzFnQ2FvYy+TuRKhawrCBQxr8xV/nIMQXyss0JktXnnwIA
I7DrCNYMS8gtO0Q9HeSjn8aFD96crnAmDEMzrheF8Kok10pZJR6ZwOD8+L+6UJZ5
1R6BozG0x3JK59NtMb2uZP8r0SBh+yYy/4U93CSu3DW40AXIOO7uz+PT8dw9zw8t
lkkgQkPaaPyJCkax7ZI9idZZ08n2YeJePsDKS/38Oz3GypMrwOIBU1z+nhwOcQoD
mnsyASiFaxBWYdii1Hcv6TnhR59LQqyjKQ7Od+jl04IsB2ti0nnzT/DtooxCyKOb
yHfQx03Z0z5iYbbOnT9xBAjMOBUIF/Xw6hs4F9RLid7jaKGDeEeCk3hsuYjF6gGt
QMWVjXaQ3ZfnqoZeB8vj2TaVYVpOPqRlN7MlQBx4Dq/Q+GD8c+4UXQ7253R1CB/M
M+GiY5u4ptWtEmLxov5tKG312Vf1rZVCGIcEj1sNpG2scq2XVkGUvTUBMpnpCZJI
HziplFYqOOl6/Y7Oj+TWJM77YY2BIOk6Pev5YfVi2oEmfDyYfLaQW00LJ7lSIKbN
Eb2hnsgFMYuUai0MEafTdcDPhyYR9vVcmrWqFKq57/U59RUr0D0cAYX+GcJ7ImTP
C2WjY3mvTGTBdG8ZDyyv62tqgQo7UbIrs1DUxpMnEdCXumq+gtH8IG5POkzY4TQH
Fx8ZAynn7pI1WVOf6SU5coNvVCN1N7nif1AGd+8Nqev+UfyenqhcuVHg05ksmTQa
xD5LkyDzI3D97icJae7I5y6A6PlBpLt66+jMOMbsl/MDat7wdFNuwX8bdGvLIwPR
Pa6xsDY8dOIujga/ANNoQ9I5GgZ1KLZ4DoUb14qtMYCyje8fMFNo3d3DqpcmpcBw
m+mYzutPkF6CIqa6fY+oLFx3XlXj2CV9/FOHfhD3SaEPO29322GRY1nwLSPv9+eL
Z+GnzRHTfpNMJai/4pA3drrMN2qlDwlK8Zw1vNyn9X0GoSXtJjmJqHXX1vd/q78X
JVp2cX9P6iUbfzVWPiFSaW+EfHgjSOQVFnv2uq1dOF2CJmx2kpaCUcT8ajy9dPFm
/pHZBTvi+caGrmaBwd8hRwFftCKl2+QyYC0n/0zNdEElf8zqorNBQ2xZnjuY7bgg
xOwyIr1DXjJF2+OTBp2F7ZbvJhGyi4YVbXEYZ9bcHuxuxXm5qFmqvxs6zPhu5IaK
fathFon4EAk2gtnGGmRnq5zMVmoTqpGgSpUWtpSWHXCxG0aKI7Ii/nlUu2jVof0w
2k4o0sT/HB1sDdDLPbZQAndZXpsVS7vKNtFS4eqvfB7J3jJcdQ7DvgOuuqAfiTSC
v/CH8qongaHksd/ivRjYVD97ML51T2c8GkXfOnVWeSsLWz5xTNbmfaORL5RSJ29r
YSAtVhK6LxZpQHwiXuzjb5Os6NEGE3GnuzELNofex8vq0D3ROlUay4ao8+q/niU3
qKLWLevK/OKAwAqqIsQB1aIgUlWcQPZ0IMh9vRQ0kATCTqSNYndQXm22o92uFoH7
pGJNt0l8cVtH0Imp8NnXLX7pkcFjktTkmpVNHB5i0zniwrlEGzVn60tKsaPrGMMT
yjHLAzMxSj1oO2Rtdyhs0KXjIK5hOlnUYF6o9iZHQk3nHl/VDVQGvUfzcV+uh0B8
FqQnXkBbkNA58M+SCO0vhEGd7iyhWm+610dhoXzYyw5ha1yAWGPNj6TAUoySWsHh
ENXOaBPDOPoLq2LtY/zSxUpZ6ILkXlOe5LB9uuN2Aq0i0CW8CQiA6KfObJYFHdpM
0sZofLTJg31civC8IDJKs6MhWjsy7dDnapdfX4KTCtwFCtSrR3BCjT3ZPeIsJneA
kaaZPdtJrKRpCHzLNH/BtHGKyUhnpzRGoXX8wXqclAhscPV1AawqURD5zvrhJZxN
GRtdjMhsL/+LO2Uv5rYrM8HVyf8aS8JMXD3Wxpkk/gJcN9Qz1fvGMfvnivftdtZE
Yf7+peVgiFRxR1GW4k1ummua2GhfpMkNM1Xz631KrehD1Ik4+xG29oR0bhr4mVB9
QOzaTJzsEFTMDiqkoFDfTRmIoPvhYJXJM22NooGfq9bLeFDxXFVp7YgnQow/rg5x
w3W3x2GeLvKl2vLzvMtqSc/9NnTNz8LWwGR/Dh5QopYGZNGtM1zx6MHiAhK+u+bM
iUJHSWq1TmkSgBwHIzX8gL+pkahS7IKXAAn3Cg2/oH4BXSENJwzwJrNe8ltr/kVc
AQgQWpds9n4Q+yD9HI4HHeR74Q0dxNg0rCc1ePUeP9x5vKvlpOj21USqnjPNTyoq
Em8td9BPTexEojy8++nyKXeOWeu6QpDof4cLLICxmlGuifIaPFIX5KXf8LRlkT0B
C2Oha6X9/Q8TqCZBJyhMZOZJibesJUM/aBjAF1QoC1exGI9fJXTlkaKs8XdM6Ugm
Spv7FM55FcGZyWznA5vDK/vuVgrajlxL8ex8tYgg8FW8iVheVqV03XFo3ro9eRti
jxO9JCfeIFeIoBdcZOWMgqujGhkHI6/LOAePZNfMrFARL1rXx3Jq1AL9NITbDQvk
1Z2FJ46a03JGv2GFRl3IQ3iD+AJuecrM649XhQuueKLGrN/ARCG3rx4Dog+9MuNP
kNe+CBNrcZDPqgCcpGQS5mBhcAQRFNJz58dlNwhzYbhKBMgZVyDYypVJAi69963w
sVWo+bgNJ7mMD9abQmFzSa9sdk0gy6JL7G8Qc3gc6Q2gHeqXL1nxjnMDMwrBUS0j
wXuQs91/LemWAb3B0AcbwnJkabgC6jHsXfqiEiGlj/LiZs4+HDZWAh3CqXfobe3e
zVLlUU4bnhhB9XO10u85RVX/5Cec4wKt5ZHnJH8AROza0v5iKa10c4LRaqgOUrKs
N+YzkiQcY0wD6SLfFD2vhq3VSl0fUCFVw204bgcsViKetTh/jgyDkY3scdoFSXP9
zeKKOYqKC+fOSqxdX3V7+HRMHcPClRP5mkkb0TDh3QwStuiDHEdl1JNU1n0Ibkya
F3JM7EgsvqAm+jiRfncD5ss5pQYaNTqRk7RcT+C9gvrOcR5eE0d5hlodPhGajUyZ
9AF0z1nFq4/H2m85jLQySZAw1slkoPmqNdNIb6eztLV775nH7HJ0+F6RdUz/IjAK
yL0WaCO15kPuJHzHrO0cjIoTS404XHtC73JXWpqSELsgS+/L9d3VefQVdAS7Z0Hh
JNcYQ6/dcvIa2FJ/L558FkA2kKgZ345Eo+u4gxigNi4c4ytilhEANvCRIXlFCwEN
9tSjCLmV7ydnMqPGCkjWL5EBBDH8iVPuqqQ0dVenuRtX5ry6bK5defG8nebBJvTt
YbYOdYTMb8QCN8VzMnIAu7+GpYEl8YV9GZwU4Q3lVUwiXqLoZOKTBqNH2rc+K7s1
/+Mr32+sA2mpwAuv6eYc4u9v7MM+mmRu3PWDamn/XuNHTEbAfB66IdLS+UZsfz3V
ZXKFjhu8htNzWHvQssllB3uc+AiNH7I/yq2/3rPl7Tb57FeDlp9Q8m5+8Nh4e5vO
xEwpghoUuzJVL8tYnA1/M1ay0j/7Z8GgbreOFwrTHamOB7srgaFDgeDAO7k9Td+K
EvXEP9F65bYH65U7LK3ig7eIryMXlKzqXAcFE43Cr1tMRyNys9P2e0ST/Yc3c9Tl
ANQPyKCTvoiprpmU9ymkn8V6mXMTQx680q7XoMWrLs0ZRZRx9Be200/hQPTLG5yL
Cl2JCR7fhMhJNh6BM/8s/VyJKSLzqg7SJUXMFGtBtLrXv47P7Sl1JCD9qwqOhZU3
Abcy77vkSvfs94DRYzrtFVcXmq+0v0W6EVqmErfvR7Dl+djwJkzsQB0IyeOa/ZZL
Sn7fjsm4AqOsbs5ztdvPp7Pu/mCDjZUj3i6L6reqOIrlqrEmMAPOkKrcbzyaBj0D
4NllPUIjeRtezPSktGeSoKDT5XQ+t7dxXAW/hG6sz1H7xJjszzp2atK7l4hrSsvP
HIQg4l+4XmucsxapO7MO3RC0uWXVaKLW7mjz/nKKopZq2ILtLaXzhIPx2oe3dNrB
GA84CilF+k8w0KUXaQzWVVwA9NjHPa0U1Kh8DJLUxbl9slTjALWr/lO2MjFE7IV0
rfmm05Ay28r85wMRUXYi8FgYaEwNK/f+uOwRXzCH5GbQdjth/9/hRvoCvcBNRQhk
TUSn9c2gSAcLNz9WZxw5Znm1K2PhTDzmD3ko1oQS/YbT2RG7Qg0UC4GqFN6sHEaB
no0sm0glhDOYUKNGmiIDkv+CCboxkxJQ/X9qr7mHkT3eq/CAJMlV8nAiGwHREWOd
K4t1mRpsH5s1S5KlOenEjyVaT0WUALTRT35mp2bZCMc9E3uSgBKWsx/ye9VpTvhx
lVmswq3D8OOyg1M/cvAv+b8CxcHYwjj7wQt0OqL0oI35djuAXi5Jlaa9lXOKOxuW
MYIuSIm6Vhwz0KjDfAKS+pzUyfRI8Fjd5eT4bzhtww5tWovXvAJxvcSFEqhKdBch
6Y+jx/kDOVzEjXqiPiQ0YZOovHJwM0b4ciQ3obqZFPePbJ2xSFSvcY9D79OTM9TS
0qmUPW88Al2QP7aTyrUfWR7KdgIeiBGG3Oat2C07xj96yf5EGSBorv26aXTx+ybh
Xl1K/bdUYDJdgWi90Qy63TUsIfXLSVC9+9neiDtfRMpYa9SPm8i2yXVtFiyb/iFy
AaaoNLZg/YFER/76i17f9jzziQvzLYylURoesdfz90ZOamz3njipPx6O4PBOgHGI
iIwInuK/80REDFjmtj0hpJfWqiskEXAw5z/zhfHkqSbAtnNdfoG8H3szSjAxDr4w
VQqi8hbLHQZgPHor1/HO/8UD8x/wzzM7d/tPTmYboxRd34dC4xw3w8KSM3UAj5xz
nFsDT6beu6mT3mPc5C5WXWwMuyFb8YrKeCMX/3DniClZfP3PcXW8cqzKVhWcY4zW
qNAUqwoE/fOzliL4YZbvv4/n4ahIvFMp4sKYKSe7koNi1TK4wqA5pRKMaWKsfhkY
2lCruq5GZCAU1EvGOmB/RpuWIfwZ+o5fq4zEkVcj/tdsklka38BRpmKAWe388D01
J8Iurb4zWkC1W6W0RLa0sQYTdCeIcYaaAwkvjE+09q8ngdi555s3lccxDF43l4jw
ZBTj6cQNKJboQvuXruHKi34p3g1QP2Wk7Rxb5Mkz2lCA0/DbOJgREdZsYh+dgjbq
TBCAsjxGA/EiTNNosuO0PYAWHbIzRtKgKTmorfRjktMkn7rMGkZmVFr6TZYwMp4a
mk7EmBD3194EnzWRHEKPkAHoGzWI/6IGOtaujPwMPwOiURrOdHI9NxKPqU/tce9l
3P0IAi5Ymgdtk5l111U7UEFE8XuZQoX+C6Hrz+E8zazz5zKrzGItdjqvSEJBH63z
I3tUq6PyxZO8Zta7UEFAKas5tAne6CH+s/NX/PR3zCbzupFyK/fRoDorN5HqfP0U
vAigi8t6Erk86N9Ly4ICG6YK+a5qgYhlvfX8I2gVK/Bt3Tf3Lm7tXhIByQbDICGS
CeJB2sCeb288LjH7Z6P8os1wHzXIEVGOjHcox5s8hn9rZ6pK03oD5Os+BhCcaiKX
69jOLrwiZu0pYlO2+dkvyVwVZfbYs31U6v/idOcSY6WY7C1QtrJLEOr6tsAemLLD
SgACSylRwL/DvIB5/+7tW9DKVAS5R8KKiRqEINdgLacQVKsQvOL0jBhzYY43CoiG
zaX3nFaKDxSOC+VwybUXD28rB3Vww0+0sII7hLZx7oFVc98psB5pcHX4AeDSmyAQ
G6oN0TTly27IJnqUctI6XIA4suLt0MQEqSGYx7BmN/v9EKExy7O4F8PqAnZuyHhW
hv7kjwGX2Bp0i+lSCeLiGVgVlaI0oEx1glKWQ6sIAHfMwRvi0ck0DyDhO3gge9s9
lUCcvX5J2C1EbjQG0fw6DWx+aQM0Vm0mwQlGlB+AbnYKXn+Dpu+lF8yzuDlOOI8M
7UywM0OnZRZ84V7BttiyNny+ioFeLMS1MCU7xQOKPQ9pMoYNZqfTfGZCJUW7xA6y
VCuVUGt/jKVLiDZjfpGk0QOoXXMdl0kQfcRyI1QUIcSyd8IcXWnphEivBdPYL6oo
E31gYaPn42i/4toUngXTw2Fn9CsYc95nVs5ow9I1ZKHkWbYzrkdLYHVmzgPn6Y8E
dunh4MHWCH+ah7uHkpdtEvPtfEbP4UBNDyfdyS27/5fSoyWeIr/IbP+zOz1sqkDz
PTBXBTbuQn1NM0Wg/jHnq/u9aU/LuTjwlZpktscgNbLNw/3HwwdA6A8YoBJQwOux
XRMJALzLSTEfFv12eNOPzyrCYK4vZO+kWyYpJTqY8J0L6rcOznuk6QJaVUW13TSs
Gbyoq1zxMY7WJAXyW3bbdGKIPJUg7CvA4hc5H4wQ+2B3KpDT5ZM179Ij+wM+2l05
Lbdwkgw8Q8vOf3J8PAZPn6/ToOHEOLr+Ro68cNuoKIYN0h1McAqpZGgHKJNP3eSd
H5Ot5zXbarn/bxGjhEedxdo7M3n5kTs3qgJtcAnHdRQbdJLj8h8XHovu+IikTlfB
skPjvc04hZBZBwYYep9QEL6X+Mnch5dQMnqfDVeFEpO7Wbf+5Ss3gh7MhpjlUFYl
QItu2/XFOJE3L67hQXd/a1p4NXpgjKURe3v7dnB0PfEyUhif1q+6JQA/7VGKilGa
gmQXPpo3agfdAxHnQKViG2/YyhjqPOf8w11oUGG1hTJ+3aqs/bJDZTMNxTTILEwT
cwEJ+vX+HiA2XBmX0mDMOPEHIfveb+qtDA6HZmDejiadN4w7uXEgirO1nXKqdRl5
jxlhHEfZwpRMpq3Vd+Q71g72qIb6HBG7S/MZUP3lTT3jO1PJ18LugvPwLRL9kfii
+fTmoReyit4qvJS/iXYppItIqLZw9fui4u2oQpgjQ3YWVOx/FXBfsSgxo5wreTEx
aoNQl3iMHQwwWk4yp0vPX7aMdeenWuhMMeSVCaaXTIkCbQF7uT5Lsp0krV/3/Xtf
4lp6k6gr5ENfCIeu3pBkY2i7fyeRSk9flSF12aMl1eKeLk5scqjvKFGxgLcW0zTO
PKvIexCt0LA985/3bKpHQGznYR2Q3H0db4LfrAhZGd3kMGfS46ZsL+593sUyTOyy
Iln0CmH5i/TpdiUrLZ9X9bc75VE+cBYN2kIM8VPzjb/PKIzLRur4Sj4+aSPx/lc+
O6/zld6OWmw3oSoDD1j2aM4+L6hjdyUixdciLURVq2S/hGlAydxLee0O28OWFu/P
iCj5f1GwUTN61rwmaC2Zy9tR70nI9GNR6B88tCd3f2U+n0BuzP5wXs09sLQrxXjS
INucttsliaX2yx34UCh27M2gwSdi7agURZ0mK96hRcjeshZ/ga72VZIs0BkHYdx/
gnZTzdfDcykeNcBZ1MN/D5xa5EEmyKKRnyoccNzzJK+noQ/KGi+T7CEOE9RX3Inq
LRFqcrN+OO7XYKAlfCOT7IuUGi6m+OnK7k7g6weUphqYCt3eyEAenscKcAeVGBEG
u66vfEq1R4cjN2AFdEL7DV7O0QWJWKjA/xdTZlAcUlcn3V430jyi/rxBkKqaHOIz
S17OhRDim43HpEG1ImkYCCh70l51NfwOVXnysjkMgRcn+jAbyI2eUI31/f7hNo5A
2A68Wigv4A5yTpmJLmqwuEm9JM2sdRvNK0n8B7K0i+uY4Q2v1Osi3QtsAp2P4WOU
Ktw6H8NfsUxqN5mWO4A3RpFT63KKkyQALqxEiyur24I8lFH7V0PLL9TsQfn/kPBN
nQ4uCRHp5UNIN7H9lpCGjYuH2hI517MLoQArwAvqmluJQrjP4IKz1sEG13xDPfER
xdCOF+t61m/3KMM48c5/pOpUA9u1qJMSg0THJNGtYwMdeZoOPuuv4IzScb1Z6hhe
gwxVceH+W8CCXCey4ccRmJFP/aXMr9LrzTi117OGiMZSns8g2+55jcNi+fQpL065
Rh9UgNTYdqL0uuxv+KFMQPk5YOCWxWAvGvLf819DMCDHQtlb5HwdOueFsrAWVw44
Tjixp01mJl8kpv1R9ep+6L9iWSazhjcoOXzlJ+YWLMYpR0YCWEqto8j8qs15UrFc
85k6J6NGaA0osahy2enzt6B11vJb5Ycr9ViMhuWKc6EyoLHKv2ObsUxc1YN3NTrq
AXjiLgkBZjJDtp4ibxYNpGMDHylK8iBGVBJS2bKu9LjuoxxYSBeS0eymJFPjF713
BkMhlQd9xxDFY2Cp4JanvPr6diPM33ZGwYblStpmtBS4fLOXeHYBG706EqAHt0a6
8z2fWSw8eqwdVq7yUmTTtBQeRDZ2cplf7+PRGErMZzoPMpeU4jPETYeotdO4XPxP
HLSqXv+pV76ipalFntG6OS4mPBf6pkFJojmVJqW5tF372LJ/pFCDJ4FczGzkg1m6
3TQMcQlfE23LBmql7grLCgyS6OHlpMuKny7MEnDECRuzizabu5cE40nl4RjYj5Eo
T19r/eh49AwdPmpe7y3jPwm/VC1TGZbES2+IyeKOh0d7/8p0VYfJJrhgbF5KbzW0
IaR/sc/PdE5xisy+u0kDUmHkk+SE/66ePZL17JEnd40vgmi8pWPZ+s/Uy6NPSfZA
nFMwnEZZmKrcXzuFkS5isBYg7UkIHLw7vsp2W07iwC8I+NAq3Rh3wPd3N7uEDodO
Iep9sQWgeCfEnQM4eH/wsa0r4LQ03XGmqaJ8cSmWbXReuDoqCQkAcYyn7cUVXfAp
xs0A46DP/PrKhsad+x7YoC9N7Ysk5KN8412no7Ap/0Q/+6Vw7E/vU38HIy7pEIhi
+MWO23Cf+f/y400M4P08a4MRb8J9AzETvZ/dmfUeDMgpWp7xpIlZQKu/mfW/v60w
nInYeygCSy9elAAIv0kSEO58hG1s9WeZgQoyqHRGQ75Jgnf03ieABMiETem42pHx
enuJ2U8SDfuR9YLMij7KVoctofcQxSDcaIXV8cruFpyDbQwHHq2nhdM8Le+miYp0
fvONnpca7MzgtnBNlVNi6m1E4niNJ65ccTNX+UYvO2mdlctkBIYh8D53zlApxlbO
wWVQ7UClZaulvmMkXl9mc6qgPIeD24fb0vJLVNLlf1A3cTyEjQHOq2FFcphdr//W
k7Usx/M3yhOZrltAl7UeutME7y9h3D5pqxvkPt2066Z0FuxCuxq+Jo77z0Lfy/lY
vrHONIVETQ3lme2HbZlKWLaFyCfeB+XzkgTa9+hTCAwtGzDQ931KAIc7LXjOCvy4
wrq5m0vJuQdPF/OXuOMXY4aVOHSy+PaJxPscwnTCVFHg1qrQ+6AcCxKfE5AZT7tQ
ZNVzLoZHoT6x/FmzrK8aDNiBkjCsp5SGMn/GOba40WO7OnWz929bifM1QPK3EAKu
mta9Xwt4Mlazo2n+snTH2GPql85CgfdBD7feYZSh5o/gKQLXu0TpAWill2IokufK
VFo2WPV+j/8zNePZ8pGCuxe8T830krojpl5CSWLwKgB4V59rdXx4F65+roKj3a7d
PVNJZL+CJlwpRgyLyKHh2XlbeHVRgZbUvcNalOQLddlPVmH96bQPwE1VvgK7Kfae
m6Q1YLnNuq9QMj7GjAq6TZaOOTS+9hF4aN6o2cfp4NXjjh/5jiT8kQxP0P183sWt
j4HOdSWXf9jwpfbK+YMVfaMsWIY7RSrAGb8u56BBlrCWoizDUMUHGW9LIQDA8lze
RBbqHwzGtrXtNOi7qeXqXNyq46Vr0krmR9cXRxuaDoE0xW3lJf9sLoc1YEYX2wnr
CLaURzlQbvo0uWHtb3HlFsKJNaWbP72ROpmQ/P55Br1siLcqyl473XnEbuLyvzMw
h0WnYJ7YXhU5f7Rp12Szx/I6UV8HOIoj0Umz/39zUfNmNgTifgsk09jr4uTihtvj
pwMI7o+NI1aI6k1toAa/FAO3GCKx8Ie+MZBLk77zFgTuims53gMuge0CrpopTs+v
dz4b0d7LS0sT9L8vOd+CFfPjSiea0pD24s/vPKhJquxVZxEFv1SBj/R00R9vnqUY
sVDNsDA/XrwwkqikJUM6Q7NBjH+K8AOxY+sdU5xqta9cFGjDt9h0FHEwekcpjZW9
ZWV8AcbM69N9qO8O9X8B6yKJF2AeRU99R9MuT3ca0PbGPxQ/gdZMhAbqNq78vQ91
1nfdfejBwWpIzrAsmOh9FZ72HAfzEz0NSQ3/O6bY/CZeN/01YlTlpR7wfsO+CHIH
5G5j6IpTe9Srt1LCFrQrbJ3+hc2kGv33jamfgESohw/UmtCtZaFM+E/w25VkNN/M
Ky3IzOm9ynELLmrEc1zXJVFKoVT03VBdhEKjL7PnqYyo4FMgYBJQDojwG7F9A8UK
rV+AtfpSrmGESXXgkTCnDlilQVnXs28rWHvYMNQWiqBbXZnfJyRP/ETt8R8I63sF
Y2leXI6N1QfH4wH0IfN7nnX+h57+SZ19TVFOcIHKw//4Y/+02Hzpomk2D9pCx0sh
8soI2gya2/pSt9LsoXvFBOdcGelWXEJ8uaC7idTtPCHn6YnUdPQnMr45Ofc7zC77
+vjCE6l58cuS8wqvrS7iUGTd3jsp+en/M45yyhiZre4f5rIQJRn5Uy/DznGNg/dt
s2fqoZpq79kqaROTxBnu4a53KokLc/vt5U7WaGBxHIXcR2BHlqPT0n97AKLF9XKg
DS1WI4C0Cz5CIceGFE+UzWmz/YgYiTZjkpA9vWG5px7ROWuPK138p4vOfExvS8rl
W6M+CTRRalqCcJ0IiJ+IrIq186m7u12Xm0005yZyTDYN6EV8w038LKXP0vZq34J9
rGIr0iT7M8RLHPPkrgIYhUhYsYld8UIqPEZmzSH3VANeIRhco/Q3btYiGpq67lQ+
IjUJ00W5cvZFOpo48XbD8cQ8XAHIZc21DFtiB3uPgt9qev83Sn1Bz9CAITltAqiB
gJOygBJwfhAzu52g7TGTCSDyzoyg08uhB8snI+kdd7V6hbA+A+khxcoLsDURnZUF
U0IK1/2RmgZAKJnovxJFzFrl81sG0mNL5sKzQZyCnXRLzrt8YUOUYUvPs8n21nFF
ShlkTC0rwxVvtqXAwOOe0ksKYS4LuYz6FZe+jH0pL1oNxNoCUGeTXzg92ep4kMkI
XKzAjFdPNx8GS2XCQxtdezJJScaeEHbnq297tzuPm7ZDAXZFVIoQYV8UztvDnzWK
3UIDm0YULlUXfv0Il3Qrcp9XLYmL4X7eVwTRmFePsXFC4+7pPEv0oOkniVo5ny4V
iSxQlhAJU7L5TYwRtx8gqR4ED/copNr2tRCYeQz0j3dXtd3jagYT32o2QXSY4dQw
Ab3kG8JpLuUSCLoAHGE7vRR5JayIZ2+aVr3jnYAhHVQaXE9Jbjc8/Lea1KraEp4+
PzIxMcyucZVfwBsMIXyabv3ZgIpUzdkH/y+o/nOf1Uju9wlQYfbek8+RwBxc2fbM
jR955R/70JgERVjjd0txgE/h1zX8UbFbhmaYHu5v4rZIF8Cvibuanf/I0BOdrLOd
kbfTAGwrnqBWjzBRQTDXRfsD0kTiv6uU6dSam7fYf6RQJusFMcDw83jldMTgRcvi
+nuFsx4xoXl/uCPb+z1EkRWmBWgCkwZHYG5/+JdIk3BFmjrsTz0pELkpLXS1oYjj
FZ26gfkt/N9qI7DP5nyJOiyxX2Myhi+XQizB6COYtT3zT2Go6NykC7rCMoL00Ak3
Ae9GKMDZ+L9qV9OAWfVYv8hGTXrNYtu1Bb0l4ht/hQWPHNhkWUOtOSDxlcho014j
dMdDYqm4kq9DdMI0XM6e9Y6vexqSflEQcyXmqN9rI5hvVoTMm9JlEjxbw60/mp4P
OeD3ynqXXzQgSTTgV6095q4vqD/NcQfkHSdk5NGwaYZWRxtWfEn8Pqq+OMct5vb8
KIj/5+WaL71LNwt3pol4nrRzPgDK/OpI+jxck6jD3stk0pxnBeH/n1jL3WxS/sdW
v1ccHxB+FvJAwCiC0coGffUj6v+Kgf2eacKJgbueBryCpP6zqdVgo1jc2e8Ic9P9
HhhvO2ZOv13L+zT0k4y9Wv/NxwllI67hu8URqNQCxhIzvXyrrvKGxcnozYuHPQDZ
3SYMv7h6VqSpFbYOxotoBo2B0QBjcnB9oDl8qFZFcUUhhYhvGsJfps7Vy12N1ERb
HmdB5y9L/Q+UrTzOgOwcwS7WQyLgylvi9mdDiq7QDEw7ebebg3sCNdtnuLN1OIHm
025AXrg4VIOimSU+EhlpJ/M5GJhTZbWbtu3aWtMwbEkNagNQaDl/38Ht4u2lGOhU
Jnw1+FT2PHSntbDgijrE3FoWYgQO2H8j8UJwohslNNTa5omOQ4sqlTx/JGVJOd0t
edaPeq2DkdVPGIVj4FJUniIqgUOc0RXfTMlcgtbBmsGlT1X7Brw9nGsDYuysYrbY
qQqkebxvuS9s6e0U/m1yV21UkzytT6fZPQWaSv4oJdca+uB5ngZNuvUnNMzPoDys
MK3+Z3bpHKaEx276EUNvtEa8yMKrnwE6QvQqiRb+ZRjUJWExZx8dK7PpYvz7cdJr
koQkByYVhHxrMni7F++5qSdTSedq+tTTgLoU6MOsOjs28dViz6G28vnD1IXan+pz
hN/ojN6d45OmQSZWLmmnDAaBjYDhRgNLNMGzzZpIRhRQFPDarjaqgZhVd+09U7xt
VXlFEVyh8/4cPqHBETaMzGhci74VPs3MjdY9ZMtRBCc/pRLTdoxCsWN7TAX/TNEd
xTAnVuWKwXKbvT8lfM+jYSlptf9P7tJoQyLT3L1DCY5GOcbtNx49qhQLhyfmphhG
0fsJugx7MmLoiW3zR0GatPSGy0ntiEsRWulCBNAQ0f3z1KLiASjRY5btA6fFjgzw
XBM+QU84/MriSz3UWqwZYqXGLAB6C5nx2OWUmTrauLTcQ5h4osMXLC15Z1qjqhBL
GaR+jcYZRgqU4rUaDUj92ANXzuThXZSi7Vx3Y77mqbT4cTe8XPi8M4fKSqTQut/H
N0nQLjpRbGeoS4RxoTjJqH7GzZnVGo//c9yI3H09YyhcO0wjGFLiPu4rNK+e2vas
xWgF4Cfh2bie3NPqjzL73thUBMWbolaJKyygCMULhyDJofjRnQCo9G44+EBC3Ow8
jrBB9YFmJYIJ7jpUJXKZz4n0ExqEEqFGDcC8jd7QimqCleJKOpIfA8N/STjMSbRu
hy13HMXiWyvQHfEKlUpy0wGu2U9JhLNOam7jNfcN4SwgdZpZGeG4SAQzRohdLmD7
ak2lP7e4VOgsT5QBkXyl1mbD6Va7rv0UT01/s9Pd4qM8NWdbEWuxdNkSxuW7sdhL
QkcW1Qp5fq6GD3k7UdYAxYujzzotn8ksawsI+xsPWsdxNa3gOBjEPP6bCevCwy7H
r/Vks89HeOxrc+RK5aXYHP+4FKw/Ouz1QOk3A4bhCHNfB2po2xTwoXfeE6TY6JvL
hkkU/Tz7F1liiGvanVwG4uWYD+CPDPjm52y1Bxl2Ay+V0KSiU9D31AecjtlixVKZ
ceAvaQZQ5QBvMmH9AQ3q9XY7a8cM5UqxEjgGU+g+9AHWqPOsOeZW7mLS/eJd5z5a
d8OtndDlK4t3gN2OfPukPycQi8Yregfdnwb+0XXu+DY/8bIAQdXLgI5E3HLg4KSR
6qmDG7tJ8YDF5GYFtrsrtO0L723bbXQAXfUhAun3An1DTFOQPkobXL3iK13EAX9O
CVNevLxwxJKiKdB8qA/y5Wzr48s8IYowNueHvr+4ZCAjdiftFTfLfu32crbME1QZ
TKuUwjYYDhq/KihRXeWvyygux8VSxn3UUzCVdTjCMs02pDQnSZ3wzetWj5+GVZHO
KTJc4zDzqWIXl5nzlW+mPsLXhOh04rwcWRM/tj8lod9tIjDJNl7lFMn4hkmyEADp
lJDneiENcxsl6XgkJIK09o0uEscaA3Tn9OlWckFT/y091M1tBH83Ac50KiVxapQM
J/Hn6jaOgeqtyeacm6fQxnIRK9EPYn1pfKEn7ZDHIxHXOvOiFA2bEXUt5kz07AFj
tFwVUa6n19kPgO0XsVZUGQYeE9wFRnKxl6qKpnaz0otj/DFCmJkPk6f7NVLHWen+
k6wSrsbQu356Z8DIKK6oAggvJBD4iCBc20X+tbX0DbBcUQLeIupjtBTdpSaxE1cM
NYMbO6rWwUrZGxtKppOs0+W5ENaSJJRUk+lD4WnEHfh8i+iPlrccay8LBmye2YYX
PZIO5qSeFslVL2/WTbjpz5BSA5VLZNi+Gl1QTSSz3XyqK5zZIQafQgrF6BQIY3w0
DOpYndITBIo5gEaSx4i5Y1PHv7lCnzXEuJ1l0aHXm02GlC69B9lcVTma145AVHmG
ILQRhktR63LDQ2v3zuqWn5a5QCbY4rdeHJosrmoh4+t+W0xYXZ5tVjuguK9SFRNJ
SfyXOOPX4NuTocFzi1dQ401R7sOst8KqU8nYOcHQaBIQDVEK3G4MNWpBo7Sn3/KD
nxFHlbSwaQr4yQEQfXZOvxjYhzlle+FBl8kwNj1gxtGDc5Pxxy//GxMjC5L2xqEp
mBEQ4mxwq589otdBcBy22SlnfKDi8nQJWUkzfS5d1WbCpsgjbayOJuHVKeSnoQPA
15bMUdC9oIXr/OQXYnFQrh3i23vpDlu8sf3xYaWZFZqwd6EsV0CdQWpwFmDgKc8t
iWj2AgcHtkOK/lBlv7KxrAIbCViLKCRhl3VKoxGrXSy8v3y1NG1BI5ZJfqVIqeVs
ocQmmlZOP+jJaZu43fKqivd+y3TDkgof0TblNQnF+3hGQ1mVLhi9LmNBLOzNpy0T
kR2FFDJEhvLMJqK3vI02r9RoQYgkctF0VUznosP2BoUCXkZQxnD6v/y60SJCS/YS
eJF0IAJvLUFcH+i9QR/gpAud812doVN4VBjaslZ7YwGItIhdneKj7Fx5qA+Erx0u
2pUxITcYDPs4oEwnRQPwRvtjd3CsbX4ikjnpesULmLb8CHx5bUT1Y9pTDRdX99yY
Pbs4sJki6TPfn2pwoUz8+1lIOduJaWM3hKQDxXYkNTiUXg+4Jk2vMwcPjJKjl5hi
uTWTLXadnMbYOTXXpM7b4eGkbncKZWkQ4sMlKeedi55h+osgOCemLIBYyyQ1qtNX
7BfYrEiEtzX8mTRsEDBSW/W+PgLaKp+7pnZ8pY72mHzgjcLWuCUXeBBXMdUhkr/8
1K+9WN1c2HOHLpnD4LbGCBEzWNWcQYW7V9wJ9gG9UPBEgOjzGhtEUfjnVODozs9v
E/i7fqyxGL82oZFvt9tI/erTphhcZDFB6Jg6htjA6C3l/ROe44fNSssmgh9uhxOp
viBPyLXzbLkrkRSpMQxXLIxZtzpKbRTVTKRc4TLIM67RdAGzUiSgIFrH0V/4HB2J
C7+YL16CEuDwlfVUbA2fx+JU2wbWq0sKpKknIAWv0beGH9jcEcwzxQtFBwzW8RhK
fjA/GWtegoxp6kGZYAoo/jkuhMk+4yEqFEd/+bsAN62cL82uZ29dcm0fcHeYH11n
J5Z2pH7JuB4wFlSCar/Sev4HStDTj2qJHkzepVc3g+KV/IDwlKTwlwncrF0/OHjb
Gsp7xuRfKdvfjLRGW3gXWldo6TG9CqFyZn6Wc6dDqigm1ytNM6LKgj7fMdJs20V5
aAe2bQwDsFpihEYJ2Q+ftukk81E9nHJe2G7Lr/uFC/sxlYDo35jKVGVEff8u+KhX
Tud0kpUzqOai+038Q/gKiwTSnbLgsE9aGHFsPgK1Eu3gCJZQdU+EpvRXqqRUMsM4
2LIlQyy35+4U0H7hdxd7VoQSMW9PNzh4JrfD2bZzKsKTubL5/jaW+Lf9lPLEPeuO
N5l1mXXOESsvM5h8MurnH4FLQ3cLlGDk9TSfonQYfk+L3wENO5d8+nvic5631Aak
cv9g/+PeVPE1u9wYgC+t1320v64m7vwOccyQrKLPdSQk0Sds2FedwrfqkzBQXtU7
AlgoQ6WlqlFyg86hNy4ceozHtLvvzbt9xUd+rLq2+4KY1Y72DEwefnWmw+iXJ4Jw
RUOF/50XlwcVDB7HsQNAex2LuuWKWZKWW/wcMGRcNa0AatncO8VDLh6Za0sWs76+
T1eboBDg97N3n4JjSilKHDTb/jwrKpXnpFpMukgZmOY1wzcL9kDgwQcUfMyhSen+
/O2VC0w6fhp4tTJlNZNWlUDh2TbG2iyt6YNaxiyfJuPgsptvmnpY6LP7Yi60msZ4
9Qiyc8FCrO+5tHrOnz2MED1m4D8oQpmkrLErnVePqNZI1AYGdWIvr5FSmrYrH0nx
TDYrtWziWxj+lNxms78LoNTDpmzoI6/76UT0AwlxHKtX2wjrexP4OgqTrVbBlkB6
oFl17jRlUokeX/r+xPYPj5piH3Cj0WaQs18DOX5DwcFU5kd2K/G9bAXaJNwSwCGL
2V5o5MIfqEFn4Im3Ya0b3fUMXY17sQC7dYzmeuvMBkpL+DjUXSqJeTPbnX0wPsSf
JQQy/E33pK2MF8oK9m79JndeA+Sdc1KGJFBNFEBxPn6VqghTXcMBVsvku+8sB3Tb
Mn0YhhkfHU8rwsJxoWjyXtt39D2iAU3bQeiR7mDzof009WX6Uc/SOhvPEQXlrCc/
kOYmjhXcwm7u0CoV3liaMx1NWMWJd9R/tnKGFvPHiUWiNZhCc0Ped4i/jY4F41dt
lWm6NrPrKANxEzw88eAQS1g3TxvCsUReQlNaSke9FWEbCC+xccWIAx06EsuCcgqN
UJZLgso3uZAR0QxcAchX6wK7ndGIgl+cjZ3ZQmTegTukuFopwVcZcYOI1vI1hYoC
dCAN4zTaawGtftL9/BMvc0tRSo5SwJuEwbC0MOie+rt2ZgRQ6RSfQNSLMs61Ys24
lTeAoBPPTQ38Or+W+w95DqUyxwNp6JAv1CO9+hQMC4b/mkiDASmBCBYKsXIGKqeR
oDAQLHQY0tqRvHxXg2Ra1HeLqC8N6Xqfsf6jXsbnVoNwmhaRMVZZFrXZwj9fLKyX
VI68hzODKwo/efDR1sgxYcqWuRohFuIIcs8x9ajLgpsiZx3BVQOvT3oQdLYPXwln
orBBq2pT44kOp9tIRG7TGEhOeGJjnJuwHlzZegCss9ZRpO/F7NkvDRmHfl2vrE7/
CXHoUjPIYSjVmaDDHEkShtF0PZYKpz/cY0SxTOfhlvvXCz7sghB/xHBb6T52FT5Y
xfObpey0RRCVMPm0qwVa6Aj7sPdWuo4iAK7+5+LCDo+v/25Ptl7vTxd94TPuJDTS
4Yb3szDlCoB4E9vy3YmEuwl7VYAGAQp4yha8O+3mLb48WXRuRJ/3YNebpFOUJSYz
i44+wy/N5xd6vMnVUQpM3VhS7bXzldCVTK7c2VV3gne4XNXFeTDcRgk1Hd64qUT6
V4M+emePwsFLB1gx3dbI0wa61MR6Peh47LGX1OL20ijEWGoKLG+mvGcjjAdQeLwr
JIwJKXjCbeqrE909F0OT+RtrVhMhyx3ZnPu0/AEr8ufNpqkHAV8F0unsDixHXK8e
sbnD6rSGGTA6YlGrdYw96liwsKHr1fpt2JRF6wOYa8l0BZlKiKVzgha7KIujveIX
0r6jyH24R2gD+28d/h4pLN2trxA+VwqKn1Umi4BflpvZ2Q80BYJqkvmXUHSxBV5s
RuXzH107euPmh61f/DI84ONKVMVl77RifvBpxfcDS6CMPojiqvKQ47j9yimJjw3o
novIvsucgpzxM/zfBinmp1j5xRpbgVdrRgBwfLSnmrv7/epFPgxVVOyDdaDYBmKm
szqQ9HrAvtMzTlz35Y5Kg5Qp/Kl9s/wozyDrUDf1qdPk8Y2vNzIvnHL6qiRcf7DB
s4p7SXgOZ8/ahJXUPJkLEJqPX6Eimtrs8K73vA7IrIrOzwdpE4G+9EuSKUZ30rTU
N3A8hV53NBxTHuu/yR1vrGQ78Yv43g1M9Kt+e2771Ho9KamEwEisOiKl8gGHLDxS
d/Q2iuJaYaT/g7cMWCX1MJcb8tpKKX8kZBXaYHN8Cdw+4RhUNaoHQUSS3D3WVI79
Wp7FqtmkjsLTtE8p6bvdwut9hCceGThCQfvfSMqF95ZRqkeoGmK+cnrHUZ46sxoS
btCf+8DoGnfiI630oQdz+yt9xp0F5V+zBcYiqUgS2pLGm43vnWHfl2eF0n0UIrqu
zx9rB4ul0LklcL4W/rqIJgf6tjNmu95JYBsFcKwzsH9CcgnZoaUdTuh3zrAY1nCt
Ef+l5uu+ZXMJRKQMXv7TRxvnRVur/Pxnh6ATdb+36YLav97C00yOgIAblJKyGMHO
rB2IuIZjIN5cfLdh7off0GrW2/6AXoxe0yxQzJJUxjccBi7hDCrlcOgyktA/YUod
gW3huc6I2OoFkUGCUKUFj+esgYYb0fkWCV+2QQhwP5UBnvoStKGPpCINmFK88nGc
hNZpbxS2+iksX3YYBT5L0I7yhdnZiljHQWOGfXMGV8tbjnNv7W2A6aDW2oMXcgYS
bcOs0LECR/TvTLoTp+BquXe/Wc7n9Zi4kGtXZv0ByziKaJC2UWv7Gx5DKNPnPvyD
Q6pa9BLlFU8Cw7amRCqeniBRG+Ic+xRMqCb4G2trIDUjrhmhq4RzkWnfM7dIV+l4
hGZjXcgKye890DXcksEIV5IwN7BuIyBMR2kVP7SGEQP2PMRYGY1ym2Mym5vWRt4N
K6DlX9lhgDKgimiJYiFKcq/Asm8y00ThKo56fJJ/WXgTEQsIrifVDHrU9+GqZm+O
ruzdWrr/rHmt4ks1xgtw7ZTrgfiCAIYGDzgMZJkQaTpKm165RJbZiwzpmBQ0NdK7
menMH4HXAwYrKGpXw2Rp5DL6WyLWEMdOffMa9GsgiApXyK+Di0xOVsAHU6dckIBK
dzQkR1zx0Vqy+k65isr1E0Et1U86i/j1mJGtLi3H1GdyfYlgc5Np8X4mz/utgl+6
m5zWyTGU8grqB5uDnJV/2PpAs62iTIiffCx9H3XGTSJr69y8CbYm6laZdRt3mjz/
2UDqXPbSc+T7SeUgIwFnk+xq9SBZSey0ce49FTAFomHtZ7f/H7Ayityk/9rbQH7g
/yo/SzImFVGSv8OOb0ivhCk5za9dWAbjSlBKWQDQrR3GZkIxtJuJ9i6aOQAH9oIH
kVIdqHxJzL/P8uX184nB3+3L8UJGJzs5VN5TajxqbS6Qg0AbY+Qbt49vP1rA8/wn
Wl7Fs5G9SB3QMt9jSGHFatYObgm1kpbi+Y9cBoJQDJNtw4h/rutbtggb9RswguvH
Xu9l/OM9glIZb8yJCCaXIHPYkEhUm5DRGBrOpSCIebtfWEM5Y0CYo8s+vstt8GR6
/tVVpgJreu2uzf/ZXMuWmSdcU20y0F6Otwhc67u5NHxWFqIiXSbV1Ph17nrLpGjb
qxUzTiB7KNj3lc0Vm1RT484y7fSnHRvvl09x8zkTAIkuRAB9eM+PbT/YJRTuDsNb
8ljMSoJw8yobv8PKc+g/xcxDUNhcM7lHbJ+lwa9RbTD/3/gAVJuE5/BipPz2fGw/
YoN1b/n6R8Fr0Kg4r5d08eO7oPlZ9I26fs89Obo3u0wquB1sN6feSZWjmHhtIERH
9erHwY4tEQe6ST3e83V/Assr7bAStL+PzLyph1pzhU8N0vYWRfCKH8i3K6uv1NsZ
t79/Mf+p4a4h22ol+eC3HqJ8IkgptGhiAgo2SHhIcNGk8FfQh6nIyLp0zePHgqFE
YzP7nLjpBrF6GtVDxsP1lMF30aNbf6Z4kNxyGMALX2dsUimLzpp+veaxjx9J69AA
E9c4XuW+ovGYJo22UCBNV0sBOLFez12L1x9ktWQ/AiaEiApnhrolPpVC+0B+C7fs
4yy47G6/dzjZpu/1beF8VYUCatUMfI72ocMpTFprE5cDo/Q75rI0uqvVTXoHTcVo
jnnz24ZkGXFlO2eu71J+2uwVYZVqWq6Je/FwszXh5kcrAw1VigEeuujejf89D1iq
juDDzQJ9FqMJjBlJroIHKEQYQIpQbPdW07vbQOta9An6D43MxCUrA1wxHm2yQ1wp
8EaHb0Z9jui0qShDaECe/yCyTpgjXtMNUrf6Mf43phP3xsaQXHfsfesNlhaC0KoS
NaPhV6FqT91XTR1wqDlPmwDWRwJDGS9xhJuDgpaSOdapPdnhElXpc7SkFXG630Jm
lYJg3DNRLX1TGj5OzMwse72x4/Z9FM2PsInmSVVWyXIBfw2lg3JwbCZUD9M3cBKh
02Zqi/kEhCbFiGlc4Ysln/Paj+8YmW7x/qWn8mYBfjPqJFgLTHHi87l/g2TNExMX
Lm66foZ9oJnaY0EBLqeuT4Ikt32sigAWtzgZoyRTKJAZw3eMHbTo2E0YrROZS6Fz
hGgGH+bNqTUZxH5SCePth6YvjRKa6c+aoJY5/5vKYhTGN+mjT9pNi/cAsxlWqw86
LFFB8+kv1lOk55xL1dr1aEldPPx8jjIE7dhrpOiEz7yR3Z6RqkajVmgST/5ss0K/
3lsM1dIzSNV4t4U3Z5wbycbHDt9oP69UngxLBQCMo27rKMaxe9+MUFNXOQP25sSp
zK3+WdB3HssnwrTBk+SgI77nAsFA+zfIBqHlTcfaZCkofBC+qGpX8Bi6mLwZUfCN
1oWJaOP7cC8COC/ArHo+n2bWrexbRTfe6YDfPlKx9iB/2I644x32uPb/sI4H5Dw+
K+FvAvD9O0r/PSCUFL9Xm1AnUCTpZfEjRQ08njv4nqtCoiJb2pjN3EA9u9kAapU6
g+Tq/W4yHrEN3b230BFQ6mm+Ph7bb1gQHlixnppbnr4n3hJ8LpBeDvicC6dffDtb
5t3o5UfQwf0rElR027MhULpp2nxRuF3Tae73yhgRHlI/fkr5ph27hAZCFU2fotOs
ZHNsTEDPCc3NF1rT7R2yju6N5OOfoQCwt9Zskwn2wEBrAaag/Vdn8y/8BVd2rs06
GbGmySgNTQN2NaRB+ri4Qrjyu7tFMSJpG1sy6i4GYLC/u1diR20f52R8LIe5tHQd
UfeBpV0t4tulIavjqXrVbzXe9CvbyT772bHKx1sxBpAOPZ4NyEz38KgtHNszPs+e
c7Mp/eOqxkxfWu6N5h2AR24LbMwjnst0HcGHNewXh7O++0JXkGrW3agBmZfI1X3L
NvbLpIVMTfYk5lqExvYq6YH6JvLafh2A3OI/7oflfx5yZXNoMa7DoYcNCer0jU+c
cWvnyNR2TEXK1Y4Mdvw8TED/AbMpRbR6hwUt8vj1eelV4tfdJsTAYPfEYk5M1/me
x+R0H4FHWKadSMSXAHdc7qspke1XKCi6qc5mkE9SuvFYetrzPeTlm8LP6pNqPho3
xIfHhzr+RdXJNP80i/tJbVm0rnocKD2L/qiyVHQOPz4TEP2Iubz7NT42y82dsW8h
+sMmXKn4Xv98d+GNfJiUfwV2aHFfLPDUnWSX/2q66EFaK9zUn+aJUVa4Tw0XRAW9
bH2+GFEQUQpZyM1MsECJ4DoafdPEqcHZ34lTxupEVdJHlkFl/QkHieTfBoxH2os5
ddoKKEMgR/GifabaOn/hjG8bzS0MxMAeUSWA+JxMvbyiD7AvKXzYEhoWibsFFc9g
hVCQJS8myGQNPtB/Ud3tEp1eTLJzi9mbqK54mMrFsXmMqJj/9AJg5NU1a7gMPIow
Xt4ZYypL8rhSodWdGYRsea4/yXKZtmnJS5MhBOI3cuu/fNdpLpqA4G//iosKzEWX
4Snlj5Kt1AEwf9jk4Ag7QM/bIlJWe3qfa7wxZ7oIWoTD+1pZGojlIsJnDp3REVnu
kMU0GE5xZIZkjAMA4leDUiU++P/H/8r3ZoQLS7UScWthfH4rILo/DHbtIRAZ1+l0
OqwuiqqXwnLeq113keBIlOcWGumajGCvF8uQ8w1AuO+Ia7QmA5GTRhn8AwnDQnEN
LSt8A8hU8r0hAfwoiwswfA/qlxOW8ve9Uh6uu4VqrKdwvvEk5vD0+4JKAS1ad9Pf
W5PbJ1ijRLzYH5F3d5KpQNb6JwNlLYkQ6ygz+evX8vtRD1lDFwqThac+IGVg1af7
ixwz7zxCsp++SVjE8tc7jQn9BxJ9FWIV8hZj7aaDkWleY8oQGScBzeY7NaWE2lbS
wxmdlob8kQG3wlbDaBtXpFzJCcOP6QpGb/cS89uPTIoXTAdljsHeIkdUyzxDz5oO
w3bRhrJWzDVQQ5FEVw/vowe7e2aJfQNWwTpkXnw4WSp7jj/jTWMnBwv1Pja95MPM
ueDpw6shxxuUgxHH+EbG0B2p3ipduOVUU+uhseXWKms8wM2qxbobr/hQNKq/h4Mf
60CpVvPvm49Ph5dns6c+LIamNJMfbXW2yV9HOSxGwCeafXjTbZKCPUOq/AkPnKy8
YxjMN+Zmy1osTye39iA0tSBJXkGb+e5LS5pZHd+589xmZiAtGjPBqT4zzpe29rA+
z6SkHHsExMQZ27usDjrc76eHcT9nALoNbkZ3Si/cea/NOzagKLwybsANk6cW7++7
kc3qqO2A5RphCLWJ29dB0Vj+G1BvbOAjWhY5riK0qRr0UDldtHrI2+DIfUZ7OSL+
IkU8/ZM94INdQM/KaKaBxm+jWn3diz6eo9a1Wl5ChJv2FU2xtezpa9/hINFRMBnt
0h+hA59JVXgcRslt6vMuEMunRsyEtiaV8+V49FLjezbTzVeKWfoJlJTVfUtUcTF1
LFEMVqsWBI+MOv/8yaQaGMXxJlE3R1n8DBKNt/+bm3BuomPLD5uunkpkgz7JbET6
jG/6i2UHlKc003kqk+XXuZtGhqSm+qARrJ1DJQH6CwzOToXmzXgR9TTRa1/1wGCq
qp6Rlyzd5OwzFuhoWGOK8einKR1oH3Hxf6iflHhwx8YBVS8sqzzun8kM2M9K1pxB
ZJRCos1a9EjBCYZynjeaVZfVnTi/F0sGTNhKrQT2ZwPMPlUYFiLfuwdcE6URUOUg
8Olq//EI+vxxj9HmeEABgnCiA/WnLa2aH2U0WKcjcKFa1juAADqJXNawc4wdkSFN
Jo7gAtYW44o1+yTVW3k7jkfMJzG+pWJoijunrSkLlGTSi24hCV1jF/yO0DDZMwTG
eYtUw5keUNlQggxRwgr65xkPfXNjbuce3PFZ7ka5Oohy+4iyhHeoTN3aVSVCrA3I
2e2zV1Szsyd3+5WbJ82CVcV6ctBUrSSNaDQTlPjxY0bHS6ZaQczKyS/uP5uG6Ohe
EF4DFo4woqKXsN8oxsH5JQxFS6jmTfjMaindmFKfgoNhPk1T8hnifwT9CME5VLcj
zln7tuMjgx2/+8tNvx0h6UW8d1AkHOOfEVaxc0a/C9xkzx9YB1op39K3x/AzDWUy
UjcqLf5WPreCiOeytPvqXSwP+kqLwTtN6ydnOjTfUEN05MIXW6T9T5hg9HmTE4yw
2ZSKGfJzo8DAgKsHivTmmLerKrq9+UNYzRvlanSwFa8utOTxOvj+v5AiU0Avx+BQ
vTmwA4C1O4yJZBOByeBW+Puf1LlhHUrCxD5ElF44l0tr2vs9SEtf1KnLKtaK2mZT
jRdQAPbSPwDZox5un3sC47muo57GI9r5MK3EPb98KcZiXSWhMy9f/FE8bU7PH6oc
xuxQ9ZrFjO+UaQKnH+RYV7NOvIGdJz0Bth6Yx+3tx9YXwByxaesyGyHAiDLURxsh
CWuXxUO1rjHaen8KWyg1z502jxxZ0HfQOPcQc9z734D4nr2oI2WBVWx0j1XPDjEB
Rpxe65ZWhsWWX9H0GlYuFZvZXWibmoepXZXhk+/q/PCxPrjQsfOetzRZbksS8qCD
PhGMg9hDMIEPLLiY9nUySJI136gHm6h7QI/5MvrCBFulbP6csw3TDNGtk1YkBQI3
74vq/s9yqY32Q8EsHkQc4HfMeB4Q2UCvgVbvE2UcZUwEfalYMs6mt1VALGX7Zm5i
m6ApBfkoqTTttADgTd3aBfx4GRJdRXFJI5g+WWqFLn0fq9jH8oSm+of6V7Rw5LNH
JatoOpvD7iXrHMtsrczj+r1g93ASLwZFAnVN95yd6GOUzfEFfxMzrXX/yhBP0kDM
EyH7n4BIBIHEreq3TqqVRpoyO/GJyj7wrxX51U/J3Mewk1KuE/KGhBOazISBZUHV
YNO8wpWYM/bO0snZcTW8BtxVhFyeperr1thTcj89uDExLMeYvOOjbKtYtAkYt8SP
82mu16OoxHoW/M/cXWJL8ANb+e4z8UafkkvIM1HrtSig+AuxgPT+uu1+7dnaT/np
clPTJw7rgL8deQ0in7E9x4y8FM34X/hiilr24+4T8yG/hFe/iW3ZgFBnbUoJg/9t
BMXBX6evtoD3JLmFnH/2lPj2eur76UFULlD3deTfmKWhjCmmPry0u8ftAcIsFJVF
zYFMX0dsDOFgeRToJOYYkWfVBNs0IJIkBaFD8OVi7YU0JWHrVi8sc63nMnRX6BCc
HK9ahoLr8jFHlsEqzhQFMfe5qKF4juFuHcGZKtb/ISkdQVbuqAhJQCR4Koq8pHsm
UOPJX0E6w0V4gCDTLjFrLty9DOBURP4B1xEQukr1/5VBuB9Yezx6yR8y4gTw4M9w
pBp7zWFAkgQeBTR8WH9H4vHU2jELCmyHjpiBM5Z5/IXX1RPgpBOKgFk5wkshlI/Q
IP8YUeRXDJ73pr6edl9ChRAEcPLTf8EL6Y9fZSmVl8ycRwcYYq3/lgwPu5yOxnKs
+Fm7jN1/vYgw3d+ZLkx3lDvNMbPmsAdF7lwcoE61clbAl3c+vFcheOwVv0NgsUIs
X/kEsd2B0hZoByyVDKetuch4NsIzyWf22wevemDzdm+/YU7/k6R4QbwHFK1cPixx
udyAeASQdYN+41YBsZqixgPavHdbo37nmam1QkFV+3IqxWlVvltyejm/rFBtD+jJ
XFScEqvwIT+/05DIQZE42N9dNxcvsgS51yWJajqE4t/HDEmMxqCGaOZnBSibuESk
XzQQb7nzD1v6bkl/c4NjKsMUp/vB024qdGlaSax2GHq3kYSe0Ougp7h/ag/lz1J4
+RnZxTkGdjZdUMJOmyIvpQKJD0aHqkjQg549QaOpqEOSZHIE+wIZu2WCO5Qwe7fC
hn46T/yjV+xlsyUsTDCmKqWdoB4vZ8+MkoAaSgDQR0nhxHCfZKy55M+gWVYTdj6/
KAZp/8Twe0miQRdPZkmesni3g1l6zVimUtWCTs+sHC7aAmRnB6YnSL/IyeJBDbQ4
A/mqXcZob3GZhYhqKHzfgKQNKkcWHAsk/QPWmPXI/okIfiUpuKlW4LamWMkb5y1U
maA2q4CKVmdDsZ7GJpYH7eaxq3Ix8WD70Wln2R3HTvTQZdt24eKYFvDrB7rVAuqi
DxN+9p5rilzFlhsg6Bt/B7HFbab9pNpwMagcfzduRJMnZ1ioo6vLcyruoK/xC3So
l5R5NLzZvNGdZZehO/9mZdugI5jpNT0HNF6gMK7q0YF0r+Owd/tr1wQ2IIbg2BdK
4ntwLVOXUBrinl+M5X2j6mRFwGbnhlNlGKJN9da9U+PfWy6jD4I164cvqolRF9v0
hnTfDTqH8vQGgGDYcJ0yYtRMrPOUYffGM4iHLOByCmmYRo6KN5Zj700Aez3svETw
wQE7JIWa9TjDqgtcZ5XrawfVma1GXAuJInhgIQY8GzH39Hf56k9C6QFnqCTRX1lR
6nFf/IUWNHhY2kUwbz9Zo0fKm71uyvGYRghPzrKmk9HA312r24I7Tirrpn/5G4Jm
kN2F7aelaZi5rJZDjeyJCLO2g6fmGSWoEcThQC1fO2MKSjtz90TfRSwG53IrP4Yb
YCf0kATErybOQFaOYYyCG7TEPQdJQzZcNj6ZOHFRU4zgMs5b98+qL4SOuHE4WI/Q
RSRNfsYZLwL0ewfiGjDaJ/716dhWnhvx+dcpDCJesAxkSyqm7oovvzDpSGHkhhxU
fujuBeu+lLUYn9QiZYOCOfnuQk5qoIz7tqLJJPPNijkfRsfT+1VRLmGZLzyg3IG5
mmmiweL6y8V33JGWPq6Mfvos5Dhs7FTbHrapSh5kD1JNGsV6sl2kYRfVUxO4G3Fr
CBFL9vSW48BUh4DzHAQTL+hRaQ2qxwTsrl3zB6gx6GTIZUhwyD6jqeoMkx6r4Jwh
KpstXYFRQLY7cPuWzaB7nLttJMG1VmnzW6BTuY/7M9h4ZfIFcVZ4nE0iy69+gMiA
gU6jHhEzjoL6CYKKs3iHm7lfkEqmQ2SuGbljgm1zGxxqYs3k0qq8VAd7hjsFNlyn
7atie1nLFssMQho9x8tloDUrRq3aFLnhbv1dQk5icDaw3KfLPQGWVM62u7idjwo5
dBISlvYRCt5YR6VrvEvbfYsxrpYx3seHqnhYmxyY3NiUkXKZCw8d1c6HrN0zb8sv
5bxOAIL/8cixgiJWltl++gJPp32kX2J//G0g1qvx/zO4lb9bgMGq3K2kxAl6RuDz
KV7hKI+NYjpEMzKi0WYBY1wnu4JsplL/eZJnPNseHpcwW0tgvPrHODJayUgo5DkO
SdRvy0FNhE4iXnv1bCdHm1csiYusOOqZPFP8SZ+FWmTMubAVzPB3dxcbPkjYBuHf
kA3n4eNmXOBjnEH9YqhBaCoFaC/NJnVKuyRdMpzZ1om4EqJJSWDusjL0AVSa5qC4
UGHbRZ0qBzptzQwqaBoGY5RiKrn4/UsbN5Abw5v0jlIe+HdMRwKLjikMmVZtX3rB
cg5R0My1s1lSk/4iZtQi/Td0yQH/ty25nsQSo47033GOW8Y+eA/1q/CFU2Dyx77r
ZK8CJYPA1qUPWEbI5pC8GC1qN//7IX+gw+xhHGqLyFNUVUsVxlxxMP+BEoSDOvzS
NcqN27+HKBdamy+/a95QRKCvfBrIfJtyrm1Jz/uri5ym3u0+nf1cNFcri7jW5o8a
6Q1W0gJ21gESahEL8pCciqIiK60Fk2cRjO7q1x6X6cW4DwgRmX/FkMFocI5Sia0E
ET21BEMT9J2yhVlpHv6MnLdQM4jDuh4nUUoYAbdnVNryZsYyQPvTgVwWKzIRRL1N
wXpjSLqb8P8+QnDNFPDv4q++zLLdk18McbdAhKExHAJYjrjqaFCtWxJErUmgNPlI
EvLhfFgVF2rxGiDyLMzPzMoX8sKUTa6Hia1ghTAldEgnR4naDw3dNxvMFDYWZ0hK
EkMVxQqXYDamvePI+81KEACN+5AihZcTZbKyrnnF6SkCvmlYsyy4n2Xo+LX6mV9L
+ybws8IAqR2oRqOTH/TOePGKJ32+8KH/7sFzl8j5Mo0UvE5htTvEh8/HAh38PKHv
ARw7eBT/H19d5/m2f3JK82b2rlay5UBc4p93OXfXS2ac8MpIRo1AKmD31EpPm3WY
ueLX9MNPhVrTF8XT/5ntTVDKDdn08/umcS/x2+T+yyjPck7tNUlgJqBb9K0hfcco
m1ESegtEK3ru+hrFHowLzphnLQ14B3QgC5B9lzPR6+TobBTsCq+aMzXfIx2iXnNu
qT4VV1WEwE8nYvkMnNz86UpzbKRgWYF5z7BAJPedZeXNVNHGaJPB+n8ajn6+4LlV
5O8iXu9yOAPuILU618QpoyaqTh4WoPqJrSM8w7/41sj5aLA6lBK73VYYa0SO5wkn
yMoBhHvAyiIRM6R/Pwo6JRW59tLpnPpmQzFvK8ytbQxspKlPPhxKIlNfvGOFlZOK
PI4ffuAYjSMmat+VEBxovcY88+fpffKcuB5qDvgdzZJisd+Jzibdnz0s+pZwQ2CN
mLn3l+RuQMubqgNjCPqcnHbKJKbjX1OZsSyxiYw6ifTrAeIMI8y9Rb3niN1ogUrD
AuNxrYrSHH+EMp74bCfg0Bx5f0wSCQK9Lof7ljtqlGYf2S07qJR0TOWydoqjUIaG
n3B8MwA3gqDxiDP8vcuteRP2Q4VeKBzdiuSQk6Q+7fyv6hCpg3Cds6iTyHD3vxHH
A15//3Nl+1ULQIcyIbZhizncW73Ulop8Q2U0S5yr6cladAJiZWXYq9Ce8Qzpz+kT
DmvLLTsct8WWpDIsxAowMzoH1rAnJD4VaTa4j7FYS2npzdiVhp5ed3tuQmz3FnVW
r/03j6u3pAywGxOlc3DxZMsEwteZT/C+z3IjC2X/T86VfxAZpQj807xGtyOv/cuy
p+dFukMjPfmQ8ec2216EGMAXu9EDC6Dm9wt7PrRVVTkvd+N8tOomXqyrS4EYR3py
LdyUfFEvD0y8rHu4D1jd1xh+B6OsnSzWGk7rL893mUuBXqm69IlpMVpP40fozcbr
w4P/2JrFL77zJPzHqqgqacIoCA9dVnXVvoHkjSbId86szAR113TLzZe/iJEgMfn6
fnahDc+1eivdymIMpfdjGOWROf5gPJbWUWV0fyOII2phJfi138xVSBzdsfF7ntI8
Iq1jC72SyW/0CiJ13GAV6jkUyXe6HXJZs3SNEv30v632GtXqF5WWSd95CgrSA3zm
acyiWSuki6dvCguJBzpjsocOKqI9o3NJPwF40EPInP72X4W73aw4sc0EWpqAB8PG
fR63aKoiyDCrep9BvwmUIBMrdtr4HrimdKH7VTv2z0x29+q8BP59Y+6RgByNmVJ1
AtHsDbABaiVT8sHb1WkGlegv3aL6sfz91dPH9OTvUTg989a5GO3iBvXI83eDkNrQ
PkhJUoTrLKA3Z+ZrQ+d0VjnbE3jwjx9hyMwkuqQ4PIuy5LUkTy7bdPhYq6aJM2zB
i+Z+06l7bj4/3xEeZH5C/6+ZAWFc7Dq6d8erWJWVXwMtCPcLKYOAhJ11R2dZ/+R2
ofdAD10kqIKOqhEhNSJP9JOPib5ojy3ZrFmvlIdDOe+tmXfdFsRV9InNqm0y2C68
OqlomCkLsiwouQ4p3g2a8bi8RibE6GB/iwePnp+49+CTCxV7Sjkap2trftQKHIyR
7Zer0UQ4es5v2jsoUNHbZArD3plZ7DaJ0QR3rRhkHV0QqP74PjIHm0xk/n2jNH0A
gt6lol0AndqyYVjO3d+6zbtBaCoxmRpEQDsx3earYFmdXHqDHm6W19mZO7krYrbq
1PxfcrTeLWDEmDwcrok7dNvuQowITpRu7KV29nCygYqLz8dgog8vzBa2+B4Jl7pf
ijHNNsWQVZPXM4l8qjZR5MC/T6mrzGUXg4ku+atttYne5InR0Lmvhn4poaD/IBET
lfJ9mG5+9Fhw4FtxJxJokK3IRqQcUyt3UAEh/RJ+uoSbNk+zjyBaUNBgzBw8FhpD
QaiVz0+E2kV7LBMpU9fAuJIF3cepB+L/GL/4yiGR/1CvFDiFAcGRn+4EC/tUXK02
dG+KGZE5397h6l57SKJGaMgZSy56sR2kp71FJAbQwXxJ2baVvJ1+WwWK1p/xrPEE
2wiNBP/O5y7rNeklPRzfxq/4BC1W25nn7IUjiesVilsxGDS3hUqGuaR3SotVhF7w
t78AmMQBOmxUjjD1BWkVZ+qYCTws/Q+vns0NYOB8sHH9R7vBGq5+wmwGWnlrG/gM
udVvY18QZv6g+DTRMIGVh8o6CUUK48e9jetiZ/QxMJjlQpJYdksOVvqT0rg49nv1
58LL3UhKlprhse0KHrFOS8hwb8Thq0XZRiuW79Vksa+ukZcKf0zbaBm7mqEoc9ZF
zh7lNYcHsReWcYQ1N7qXLzGfoncMlrjPNBpx13zbA+U7c+1N8Yhbu74taxQ1GvHC
0PUkEpFFyWfqV9qctUwpEXo/yYay/SvLfbCkrAlp2KlVGL+RZrlmF0R/uGsAQZfi
8GkAvssme02sojgCvHOVB9UMN+euzFcqvmmJUgylN058Rwnh/ffpcunpmv8UW65z
W66lycDA++452myoPTZReEGcASkFwNG7VDaJy/IkYflpkzUKRs756aVUW3kr+RfC
NS9Yo7ykCb4HaVJFSbDuNMv7XlTGdo/55tfBlFoZ+Szj3qTdirP7rp8WLfEXaBvw
N/6Qqh89a7pOpT0u4WyuCuCOUWqUcTW40KfwuPsACSJCeZ77uBbHKU7wpmOhjeIF
ZrNxAH9j4sJvEREIzeYqu5Zt98PNwOJOS5MdY3YTeY5ECmo5OmEQQLoDG3q3B4T5
Rq0jg7zs0lg87+iZmrNQL6WMWRuP6lTDJFCBXqGf390/J+PB9/WzpAzglSF0EQrB
4sCTkCs+fN/+r6ZY2CAFVnVzZfynwWWuXfB/s6Ss3Ez24UTpkvD5bGwUZmwWRhUI
9YvDotP18DflGzbcXc6tuDCZDTjCLG7c0YxGYfH/eZG51t9Tp2osG+EfPREHP+fg
8deSbl2urqc2gYHx8C03emru3aJ0JRaHaxI4OrCrSR/0ScbRBNiBZrGgcNX5sOWy
nOwd0+el9RonZpl66BLY+xhKTu/rXhQjNhXDQX/jnVN+9d+CGh60x/5+Vmo6mX51
EHW2PWwWUbZCFrBei2Q/RVsAFoSUKDWhCkEPFkuXL0FzxaeHCkwO7TfbYytNl6Cu
Sg5ouPWVergNJgAjWJ2FzZMyP2E1EvuYbSKhZsb4hJlkJh3exGGbP79apIZHrL8L
2j2M+EaVQf2x/d6U1cOiknWdRucqXkc41rvAD4BW8tfj38HTvEWEverBr8k4lCZ7
iB0HctAB/eKDzORiJbWImXB5oF9GKkL1YwLLJf+IM0aIFLfjX3Mnkvr348nc77bv
YrLP/JnkGrfU9v92mj59n8j8z1pRCrp0joZs+879rGvIQbLhVm6P2gATx+aq4b3T
QDUKqLuzoSApV+BhrdK/SfnbA/X9U7RBG6Hb6vwbHsAbx02/C5hK6uEidigScWUm
Uzs1DpS6jJcZjcU3Rd7nN2Rjao2E26DNI+WYtgZexdxmmXOjZpPl/ClJnml6nIb7
fO+bxxf6qqxBB2KQ45qzSY3WwiJ4eAL29goXDTgRgbdqXNufMpR5cDzsZ19pE/iJ
MpP/GjdbQyp8DY6MuGYvT2JhxHFrBJaEC4sllenF7ROylTOtgew435wnDtFEgtrE
HCIvMzhBLvP1zTtgJz6w/ovKVN0KNbwFuqtXTai0LjYiwED1TAfD96zp+pipmyj8
qlX//GYaBaCsQ+eWtoZlSjzi4XzEsPFKbV6UwSEBOIeGc4GLdvJOED6OhOme5z3V
UBNCLB5sw215wPYhdVWtt5mg+Vq7UATvVcjZP5W7bk3vjxApX8nCLQ2v8f/K166P
3ateGLwRrfrjmHerlEsxbW7+L1HNxKmvezFCMMK/hoeDfJznPzgLaMEtlYlBJLJ/
0PZEdn0di+Nr5waEDvTRyVbuViYMr57b69K/ABhQus1DO71TGBjWavIKSlFQEw6u
sEsBAqyg9qu21YNcchGEBGolkCzKexVfJpbqlRaulCKmljJSeu0OLBO//xfUroUX
cStXc+esFtJdSJd345gx0k0VCpfKSPB5wC1eEm9Di54PSrz4+Nv46ULtc+ZOUfUy
9oco0N1N0OapNdZahI71MRjO3q+VjwBckgqtBelx4NrxHJeiA9FXWP9MfCbC7vW3
ZoBpxdam1Xdd9o2EQ1c5UohpvWNNUKBizwuJfM5ugdpBPHs/MU//qeSDnfl64TcG
1Tvmh/6EHnYAfPmYqtbaWpovR/aoWyNSWuX6TXyQVBiFPVmEuh4JA9od3+qyRkzW
KsQr7zKuagowkWAliplAVSIfOKg50TRtkavDtndf23nRQ9wx/wavIsPhpPWy4cAD
6bA2GLkMkyxuD2m3rQhfxLD/e+EkoqdxlPpcUHPoa01KI6vE2IXJZp7kPSy4815I
25dfV7MXAS8m698lrSWOIkbsq/PYXYaFFvKnx+9J9QHITS6UBIKNMJR8TtN8GOqZ
tX5DNvsV2aTPuQn3E3C4O3/B5iMu1tKDXD39y27v7NrO1M6blVuRZ37EsXjc0OhB
eB5Rn3MfnJu8nBjo3fySMlpaRd5EMZNDvOqSh3ditbIyy369yAslAusSbESD4sEy
RZF3aNje8k+nw7y0xhyaqKe1CT+OogxpAgSJt7t3N7OIyPviUJW0v+bIYnDW7Mh4
UgpA9jAzdRtdu0Nj6w04QD0lRlkikC7zUglVM3Qhip1obADKxITc04Ro0bhZkUJn
v6RrmIf7PO5L2EtJ857GPVpFisNZUMBAkZSAoMQRq3+lAz9G1Z6MYGrdytRy0GHl
E6+DnDwuXPM/4Sk9bDZy2rc4n/bvZK+oUkIAOkP/wWA4/+9aJUXi/eyWUsJZo2bM
IMMDX3CdwroRhifuURmqwToVgzD47yPQ5wQMX0bb9gRfgiL3S0vuPwTTFXol+5B9
MtFOhGX1pwBwzDeePZOghC/e0WrS6+VC7nThlUv8iDwIuUhjjH8bipInlDCdIEXh
9OGU67ovCEPi62LxMbjjKUJ2F3RGch/5MLeYYVYsU0QtSlee4VeZVE7sepvKxxGQ
oRpWkAPrIIvpIslKsqG3q31Qi+U8SLRwuuF5gOkffcanY7CWeqoJSwWv/qBWhSw0
ubcX4rZdRK+kfKBTJfCrjbv0kd+fPLgzM6BtkANJ6GDDcTkdEozeUejg2wjUOvTx
Q+9dgD/sfVPriQA169H1kxGyw0WCIIjUqHsqh7HP6yijthX2mQIebnHRhhQlL2O0
B+VyA539DYbCmR9GE3hcvAbgV0uET4NKCMzmwPZ26Pja+hdqhgK1xyUtx3u6JI1N
4gJnGEz/kUggwlQXU/134nw8ZSx6VGiItO4KOV2bR6NVGRoz9Of/W3RUpXehKW6j
pFUJP5hSkcIZL2cYPPUPn4Ug0ycp6GkRx/CKcTH+w78S07XbG0eU2jBtvypybEBl
TPpxJnKbq4gzuYf16P7SiPW0mzEliVki0IjfzS3rS1EKhbfufGT1T5pnpPD+TdYn
dM90hW2BzXOrRafjF524wawvZA/8aDpye7Zoc/frKNtptFoje3DLhKy572ULtuGz
AoCHcOvVETi6Aiyjf/BB9eoML5VqpAiM03XPJW7FpJMivuaBPgtU5EqRaG96fQka
Hga7s73a91G8RCdPPtb0A8IgmwDD3VDY2O828ivnqjZwi25P2GwL0BBycN+TegcQ
g3cpUaEWZsw676ukQdfRFasvnrutf0kLz6HkfwOViL0QnUwkjFkcIM+KGGOQ5xdk
8WOS2IaorS7V3v1JJfthq8R+xmw+qFm+DM2B7Wt+uShghZin0Bn31y663aKSb3CH
QMP32xIFTrfVlwOf3nFz3o4s/S/So/uBI5a0a+d49sggT7pr/0TuVLBX+RC4BwSn
D7lS/nbefDKIWhqSQ5Bu/HVFIwu16vg5o6eqPOiHrYQIEx3OGL4caLZa+Uby5VQi
f80zRygSFEtxTwfToVbaj1j6U2A+e8afB/pjycdxc3VVxqTnMRCccIyh8zJmZho/
TwRs2gi2OwlxjTS5E9dPXn78pmOpySxdIcloIGgxKIVABTJW+FC4aNQZ41r/BXLo
wgGa9X0BF1GlLVnHcZeOKe1fVHg2s20ou8CiR4yaytsBGjuQnUNZfN0SNpknJ72S
mvCtrBxT+IMo6xxgm12IMWBr+k7RcNQq8zfp8NWFnh8sNaT0PR2KOgaHGeLVG5bj
dcOIDQ0h0idtD1o+wPMrc94sBmmBpTwPoV0SKETstOamesMF027Z5v3HRf1CqalV
TxRs4MDZPOfX3OwUuRMysOjEXySjG0Vcp+uH6sgDG1MICTnufshYfAlF4PU5mOTq
FAFfCGINXA3WvJEJivft2XP6UUC0UjbS3vxWvYD8GFTRtCNzHB8tTF8C6yr+CXoW
lX4OEAOBZfKeuLrOiWzJVuk3QyFL3BdjTYhxTl4fXsym9UEiu2mYOTUAZgEhVFCP
WSwjrzlfC6WiOiMCkTONGWAW+9T3B9UwNcBY7GS8vMr4oH71bJK5xKJBc9Q+EX3z
6Ou66SDG0lqKI4n5wiXE3bfEjc5Q+y0j19V8WOY+Yl20PUbyvl9F+XJd8ufnmq0v
n+3p7rudxJrnVXHA1QxmXXnQ6vy0fIb1ea0ibrW+bSfHshkWOAiKXbG+Ue9miN9L
VOYe5NPkUBS8+XujfRw+nGeSK5lMXADYW7II8qFoKKl7icI2iNFFJrWQZr0b+4ET
vh7R6sIgo+xQmAeriHfnWFTnZmnMIAEQi5yw+NQ7v/iOyJxlpKbK8HARt2VlS17n
Eisl6dIQwyS85kyPlaqEpOJu2U/UdrwMRWzwKOG8y4+g05zwgjrX3nJY97zCU7tP
6aGVScx+14x9Fb+qcZ0b0W1KzF1WfLXv7DpJHeLKHH5YrJ1iId+D5eROSCkAkXlY
T2/TcEfdsgeJD1iPh/jlNuDlMkUoRGi7SUTfu8mPlfW1LJh6LgvmmlnnZXf0MBEK
oUt15pFDrhpsnQb6FvWwnYOnfaNt8zzgyA+M5DCjFxLMV81NUKqqeByhX13v1W0Y
f4bg/LBnkcRzOBY2O+C4FL6rzIzQJczkW68B+6fuF8V4cQ03Rk+pkso6NOyAJpIC
J3/U2Vq/fcg/aBBu8NesfsyqxqRhYzWB+SudsWU9xErC3CGEwacPmX5KtkkFrcqU
XkmlZrxQwrH0YVkg0wQB2P3Sk6Cu5ptYASMVMPY7A/YmSCKXpyFDTLWVarLs/Nur
N85QTpdi8gUPv3fAuvyr/dEtEK+4BcA0SkLxUbUa0jkMltgD7BbvhGnFpZbfVHlI
z2XpiYoGNlidW7LA4Ok9+s0bkJmyuSXbXHOJ05naDcT2mqtts7FX1fVCEKE479N0
Ko0ZO5/sfIlhLpPmAmpw6Eh0mf2WifGOTSFUaVsZ5+RYbVoClWkGXCNS7nvxlsCu
Bki5KWgO6mssiLIjDu+20UjIDhK3rrIYay11XoQpGY8ADMFCz6qWvdUuzqvzh28W
SBoRJPA2OntrgQUGlGnbwXi1zBCXPvul8rlPn4/f97TOZP+dB6Xy+hFmlEgXtum8
i6rytL21Jj/XEAir2XaZpLfMqMTkH8Tfr3oqnSiruVdQOEcPViu5zi91SPYWjARm
u+MLLSVU74eRA9fQS680K/lk0krGAOSqfQ+FIVLeOEN0pFvs/rKJH8PmZFW3RGls
XzAg6MIeRf9HY3QSGRc+SParvrjVvUETezQm9zlDCrE1BjDvIC2fLpcsgRWZvAzU
hXITf4SsCG69Kl489DZsJeJ2I/sjk1SamgtNSFU/64ZtWnXGlBTDbhhh4TXb1Gx3
TzZU22H7NbKuso1MAqdLcf5QV1CYtvwNoTfWvlJAl7/JBDS5IN6Rh6oRaTMWPgch
2I+FvE9Ok8g16RFZ0irwTThXxpqRJ4Ssxc5YE5HrB1dI8zJKhm92oZdU/l2FiPV4
VIHrdIDjg0PWC0Pz73N5hY+CUUDNMttVSEcW4dpF0CSXqCVTJF1cyXXqnILZjlJa
3Gz/D/x9No6h+nYpwLn35gYOWOSHmR2fPinlxU6qCICz7RUOadWNwoPfNqxwbHYu
Mraz9dDSFFiJaEvcVVEzB2FR1h+rbYtNww8NaKQXTzEE8pwIruYeTdN/ynGgSdZB
8km996HkRK7/WqgXwGHl4CUSiVs1JTEkK/YMJyfejn8J+lGcSUF/mRq4NPnJhkUq
3KMrKHzQi4QHgwLpwL8TJyYdfMKhXUxvezBtLbUe0cOzgrSozPIpFthTY+gRAedy
Qo39aFubfOOId+iiC4f/tM2vulexUj7VNmbBeohkpCPHbyaiExqMNyWnIEt47HvA
Kp8gKIP2i8kKCW3Pf834YA3U6Ret117eCAGIP4HxmAOtYvyrdKz7dHg15KpVu6eH
VvG0QiWqDTdARbThv3PjTw9zQZN2WnnSEt6FbvxKiZaX2DCXqdzXLQcKWkN18IbW
PaxhUp+mfbvwcr+ftqtOGyKQliLmjvSTwGe7xMr/izP4EAer4W9Rq4zPTS/iclPQ
tPJfF8lsyp8jF2+3o+yNLttW4wOBSkTQWVhLd1wVIy1+UJK4dPbqVIVzcGbQhSsc
LNwbiiwGGYPFpPRGEg9InvMCSQZL5L8OTpJkZ8HSdLhl/7GKVDyPwGX5h/Zygte2
jYo30NMMqNr4GtuvQi9SkN6EAXLArmB2HiBdTr0fLqpE7V2nfrW6YZRcIRIUkrpC
iz6ekOkECUotyVwQNojXvujgARvmrBQVBEz4cVlOIqKaPAQs34NMbDR4f2K/vt8P
1DSm+Rgau0szM4K3u26l1CGHQ22gXiPtx7Byv8GXuS67lnAhZHGjGPqNxnnV5yjN
aKSzIW+P03l48PzSkaq/Pls55tIgD6LLURN4DMNPDX+FLfmzCDmNb2NV545ThcvT
OUBx7VHOKXnthYfIHPtu8jCCu36+XJV4DBJ6VgLrDuSTzMBFyQM+VsxtRJFE2gF0
RwpEmvH+8IjVdTXYQZdNUNPvy9lrgNReGYQhwzCuFjVeChubbSnipAheeM7CfoNK
lLOK9B0RGhvtTTCTc+50czfaU1dBmbqBFQpTHdizyqOIz0RMwrhlZ9AkmhdyVK4o
T4u8Pd8GPUm9Wh+rJic37F9rgMbkE0uQVSl8fEyLb1Mh8UrYdYAO0mFiKXaZTNPb
4S6HACCgG5gK+ewulZE/QKm//y27xj2IObGJDJQ1W0+VAIVXILDCbPlpvDmUTcBq
H2pb1f7DFlkUJvzl5j45UhQ9S6ZT+QP93/DvMSjBU1oiPzJbXHmX9/s+w4RDvB9h
qt9Pfxg/lGOcCHGupvOShb4STTjwhSCJFMXFFtsst2LSoD/rtFr0nZ+KeE+Onnsl
NwV65gTESDRxqKq7PtrTHKd7dOsEizYbs81+WcwKdyUBz9hMjStIKwWN6WydPuV5
k+zQgZmQ6IF2xnVGWzD65phs+k6b8v5rKt15CsAGWj1m7UKLsGAjC8bwjC354E6R
xH3ek2FH6sLeDz4ir3UsIrh3ta7kCnSwmMlMHpQ5vWRA1vqf2tFS9dMqROoLnMPN
L5kXtpzgUUkpxQCtVBUe7juKRzMN28Q3rHEi1sMWXnNHa4yf9t6xCf8n+nnIJ76m
WsWObVJSrVRzaYiOBmDLf2stHDkkQGO8Vq7Uy5Yqb55XXSer39opIe/IEikfZZJn
SB2R0yxdlePLxmpKaTX00pM6c1CeMNf6ehYSzldB940ltPdbqV7QUP43vwHfZP51
GmrOCqc99SvnUJbjjx0DkKZdxoYYIZauNx89spQ+e9GWEE218I+wdNv6HP+Mq9ba
frx5ZqrA2tX6x54C9EJfezzzzAXrXtqFfUC3SDR+c9DYpkCcjvYGpt1A1cSFTMcC
yEnXk/gmQHATkuPy0OwzhQPp34MVN/lbX3GcIqeQESO8Gc9jzTJWZ41mkvVgWaJP
JTjBtOGOhP0pEd3pOfzTirMxTpdgTCMR5qOgc399RzoGVHsDeXtq2Tx2ng1WR561
v3srJL22LaofBlH1Q1w5TO81MeaVKA5ESDSnpBtu39b9krp8O0EpR14uDgEUnpIw
iENR13WesxPteza9SFX+yOTt7tPj03CtJcxCuJDAnCM0oGEQ2NCvAsStSbYAtggm
my5f3Ue4MXoh/dWPJlY+5KglV17Ld4MdGgZqFAaQ8dV/Sfj+7/aD3pS90TRnK9l9
WEttcm5JrOnYubSC3lj5UHDpgJkL86/DD2UpVRcFwiQjx8DkYpGF1eGN1a9kvSgA
tGHXAzWyp+7YRtEL3T3q92Y2UncMdp1fmR4xKYDPNJdSnIKAwKi7dQyPxirG3kdd
+BRVPrvWRAoc6AzEtTqpp4wyXUlztfF6hxJ2S8keJp1kJUIY8UlpvvJ+UJ4HAyfF
SkflajKCsJqSwcAWwsidYeR4rD1Oekigjhr+X10lkAAidZ8wY3aopc0UykiTCksP
AT9LIKaELB7eKQbIGbtS7AWWOSAhYoVcR5GVyeyxZfAww16r4xMbU/b9g5IvMYYW
zelVxrwR51cvEte08S7y4cxEabBIphG6lVQgUuwMFWXyi3eRjZfLKfG3sLTvbYmo
P4ClFnhBJ/lB0gf15IBLsMuQHkJTsuI+VloQacR/cZ7AZucmk2kbs5/hRlMiSAWH
WMPKTAag1OimTQYO2f2DzRaiZSadKdMkhHQvx9YclbfzF4ij1d0eyioEgLcEOlrm
1sZbKP7PasI334MItfTjZbumd6hdvKY8Oy6FIKGf6YYvhY+Gv29QuIG1IUDwfcWW
w6QaKD3P5fYmac4QiKRIOCWCgCDYevgexWtUfvx31SA3UxcDkXDNRLZ8Kmf+qEjn
I6jutrA5kldIgPMPb6/QC5FiScGPcfX/Cyi34Tis58l1ZBky2YNJgJE8HfOzJpDA
UINKne4AIqQCE3Ts+03VvDas5RMVPVdZPyk2ds+dTOmfTTX99dAOkDzxkN9z/pr0
e5rbD+EMUNDoHQS9c3REFcHOjp/Ms5LiWbTe3fRSBnmCCiPQHNkm/a00YHgtT1ql
sRxyPdYYEOv2M4suJqYFppcqsznC9Ci0gHUtg0iUmAVArvVnaSoQGrFTN+DZg6Gq
+lA7M3TPIQb/yhCiXXzi7cPY4mh7YBx53a2W+axBqZd/TUiLi19Vl3sdubpTVmCS
uM0EntyZJ9BOnd1sWBjQISEApNM/sVdDrNoXDN3XD0gOK3qkVsCeF2voWvC+QHIq
jpSzrpGJJGnmbLT99gRh2NWvkNWNXKVnuqTGND+ZRVvOywAIiakU7LEH0iuvCMpR
jvS4jTzESYw4mMNIoMPoRpFlrzM3BW4ZgR0xSTDca9cHTA9WA8ATlZgLriCj4LeH
5Sjtb7qahk8O5sZuJRs28adFNBaqVYOA9wsZ9qRx+lJu/eBKsVQSkN+6vXC8AE7i
6AZE66LROBepWQh/4RITl2quTE61ZPJ6534cZ7/WoTZfGyKfaG5fJKpssv/BUTtu
l29pXjhL4j3jRqk5a4JExSPlVu8cOdUKij7z8Ur7m7GlJxBHDUEzRTy13s99OvnE
RZPbfC3xpna2fdOn1nal8j4nPATn0Ev6tLaGFwJ8Keal/3Ec+/EerROf6PZmiYSv
3fJHFjhKCD5nx6+beRoTR6qgLs89n02EQke3PvhE+ya59w9AztiZ+AKo51LDT85x
2ru6jYqjSvNZwq7P1ZrsxX9zIyZel0n0jNgXYJeo1kHiWZSJigxinJIm672Jo95P
Feirc1RF8WaSj1lAczYKkHTq1Vw3EIYXl9huHGoWEUrC+hZj60cIJ3JoBXUsDnJ3
hCFsx0sMgqk62OyP3PsIwUR7wDC/a9b/qXAqnzQwsIQyIEN4biH0HWlCvJlqW0Pq
nmcM0GXV8jNDhTr5CRKhX7+B28tDUHNNNwvTMv9S5syNrgLWYK30J43rop8mJkL0
tYYGJSH7uFOVI5pcJewOBWSF+M/lav6sFYDYsJeB/mDB9RXLkzcsvaVljm2EycS0
bgtSLYswDFaVvOE/Y2hS1s1+XOMeKQlnxZ+KFddboHmPiwP09odAD5Fk7nn6FmRU
E/tTUScIMIaStRX2/gp8z9X2G9sJGVW2KpBmRCDLztuJrJSLM10pph8j5zgL38dG
/hXwkIIQmKfQUPJe4elSDCTswV3DkUVvGrgtBhtNwAN4B80/1CKK9JuRANKOjaVe
53UPiCFO2gpgm45TUKx6br688laVxCcNWNJlqPEya+/2qlI5DapL3VrTRhNpPnvE
ZfyOOaNB4AkYHSatqiB5d+moqxz1qob3d/h+hRuMgRrBdkzzeG3F3RHsVJmxF+4I
WtwwtXqXTJ0pQ4PTJNg9ZsZy2UnTupDWrDK06ZkrDnhzNnCX8Qwovo90Q/a/6390
HpWCQ88sD2qEjD1gLOiAAcsh92b873ssFQ9WGgSNHVwa5jF0cDFSCLfqYIM8cTke
dNG87hwTTBu1fU4x0JItqNDHUexkgcwEf1WP4jj87e/qXbrXZt0bBZALjkUL+vJI
J5H1yg+tINQGxDKA+O2UkNI0pj6ZcAPU8Xs2gk5PKrOrBtRTI2QnTFwwrmcN9u1M
hCzda0qWSxSOIDvWWX6lY6UtutI+HKfi0V51REskx75x4ONBiaT3MaCXIDyco04n
GwyuAUbU6wTwN6zCIkWkttBVhNeDc0CRn5Crndkyk8DBILICc0kRztRgYV0txRz4
MngBGSr3RNzJUQaEVHiIpSFvBe7aiqahDZy0A0ZsPT8SztAeqaxIaBU1VDnxGV4+
h3/ly3BPPcKJGxJdxu2fTmsaLNXkYOr5yP/XVW4XCrpf00edqCHI8NJco0aRClmL
hHV7/2qTqk/RJERLN/bDBZYB4SIka1lIj8p0/kukGCMgnmg8LSLUrPOmaHcG8zta
TqC3r1N7m4HeKYgO5yx26ZrF3cMg7QRhdxOLDK3F8x9svGuFc7EuwZAR1IT8CII4
YTzYST0RLHyawG2jEiT7wLN2Jy5tPGcvrJRT6uI8KUUdrTdpIG9zzcrRlHXHXScK
K3rymLEpyYt30mXzUZv61yoDD9jxyhnQNqtkYzEIIVmWvcE4frBvHs8ePwMQ7eOI
xnngJkRZsb08i1bJebP4qMedeYQ79FK1zSJmwww8pkGk5OgwUSPm94/LjgxopYbi
omdONO9EcNiDcdWYSBCHnUypAlVLzURP35qTxcM2LS/B0DzD3+UZatiKoss6v7ju
U5BKro44bZXlHpwVb23W0P6sACa6wW5itXDF2dqYGr/F6tEJnEtOk49PAZM0+8YE
hh2H8V8zbA0QJR90IPPMxom9KzNqnurlfbVC30JJAgIUs0wb8KH6K17z/9zevWkp
WaMgs/+gMwBKAKHE9Y4BUxPEznWI0tCQFh0rmKQYp5pgEjscso1zTgS9ybIpU2bu
z8Q+nGmolDg11QR+zZZLAOp8bbxDv6D2lOjTFGNYwi81mQoIUJ8hvpdkR9Qb+XLc
7LdneF0dtJ53hpQxSrtYSN7cJvgp1Grq/hN+v6JpyLzs6qDue4a/7KRDvxMsjsKx
Xem5ZivasvkIfwgPPJqClyDTqabvh0njcq/CDIdvVAlBtVkKMZQDOInbB2JssoQ6
BivlXtreUDKsUxsRXD7biG5zF3pEgmTUMg+4JnHpXqahd1cnvdLU6EQ/+OTSkbDa
jS4yYF5HYpBMd4eB1VC+i6+Gw8OtOKzOm/U62toYPI4wnZhbesLPDGDw2Le+HeBn
jnJ8hwbYCRd40pzrrdI7cHTFfTfjaaSJ4h+XjLv7wZuLvn2UdjrQLhfFhOdRVFPO
dX5n7R5nBNByj6N585mcVu3Q1FqSBJPmuzJheC3ucQmVI5p3nSLqGEfXnj7w/aeQ
fQIXf9UpsEzO0/COlh7844fNEAZdZFlvq3Mhs5tin/HwRiFIPlBdaEmMEHkyGZ2i
ag2hYcu0ENBG14Toq4ktfrR9BwrRhlZbMuasBdlYxjN5PYV84gTvUUp0Y+1+Wn3v
pdLNUlIvUG+NpxA9SDt/zDfJskX/LpMiENFtk7G6bcgCdWeXlW7R1D+A9FKf6vur
Pb7xG4WWN8isdUxn6XeV/EaTF6ZUb7NFnllImlagi+vkzoZ5uqhyJFxwP9+nee9F
6cheWzsA0PCWJrFEYCXbtH4LplaMsqYAh4tB+bLay/HwK/34/glO5wyihzKxzCek
1I5pnEXExscON81bZ+cecrrCdzFGlk9M17EnJSzd5kv59FAfbIdC+OcYeGacJJHV
s5mX6POzEXAXfeDG5gEPqeuZcXjunxamsEQkFRTuVBEOQ+DEgauFxAS2RUFksqLc
T2fDF0fBK70VbcUkxpTX9B2h2hAXFyIxxkrMSzlVfma1WdwpY21YAWdnYzNHDA2j
0pJ9DJZtM1gD4XICTqRJ9xNDFcjAgvlBzzSIeyHsvBds5yRtj20m3emLUA4cpIol
CMwIhw1dLVKohGnOZgRARGy9ufCCyu73gyaURd3FfumVJlnQ8Yq2+JqUGPzTO2Ch
ye/8FDF8QrSXAi1a3mZvDUOqGW5Zs0Q29zvZzcyCRo2UoAT+SpgCJvibYRst5w1R
TkbWYUON5q0ix02eBnl2o4K8swhoSmSihCRr2rlhByPRfAPD3dv5FQJvBzhmJgRq
TAtmc/rI5rzdA7QsUszsPTvo+qz4A8CXqR9d/T9FJe/dTAJ+MVexI39+89EPS87r
1rxgzzDr7kmNnEMz0jyc5lerIdUGMq7tTagop/bFOX3S9KllYjO5abpK7ybhZgcn
XX+oOwZOSru0xSu1pkFDxntm4LTJy5t+xGVQiHYJuKA2bVO/te7RCEkyguzZQuZc
O4meW7xETC/EY7yY7skaQbHZlI273oFaE5qAJg3L3JnNXHu7lyMEDdPwsShVNv8y
Q/HFmjnYBV3rVUkIv61rBFV68EmKZNR9wZNRHeijTPFfAXLhu9qnBbAKg1K41jbQ
eKzIbzEiAkHWjnwTF+5LH52iYNZeUXvvTt8wqs6XqsVsnwHAiTy35GA/B+d/PWNY
ddZPPr48/LFf//S9JfzxZn3vav7ChW7tjCl8tRNHDnNvv0lCYNDX2PB4wJuzU1Hx
SchnBpRRbh7HGu94wLdZwNF/nyVmgqYYwrdnnM/gsr9S6gzZfZ4ce+HY3nb4JsGl
5QnRhBelYRzMOYU/L+DmErvAjU0os2qUfKcE72EWKgWRNXH8+4xEr9gAFA7pGKez
uNx0/7/AlAGAJwnb5aJ4tYI9Z1lMB1dt+9Igbgl4FC2+sxhFd4xAZfNrQ1yw4tVH
F1XcHfo8U2HmsdWjFaVd5TCEbEo7vQH8t+uZPvn9WrOjbT4Ru+5eXPEKjjcDwYZX
Xiv5ij6sN1Fta7QU4kbgWElmQ3SvysXGLEsj37ccJ/fKYkOkP70Enmm1h47Phvka
2yd1DXsHtgbPM327vKWswrxmecsoyp45YLihHyLDWTQodvyx6KTkv6kd5yhYn/P2
eQWo2/4lPFpg2RBoI09gI7h7K0+gl6CJOFPmIX/msrevnq2mXE3W/6kYCkJRCGN7
ZGyMv3PAg1rIU2Ev82QKCpSdm483jcm2AgjcOFFACvn35oYNAvfFQKKw96sUw2zN
1y58r9RUIh8GHnGU4v4dckka6g/mDxvcRWkCDAhyVXH9vO488OIrjov/Ppw209sL
W4dWQ4WWCscUlRv4ummmcnOnBWA7kvFyzliiKAM1rd+JoR0x+ab5IEk9E+qLobMg
t5Yb8b0mFRKpAu3Rm5LBDxVGEBjTsLM3QPgCAiQLcJUNXSWm7IL7ZriWT3WOQrL3
pMiXTb920iaaJkzRF3tp5wCmUMCCv69ZXDfQctCrPtyogADdlj6jqr/pnPSqdOPG
alJWyQOYzNv8GBFF8KrPUIPKhevbydNptOu366xodZnmAMj1TPzQVhTeTuq0gkSw
m9foc6ZeVHe2PhdDT1OkSMaa/ka/82dnVEPrutXzrKzcKz361HF5+gVyQZWRi52e
Wz0SrbVy0ujlgDALhDsJga1XIVCXcsQ4/5+wYdQD8jENfeW33J0BIR1fTQ4HAgJQ
TIBSHiyBiFPFD0nc5K8S+ZHAEj7MGsChqOuhP7WhRIuGl5CoubvrGo6KUqX9dsa2
uyqSVIqEMZxxflUqOuF9p/eCNH8aFpnk1HZX/toktj1l3ObcYbt8pYu4t0147s+f
aUcDIo2D0bQc/AJVTevOzKDmp+lesyNt7HrTbM2zYMF+gFJ2laopNjDdeKZxwVHh
ze43svzNRAXKm08GytCuogQVAs6TYfflKCWxPllXFgYvIlXUCiRp7agfcEUr13h9
tXtclk2pWNv/kWhPyFKX5Fmxe64hXQZUKtEZUTeL8zBCgcGzp6dNMG488WC0EME/
w5kgtwrV2q9dRAXmhHavvf3qALdOkDUzQdGP7PcoEyuAngVk8y0rjg8rLKvZcoml
2F2clugPok5cSLS6H0d29q3STeTfhLHwNDpvcwB5F2SBr9KOclaHdNOO2SLWj2uh
Yqvx0x730OP2wre+VYX5vLm9LYVQ9YD9YaHe7UXMggfKkalYJqhvRJKh+E/vaUQ8
2wfdv75Ii7jQEgF4oltA4loFTVGVPKG4TDdI/lrL5UOX8uQaVHbixxgZdnHGOtMw
O4wanMSfM6LCKczA3BvAl7HQvbKsw+A2cCm11ORGHA2zyvpmw4LGIL4Xi1LtRv/+
40RjeOLittCKQ5KQnJeaAxztOYr3G71KMXk2vbXpUoHJal6aNJTDmGDmMz36XENU
CeYp5RlKGFDwx3NsTixLG0gc6eQyhlFsJTSOxArqwti81hWJ1PQ7GMVonPCwDGDz
oAjGjcky4ipAFemEI+JCVTnTQxqC9q+No5il3+DwMLTCzxv6715HNtgkjNLjeEaK
S5tlfha2bhIo8gT6+J+EUZLiqia39YImYDA49a/SwdaW9dWi5n47vTvh6FMKUQFg
DXYLFBjxqHEffiFl9WNwqmw8LhSKDRDWnSHeyyP6NoqA1tW4zZP8tGXA+MIc5uEE
EtgqTOZNeu+dQ3/c2emE0eddLE1uYjy806vbJ3iNvPzP1LZm7fTvWMJYjuoRgPkC
qNWLE5pSIkZIesbcmsr2EawDiH4nfdQKmagSXFxNmFup4vLmGT1dkfjcoSyzGJIn
SAo6i+zwLylJkqL0zAn62Ym+EKXRSD2gwVqDlXZD1yBVsVs1KkIRe9mEuSllxoOA
qzJk54U73afJasGxcNTwyyf7oOGOqbxeNM7Min6gA47T2HvA2UQvA727PSRwMyZd
2lQL3leF9J+q+HkE3ELvTJ3/WZaLsUYhIQUCEAVw20uT4oYJteN2m10pu6Y4zbWg
JM+L9OjyV8HGC3mNXrBpFY8AYcVfq7qwL9DKCnyzU66J5QoTJS3oNLoudtpzGert
7Gtmk7WjbxOpez9+4ltd3drkFWLUkd5F9DU6alDM3TEoogXSV4fhvVu5Kv2cQPLP
wKAwl1VadNjlGosJb4p1FEGpBbqITvaVFx4Gso8vbp6R7EtgHgHw88cRCbNNRByj
g3tAKmy5OszsTB18AstNzMbJduc8IMYKy/VK2JSqKjSPHnByOauIGRtPMjcqjYaQ
y8NS/op7aJVOQ1UPVAb6YXhqHwFy49YCi1eveLllivZa04xgEsnhHU9iQPUW36Py
qlriTrSFaTaOe/gZEknnXNSzuulioAHceOfgxjeBy11i3rahgO4NXLhLv/ujvUoU
UaBvcJMYrX+Rb4Z6/pnvCORi9DOdJea3HjtnTEZtr/CYKsxciXU8Hgsx1KsH0Pl7
s3IE1zEz4KgU2JXR2PB8Jm53ERRrTZDDLqVYS03hpcn4uOrxC25VFkFbDZ1GbS7A
/EfRBYI8sEZpLw7JFf/qLa5fPbTxAgGdVB0fSRLJnqwlss9rsBocGIHpg73aWfKT
LtDWY8os5AuR9yqoXIrmyYnwGbqZZzbUaLOVEqjjJgzg/xs2U43Q3Usp9htrwHEQ
N5YayT6n4O7qb/Y4DN/7NePH0LLZ9vGmFNaQzdGw5vIyPgCUYRJMutyFe6qU087B
BAuqdDJ7H7M91292UWztljRe1LezfgxovxSet37m1VBEeb/ODM5q9iZEc0645fln
iJqpWzjfkbZFcdHuJHqjR0GKoGc9rb0vesTTdeAoq0ieJCuogwJYVQH6ekadAfAX
t+DqVoWLS2hIZp4inb6z0JDU8M4vZThfY0ZjzbxIXM4sVx9qitqnyJeLt7Xh5TMH
5Z3F8wq23dvdGGuKSj28UNZhULNurUAsDP/WMstjuFwYVVc0RFqDyNzEONnXCcHr
6O59JQEDDk48c5b08Kotcv6J2IF83hrNCh2rywro0GV5faojPxNWUk/fyIWmbLto
f5yS4igi72XCrfSAgWRba9wTz3eHxaFsa6FBuIU8tROpYfrPFDc4cBzs8rVqouk4
5B90HnKi34vSlT1+oulcQqNItLJrH48ILrGJi7d5q94P++JraKEr2ZvSYl7pc31H
iQtl1eTK7Y/cBIRFFcCdjGwW4zI4jyfDrUIifsk5aQHa/mCqsJao2mHlcnzTeKes
N0nrnV9PSyfiosYqPOktc37A1ykAglE0a5K+jHTlY4/ghg7rEm0Qf4LKqgj/ibhf
bsqlUAn6+30PRRGbQwbb+FD4O3ztunbcxUU9G7bsYaB26rQRhLhQsfyj6DGh53og
bpHPUUjlTauDcfqtAE169Xuq6xcPnBQp7/U6Npjkh8G0/GWhPjADidmA76QiDxrU
njJebajwSuO8oH25xbkNapC1xbYCepDfkEjkrC1ex8hja/wsRCRG3WrhH8F/gk8T
OZUVfQfaCYnr+YJe44xRQsnB+qECJX6qFlAOMzRr5fwDBVFiHWN3/QDy9QqfQ2AO
bREs0fZBUm8aLfjpDIEhIi3x+cAt09mr1r+g2IYMCSKdwP2eEDCJcQjQzEbF/DK0
Vke9Gyk6OwSGMCbkHQ9IJDbeeb18Ye6frHfLHvruM2S969bHqvKHK6ml0OxjtKbj
AaSXEH7A0HVrudMUa0lNeWp35thJ/0z5SYV++CCUgl8tnHxLjto1o5CLHsRCNkgH
eKeDG3CA/Jfn4bjiyBrItJGHUo5zDNuh/X8eI3es3xxtm3FJHb3bV1SDQ4N0hODQ
FmiWA0qEFc0Do3NxNbynHCbiZIviRVLuVSVFkzpruewQ8qDaceWM1yCG/JNNTHlq
KRayE0iR4Qrt0ILaFUa6nDBOd9HH1nD8X7dmoe2gkJe8b+h68O91vad7fdfYDSKU
xMIChDRrWrG2q7D9GjmXbOXF2Bo41MSrBgzCp1AlyzAp11Ve2VlGQ/YGp2YV8r/Z
2azJLzP9ataYJ26JqgWYvuTp+GMaVjiwm46ekX6UJDwSKd+UfKB7vMcSjW9ozKYW
ENruF63En4pAwYJE/kik1mDvYsFibYNbRo/J0KkHfpLF9af4Crw1keqWLXp9/1Dv
loOFPJX55rTdIYoElMAUzG0PCFJygKEkVChgw4N7grQC9gSWq+Ok72VJqkKSeCJa
DSkWR4AwsOA8JF5FNobo+iquK2e7ReGyoJxZxes/CWIayMn095K4NugkGynETSFn
OGE51/YpM0cD13P4lud6RpKIilKe4BUqSn27MLro/lTbDXvwJsb1qgz/Aq9QwSpI
uHsRuSQKTVsWIUQZSe/32kCvJf5oaLc3I66nhUi+NVmQMI/qIU47PZucRwOLURZY
v/bCRFYQL5f91VTkU2tv/GTKVwhtk6K0V4keN2B2rNmL+OBBibzHbvXP1gU9OHNb
NW+Y50NzTKfQfqTifotx9nNjHymcwRmuLDlDfm1P2OS9ApuYC/k4T3dDcavCHFgf
DFu5LS7IRVvuc1giTUDUOiHDHTCw8D/JL7NeTF3zNbxpn9MDFWrMfStoL17n7bmG
D8fkm2axvNQtiDdvBKYVT2vCX2TW96uAPl8H5/uJOXRHnrbo//6moCQNem0656la
cos5uItZdwvUmsJttBfd0TZmSk9xI8DuxL71b8iCa0uhtna2qjl2/2kvDeto6d58
qB2ZJziF0losCpMBDWLfVhHTAH7BzKlAPM7pxvZsGmAxIbzUUKyNe1Ox4mjJ4dzf
f37UfC/Gl2YLPn64fPLA8DnCtYOEPLxjH7fSkqezPOxqnLXB6c+UqDycgfBqez7q
gfVidlKrbIHaAH9NU57m/e7QKfwcMkc5lq5cB+GgnGnb5qM+QTYxSnerjeHv3CRM
whHfOKjeBhdroZDWFnt5xSMmbdbgJpGbBvatG/YKm7+9lDCkEaTMCqdcR4dVE8HG
BIDnt764O0E3fEIo+/79SfbbWt308iOA0TccFFX4S9TQTiST5qvrccvl6FPFMhtU
tl9z9hPEojb8puNMFAXj9hOlyvYzxmxmnf/YH7ULvW1tgyGsh1Am1oKAuD/H1G+I
fxPnSSCOu2vfUsPAGIfloCKqLanwaoANzBTnuoRJetSNa9DQMc4dBtqvkihld4QM
LpH5VBhBeQn1R/duz1kakoKvyot4+XweNPmfoRyUqb8IBkcG8OTTlx2yu9l1YN3v
z8rtByu1+Bw+dJIcFwBo6NAkFJejdbLfnMkUrvW0KbxnUmEH0PGg/FPPivO4vmsN
V1+kUKrzKlsNi8/k9CehWOtDZwn4aJnkd1G2tFglVXKXcPLfX4F/yZG2uUQg0iTx
kkR6j/8yTBVPhpzonP6zYEOcgqzmFc9HCFRpc+2fa2v/mNlqinvPkH4rljjOQENm
pmHrGuFOW56yG6UnIhkOqbqegzNiDO0DM+qryNYo0owhP6NPKbvkAQABFRoabL8R
3RiznaGVlMzMJOn2/ZwY3eT7DP/Mde/z1dTJXt9HCwlmtIWDmrnAS5MBBVNrG5AM
mgVAm/K8R+nnULCrDF5XC/ZTXacAz+9UiLR/UFJ6FkVAwjbUIqfOdziGvQjq9AlW
BqIxd0od8yBc7FeBr7zliH5lUNVmE8Ds1xNv1aPZHiKWgC2exbTQKE1WzLqGYlc0
ud3zfOVc9SkbqBhdWZpgz1HFcaO+y//q+1zbdMA7myHzrlcKRT+97Q3mTzjWfc+Z
7TCC0dfC8RdVqwZ3qk/AkFjPJQQTwRZ9dSoUhgxmMbEBiU2ZtC7NGWuCPaejtR6/
QKWia555CBqtwxEkM8t6yMjFqEtrrWtoY31KxqfdmC0aSQj5O4tkG+KFwhzJskSa
t3y5VurkGrRKgWjFriy6T56ZzcfEazd5sWWy8G04XXsrmf1IxZEEQCV+8DoCMvDL
914Tz6KXy4kK6cC9t+8aiUToP+2mZF7WdzSunOXv2182P11VbX43SZ2IiihlaWvW
pHHzB4QUjoq/DqsQBo/5O0nWLtmmgd+zCYMqOh1cULkKMf6zLJr2wEftsZ3kRZKB
ngP3Bj2Rl6lIGIn6T+qpqwMVTT2RI6BIOkccQFkN45FdkFoGv0PQ5N1O+XD5L/n9
UsnLr/0DbJ8oYN8JDa38PMJOcruu1KdgkrgeG5fKleFHLTzK+8qGasNdusCozHJP
7WxfV5pMgWeDL4jNlnbsGk0X29NwEXymBd5oUN5dqwefpLuDyzUx/LKHKtwvJWq8
8HVWanDNZUkGj3EpURPKxOhxSUErlEFQw2uJL46SO04mrH92ZCCFJV9sjj6TkU7A
gJE0umG4eqlMk9ow8Lo+KEUl8jhvwS5yeObkElw9/cWkXwKUrSj7MEpwiXK9scZP
MD4f/9mNeOol4w6HlsHd3RILVHZXC1aaQbe0U2C4dZorrpvVfA47QrWt5O+1FytG
h5gcjoRo/URqJUTRw1GQhWVVbLT+S82ZZ53sL9kZGpsvCrBJmcIsdnb83uqy4jRk
reSn8/pVulcN0riLJ1JcsmdlKI/VU1rRgOHFDFWmmH/nBmz4t0J2XIeuvs0UAkBu
Sqyt60xZ9fOWxDzowRKCFeo6J2C0q2StK4JTqJ8rM2W0cn46GZv2mhSpUbdD48Og
uvQGuMBaheizJAorGMpuA78cGZLywQ9DGufmR5Se3zXEw8lLUIR7yi0yDBRW6sJ2
HGCf0uMz8zbchZMjlvXsZea/HH/M5cljcWxi8i3q48AvPklXVz1yZSbOdyGyn4o/
WXwa39YY/DfAvFm4EOUBmPNMIwP6mPI03EE+jFt6CFXk1oM26FoTdAVlKR/G7fgt
W9id55ZhAW6qKOYGS3YuhYDA6Eo4Vl8TwSjHyarbC/jq9SHeqLgSphZVROClqIcx
huwAH7ciBdn+TYonw8UMsCYSWpMxTbJPAOA1/KBK/85nvy5ekXw7PF0wgRXxQEIr
CENbj16DRfuLkZoPlVicsVpvxcraq125HThyvJ3G5lbEX2WP0qwNnPU8Y47s9qVG
yoyORRUBM1tloG8XigTKhlwLS3y8YkNlwJ9+jfdwZBWBmCka62XOJdMr9WQQRpFH
m+n5G7JZ6MA+Zo76CmHPdfsgp1Shr5D5N0tvTx2y4f/MfzG1avLHiVVLjn/g0V10
EN659RB7H+y/1/sTxM6QBx5lokTb0INEZJichJqaLzUPt75zLc1hlocjL0cVWAF0
QfwL16e/9NkZC/4V0L1xGjT63m9B0wys6cHpJExHHPhFtbK3Ec8BRRLqSTuXe0Mo
lWEAhf5AwocaCfSbu5L8ZJJ48Tk5lZItEnpXxIMFZQBNOEyZn11wxBdHmS2ANxjf
houRg2i64nVz6KvhEAZkig3uk6VpqL725hHsfUdQ7Deg3VVJ7o8RpHCs5N0jI9C9
ExGMBXnCFr2AzqK60/dvtP6Wy7MrcfbuiA85Gm98JhgBOPOC+SMTQuLqfz4OIkYn
HwX6I0Sfxu8U4HRiz84ALigRtn2MfeU9IHZJH3wqFgZ3btfR9Yxy9zEVa/tVUMu5
i7+/maZ7VDMuVh1hKpU0O8JtcX1zi0etmVDgZk7F5alJ/sA7Y62lvM7upb/suzMw
eSa44VJarACiZlAkoG7wFr+kRrPIMHKkaBJ4DavluTQuFgDDqwl5tx4V+wLmANpF
GjtB+6yrS+bkq2EIfWiRoBzI5nnoqIdkxxvEQwMddmieHsBUqA6y082P2zy50tXm
IYUgUK/obd0VkR/JqP7inT+d9b5FfS39OWfIu4PAloCXLxIV60P+c3VgZOguxzSJ
28D/MfL8lc5c/KIrHCAjZo/yrApOb57XD1HcfQ/aDlwN83lMy2KyrXUfGErhb2X5
qhMvjUzE7hcHpUVGK9Hk2k2bjxbadzLtO8HOz31kj4+fV6eVtHU+5SW6B90Jw9RE
N47WaRcN2tmGZ2Q4YZoXS2np2sHa54c4mu0poElDaqBObEXRNUrcxbmU7yAehL3o
3OGrqzeuU/j4nn35u04lFPsXDEM2P2dgYpaEgupn3TwXiDH81BQpYsH4EBs8tVQ4
ZfgUtG9Ugtd/DlU3KxcHGd26Isd1BCuSkxcPG86QbDD9SFi+eUlrVk7hwa7O2SMy
Z+gNHoS8Wb+pBKWcTtQ4n6kf1z6FTvGL/Y8R8aIy+sbVXgSsHH9KhMLtm+ojnlm4
w3BjFTVNJxEoRkZMh2BGkPrdq4GDgIsT3P1Ty+DDmAnlsCn5TWBobJ2rv2waOMwp
hv7AWDE6gPBn+7QJJg7Sdms7knyte+hj+NYsHGMtIWUCuXf3J/I81c+GTUGVv2UR
EH374Wu8tJYHVOCN/40f//cE8Aj86mpEaMjf/FeAaR544111QFo9oiDEuaYtY8xq
/RlD/47+eZGW+FB8f7TEp1/c1GrtS6c7FP//9+JWcY4vc+hI2MwIUieypgO9e26H
EPdmdwJQxx59f7c9cFmkJlxHcg4d4qF6ARkWZSUeSKl8HpqkAwlN3rqlQ8kP7+mA
ZTOwXx1FC3n3h3aHxigOJ7hzxlbYWLPfpdb5ocxff7HPpf3NFRFqArIrr4Rq6y7F
11KuFAe0d/2bKYnY92frZML2Qa2C5zF2q+Lv5HaIMm3uk7/ofqYNAKjeifjBF3cb
1K8oWkm7HHwH4kKR+ytldDsThmoTKwtPbIZY6m0pO0XZw9hJHiY6qlw+cO+mJ5PU
85QVXwMSwxdeaE6mGK2MmZIo359ckkFOefz2lkpE+9rTTMOshHM0omsu8U8V+n4d
bXqvWmXhOa+DT9ImEPZaL9HD5f5DjaCNitMaSb6KTFL9Rlig20iNLYecI8ItjbXn
ZWQkk1Ixx6hMwAlXlcyQ/AGCQhoPHULgDfhGwEKEVZNbMxgrw6xXBxMrHkOBjd2B
1hYX55DSsAC31DCP1z5gPCVRJMYimu0d8/SkvZ6Ojr5cqDhiv7WYRfpyabYDdbnV
mM8OffI9F3z54Y65vyiQfSG6QBlezo59Z4nFa86STqA388BWg33ybMKxrD9cBpS1
NNZOk0mEEgOp46rg0RLPmUfGK6EbP9aMT7+J+IM7Wemd+7+R06wz0d7ovMz4rgZT
JCdYMKIZt73GY/md8KOaE1JnRpPKLGrs2CgTNs1mOxmIejoIDXEqDfzX2BzYYqvj
9+MAoHE//3uw9AmbN/XqXfrICL2JES6Cl4eULy2adKUsNRIrrwlajV2fl7/s0ZP0
QvGU6oqSCest61eRR4b88lVW0eagfBl4ydTZ3TIGzUGZgzOSnyjQS46Y9w0aBuTX
+TtgUkZP9IKb1Mm9GLmMmjrfqh+o0FWBToq/gLAU+/fRers4Ri0EHGeRaX4RNwpS
o3zwuOxnZEoad8Z/AwQw9oLXpk7nEi29AFj2m+GuKVSQO7FvECurBP3oQuW34GV6
zGMLv8Tu6xm1Ahobs1NGwSrsz4cMXULA/4m/HuKmLLzC4GoqcbcxcRxMLeppj/iZ
CmtR2FQEtgjjKINDbi5V+UQI7uaLbMmZPUfIRSou4hiWCjVefTF/aLI4lRx9i+jj
ZEqYU1+XPN182SK+OAhWl0mHWdzu/tcno8IdvMTAqrKRYL3Z+8oWOs2ZlVXMIcyt
xayWriZXV+BRObiVWTfAPrvdQum1m7c3eaeEyFQSXwopzg7ZeNW7WsaacTYUD/CM
PTuIwxgi1xXh8psaTHzKEwEaz9druq04XTLXUxnd1rFZbh+LLEmGLSAow6+M0VFf
OXM6OpVFnMi2kRBBXpbJ12DieCiOA3fQNsc0By4EJ1QX9nj4b+vBLyK/vssmzjKD
cmQ4abO+8YSy5aCVlI2bDzHrw3+rZ91/7qWey1oMy9jc1wFiEFrID48Wearm+B9m
xVsJlYQYMbLwVHQS+qwmSHFNc1hO253qyH1MTSPn1uWygXguqwNcg3Thyg6DHMgt
aEepNjo/EBwncQFzK58EewzFfachvWRuhXOFlI5n5ofbUQ2R2BQO/Gy3oFoAKlx2
/eZ4MRYR6rPFnB0r9hcTGIdvVJjSjWdhDTYbVlJoth93VCLFGrOoLxiTyAjTWkqk
jBNP96WbC2ZlddKPw/fwPcwD17ZB/7NZiqlppd4bKf99GZCDa/QsS3obvrjy3qzG
jSpor7lX23usr/d3kWhoo8qq47PNZgXe5rGKtdZgBAXFUwx/UCJsejoWVEvubxZP
okXer0+ZRY4tdqX23yNT2rrVU7682s3UA7R1X9nmbcxMde7um8u4KgeRsyaf53Di
bILuBcgGQMIBdDyfCfpJBqIgNSwkvPtjvIkHLRkW1PrmYAxmEyQZ++Y08ih9S+kn
b6nJIdGAbNgv4LHXlMDkcmgfPFjVRAGi22PeFzpawXWdhVdXCiAsm8dkxgsCKZK0
EIGZXWSJgaWA8N90UhsSiCGhy5xN55WPsM8qUFuBPm/+zOcQaAS2b0Sd2GpvWL5n
4ncIdfdI2swHtgYHwEFmQqpcB566s0dViE5QImZBv9IZBCrGa4krOLcOotzJN8XB
YERwyNKhlpI0fSpBdyJk+VW8u99tGVQjuLzjNsBKGQku2WO5Z0N2fCZbhXagB82p
H0bwxgeGO+4UdpIcTowExt59c+TCk4cvrMbYv/V37OdvYsbcnryP9KIS0E03HrsC
XoKxwa9dh80UhYZY8ypkfTrF7rMwtfL1FFmZT5GAJKy/J8nxdPpidDff8Fxr+ID9
nOpJ+t4dURoWZEy+5ER7U/tTokSrBBz0n/pOY5b5+j9/c/CvDCo4EP7C2RIJFKMk
+Yi0tUpquyunL6NP1v2hXt/8uw7wE65jA2uxjQuCCcFhUS3HbB5dr8qTfZ1/JlFo
a3vlU41JRqvIaK5SnzARbHS/38J/TcbqVKfHx/GXPKu7R78nJLw1G+pdfzsumrJg
eBA0uqvUv7WYMhvxcfp2X2cSoLvJyzE1JLMR6GEofi76MNpF6C80Rbh3rAGUxes1
d/0yxu7b8Jdw6tsuGiabh42kRev0t1nlN6RkxM2G3+Ak6feZX9pUrAZXsjkbpNhq
Js3xcIWpxu+0ovjRbGwN3ynMETxih1uDvwDqXoDhJ0wxDEKLzGwEcCf1M+8IUN3g
VxsxEEUfEcqEpeRusyj7JZheMXVcpH9++LQlhCKWPyKNACY5eWayACNe1llJo10f
H0rOzu01byS2TNXMczxm2s6dhTviYrD6TkTbWSkkkgRh85z6QVx/z9y9CMJ5CmaT
jMzy2JeXxvf0oQKa/pKjFN9J3f0FEeFV1LG3PBR8gdGCetbcl47pczT1GzWpvxOK
ZAYMyzeICgsh4PenftoeoOEFMo9NA+goBJOeBqnI0OivR0syfq1KsWZEgdsD9jL3
eEAn2p0f/2imlDloju05fQ8pGYLQ6NUAmFVVAIctTraj3/Le6kcGA9Et+8Rp1arX
+G7GnE2/RvIuXe5KsA5odQsc4Ndvydq8nBPswgidnaCr4ANHxYAqn/0Ss0StWIHc
C5xPuX2dncPD3R1wPDmQDLJdQGoMiKDCFPlB5qOy1sq97RYFbgsod6AYK3LCde7o
Qr7gJiWjlIPG4g0T+mvmnyfM7jRFK8YXcjfyZx1faUgjUoIrGC77yJ9yjoGWaf+w
2Zf8EM1qMdzyut0y3jw309+RQwDqN54Sn2cfgPRDWnkl0FviphWpsiXNYwwgEbYj
RgqcMd1nzn6h5usO8pa7qYC8K46aeN1g4W2/AKKIjbp/rm3Nl51WR1xjx2TCAZZP
kAPDCAPOl0KxjKDpxWBiZO00Jvddaa63cPdcl1w8qVhNl9TbuRlAZ0iotlJKV+tK
jfrwo9F0wWTCH5B61uNv9jt5ZRxgVJsacX7ciASHaBdGrBeTy/l1idCbr45e/vA0
jq3lyVGnzQcJyUtqla7/dmHkGtQApVuSf+Rt8Wpr20VZAeSaSbJswJlKfgtzxf3E
t89UN3R+suF3HUpE2VMzGDao7/8S+Szm/HW+909uQh7vDhlKmJrWzlIgeo9g03Le
U1igg2DSKZhTdZwOjPS1jdvZ5m/WM0fMkk1ykMVinKntnDJsNt1dmJKS7gsqb6J5
QbtipaGOijdng7a6A+OAQK3gBSKgjJ9KBr+R1gppnxNyKyzw8ov9mx1SyCy1mbaJ
Y5oGA0y7LckOOsNb16MosJ37inqMbw79lbZ3ikUmOOgMdRagVx6lUTZKxHGbh50S
bVvnOWfZxSYXu1rLtZPIuRVCIw2NC84ovhb9RADjmfz14ytTEqIPFeiGVbjQ0N+T
bCenX3/kM46diohfzV1a67lKu20uHm4/uIR2xB35OSPL0m/Zoi1RBmHuMBfC6NLl
YQiUH6iyfFRqIsAdYURqzDgQqBdD9Df0kMZXo+YWUVyg6O4hddicS9wU5USgstTM
gfBYKBMtTzgm52YSJqo0jGhd6v1s4NxPp1VX1+XlTt0LgDTYUvJNNStALAHPmj66
v93OWB0kOit8M/Op9GBZMV1JAZKXN/Gi0sjnhFWO/YRElmNA4am/3N5udUXXGt8v
rAdGPOmI81RcnDydMwezAvow/jz13uRGG6WyBeXHPezn2+8D/FZC9fTTVFdDLxmQ
v8VBAMzPEfc4wTBZiubMCRG3FBFnqeeY/Cm1p97l+144oW+E7TYtCxbs6VM782Vq
QDIIPHf/SRixh+hKqu1MWYnf5oVHKzkjoRM1ke1n4uh1/8siUH4HJ/DzvHxCJVSs
n1FvkLmi0hTYqJ19ZANAGNjcrKdiK2ivEXiH9Id1kCTj5xTks/kKrHqPGtPqKXnF
zqQcTTd8Fanya5I7dNW4YaJZsmZxsM6WZFT/otWgJ0EmFxMMI1KQIJ08vHPS6vCs
GuJhjLVfWZeHJnD8S1HFtRETKoO1Bvyp1YsgGjJWEXss14sM8kkMGkgnOg0Miadf
TJkSUYZJBKnZrVC9zRvs2eaKpuCU/Fgfyiokh4K6DOirFVEKhnoN34js3AQoqfUd
Vn5MxxxrqXmG2vpqpnj1BMwrqM8GV0WIlwH7PwIiz+8WzxpqyxtOjZPfRxPQlTWp
RExCUkg1Vv+k+v4DBjhvvG1PcJnX+MEXQlpBxEGInQpu1nvpJvQds0aurIb1hDo+
D7qKh9S/qTVO+Bbvy9GSzG9kjGpuf583ajEnWOiNGJNbnYqNrKp1R1J4PLtSZgke
i409LjoO38s1dkQ+6qw8720kGev6Z9SqOG756pD6I411C2R+3fhvSA0DR6Y1jEl1
7Kt2HnBhptYcaBlWmfIRDmq4iFrLOD2ev5WRrhHyfYSXBteSn+C5zqERrYZ3zvfl
fo7OaOI6dCeiW4B8eoHlapCxZvG7CEwyV9C2gyG9g1zrs6JSz/qrpP/XrgMRSh5E
lsrmXdb3pM+28v1d4uXmXoR7jycIfjQDkO/cwxtsRHdRu8w39OD4rWnIywB+csW5
mT0Q53NKCSwEkzswPFG8IrwtBPMUAwqgpb7Tgq2CwfJY2k0UaKIJAinSX4tsujyx
POVism81EOT/EIW+xV6csF2LE+PoGFAfTVcccREolqyWFUihev0XtiNjSGfgxE4n
l63JDBNRcWogcNJMhqSFOSsXnjio2LVo21EL5kqtxo2rneXCnloNy0F8GH+QL9fH
f2VVMXBFeKCs9axeoKHhEAepX9/F2h2Ylw5jEPml7V24kIjswoqrs/rh3u7E9LPA
xxjAJjWZunSZfDdYA56gcFMcak0B2tLmOvswxmgBJnUOMJCDSkPhEL6GBH10ufzF
c/C4v0DRyAKjq9p1FDITmX/+j9kJa8kvPxLvuhP7fQ7pKauJ+OQ6u7XcPElALG1i
co8vXAeFcvYas3kh8k5XopEinTLIx35FpJwX7Vb4qfUPLwkXLliEdDRytAe95Gma
H3RRdq4uMyMFo2J8lM1QGZ2g74iMQrIn3H18fNvHZsaZSmsgW+36/1DyqwzKvM+v
ctfpscs0mYCENsG+901B7h7pl9D6eK5B8/A6ia7eLLVQ3XB7ONaiGffJDNgmfFUp
gusdjIbv8w9mCZG8OjuikYBqxsRpyvBp1KvU6POb8QrgCLzw3tmg6Gp26k2LKP0J
eL3jZEoYH3T3SKcMrCxIb27Qs2WvFygMFYqM+nL13rx/E7V+TmdT09KFoInPeTMj
JQt/nJ/2zhaumGWjXp4AscjoOyyWMVSGvXE1I/ws2gsGNfy+lSmET7Zom1JcrEPN
0WRXZHmiTgRKLMGL9xajZ3kjsD6u3GON5Ms+MlzOYRN2+yljJGRyflIo9OnjiwBK
OPNiY7x74XT5dEog1adLpbgte4uj1CbcT65KFGZTlbz+eCJNNcr+BGH1XweII6OP
yxGcm4qmuEb6CNLhg1ltUoZ3O8w1kxz2fhrsb5Jc3KZmesNE6Y/HlxQmq/UQ3s1N
XoDbOnW2FAbfSTjRB9kDrQVh/mM2kigm96zbX2Ha44xcVWX1mIQEFT25KDSiedwc
9qu+znqI0B+J8lwq/Kwqrl8iR4KqHLk2ZFRwZ0K2HsCGli3r8RGEcNAkbDt3rXYO
HIPA7nEfsPtA2Dm5ZoUSCaqXpvzQ95Ld3wwjq4ZI3SK9Mw85BjB+e2L7UGKs4WHg
YielB0QIU6eH9k72IwdXDsshx4aRtA4mIp8ICVFmKN3VnuWsGwRHEiKBCnKG/7be
ep23JYUo5xrSWEivzaebv4lvui74qs1y1QL+4UJ/caO8J9289IR1NEklrPFXkngv
GiDnJIvMGXBx+pnbdrvF0QmsrF9Ns27FPkxTepQxnJv/WSA21HCDYe6q4b2Aqvjj
wWDaocDv7nGu1WFMIVP1eg+F5Fiy1KDuYBb6RVsOpdbIiIHXQGQFL9Ppg6jw1P3R
A4ViMPg8PQ6nwzKAnbaQztpDNYWWOxAqdth/MPh3HrXGkS0d4BXvyLvs2uEQZRdv
yLnf23kHIc3Cneh5XLR30LrLbkaQHcpDLuOrja+h438IYwSKRJtcPIIhMWKXke5U
PfeX7HtQetlMgCGAv6hHxQ4O+9jrJEkz2bKsGzbIzMDyxL+Joql4E1TG2zyDtjDH
R+dCe4119LvyyIPVOhsZyUhtXpMePePvslNpb3xRe2Uqp7v6ErqvQRkb6IiW2O0F
bRiw5DjkOMoi6MixRSsXTUaPFOa8gY8jqVdGtiq3umVf5XSo+IHbcuE2eDMR/Fab
Byw9/6nudsiQQ9yypSD6w9m68HHnwmmKlTB4NBkmlJ/YnUuDLkIZJkyu4E3fu5dU
sSm3pJdpXSxPco9HWY43UIfdSn6smVboZrEoQmh7B1ZuqXK3tclvwJaCScMIEY5V
CpBo8Iahq6v88y9yZqQRawy3jEIb/HkL7bC3ERAsBnJYRJyx6vIfq57LInpWvD1p
K53I+oPy/1YRMPuQGTqVVc0d2JaFOH3/V1LGvbPWilWH8DM9H1o3Hs2mFF1gcH5z
AqDN3Y3/V/gNhENKENcxwanuy2qlaMpozhQIqTsPcfonlwEvH0s4bN0lpPVqSI5Z
K/VeqapLu2udzM1oRqMg+HI01tc9gaYUb9DjQ+YoerKjH+GJkrrQ369qKiCOgLRj
h/1tl61sePBa381s1FUezJKKjIZD+6hCoN8r35r2LHA+bcx3IqLnTG7XvYOayQ9v
tX/s0pOYEE/q68vy93B2WYX1kaTgHGFazM7xfbvO7hnXmEki/yK2SBq4OLcAeNwY
Lh21jg/tKa5CS4KlPnTa6WFlzmkslPZ5O0J81a0rPMg1m05rpKPN1OTm5I42KJkT
zf7JFyxLo5VNE+OBPfCCD+MMrqJ/tuIPHm1moFxkiMVR2qCiG11aRL68jZQfZec8
rHTHFOh6WUBgdG+F4myb5ea0nKBJGIQ5Doutw3kSgFYlRSBdQpZ6kMkFgDirEJV3
n9f87+2yiCKP4zG7Ey5Yx/YcTi2LcQ6oblA1W8XKFPlyMmzCRWJBl6LlEwsPYoHu
8vhitXzKSpevfA/CdIHfJAojMSgBFN0ZzjQLC76/BvXG56xZgWtsgJjPEvTA335U
IalaCtj5ntV3NlL8/SI45NvVr9O25ZKZ//N5eCUE9Y9XRWSzaIme6fOOcmaLAIIF
WMO3q5PSIZng3TL/1GhIQFT27mZxGAvw/uqz+ViFYyEtT1IcAtksmDTtX5q10TYW
SQOT1qvPdrvDUjpJX8lLf7Jc2rlCooCUxm9wSQIBroUUxoXmBEfCDnTVk2Kn/oHK
FfLHcaWilEKVAXxBTqU/jp3rqo5MX7SabLL6eUtBh0ffguVS6PvNS9703sQevxVr
I0aQNR9w0lglJV2f19KaGMDtMpRMeMomf9EBf5vqY5AkyEtPPehRKqHb2WcVVbvn
wpxoWpmzVDrRwF1V3Cki7RO9XOaknT7cbFRgtUrVYY6f2UvAhSZvN9Pvf5LUuL8F
ydC2CwDifYvKfJF+ziviiAFvjlOsxq2iXREh1gb0zqDSqWewEztjLw2CpfGCcfYh
YHxeYduQF54sJpeEehog2lJGeiMq72IEK62VraOULZPrdXLfs900nYFvUplcs4WL
xaTULAGx1D0ERRoIn72ic7hVBJK25YQChknYmvVe28TuslZdYUkXRtummMg3ZSLm
8Ws30Wd0c9bK4xplRV5z8FP0WyaIKaUh9FZbtCjCtiNblQcN+JZfM6JlVpgNJKwg
sXMzgqfSPGi4pGgjYuCmJhbvBXTpTuEEE29G/LW4RbE4j+yimGNxqthcfnOTPT2h
RxCm6z65EfH5YP9uO7grv3HSA6x/gABbFgXFTUU+vHZ7S7Ou43mDOOnH2vXP8ulO
/EWMKHtCUvzPmfh5kvyiOOFUlTHDHLIudYnL5uHTkw8t92/qdn+jpodiVSV+/cfl
T2zdr8rrvN6kClchzOKotydfOcveiwUC7yO0aotI93BYkbwfsIgxlUxcmd+HJfSH
LdLXQbuqcJXYSdMLytYyAA4gNJYozrU6PegNw/W1BDBO4zXszGohO8qxNaBuSHtk
ynV10DjbaxZcI83PCYwAOxqqjQKL/mZF6EDqlvAbSPDzteNPLhc8P0LyUT50BB6o
VOkPnTBUR22BCDVRshwWCRUFpAMUPLEn81Y3v7qZBEHwituiqA2lUGc+FDtdosg/
snzqcXjE1+zZouAyCuD24kBm0xC0w9cIUOIf1z3C9La7LxYprw3pmwTLLb2pLi6d
oujn0o7vQL/ep1zKq0W7ypwIV/wk412ksQl0QO4Q0ssZ3kTPtv1YHJOuHp3u18hU
qSYoLcQWOFbn1G215UZyYXYbn5XB7ndWTNIdHd9A3j/hel22KGQv7L9B1cp2/HN7
bslRSbCv5915jIrDRo07Olv+jOzQO1jjuX37FUI4KbXSx+E0r1MzXSLqskKEAfyC
BYLRztGzmICV6FNpYl+zEb40KnBfnFYHI7uvGjdPWERYWMUliI5REpUce4307gcm
nGRhyRXcNEtWlI5sKohFnTx9YXicXbTTTlSELJy+DnG19CunOUbHdejgeeYRAQND
8NnUuBcnAlCLJ0/Xb2oHKIvccYpGTfh0eSDAQqgIxjBYQv82fhQ9LkjYgauFWLLp
kdFTIdZhNTkBRPbxNVsWC+uJGFSmkXo+/dP8Lp0+MJFuQ1gQa8762O2h2HmcF/8u
u/INuSnaYgG8gMSgy7PaMJ6sj0GFAZobvFmBFMkd4yu/68LLpG5XdEW8DYVN2k3w
m8BPjHIZ7AaSZxxuaXHFD29zTfia38MHct93/ELxEa7N0tNxI+bwU9To5IYPdywX
W+ZzmZ9C/nuRjIIo3Ohy0myd5X5Y7g5KNuAM9kmHC8KB7pTjU1RLLAkn4nAm2XVs
tFVCNdXaSnJA32toJG5o98rAC8gGdexM7YuVSPZoOS1VEncjwdlKW7zcaNDY82Mp
LeKqM9p0pYgWHu0U9VgSQP3yKHMw3csFh4LEWz6w0uf4mziFFNW08Nq4KL9X4vIo
z4eX819dlSkIj+cnrpfbmAA7LV+RlP25uv47hiq10TkdF6Pm5OlFBWHf42ktByJp
YhC/hFJI12dQQBY4KlD/xHlOYV+GS2wkV9AnD2N7tAEJR9QXzO0KuHqlegsr+iFj
IIO/7aFbwm8Q/bJL3k9iqHl+NJQ3VOAJZQBA3PV4ekPls2tWpSXPxNVl7wDdL5C7
Kp6ZTFiLSKzLKxhjO74A3n6P8rkH/kGvad19SVRL1DjesAZcsudY/g1DdMIXsrG1
pkcxB3Pxvlm5bNie3tWcYmLvmPET/+jTZ3XnM1eW1bpf4VrqD5+HR6u7psBmf2tk
eFeVquP+NDy30g4lRGTn3mPdK9R9MvOijOhgwQ+FN+iPCUxFGzJUMsxYadR5Weyf
vNJ94vkra09UaMyzSdbdMlk+vwqnd3yaUevMR3peU5BX0memVVt1/tj3zFBYltAn
10urQQhjOcuuJK8W0hdLK7TU1lfwG3/sbCfvphDDkObSn2GE29ymYopb0Qdxv0ha
lBmI89N5owrxl9DJxvrmv9JbQyHpli84hH6+cgsrqrmVTQhKMuhTg5P7QEsSXO1L
khbjx4yU143ixPb5M9rd1i4vIcXJ9fP8a+hiZAU1Y/spxw0z5sxsNnLIsZg2U1ZD
sUfC2mRi5lsA88SRRplWXmolz0fzXn1DHPxZq8VLgsvonMI1RJGzH8wFyg/EuMG4
zJanHMI2pcKaTxmVu6CXU4j2gorxDz1NuXcI8wvqeBBPEtyqulecItWDEFWd6DRI
dD0482Vmtag+OnKGbgLflrAhESirW0rLUDqJx01dtkEAWs/4jQU3YAXuhRMY/W4F
YGfYzDiAvdCkb9Hjabdg2VkEb5Cj0JMaUGiONGKsAHtISWICpAuwZlbEK+HT5kru
d5y/loiZBwutbQFFCb0wY1lfTs5c3pHzB709M29dJC2QQNizspeu9OEuIiHxYBNk
rsoHxgrCeKDwGI5dnYddAmNsAsSoaMrtt9RV1/hYNDz4EdpoEDV2158r+Hp9IwSy
ZywHRyVQl855+hiYouRCIaFGyCIHSANa9iiCzNI6SQOgOHMEGSjRQFkINnN5ociU
HQWAjXRULySbSEGCYSBpdNtTtl3m8is9dMUkwPF8Uxd3FLfdH6G18bNQQlCTCOws
+HLMaz7ZiGtOfIRVhQ5GhexzkuBWLUPw6ZJ8eTUBU283v0jCmbDRn1qqpAnX06c+
Ji70eneWz9S075XxPVd028P0esyQrrjpuAyD9JQYlQkx80+fx3qlYuZd365m2X0O
oH3U6iLfReQMsWWysPhYwVWQx68agOn2kJ9hJ9rP/zBSgN66SZxTcaDuUxakxvAM
BBPC0o9QvmMsGpeJvPKF3TWKmRa3UK6LEDsb3a/Tm6C1IBebAPpxJG3mICPRxjrT
FmF/h36V2sgN3NVrQqDgtqCjl3OtlJFEssEjvUnMc7wPA+fekVLZ34AMpQiJbT+1
4e9FA+xzJ/TVNg2ZnvCT8k0wpwBM6jnVLzoD7O59loGID450GdtH+KEjAR0qNDFO
EC37N/Xj4uMm+q5ztNra+iRAqsFquE6em40Cr9PPRCYrCIYf4lKERbwK3wUu6vGI
AZJ4qXN//XdYHr6cJ0cT2c8vjSnj4qLMdlSoyv7TB/jvcBozbub9ZYnq+9JJUk+7
gFxmGCoL1fWTLroO995UlzMLkonsu/3M4Uu/clo0bKVaEMV5MCKY1clqXEn9wSzZ
ns/TTxxgXxv8bG9wHHuAbMd3zm6uAxjYJ7pvIqIao7mCD+tjf5glQ0Tt0cBDeJw1
NeqTb9YWjnSVtZuCTS8Xis38t1u4qtl30MS0YBOuaMKoHGN1LSPCq/myizpCun8V
h1FGtJR0IxZt6XHmEpCRf7sKOzdTPjJTeu09QQEQG708M9g/P+y/utw5eaRTd53C
8ibGOFwJvRAm5VFsB1PiqBvhHdsoZDyWby3A5f+vuIcGRVcGtMZay1MN/VMQwmL2
FQI/gsZJX2jQAOQKskkAZFytNhjExUFyOMxd2YjT1qupZXRJaB/9JOeUa1Q68vuH
tj4yCzao2+pDZPUvWL7tyAwmeaqYYrmZZMJDGX3k7cuB66m/ZAt71KugAbU3mkCB
n/VYqxom8gisOmkLvMxeLKFBJn1qF4Aelz2a8ByII71YnO3cmIy50wnChsS1U8PX
qKa3Htj8KQuvf3FPGD8ZxqI/ewoSIFo5bmEhL3fzfsFEv110xnV6mke32X9UiIB/
DVgqXbiDq6Bhy6dIyMierOfHV6crObL2Gz9ipSuGhPDoVvgb8zjNtBZ1pkEAYisF
WKVa9Do1ou2E2g/mXnUGH8h8RKAZRjmkdyb3FKOpXUBL7awiqbkDgJDiz3oUqkwp
8cfcxy3JdlviuXbEpMCJiJ1H5SSB0JrQVKrZSl2gfnj1o3tANkkmgT34H7g/AxuC
A9r3cv8Z/BMBelm8mT6V0BkViATepW5VNZLrJg85q0eeMakEDb5L8wZ+O4obLgV+
9ahfjTDUcBddlgwJg5njGheJcZ9C63MSlCGPunCC9dD2uSBVbIGuBjCJ3zRg3/h1
rlCCqZDOFLv+lTXRWEEXf+hO4NwsSVrbr8XOTFYcxJnrVsxxZfsZCjFRnOcaV+pm
IcN+0+R7FjhQnDoyedzQd7uViw6GJw7zQKlFkqAoUoTfeb+ofDo0fu2fPfIJQO6m
DIAHFxjV8RHL0N4AiBItZD1j2txpOcFWLDWwJKOP5hElHywh8NO4zDMItn5NjZv+
gH9KG/6ICGxjQBkPbMTsLW6mLph6P6NqN/1BJCNRZl8o+8b5AkFXb3p/z8ebLwRj
lV878XM+IhvQyQ1HVx6BIame6AbPDFUQMmbIUliJ9MqId7ZWAOKHv/6pBbi+7SvV
dLNF1NybdksC+Hw6e9f5OBdfhoUrC1NgrbpTEulri8VFjklJFoUxUGU3NCoQOJqb
XIlf058mEiaw5RlGzKCrbI2FyWfM0wGsBs0LLZ0b+1XYePop9znhq/hHB/qKvsJX
Bhe6HxrOXQXJNnfpmAdPrszD5Q7EIhmTQt9HGPLSEorC63QwwmB+VX9ShNvvxJiD
SIjfwF6a0Pfn1Ekx3koFq/2MrtUZAy9q5DXKs2OpvT6KZL9l+pVqY9lAwlm4juPZ
GEcALNE2DsymhoV8Ms2tSXKxpPQO19YIPZQJmz4DdnJbDnEHiyEFDYZOjiRkvZLS
ggjthni2X2mxfKnd+SLGWE4lvKuvfU3/Yd8MGpT3XTqHfgFY69pF73TIN0ReQwnN
NZRGAPDeBboLn4rMHB0zp3gl8TQ+78853Zy1zDUSetVk2OtS3oS7G6I7FMKHB5Y9
fpliimugA10jYXtgzMq2TusUJJ8uhlaho2oYrUJNYRd+sWeoYX7CS4oQkapueXb3
lzeNLE5ZvcGUlnjtvBkcV2olyrbiQh04krvyaoOsihUK0GIln+S0kAJzpVAiqJy1
rpsrdu3fv8yBpVoE+tbqC45zhyWPrKtAk/ndVC0ThzBQueMABe+ml0CF35KJ12E3
x4xbZIWCjW7DMllaQwCdAN3hb77PaAAuYQfx07JKbSQkeuVMo9YXsQQpPijGVVjt
uZSQ1vjcB4nSEI4/v6ykx7tTsJJxHOuDtxuas5aoB90+vivaRZk7CGQdHroEAROu
EAHxvHKWWhWQpLFEJzBX5BpBc37fmA5pmZIOYdzTfM7g7rRXCC8762YJuooOayFr
yWM2MnVtd699wYP5YmrSBM+nvGGBveCr7BN7eQPOse64FFkNmqT15Qwp5QLU4zEL
bu9kkRUT58UIq+a3aMgj+VUhioyLHtaJ5q7mLHedswr2zSTKSGS0r0pvpVKwAcgn
CSaMCav1fRl0pD/kQvhHqzHd5ooAmb6MrVZIXHz9R5TmEK4klIiD+k6k8OJlpq1M
HCiknnRLu4sqLfOHezPG6JjB5HIspVO5meL1B1ayV1rD7nBBxiBZHCoClBW/6LGb
lcdiUTg7SAM8dj5ZGPA5qsY6bMDpMKe/j5kmKzZYb4DRbyI4eTTmiR51RDJ/xi7i
7nLqq+pD2mL3kftKRi4P9wHPVkJWiYXVSB8cpJhp+Br+Nuh5S6FjLb9TBPVbFhPZ
0uMvke2v51So+6/DJ3nXl7/lmCfZxlb+hoMxeLyejwu38NxXT3pPrZrEvJK1M+2/
JxaoSG3QeDh1aYdadKhfK8DNJr3m9mJ0IJfuzO/hO/vPaVOpLog7MdRD4yY033dR
+hBf6lXA3oOa+EwDJumxblMZwCfSj1EFv6OCN9EMeGF3zRebsQRLW/GI8xX3poG5
qv8z/brrvCjX48aXbif5wW7T8hU89Nsd9iiEPqIP8KBAsFhlNLyTJu3UVpddbcf7
AsM+xrjjmqb3ffaEufTJQYNr5/ylziv3uatpLWnQsnswqAK8MIw65DL9u8JRaWXw
3JURe06zaY/A1hZVJOVatrUFWBU8LDcwMfnfzqS4A3HAXekd7RWopSK7Mdj8/JOT
ifyE1giZbldlGJKRw2JXr3Po/lw5PEc38u19lcGjxlAKhtJFF+koD5g8lgHCXDs1
VYWmVaOJRLtztOsb8KJzHFr9jFD0iYLMNDOdC2jVf9lr3baxKrjbhTxmlfCOPIuD
t9D1UEQ6wp+8g33IrTHUxMrz3wbbCeDN6gBTPhCvSu2NJKxZMrgbzFomGRqm9r3W
08HzsqXTALc55FldrBJ+PYMlPCzrzUE5uUwlCKmsjgZsuQ+W3MhNeD1fzffzb0++
9UVVpgHviagbu6P1E8ynx2F85kgMXdlXBRdKLjZG66vDejcQJjoriTV70iOol7tt
44IPrs4FzoceqzABj2RL3pQJ0yb9P12bX0/TwkZRV15P36z909NMBg8uFeqCplmL
pmp3EExrzrGkPayeCnJucDqqBPy15sVMOj51PHsMGgydECDNZWra5MnPWnBq46mO
NgvlMnY++X0DnWstN3kGcXzZTbraj/matm0eO6umwUew81Ho+gaG33qxzHgacpbV
d+It9kUuSKwWaVtsDweueNTOKQOgJPR2KmMeUqUChAp9IdbVLCqg0Dg8k1wuH0o1
MYNDjVrX/Vz2KIOiPPIeYNXMsBnYVts7MGK1W7k/DB+400Ao7yrmEmYhPZCMYp/R
v9JGh4OfTTxYDU2PqM5wzrumew/WyxAd4A5uDAuJpFlnOKqlozvgfcNYosFP87Cg
54ejRLtWO+bC1VdoA/Pc7yFSAfWqWgkSNSyzFBjwiM6VDwPmXeSpo7wR62InreZa
SwTA9gb5nSAZkEmW966HP8TGSqwx+5OvKMNuCsmxWwf2fVHNyaKsFiMh8Revw8jm
qOtguH9fNJtfhY4jJWFJwiFIW/y0SGpKVRsLsWPTgcfw/1OoGimMsGE4Yc2q1+ii
VIBWFB08nj6Gr2HsoP+xXGLs1QhfoAyw9g2pJp6+pto7xfs14fww5xv6CHlI8BDU
0o7IOoQux3FYYs/1iDUjWRQ2VLxKePCnc3Lx8r6ClBAWSb9gDrgxzj6YyhACqsTe
WlhCpHXzm3fBFLpLa13E6a/i9TN8DAvTtPDdr8s55HcABMLF5qL9yTcxZiZCEK7a
GNgoszzQHxrB/6YoyVSZXsaB9fDzfqgjAei+2q2Q9xFTXVvMXLfCFhHUGvjKE7+F
MMUp4JMrlSnR6JwikeeGmnPeQEACZ0c6/+P4P0xIA1w8JG/Qqv/R566jxjtMfIT0
O4C0WZC64c29VwouRhc9TBNfzwfKbVS196N9qys1khDhEmgKCGvT+bTPatvMBlo9
iHn1vjpmCHCLsJUTMcROTxAiez6unyZ5QBO7MSeuhlOuPu0BNPopv627WFpCwTEu
a35ioMGiuIwPmCrzNozaH6+R9ewDLPElHmZUwVFrj2yLk2CZRmBv3O3fYqY1D4Iy
QYEfdeafcQr4EYOrCt1kwEbnRti/SmVNXsthEk0X9TvnMLzBsFIL9gYNjnPQkBXL
fWPf4Ql1Pv1P5NSk7QHSXZTtbS2UOKtFm8bRaQOCCbctdcFu0zc8MqP4gjMQ2DD7
Y0f8sfBh+gJr1+2i229mAz8/d2scEweOpJwPOTCl3mwWzJMl+PcBVotwr9gZSREc
LE3sXd1AigwV3CHc3aGu+qbLqCKNxP5CL/R4Z4553wKm4qIIgR9bCt8fbjbIUMzK
22FbAhFsrOpzHCiRFO7SUjN+XQdH9gX6Eff1wstmbtTQU2TCK6kBkLUGGgXzkcc1
+43RKh+wmdmD3cfxWZuNIQQcNbmFBh/LhGg9BsrhNQ7idsjNK66kstNV/KtiIj4W
DTXchR6fpPT31pu01w3+VklIFXdwemWBwJF44sJ0slBD+Q74hCo+7nqDsbU4zfR1
jl58lkm32lWLRWx6T60+iRBHhUZKLEA+DZ/n3QrEr4QAobRAmu8430M6UnnlRzf8
86ouYGClGZPCt1YdCoYeRCjhig2mEmyTRMYEInVkczzY4nHEJEq933rxh1xdKRjf
OMa1FndQ/ZbTAp3gUkkkFxS8o4pEJR2EKg2T8ZDWhF5269h6sO5DeRHVXLUPWWnF
H6EsKtZuAUrrJ0903CsbXp/s+DDwl4O7sm143rnmcyY1A82vJk2LX07YUDDo8z0e
+NWFzcl5SLXGTbnlKAq51sSja6VLN1j7oBq2ke6AwKFCEKeQEIe7vly6w4ywF3pp
n6GeRa/NM3NOaNRuAF+kbKqgD8kFbX3PntGsFj5nbcVCTmFAPVomK4jO8C/6sTab
aqFclztvOr+XgqTu5wcRvde8CJajSZdSN3BctMkpyqDv5x+UfMsoJLRUt6KMz2oh
gff84Rcjn2IxvnazG5JOGEc+tInye8jggfT3ks1vEycc4Q8JVl3D2B1BTzjpgZcg
3LE5m++VQ0LsKqrlQiINcRJVfa7mne8nvt/hjcJdEydGUYEA5KTsANTL0HeRfb7u
TFxCPunSeyNQUSQCayZXN3ZIV8EM8iwLiHgwjZ9KfOP+oDowKZkv893QGzALrfBe
30XnpOc+cJwmyRZhMjk80jXUNT0hflXectBYDrtXN9gmuTnObAPhABvAnY8cImtf
Q03zEsixIRYtNP71RUjvUVCrVQJ/U8AkgZfjYTOO//eKGjBb4v0Z8RgLLe6uPquW
D8yLGqA0fABb6Vlqc70hyvWJXymV3xi2ZdktNop4iWclr63OOxSCrfLIV2dhA9x8
b/FKL9aU7A7qyc7ElB8bwYj8eejPGZEep8eRloXu1FpZG+e54+3GckgvqM1ldL7x
sYHEL2Ko/3g6jnTnQ70AfsWMyeb1Pywgy88+alSBfmFbI1oWRV3bwYRCObMKRpMH
k0RRoBvTQY0L3oRC6IuxscuOM08gSXcF1YIXpLZfejA+WumqBID9N4hw9OXUZFp7
bKMKR+IbiRYBQAo5RdCy8lnDS2KiI5KflMYt8/KzEayPni/kKGp36YR048CRHi6U
BuMkFVvInIHTSLNkUf9rVK1ZtnBYy9HGroNhiX6UkYTy8lVXO53RIArqxzIK7WVC
48Z+qmtTKgMXHwvoqs1ucSnnb6TUjYFkdZPkMvU7vYiF1I5Wxj/uVGFXmpZmOUmd
cbFhK4PY6v0PinO+XjmBKSULhES5VGfqoORGReh/zc+jDohwMr7tDEsykM1noDoi
gEVswAcnbeRCSawNMMJFvFi5X//VX+gVlIntfSDnQvIkmKwXgWnlQGmLBc4CpeFk
UI0ul+NoPo5lQbHh5GCvRUE2Y9qOWehRKR0eH1jj0xgDJ7bFzuxnAI4nzV2GPn+k
z4rlxUr4ZxyPa7zgiUkTtJik4AipwNN+cP2o7pZR9LNGXtUKdJXskwK6p7M16/oG
dCzcLQ46N8fS3VbILjinvD1k+hnWsDXUnrFk1i1B2NACvqKA/dDjuaQ8P0Y4YpQv
wbZJzAB38MdLKx3a3ynXyt4e9BtPTSWYN7M8Y9ifOPhKqEbByX3CnF+qHnNlFS4/
RqHZLsj9iPTLwOMrV7CfYbly2px5WnxSUwbMyOfZg9MKB07A5GV0lEKeDmMV+DpV
Mtd49iiaIc+LKCj4gavnxknPuF07UcGGWNtIIqdgc99KdZr6YA5Qt3npzLbfDNgF
Eqjj0bNmDGUQ85VDPC4oz/g49jTqBeHqVybSr8xq+RLFBPkdzj0JK+D2uek/8mQ0
gA33aBYHn7+KwH+mMOD+Jfgn64qzIfXZWWqA0q5r9+MskeN8xYbhtHUmyUmnWj2G
F77R/Sx+vEMJe84BqtnmifDQaV1JhKunI7HkrAeJf+Gsxb8Aalx8rX7eLcL+GmuJ
xi1dh8txmRgciT28e35T3ETW6LkJ4jXVSWqOOycrySlYb3/vcAFnc1eSttmCmlMu
1vi0VpDyhjju0lCCV1ZZUcMJazqW7gzy7QvA814IyHTSCYzq1gy7av3FQEd86Jlj
fDM0HFm9LwPX5G5Bcdt2uJDgPJjvhpwLEhU7R3t51AagHxNJyO4kQ6Rr7H0P6Oe2
QOmp1hKxKNUJdYguv19rUzBD1+ZZfX/XLEe4nJwtRz4EufEnr2vpgGl2amWQdyD0
nvN+sxwsWFjq39EGx2/XSh0o/QzWLassGmtDoOpDdskk0qn8NzGpdYUE4j6Vs3IK
qU4i4H+a0Om8alClM0GsvoEnn1E5nC8JQYkivxuMx4hfxXRoQER77Fwk6OoR8cuj
+qRdisaG8fV4OZHPfZKIXK2ALsYGYfk9his2ErQVHS62hiAeAxJg1x3FOQZfL2z+
xLQCdsGD0AlLl33KrGWuHn+ZNWc5dpxInDJdA0DWprddjkrKiU7RtPUCHBUUFVka
+gFqNmRi1JAbegHlIbzkxL1vEGRZjoifYg+HY8ktft//yys4HBuTtuSwtyQQXble
XN5Ex/F9wNRI5EituMpcSLvmzq8I8CT6YRpcJZICxMCg+iexRnK36w/OhRTqA7dc
rqnpDIAYb+6OkzFwco68kLPcxCyla7E67DMS/t0GwScScrHibjnVVMM+LZUVdlVd
8qFRRXxi8R3jX2y0APeDwsgGeKdudp7zWId+f1h3BAdJszrL7KGsiJPDXHacIsKC
0K7i/dRnWBF2+oQQFpjUtyQBj7PYbsMYLdZxJdMZnsBmynyY94j3pnSIq1GOnY/0
7tvWWMfuZP4ZC2F8RMhhdwM7q1pc0d7wmt9qMJ/l6CLJutq+3v2OVfCN90BqDzx+
Z4xajIkMGceBli4R1kmCb+xXF9jRL/DHZmiDBsOmR237zI2S6j/OWH6f7AYdZrue
p/rfYBIkbkA/X65hMinnPOly3ebYetLRd/sFaAzGnVGsuFMttN1ydUzf+5kTvfHR
HMhG0XRIsalKDexImFN8cohInnxwHKCjnVpudhK8ncqk8uFg3R5MqeQ3VemdhsJn
ITeSAXGVyqBhpwvNLfZRiQOSmfJxrjJ7mGU6KiV+HWUDOaiPOOHJQVEsFgzfHujp
NNyI+Ru+7qwYl9xEL18IqHFMhxu4aZ/BRY6Rw6H/Gp/v08oza2bSysz3n7MaKPja
8a0b9GfdfVPJUDvvJXUPIG/r+qQnNzVF+fVR9Uaos30zeLANKlNhijRETxV5x+2w
ALqgQbqNOMYn4fUdVgiTSx4d0Qj/lBCma2Ant7NhVaB2R4zeo8/U/9+9WhfNgNaq
Wr+q6T17kyekF3kKQic+kg7drzWwULoQPDGfkwb4NYqkKeUAwdDe/f8s+yWDWq2p
iPD//ayxhZVT8pG6YHBrIbqJ6oXFSlIdYIjqIrlY9ZtBNdJ/jLh3OqtSYC8FTXIQ
ZcEsYyaLcQUdMaPLIyWhS4P+JhOy+t9l/iljbZZjOsRVByddsAmtYgvk3e7LMepp
EPAxOm90m8A9AtQHomzdEZ6GFa0751VwXytqRSrQOn0iQzuk5kppHTEgbo8Gwkmo
70YMwetxtF8q15Ib/voZqQYhxIyZny0r1L9iK3cYh6HJEVJjyOxhHAJJ719EzAsH
T0cG2DGW+hshYiJZObDjEpoHNXwk8xNWCUiU5CQGb4FtlhWzhV/TM0etZcI6OJpc
ma8HQVXVtHGac8NqD0u7LhI+o4cyHY/sGczbCBSiDQNbWJTktu7CWcJezxnqW775
U1kcQvSWue/UIHEFbuGmqm/wb8efw9BSoFXAN8i+NydYLEVkYL9galY5DdpSCXXm
u7zTj1t1KJNpzCIByGLpliMxP/0g7uPWNu7KX4Zo2QSFXjKplNtgy1CeO5iMbGOk
CJEmBeVlAHDIaruehzxtjqOrtbW8aFOcnfGNCqorZ5pjgt9278XXwt56xWZ+P2cK
NWxFQgIePwGOg+o9qYDeOYa2uSrSrT45PkutJse0fwMKmgvMbaYW2bFreWiDUcdQ
1v3cJsmVDGy/n1uG+KkSK6svky6DC0xRarYsFJJZsokh4Y+p1hWNnaHj3dUTSk4l
yC3PSHCD/93nI3yCKiG5lur/S6cG8eHPvrgfpJGxeyfoZlSIGJwULW3XMpSLEn3J
t+KPUda6V3UHQuN84YcMsRmwAkjJJbtKTq0nO5P/KavZXZRrQRXV2ujxO4aNybw4
3hq5NJH+/GHPABFFQc5cuvXiagp2aY2bttYECKPLMXfvm2yOde7Hcv5Jp6DULKG0
E2up73olPl9nj4j6OteSjro5KBYOJakiq4E0CNV9kkXVewSzi/U0ZM2EZQs5PXHv
RtDE+CbcuwTNrPqJOjXdMSAAnymXaqumaUoYt1YFJ5Y+ewZk2/X1I0d8Y2ZMa7jm
tTK5GNTibVRim3Yd/zkXo1PlbFGeoQgyMIHt//RYU5FrLodIYkUBiMSjmsYeemh+
LQcDp71nbfaSvqYrSMpIxb3Q+BS51kXPohkOrkhl/56XhI54soI1ym86Wfp7n+Ql
84XKJemx1s7jjBpHmO4Xryhy8f5X/FsUwIsn/gQ7iEGEGM7vuO+M+6x+Snkb1hsL
GHkw0gtSGPACbe8Rr1QG7pzdkbzIju/C/t6xTuxif2D1ou2oYA+MZeTPOD9uzvel
i8tUlcfLJJ1MLkwLosnEMpjd6fACDeik5wR8soALFU8bu+qahrDPmkyXq7SNcYMi
y3QrlqUrQCzLpvKzXzp3H9TibfFnTH1wafIJPubOWQ+OprBXZskrQSCn0Rj5Rkyq
zTdkxaQqtz8rS4/1oxIo0MC5ix7uR3tYigIZj1crnqX0HvREpFnWUCUlKOWu/Kwh
vPAMJZbzMGdSowtoAu9hlUSxItA0o1iINSnqpI1iiqmwXwh/ylzmK/hvuD/PwBDN
RFJQA0wY8fsO1vcWntjT9if5VTdz0LN1hfAuGyn4/65rEaFf9L81tevU2AlGzGbD
7Vs4GfOk8ssbWSK1VgzkSrHegu1KPDik5ehK+zRv32eFoUWEpVF1MafEQ/sBPupM
fSAycQcRxncMc1H+f8J99S6i1iLlJZE/l+0XdoPM5n8uqBZOGHp5tpBMamzKHZeE
oxNftIVe+eG9gqxNXCMDSSOgEXZ87CqsPjPzPplpC1H+L9VpvczP4IAYE0IvkBF3
hPHFcYhboFik+rtUsDc2lejfQJSoVDldzHlRKMzEOybUv2V5CYIBDs0yAsBwqmGC
ozwsxw3qBG50upDNMTDIklyT01o5UfWCYp0ZqK8tU+jaznrk2vFpo1bM1q3dx41b
7ztbTBx2mY1PnkOqb765dsAyYMPGQABgalbl9xIXMB6jBF3a7NPzDI6nFdZH5nm1
/4KVJRtO1hqpLvHA6kXQxSO0JvQxjWoXhmBmPWFpjdrSmRiT33e9yp9HRU+z8DVA
xZIfP+PptZWmdcg7YbNDi48y+iuBRCzurmXANPZ4wV4SLmizROc7B6Y1vh2XSWwZ
N0XDpPqG6dAmtG5VP9Qns534auIB2kKgRoGMb1LGr7iIXBpS7oKJJnAnsZ+CRoKP
2DdlQom2DFktzqm6JXCwVKI5acExt+NLfrzSLzpWT1xvpx1GWr9M9HoVzn4XHQei
DHWhbYEpAv0D5een4M1znelwWBoYvXEKKZ3N1Koe92eRyYeXR836U6KUlHpvUywo
NQu3kEj1xVQ1NG4Zc8WKFC9SZcgAG12JjQyZMDfRuMlVW5lTrjZOcdg0KjAuS7eP
lQDnZ1IYhRTebU/WDfAcC2dNGzYYfW0Ks/ArtFzi9Vw61nLUAHrhUQS2saFvDxRk
pKJ4SKFfRDrDpF5UxVlOHJE5KXL+ZI1WxGmhZiDZpADOI5rrbSe75maq7HhZX5t0
/314ygfaDhDKqRpY7S5RpgBVHx1soeXE0rqJoiA6UmfimLhsclB8GTku2PHqHy8M
WCdebaq+SusVrif0Um4lcJBU/DsI83JTgi4K/VYkwof2TMIDLLNHm43TF39liUAZ
tsqmCUWpqtDZCFUw1GyT+QT39idZRI7y/zmL0okRgt9b9ej3O4AsXqXvTX3F5lPR
LUHh/tIN4MNt07SpUVfqcCINhCSxufMEViu0uehoPTZkg9wMcrohA61m8H/KgIgB
C+I1EMCMd/McdKdosAobChDsckBzoS82vvuBMEfeTo1ux3O/ZzVVpNq1g4l/s9yK
pSGJtl4XXL9pNputD74z+vQnbEqHuuGRBTEx1CXqniYREiLUic9S0e3kqwHbojJQ
+yArD0xzzTSwakoP84q0IDwqHWOqsY1x69Mu3GoaeLUyL4nw6fr0yaWGsSbsnptV
FMeb6kqDRLAUfAN56BQa2l4o83eAlDVzA0OJUyOxsx+Ugoz6dQ2vDSzuQG6mppoL
zQ5bvqrtVC7CZjUqEK8AoS/jIZZedm1tCaG4rNEKcDBa4pfJoj83Ey0znnwehZgE
ZpSl9lwf3TVJRLfFjINx++U0K7JmQoELVmheQctrHZIdZ3HJiRxqaEInrMY1+j6f
uAZI9rqNSan7MYhMaB3/gkS9mHO4rKpcaFehyXtpQ9gFF7sPd11d1uCSx/XYH/dx
YVo8M9ns3kAUmM4p3fRY5ZollZuaUWKU6pPg+qXXK/CRssjQOB7FFZ1dB5PAcfiM
Ao2eFUwbkUOb1/nk8cslX2xJEPW5klJSOE+BDCJaZs1FZk07RmHuwqvMR+LDHvi0
lugNr0Cfce7sTYoHCgTI1EYYaK/ahLHwW16cHPmzjoOwCsB3P9UYAiMfyyuFeVTa
VOIfLP39AFBcsNs0S093wQHNPG3SIpF5q6+q0jJG1Qd+XgW6/wbNdjDtpv3+Odnp
1SsfsKJVNfHnk/WG/Wv6Q6qF8zjqUKUX2sEm4Zi05HkcurIcx1bs8IsfufxOJOsj
ow0t+IKcpEXYnBmnGZgsRo+KDBC3fcpLzjEhvNdJ6N3D3UllK6nmaJMWRm0bqvNf
hMBwdh5+RYZawIQ+xR1TYoX8E9G8SlIMtOwIlAIsWvDUeD9ZWtFeu6hZADY7j5ii
hgtc5SqbzQvjsQn8CzQkFefI/ZLePtCgmoHf9goak2ysHwiz71SQozfsNQBxWDJJ
3vKuXicfdccc1hptiQ3djDUTIMStmWyrG9UYuMb4L3ZsizbkFGG2fFvj+sya8DQc
dpwRTAe3CzmiT46VkE9zg7Z2zRBn6ABhrojm31GgSy/bjTkN/kmrA62PUzZ83wcU
N8XGHD+VBAAEctZOPjTIYRXPpNAaHWlhWfwSVBIQMTHoCYBLmb70KxCz4r/3U72R
Oa+mevFxUA9V7pqfAwraI5JP/H8x3bMHanLDrlE/N/zVbof4WK/bne3/KsV1aOAx
9DnAPocy+jarRRlO6PRx7O/2W3H5cSUaLGIbLJsqoU9aGg4EB5B7Aw0GnzU28FrA
3c0RyYFsGrAofeGM8wpY2ld8r11bUOnY32MO4QMBjDPCiSkf4LsHBPozpebczvRg
Nw9N3q6nJWqEyVtloiGHKFKPn6hm67KDM+IAe2HxKtljPX0uRnJp+C9H0pO35rfA
aETK1Jp/vbiio396q/HG7YdwBFqO9Flt/nGFUfSzsf8r5+DVvYKfHZxuG3mzVjL0
ekLq816AkzVx+9Q7Nx7KG5kpg01a6BPdqGQ+fFlvPr8r/S4iXKRbKwzECJ2CVQR8
uDTiIHNC3O1pt9VdZ5JaWJ4GbJPNEMI9Afb2ZRJlBkk391sEmeeYurSiVjUpj+HN
RJ6RPUogis9oNivOVO0uNSjc0GFv92NOLCFD6wCz/5V63YOASmb08gvGP0u59x73
qCbdcYeOQXC7shs/nf5XRgP7nuij3pvMq6Mw0w0vDAvZNaNMMz4z9vFxmN/96X2p
TtG8IpdU0DrnMoa2kzdly0VN8lWEKZDGusQ6BxJvt/0kav31K7gGHnIKDX0cP3ZS
GKZKcusdYMPB7GUfe2+h2KH1Ug1M1ZzcJG+8GjTkvJBBzFrk3Xr5serXpt/Dnu20
S2w6NuAK8hz5P/V/GECwnkGfZOaaUjef/dB+pUOdIA9iDjbdN3TAAya8qpXa/9eG
6lW7dilaCNESw3ypMgHFQ/c1ibQkylZeobCNi7z1C13KFaDaiZG7UmCypOiYMNwk
LxvvTzfT/UKtLxqFaHH/+D515Z9N4lpbRzhiKdmnhuV+AFTdc2AYfl9dp4+awiia
+HveCrNEktdWVowlbk+yO9PP1PVz6A8i3KfBCFKBo4TgG60ZO+cAojJP+yywBnV8
/HCW0YfCR4tSAvZVDYSWLA99x9ljRc18dOfa2vvAzMQ/uE+8Lbd6tUn2kMRkj/t1
hHgd3i+ZQFA//VRMqJ7KXHP2YFvZmOyCHD9InEtFfBbrTR6WwznVkDaJZLj/IaNx
ncpaiFvE9nT/LH4Iei1AEdksfKPG83ZK4m7zMLPvgzs7WLPNE7MhPexCzZeRVMMw
3nhCxCfihZOIk6MpEmq2qG07aGiF53Esd1fXd1L6XN75sOZGz8TzcQMUbcPjxGeR
IQZxUOB2DsMFXXIzrjkmMcz0VadkTql+UhZt2zUg/cccDKqVM89pJSgvMcTwIl1M
x5SEIxIg9A2w+0B2EljhZUrch8mkqLj6OAyqgfD/6g0zFQyg+KuUwG4dkxR+suD7
m/rswWf4QT6JKQK9IpOz1mJ/qm6GBxHwnzi7JjO4JX+gra8AkUA1HDV9F9cgMUhb
mNEQjh6tLsRMcWgci2wwFN2VtkWyGJAhY1oz46mRMgvpZ+HnmH28JbsFPAgmpHx9
LrNM6a2DTfMDxwTJLo2ZDRyf6Pxgfx+Kzl81jjYX7vIXmDu7tuY8MwLohSokCLev
dq9j+ljd77nBuHj3hSMDMdAMseXtyrypzPR2tAspiWj3LilJGUTETQrbOUxwszGL
VcyUiTJLR+Y9AQ/kSkAzBfTeM0kIhItR+OTk89V6nI2+PRIfdLL3fL8Ar6c84ilN
jwfmWHRdDL6nXuxL4ewLQdIrN7x+97ruHjhZt25C2xaDQZEdg9WlXJ//s4B6hhoy
5on47Nqk9IRtkDYpVteGnAwk/yNNjNCMKZb1ocyzvS3Xe7Th8HwilY5ugkkYIkwv
qxUuxo8IJCTNj1xykpWIA+dg3HkfV5sHN0vsKwNfvW+1WPeFBwl4fZOC7zToTRLg
iIfX4ERDn0qTqvkcKbxR0Y+kxxAOyFghLi0SKXXYgInbtIXeXFZDZiUmbPbd/hxh
h77MMuR3cX3Bp7y4iAUvI/DZch4wxUPjrWWi4WVV7OdnS2XapRufWOFSW2wqik0N
DLSHpiLoxgffww8YyERYQvItNyiGDB8PMwxB1bsIw2z0nJGa+OehgUw4wsNSub5B
pq4IM6NqBNbwCXIYYLXFl3REb2fSgm0ILjlSkmEWFS1nxUz1805JXPoYuzN7ORE+
tH0JIo4SoXYbWTxHZAtaTImlORp4VMOM5Has/6Cnbo3KvgkiPGqTU433sLm0AXGV
eKExwK0TYIWDLCc8M0Po4JX9dPvBBOvblGo2MAISMp0xhnaBHU1n0cbjiJffF46a
nTt5fJwzG3Qc+FzX00zVDbmqb0f74YfLf2/xek5y2eQOvyCWihwoiWif97T60pHP
24wLqb0XCtik38lrqjVIU/nyUg0ouB8vI8jiRk0f/DXQm78QQTaIXZW9HNeyxDGp
qkQ1v0Ji/12uNsgYdPDSlwTE8d2nXayqNt4poBzzyIjTrjwvHue5rHa0ohiI+2/h
bsCIV7OgXtIbo4vjfott/S7N61Tbdsjn0ii2wsVy9bPAvdhbYmS1Fo5fQg3ub+t6
vHdHxa+xchVLi1dDtPZRXcUtPVAH+vkkJHKbklAxgTC/f0imvjJMYYEx9qJccUAA
5vLtSOss1ynB9j9RaxAJEy3PkIHPqt3KEc4bCjORqYE9aOm2MDRSC+3e/Tqrenh+
ErF9274U17Zq7HPR1QXkYiTV5yrsbOUgwUqzGI+PHI/mjKjI18ffbhTBQ0YGOUYI
E3nb9omCtsA37heUy6fHBupQ8zmQEMMLoHM8S/V4WBpJZwtk4TJkybcaocOpeCyr
UTA5sSpRORaS7mB81QQnRKmVEwL5803W83cmq4V6NpziIxiesHYe/S0ITCmYCkTe
egwV0psZWNwYwQohJYpzHaXhG8D2JaQF8zpVz9fFTIWsR0elFpYzesZtBXsoGMfe
xaVftVvgW2B5Z3kUCanQtt40arwCMCSNBDUVJq0WhlDC5ZklrpXziDKKapiwIUHb
SotVQMeZ8Vhht9+Lqh3HnJPLk+h0TrjMQcOdi2bdiRLKidUeMurN7PGtj5NxI7v1
qB0yoAFR2U6duwfQ07HgobPxPIdyHf3QKI7+uUXZBDAnqF63d6pj/Yc2Kfj/wl0w
hGaBT+XKWzJotKMxMB+Dd7HGvgNMFt3J/aywfgpJoaMjmSZwTBqNbeDeIEWJx1T+
gRtO5p7UOz9ZuH3oVAXCsb0LPaTaKiQuBPz+IkU9dUcwUgKTzwcjOr6CbmY5P9zy
PiVAMIZYqH8wG+kvgiMSEzRx9j939CA3g7xbKy6iyhBtGLrqexb2w564Gfq5O+jD
Wz2ynkjP4CS05W7CCE1ZmGY1w5JaD2QhyW1ZxkbdADYFv7YhYXb+dvK8wcMBsrLj
fIePK2ilcZdoZPm00vWF0BO8WLEgmRKSI+wMilnCikJHcCPEitjsT80VXoK5zNPx
QPNqubLiLFXoqxoGUtRkS4qp1VcYrRqil5JXUiBuVA/ZHQCkgLJQ++iQPiqdTDna
XXsObRLnsjgu+DP0fnx2DE6Vo1tddBQEC63zm85qchoWTERvVHNc4tD7AwMNgb8P
SK2184rsmvX2SCGc6u3LtjClOKzpQgN407yr/IYtwpU8+2RuUWTCNtpniM6ANXRD
99Hto4cM30KT2KLL/BXRBQjhQjtFE5oKcopPBGwoLn7LZKGWBk/HFd+tDIYqoVXl
utVI5i0zDo3KrInzdkzqIWhTQZVDaalbDLsXqtsrAkScpO+1Vox0NaQbF0Ex4fy2
iXmDdd+3wTAKxu8i6MLw6gFANqpThODHCetTOely/WFUPJoxCz7F1oJTKLvL4aPt
euGTcqQDsD41SsB3GaRg9v3cZRWsetJo1ArT2/U5PhHKBdc4NhwUqjzGkxMavsUb
9DUaH05xwoy60S5X3YwpKzoXGQYHVXsus/Up1TF69klZWdguSCnYEch2UaoauMlf
ANTaJp50NDHO81ckrtwLVZ35VfjMcOnylLYNSSLBUxodacpp+4l6KesPAsEfNLim
L8V+1W5Lr2ZL1r58oZKPP0n2zcbcAaq6kk1JHDJBS3nG8kdIOzU6HrzHaENFM4Mu
vNJbVYvbFrE+oI4YPujNrpeYb5SFhtw7LKosBwsyElxvcXr5mm+wwbD44B+L/MFe
fAY7BJFT0gDvPyhUsV1b2VVYD7HsUcvKNLMqRP6UeWE6qRM87BgVOpg4KCJhmzxB
6R0OPaAbXD/4dv69UoVtYGtPvf46AbeHFcGJ0+S+VfgCHRwlvdjhpu+zE9ajQN2p
RkPSkIyjJyEQqH9Nf/+i6eKt1JREfJkSqsqaXKTdMRXj/Augoob6xsjL6eh7CMcy
wx3fHIF9yVkMDftr8VW4rzktAbZ3CwknGAav9/590L8=
`pragma protect end_protected
