`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WhgG52taTU0im8a7ngJGiXpeMD2sxRuq2gzM8xUPl8TupAWIeJFPAt1VKSzDGUeG
KxerH6uvrjlQrqln1+QCsvRy8zgeQ3eZvtOqaguQ8tLTzboi6EaeT286ugfLxIMo
I5ZNijsjwuez2KsNCRTw/QgkYHtdcXKOqg5fYZ78DoU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 98768)
TuO2uUWbqaXQH/wK2dEuLCLNC8TraJR6JtRMe1/iSzKILSInZSwyOnIhYkgEfH/Z
QkaJm67Iyhkwz2q+FlqZ28herNO+x2+Ez+f96K4RlDQMQNcK2wx0bx+mUmxJT7q7
LTaNP/1VcdzmFjT0jDVavxlTXtA8kDhvOIUX3MLLXagvVSTEq42IkgWJSg+EUz+M
d/2BtrK+SravM1naX9zrwpvjUdAQFi93gHIYa5xipvqotx8MClyFqYhpj0m9oB/D
O1if2fTmdQpph+bybR9+G1ZsjpDBoNDbXOCum1vH5qjq7O4xLQV97WsjsH8ZBztE
H7HTFHIB6k7MuShAKnFi4IVFr/bPjWACyZe8kz4Fk1bxA4X5OuT0/cJ2UlsXE8qd
NHOc4sFuY6+z/4wiDS1Ovrjqehn4S0hdGuNiUdKRGLLG8smJosawh07itbTjQqlc
Njzg//hgqhuOORsnXQsmNIFw2AglgTIZYrsOKtyo36R1ev4xz2I8Qi3szufnh8+E
H5F+mAWmJcMH5yUTXd1M2IcfcNpTmauQtA+xxjKJQsc5d1liGbJ1KbFiYH1N/QVM
XyLdZiic4eTvK5i7fOkvju6GnFvAN/OmGayvBazelpogtFgDRg6FbujvUJ05ZJBt
MTS41laA2yISjt29deQ5lAW81FYvE8DYc90Gmm6Z71zn7DucNNyoH4IapioO/hkZ
SpGIsaRaPcGlzGYauTBipHRpwXuhHiXqfQZbbs8T6TR7t+Kx3hLxoiW1X+efRo0M
NvZ8tb5VwLZqJkz/VnoyU/jRWkEL1hVCW3lcmtyyEGOUJNAmKqtExAuD0VWV39dG
8FUTKmLj5vYmkMgts4ayFdgVrTySB4CtsS5cE9t5dpYw49lyShS8x2d5qwt6Dt+3
1y/+H3ia0vvH8buwn65hG3zwBUsaUUPvVpK+EEMR1vbApwaMiMRtSR6SkfMOc76D
E8GYZXpzBphE6A9RqM3ny+l/72Ar+jDqxC6lrYYlzNG+hV+J/PV7bio/4Uq622Wm
qKOaDm0EfYV6BXPvBvgsOB+PVvP4LgroicRBbG0qCB+SrKEo3vwf6ZU+riGEi9UP
7x6L5rRnjxOj1mz7CA5sRLroySBhsEpaQp1DC3FXge+x4fHNDPYPPbyQvOcjx3A9
39NJzTut1CQUSg6cTaXGbAl4t8xpUkPU6WCMTjXymjg5w5s4tlE2GEA8RZ4LvAht
XICIljm/GEQQCJOGGLOyobGXHKFk4K+ML7Sk7AKLABpI7ala88v2aI1whhAvRMon
FuRlI5LHHTdP06gzrLUyy1m0lJN9eWah0bBOJ7wOwRZNrh4OoWx1bSQv6lyogTA6
hnnDanQEYPiWcyv24mMum8audAMW0EqFX/tWI1bHs3x8/DIR/6OgyJx+Q7pBjNMQ
Uyax5M9jgViCG5yztwbO8aHGbPe3xypx0LQyTHPTZQp762us+T+zK06sAUtIS1zh
IviJRQJvlx6pk9NnZO5pLN/qyhQvUA4K95Lw1rZHAc+m8c3hhsVnytaJMxopPRQd
T8UuM1p4w76KNg/j8v6TTsoCZDG5qeVzZoJG71axQKj4XwWh9oOZqlz6idaPhjq5
a9TGsZWrquFF1uztkl4oaD6HaoAEeqNZfkQIVmEbVehjpbkCbambEkEaoBE3aa12
V8atIi+kIbnZ6OhKw1KsXx8OI3pFa+r8SFkoV5APscln5roKAlcHk3xb7OUHrcH9
8kLjcNJ68d1VIveMSYrYU0Yxf6aY76GML5cLySu0yl+rCuTpHH/wwmCWbl1sKMFc
HhT9gUNAXOhp9wrLFgxHKr1DnsOGFNpzzVzM1Z2TjV4wYHWPNfK/TI5FswB95Yad
abkoiFq6zDptjj9H1ryhvujC5+6WnGVE17M5dVgwSDueE/RispnfveZyEVAKkMpo
qgJb67bCZgdjp5qiKdIOL0yUyO9994Gll1pMMQOqyKR60FdpJd6Q68Xfye3XYuXM
4BkvtUe1yO0JJiNGNqCsnIyi+OGJfVgJTP1gIX29BkLp3BOHqz5vB51e+FEcNziq
lrIXvpYRrjR+8LeKBcGGmPAqL0rrcEiM4ISeVKe+2XPOlGn6WoNrIaak9dDyGqKx
MiH9fGJCOtgw6CB+wHuTFo1N3TZG3HG/rfNg/ruAJmrNJ0SUrFgkIWIRynbIUC30
kcrl0A1U8La0MBpZKvOUt5KigW5d3plnoogfZQ9PSW03pXf7mp+am3EFq6FH7hPU
h0h+Chgcu4smz8bXdsrQTx8OadD0R+tD3uIrSjpC/VFZ0iKXXPVFENomYQy8/qNS
Lb3nF/OPIAMF9BKS9+nVJT9E6xN2l+2QlqMMlxunpUV8CkwxbETHwmPkHFOokFkF
LJeRBeRcGb1uHFvO8eC38/6rwY40YbI6628QGFDP0zfdjoGAsD6HcbCEakbNvv8m
ULbJMg6aeupNuy1zUplIKjLGoReGJhUluH/iePNqaN2RTPClcDswsJccncxjIw5x
fpnFKXPH7ktv4axOqPwHUjpxU+LzlqCxJJHxSz+O07yDe7hz/tmTC/p/oR/Mqc4a
/caTV3KB2IquIRciYPCC5A/wFM0Jh62WQ3oYccdukT2k7/tADm9xHvwahw0JFej+
J0c53HM4OirXDDHwsUlZKFJLgDE9ZcLsxhba1ZeoD7Whnh3rqPE8toZUJBv+JRa6
sGwn21RQZbG2i1kdr+tAtqgQlfZB0CEjfYp8SFref+/2wgOsFU9N63FQpxZNBQgh
6k0iSOQ1NRW4yt2BxUEbYNzi+VlBhnG+cIhTpsDZ0tFAU3wW7eEYaZaCsDIRh+eg
KEfr0Yjfcbzt49LIrp+IBMjPUJkGmjZt0CXOtUvWFdqloGy6nVx/G3jefBmfhowj
iVyCZF6LIZyc8FiKg/tTZ8PUPurjBJ/ItnFrUiNbVSENOhobEEbdePnXAun3EDug
rH4YIBi4duMZw3TXZM1M1CPnhXUd/QmVoIuSMN6ea+oXSYAESzuhTNEIOuz4EtSV
c+0LnMdq/Iuqc4VsknvtIK7GJZR8eCNfroKEAoAlhcyP2tcKf+rnWcjW/u6Yz9ll
UMYN2jpQp67mvpUUUr2UbJ5EpTnPogtPTw96qZtbeKuuixBTF+AlRU5ExthNDf6Y
skRne+pJFrt+UDY/hFHPVhtKnyyUzQ0Japfvem8wWI8AC1+mvMM3++VZyFA39AAP
v+U6PgNVkD7dyRTKHdCEqViUmNgbvNRRTxT+4phSxbTMdOWnRCbYQH/LG2x1sgQQ
Vs1Rw1ENUL3VSXmWbBl5S9PcHCQW6TX4Ei2JdauA5azzsWE6i9ehZzVGhIIy51qC
ZnzNmJkaIPeD+w41/prf2ZWWpVz6uqtVA6opRCQ5Uguxs6sHplQVo3iNWRsk0iRz
S/iluwfF/WC2uU4zkZFTkDtBWbwE3ss/7HZ6UFpPaa8eJAnOYdBTX3mYR4OIDBNQ
gGGaZZUV9gs7oU5eG9b0es+c81sfDIfSrThRwNPm5s1Zg3PblCE1t4oqbxA9Qyu2
cHUZ/X2ZlYg+X6iITJYROytnS4H2EDI03O0J/FrAaC6rn7ervxLt8oGs59uU6b/5
to+FDFc6ehn57jqeKPrc9O5O19yC5NnLPj9xjJ+P+E1ctXQHeYR8TqmRQ5ksd2Jr
BnyGG3cmeumuuuw9Xg0ZO2tXdcnB5ZERBQjY0JHitf9cNHScRIvbsqaJ+3obF3Pz
ifg25mC9sruf/FxKHjwIh8G8MFQgWeFL8jHGh9d26eFic3tOGJyr6M9p739Xg5r4
ynjSMl6b2jTUvghLr7wYhcdtD1nN4jf1a/46Zqv+WsTCz9pxR4caKY7GYZAtK6YZ
YLW2sU85ntt8kR1ZFcFcwmifS85q7/5Zx6ox5O/pgTIGYkAMluirvTEw/68Phg+7
N/bh461ZrBjZkzJyAw9fx23JrUmX3ZXs//oI7xDLZbyhKDfhHQghI/hzHyz2H6o0
BY7tqcISzq8p/V+zYrQt3OWGusVmpa4qFfZn5brq1Iq/Ju7nNGoAJl3BRdHc3/cp
WwIaBlkO2TKuZiKDrqbcb32mW7UgSkKeqa65G7Gl486TmmAKs2r37bTyVrixCiMD
QJQEEDtLvrH6kZ38XkrEXL6p5IOFzzb4djl8eUxZQwsuAvZ6CSlCOIdNO0Se6cKf
0dBLHD+0davOgwXU3oUTum0IEWc3XrOkpAhxbK5L9Uo8DNBOx1p5VURZwrKKZpmW
/UvbiSsrr9O5+aahRQlmDrdr+oA7Lv5/4cg7m1QxpNKjxMvp+wN8R9zKBjPg+ooh
RXO3dbTrFAKEvMkM2Xz9Al3khYzxQDk9ZqXxid1FuTbMfIDjj2XZ9czLFAvTRYv+
dya2FxPK//AMQGDfDxqtNblN4jmu4rsSZ440aQbjGg/vyrS50inHBgMaSiadfG7x
9znXTEYAgEdVHpx5c0XcQxjqk2cWj6LL1LDoqf0BP8wGSbGhnMV7vhg4XGOTJdKD
KxxhhVLqu098u2jFWZgGnYLdAAL4n0NHrLwo9V6XKf4j5UJf8JPD3jzUSDSuh8nr
RguqscGmkNEnzESuA/XWAsOpWooGj71mBVJa00JCxF9UpOg2J/XeqYbr/CN7yf8f
qZpkCt/NcAXfcfIXZ7XvKdtuspzRFUnBEZ/lOvWauq7XH7DVq5m9o+hZ24hORwJf
aiQjEuCNVsd+K21GnRbEMKFXkmnVHXrFPlkQFbYuYOzgEIbhJZF7qu2xZPv71mWv
EqKeY6zzQBWbD0Z3FSDBco84jgDLX5wPx/VZ7Y19ZGupl1RkOTBtjQvNobZDP3PU
o3KNzGvFPD9KUVBkeNOjvCYkKAeW8hrlRSUxGkDXOM4IEva46bglj44nM/o4RMrL
6wI7pzWVVovchClrkD0XWIsAmVLIkaeJvL+vkGNnMxQ1eJwEi/bmVWHSq++K5Vzv
97f+/PKYHs+dF7hYr2lfV2CdfZPOBTE7y8VkEp3m+c0/pleMRTtzs9Bcvipvt3X6
/R+R8VIuC8NOSyYOTq7KSxXndWoG3m6OoIZspbYrDHjA128Q9BmgC+b/Wsxtre6I
Xd0i0wZlh0YU6X+Y5IRjmJq1W5zDJq6p3vBXwTpzsfr7cbUzTavwlDyftSr60geA
w0GUX+K0iLv1YI3ak+iKmoQjWL/RI4nQG0EXCJ9aVLyzUCuxf7tlyjeArV5iNcnl
KqI6MWWWxYdCRbDP8pBSRdjs5wBKI6Asvjou0Ds5J0sWMT8BSnoOJnA6jYCOGVvU
vL7lhzRI5vbHcHgDTYCTArUK4YPqYUbPSetQU2AuZ+ZlBOWvlLijFXfbUtb9E4mo
4JdXP+Kgwfvyo5QgePvZZMO0iExiZ4T92AuuCdMTIa+qCFdUf+b4WoMzjAFhygih
J7j7darhw10ul4a/C9iNg3RYxy8wfsrVujqPMlu+SNxwtKc2Zddd2B4IiowNgT9j
lzopAKYzYb+sveEyAAlhbYB5Cy3tpsgGTZli4HmEGsKsYbvfJxi4t5iqQr0ZZGh6
yFKoip74hI7z8cASLG6TIQMu0adNBfRcucBtt/2eZ5Y7F+9q3LBI1rXwB2X/kZ6k
YLP/bX6vswkuTG4uuy6yIqfcNwgMcTmszM9Phskr36VDtSAumuzAzqaRfnMmKQro
caWy2wIfr7GmLfSl0IpkjZie8GpHbMuC6LYfi2VvNeO8Z0HSN1s8ArE5uGnbxxo3
YSr0Yc8BP7qNffS7rHThDYgVAgZbBT6YrXeVpfoJ+JE8+9rtzrDBRBj99ESNSGIQ
Z0TOwfMpnvnUsh2S1Cs0wzO/mvM/haguv0XFWfb8vCte6Po3iS8neCjZzMlwymwT
lIyzbqeTO02NkgMLAKm9cC8liEeslROfYgjrtQrqxTaNYw5XtFfa3A395ptgTIAI
CIzMdDGT4puouJNUdBm4huP6/D1MKAxgHovSPh1H4vrIquiVtDk5nRU5do6Spqnd
KPFExhagNuHhgaeldroP2CnAUz1EPSIw9I6pKBk35BJ1l5EUHUx+YYUPwxsHc+Bv
Y2AHG9v5TJ2aILyV1Om7xL1HqQuWU8JHJiYTeKGAcBlM2ApiRdV+p9uDM01793hO
UJ6Zv67U+CCT18XVL1ukNIbF1b+0W80IjX0RWRKAKmENJDm2NIOaKTgv+p6vxGtm
iBv/scUoMYlyh98tKpK26U1oEtc7KKmWM0HTrPS+JAPLsWgnvrJradEW2UHQzJe2
dBNAmhkTxrElG/oZlSkoaS0KUW2lqU++i8WYwegh84XRj0RMWUAy/zLMSJoAT6Ai
4i0N5AOfcLX4xoyMdi89xjRLbNiEtQEI3Dw8zXwXQZdn3qIX6GNlhsrpVz+26U2O
d4ubFzhXubcemFBQAMBIDm8wWdeDbNtVne/8NGtwuQTTCMQBsxEaH9SqD53VVIhe
yQAzDDJHOL7uQSumObKqhZdcm6avizF64jQW2g6BB3Kv+hsuvnu2PWlrRFYzxvKZ
875rLMBcvlem5eoQwrbzLtLsDYGeqLBHimNBXlqDmmt4HOGZxfK5UlYGiisMur1x
x/GyDy7rEtkhs26/iAyXS2PevVdxrQCyievpH4Cz7O1WA18FVSprxIyVhlVgj0jv
zbYJQvT0whlA3QWe0fg7rXuBRdRg+x1wZ2t2S8cE4LH6a0QPe4Qv11wwtgRjTBIR
vGYejj9fzvpHry19ucOzauQY8bJ69y25oN7NhsAWhDq1+xGzVd4JRI17bkIDaEX5
4UJ8UIVbIZJ0+kkB5DpQyph+zFm3yOR/VfZm6CoVhCtOgYawJiJ2rA4p5uw8WEIl
4WgbX9zUz5NSKGXQVpUk2w/lm0/5vHvXsmwHW1vEDG4I2ZluJJT4njanK+bbC8ZQ
cQ057G61oITVViA8cupJPTYTsSBzXHaoRob+8czjzCCj9j7cqb/erO/NT62ZieLP
/QQMmlSGiwG0i+oaERPJlVlB9ajNy/FPepuifk5MHt7QshlV+sE5YLSf8GANwvXZ
X6dhxrlO3TBJXgmPUXueu/a5cTCXqxYaKFYJ5eIm1EKXuAbORtWuix5IxarHhW9I
zxMmA7SfaKRHrQ2uv/+8xHq+FNiijMBxO4EkCzG8+ylsxJgrtA7nLcD5aYz45iho
6060bYyHpPEDcPrTKe+6vB9i76byihKz2FTO3N8Tinwfc7qvRDB1MElQRJL+ekgG
q7laUmSE1ljgvbgiH1ae+U1oIhOIlKTJS19iCwEDwY3l4S436TxLNhMltf/YQyWE
aR9CvLgnA7ebyQIOLY4ufIbZLzi8dQU1+yBXgWkwyGYJ16fQGOwqJwUExap8nGDr
HBd8vH/u/dfGbEiP0cRSC7h/v8JsRx2g98rLqNa6UX4yHWRfozJipktnkrvbA61K
jN5+YrKzzfJr29g723g1Xu3TD62UVCGpcUSXJPRT9n2RQurstHqvVqgAGCIVeFcs
oj/Z3c5gO6FSDA8QY3fIUTYzfzwoXIPYV5t+oYtuXILkWqv1ctSHwFqVyQ30DIcH
da1U3Nh/azpdul9N4JnLkcDK0zdStFfJG9f74yEbjotE1qgyVocbeBTp8ZGITqI/
FXjdrzQkHTZNwwAj+UJqla/UdWF9hKNrXjbbyP+d5qDVl8bFSW0FKKtdMJKQGT4I
mFYJnIFdOn4PqJ4uEmZyvg5/6od5lMyzRX1R0IvV9KFfxNN7CpfjfHI9MbV/0sLN
jWiYJIYAC/BxXfg/uG96CJ3kH3pOmAruGJYsHr+/ySFhyT6PxMf511AmvQ+R8fUg
5a/0McQeVG7nt/wNojzC+HtOkSO39r4L4sDj+v0EWqKUYlRBKERJbzd3HI6RmrTy
cd2zEV37kHX9qUf9Ui88sT9slwHZQAIfFcWaIAHGHAAhf+baBjRpen9nzE35FuOV
u/s9FD2NQT1A9N02MxkiEOnJYrmj4t4oq8UeGRyfna2bACzD/4kbyUiNBzpufVzh
jQHLCSQ/buqlNRnkcNOlbAq+XSS9QmXb+wD7kC/9GfneFqHK8KvIseSB/6KCVAIm
P6VNv/AW9BQt38Gkb4hbtdm0rKKQ7gSk3kvW2B0CLPhVumlNucxN52QSQL5yRbLx
be3G04BlCr8yV4uQEAzhLDcjLDOU8YQd9NJycVcdSZNG7WE3umgMM9jd7NMepIPR
oI+y8jbsDGtZUomM+mYybhUhJZ9QDkWXnKSRo6jmqBw1NGZ+uME91a8UW2KvyeE4
SqNitErhOH/biwbtYxr4/bRhaUj4PNfEKedAIvJa9Nuzz1w3JwkhoDmJx0g/15gY
4/pV8F2QbRvv+Pzar361tJvXx/mNWvjj0TCy5IyFDzKiC9322lBO3j7GIfdsXYlb
ENXR4VbvWG7YDlOZWXzPuT4PXOyANhqruqrwWcztNN9z/NOVexd3ADpcbsGTOmYJ
uMim0TDAHLUC3OHhXz+VW6yOUjBC8436b7fCx4aJdbP0qJbZDTVu2hBoZYF9Nhok
IRXHG4btmJn77l/TAf1ZHIOvmT0lvncVHgdPEnPGmxCEXuLeHdHMhKST7Lg5KOe4
H0jhGX0SK1fT+WCUXteR0YQpWo5dQRAyKbcDduLt8rwNIiUiJtVs+/5EIj+1cm3l
dwbzZwqWpmBjGUDFRU5po9YHhAKZbLfT0vUbGNwEc77yu1Kv2iUqFONZOyPE9eMv
LJQnUS+1W/0lMLCZoHpBubcPCODPWRBffr5l5yaeYNdlW+K1T+ZYJNuEXheP5X5R
teXdT7J4qygMFDsQBMlOAuLZ2ND9avEQhcLllDkggHeBRK/1c1tt6eqgn1p0B0Sv
O5X+JC8uTV72rjwZ6UjlKmdQR0wXpW1dUE6FceSUvTvXR/YsJliOkTLDbuKnwMxB
wJMSIav3HAFV3ALvU+2Pwi2Sg/ZObBnXKPFhbF9c2BJO6wbFuxqOnoD3PbW5PEWc
28dzAwaGG7ftHR6RoaZIskh2Tj4+q5EfCo6Hl6s/tZiU96+HkpkJCZ0YQVNZU6us
FuKuEA0+KhvKTRvzCYEx+G2z9FmrCsURWluVSAw2Nk6hbtl/0fxCKuhDGEsXH+8U
CDnKALajU3HYMaviC0pOY0jqmXZLzG3zrg5dta3M7tK742TZD8bI2wH3ZOahuS4e
LLeMp0y7BEb1C4l0ww2Aan0HlwJEE7dlTvYo+biys2ltdZI+80er5WeQloUtVQPF
+4qa3vTkoL5XKjj38CdoyDtnXvTQ8Wfwpqi/arjVM019t5fMmo1iEf5E2TpA+bIk
6lw+EO1nlzUsVO/MVjQoLGkeUecHX/dzklYuCvfR92RYZBNJPm2h9WZ2UFYi25bY
KWQHhTUzHw0r2hn5Uevfc3mEZRfGUXcxbSEeH/NCeQknxaHZNWk9QaMon9X+KQvb
EVbuxFZ+22GceBB4ZSMVotRutFnPpnGUUVfvbt255uUNLE+lIqM8ngwM0Z951oEc
nhZS9Zks1EKF5Ml7SiflOKRv1x9aLUmz8WTcmFiLxDJtZ1Rgmk5t7HIlcpNT3eBg
V5/7yUOFy6ffTW+Fl/Z9s5XFBLyxIg8N8vjCAB0CSzDonX3bB2JS/Lm4lCHWAfSi
NdBQo+SCBOYZUc7t45xx3lyCfU0MKCEPxgHCE6rfELCocI6iUgHbrPKdn5vho91d
Qx17cChKMfr+5eZgYlA2zz+LRwxJ0E6FRMmdXVeBN7pKTOplRmzv1vIEN8VVHTsA
uazV630Ei7w5EqCD8CnynHfFfoivOc6AoyWrVdzurfxcTkcvYAKPMcdQXgql9Pfi
bjk2d2jPzNIhTBMsbv05SIJfFoDswzvqezn/9dn6j1U+dRDVyYCSgy4xEvIsvjOD
qpMfqh/ffLBnuMEsk5wCdv659DQMVRkctKxCZO4DkIIj7DG3eRSKsF6K7BhtHYbi
4YkusYn4pr3L9Ah6D+NIrnsDQbiBabKMAfx13eYXNMhYsrs5mnYcZSrziclBfcMD
r28K89PJHC8Md+Ne6Ee8MhqePNqKZ7UPaGd1rs2uKXpF/efgXX6FUm3gX9X2xBOP
EzWAN8i//KAD/7tiFJZZsD8xg4Yv5D4cwaXgl7GCo5mJ8DvjrDr2MxYe0ki2Hu1A
1h+zhDJ6qmulcNDd1I+0t0Q0pL3OoCe9RYEN0joZQbPRP+QNDtblO0179yQ+y0RF
iZjmG5vMxCkS2L9p5jGwX1N+6j0z5A2XmWIfggab+OYf+kwJmb3tJXlAd2ogy+MX
BkCCQDfS4Q08gm3kSVirF9Ildf89FU2hpMus4nMayxqQO4Yjbzx2x++ymD7xvNnb
0mTP+qzsck+lzIlpDlrmQJg12rRTBViNGkh7jJVYO2yN/Ydxcw/awaXtlJ6frTl1
vZs1fdW8lWiapWJ/KQIL+x4HE5k7nogNyJZx+oRAmOqr+5Bcqj9laUD/hDe3FdEF
vJCDdFwx6R/qJ60IzpCx54PQFu2usXbmymlkDrGIAu2gqNNrrJA9njtZ/pOID9bi
Pooacg89xNvu90cnALR+ioSvZjkxfuHgtCgfKYfV7QOIX0zobiHmnvyPbazZPTpB
/3opFLi8eb+9oAyJIGDRUQlZ5AT7BGUEB/hTxZ8C8eMe+xgFhJVMA/NCDRTTkWXC
NcTBuVtrWJNyTY9dNNGWUCW6VT6TMttg9AI5/sZ1kjqI211bGPqXm4FBiyVQsm4O
q/OGE55rggdPJzqRWg39RT9W1kP67wu4cvI55VVHMoQECtW4WmUqlKZPid9ky8dG
BNCDWjhFasDvpJ3otUUF8i4yx9Hp8OSYUn+NZwk5rc7Nx6c3bKm3lw47GJA/4aiw
I+7jiq6KvVTl4C1XMCQKgzH/+5mfTCIGuLVK1X+W3Rt7co0vSwY9EqHPLcOno1KQ
Vz6z+X4rp4QNOSEn470Dt96Js3BugpejwOu4OOkwvuilwZR3p7Jt99pXDHfDdmhn
4Fa/YbmrXhBPRMM/UcwZSHwu8TlD3A6ETcwlmEWL9DH0nJ5jBm5uWz/wgXcFHbTp
ve9rCZXeTeL+eTt/+mQuyVK9eDx8+VtHuswKtJwvf3MloPGYA3bhJkN7p/pSvDzf
piAbt0/ehzWt1USOD1wGGWBEytlgXWkYe1DDZ0tezRVvch28fiifufFXHWWMyOt9
VTelrCxUemXgzl+GUwV7eX6FE4DjkSz6tXn2mesTp1ndEEOQqSfRqIZxXNyB2DWZ
oolcx4hLAb4LcqcJSNZJmGcUM6cDUsxiJqMA+s2IHeSW7cbppfektC8QZ0ByLNuC
znxCFRzF4YaK411okhqCt+YWD+5COGrnQIPrxE9/SS56op7fZkaRJhGorFD+jpWZ
0BT2UVWBWDGJ2Q6uMgM/SfqVizJaT9pryropmGtCejiA2nMZmkIc6WhsQYoXqSqm
vlcJXdWZN4cKt6vjz8Dt0hZSh0fXP0UqA8R/be+w9bNlm2hTzohrFXXv487Ia6xJ
bHDCYKWbxBHBykeOR33v5Sk+/w88HlZEyszbhOK4doHypyvdOzM3lZyb5nU1qjxT
I2iibUsTA3fhLiO6VMktICRz+Tu/w+979wFA1FLYj4I8WhPlsza54Qit5P3M2Kss
/2H+jzRh5dOcMyWNmK2hQsd8mxD9wiHpZ7rL/3kbMVDPCEIaWnhmvmj+UcALi9qb
cMnGUxBMItcsiiq2laXeNfVDUFYlNJrdU6YhbVPZw/sZ4zLVbbeiLwb6vAdbPQUs
8r1FSK8gLaChd3la27pwk22Gzl9DoY0UpIpAZi+XRLKj0X7RDdRJ9LKyAflfhxiq
jJ/2YI5WJI4ugaAb8QiCcP5Wff2HAMclEzg9GG9ulliq2ZovTsEQAgV+13C7sJCo
trCiW6u2loC4M1z3fml3AcbGNf9qkbuBP5p3CSSO4VKmZPdQJZ1DYOGCq/PTGsWp
eKr/3f5pyhSn3sA8YKR1serB+BQLKT/0QxRj0c5saFKTX2pEL+XLnd774TrH2BhC
5SX2PDrcNHDvwJMglBzi4rwIKiS1gIwLHHpZbrX64opbd6f3+e/PRsd+cM0LBxDv
ekh6cpXIW7d+wp0LXVjV8DdQ7xWpi5wTV9vDJ+piFzarzlHbzgxFRUVwtHIQ+3yT
vnO0eIoqtxKrj13yF5b/et4f2ZOE9Uva2PxfGHVY8/uSlVw2fetnZ2Qo6NuuMVtJ
EzfckWc5y49fhT4T3ROorMdyQFuvWPIwy3LmtxAeGfMA6sThUW4Z+VGnIFjeALUF
MMrA9U0Q8EjHiIN/eXin9Xtm6bag1plMb7nmYNODiVuwndMpBg2TJBugvfYhnrYq
vP2gilodpivY9Vh8S6W/eIe1WJ0W9PernwTAAtISDrbP1RHXKikrxPV0qFL1jNgn
WxiGliscRr2H4BXLjkSPJtzoq9QHON9cO2JKkItXpqGMQfZZ99EJLLz+0/2mCYpH
h39wbI17ETYnEAtFcLiB0Ia6p4Akd/3G5y6sftO+UblisWiEA7KfmVqBwCBhHMyF
xtmeWGOK+J+nBTiugSM+jJGTdKOhFZukKCO6a4D16E1cvAL1cToDxODnHew9/X5u
w8GWhPKoOpcAHbMI957qHekx4t0M3pAi//51CNvvV8kAzMuUZ3N9bSGnt8g0hJQh
Gv30akuUdQAGtH7GjMUDaubyOCmV0kE6YagLoIWIpigosENDyIcySWb7Yy7DncqR
LIS4IL4u12ISU1E2f/wLSips4UzR2KX9vvQv2PKuJxwaM1EMqie8uhlg8vQE7qyM
twImfhB/W5Q1iWl/CSPgrV3lqX0tvy09foV6TbJ64qFAgkN6j2IBEJEUiet1dRbF
XERueo5fiz7bDYir4eB1tt4LxYNlamit7phN6M0ST/jw1hQ7WrJ0mrJAr92TdyMA
rlP4P26qLBSXiMHiTAMe72Um48y9tO35ApFY3aVhQPN11mapG97Nv7g3lD/KB/c2
9PxAwZqbCirk4qCMWvfaAVmU9FjOLNxIqUqv4eOh5G1I4NwFUvHqiFLiAPcuPFL5
JlNt0AsGIEegUE7yo30J5ZhwCXwxWz1sELplIJHVYmLAG20jfJTg3CrRJSb7gL6U
ha5+fBUi7SyyWq/Fbr89JnHS15waMUM3GCKcsaQVHuF7ljZggEVxieXD0PoJGCw9
JzZtcAR2+vATWatsvI3G7/sWl0YtObfjYH6fB3bzPAqle6PRHyfAhfTnBIuod99M
m2YKIwc0jTTDwIUTqixoiNQ6JfidChm2H9qvqGfp13AJ1TlHOIIVhj5Aev/cJNGU
LoYlIoxIxMbpKe0903vf5CbJN4hscLLc9xiC8qF4mGiDZTyvK46UEutAcmEs+gSG
0xXTVl06CmfXuNAXruyDuTP3xIYBPFb9XvyyOO0Pq0bpY+8DlNaWN8PS0tBXd1XE
6r1Rke6mlkEZ/zr6YfkcRnKV+UNcJ85AoRJr3fVl304Q4wFDv+OnYN+b2grkVPVP
9/Kqn6Ot14Am0lohCsnDPly6tySaHWOMU6mOC7/0bEAINiinGfGOPkAf5fqST/58
In51kJWCh3TjPftKszbYq1xAiDBIwqi5BFd2kKIhgvHU/CcLurMM+Sq4AQ1hZRTG
Z3aRlqhEuLqzOGMhen94YRVNi0Egxo6c5/V3Tk0v7f8Mjw4t3zAhh7YAFZXSHjg8
sx0WdiMCXb2lpg+7N0c+T0Q/XxlF+zpcIsltlwMgfDIhJ7dHAHp7uJ1Tc1/zovGV
TSGZ9VFv0eviNhD/KQJp9TiMjQWi8SnsHdS7sT05yUPDnFue9f9GCqbWlpb5kDtw
Hxhl5l0iW8IaYAldo0+3m8bcOWLHwbPgOpOh2wceKnoTx+zd4TedyFBtnFIofzsj
Uh2QgVgfAfyI2t58pGUZDkddYK6EQjU1lxtdnP0nCMDk4b1VnFLtSr4cueqcNVT+
psKeoSM5Tx15j+4iqAF63GvId7m847pVCeuK5QnZs8SsYuSaYFK/3UcU+cr2a3t8
NUjS1aZH9p5kaz7MwJmg9bmJC7W5FRvPFzRzz1JVrHN8sqXF4ueRecxBKjX7Bkev
yNEPX7SzB+LAt3SJq12uyXFvBWjGaUUzWpBueAViszyiWFmFk5T+DkbgJjpG1lSk
oM5DFGjRPJ9MfE84c/Y4s097jlQsaojPVhK16aznB0TFWIwEBEPbTHcqJD/yEE0B
+gr7oiBOyfzawnVVvl38GJRrSvj7i1l+axXOGyM4G1YFUmS7zkNJJX73cLiA9kZt
owzYs6goVGZi4c6L7pni2n8tfHsCTQoI09HUMGsozsAov8D+dIraOhl0azRrlzlw
UuniAj/xY+Jw7IPCZp/bfZn7X0YaqVKBOCOu66SKJOwvRatYZCOmNnDIC8tJj99u
XRqglELzTevoHJo5zR0TOUkRsZBv4wmS70u6wwBy+c1KCCyQjgd/7/TXLoPek0Z8
zaaJDoeF51Fa2cfPlynXag7kBl52yRQ8YrTfDAdNi0Fm+RwsT6TEFDJif7X2keEq
sfAUegX2zTYWI0zQSaD4Eti0c8O82qnFaJFxJdzv1HiwkJDpo99ozRgvgGd28n5T
33fU1g8dEjsIhyLzXTQjGO9+onI/CYZrbBaPwRbDiVbNVIFK2/QGIuow4/2xXAcf
JxWmwt7qqNq2icpiIL/Y35NLZQLsU8I1Sw/R199TgBALaHR4+Fzi61tNEIqRlC6F
d8QEKC9jMp06HuHiJzH4X80k1Et6k8VjZ79obRYZ5iaw/hnZ0ZtaCc3ZPbbwSX4w
216KiPcWbot6+ADeSh21rHgDcYqWzNGnIGtUCG4ENV1JYtupP7GLzT57vJmyIzpX
TDWKV/MWxKmqIXddJoc3wmEPVUNe7+r65AzAF54wDJ2UMQQ58p14QwntkpaW+SiW
j7vJ8UFGuMNqxZGkqAeXG+mXOPPv5dmi6igmj1cEjv6iEJtL28Qzx52sK2GF/ot9
YexwFr7zd0OlbJpUjKdp6efnx9pUK4M2sqUl5es4KOzz8dzJ4+tkwot0HY387OCc
oEjC3Z48oHj7maueprvIFvsk0uIjSVq2YTUtCTSNEzfQSIGHoH+E6bSuMFfK9BmY
mTOlNTGGt696h80NxOU/TfbLqDAToJNpb0vjpzHudQQzXP1pYDjI7MmprGrF9S57
dXgUlrXW4Bbc7ZGJ0r3z/60EYiayZIaFi9VOYSyaXFoh9ky72fG7B9ptIP7rfNO/
8HOEPGD6igkpyKbWqdOSSYp7poc1o2MxrZCf9PmLkHTmjJU7Pxy0nUZXUGBJ277k
AoRCIR74GeKeZ7cFCb15RUdObJ2+S2N0cH38GjlgJZJO7b+Yv6dsMVb7igc89jEe
Ulhww/NdSuAgkoYGeH2S3cBx/H9B3IUaOx/X6sD5AS5UK5xfqLZMQu+t53WkOVl6
tTgQ5ob/k04Si4wiKnjkYerXzvFN4jZKUKmwVdJXuOHSib6/ZCMvVt8iRIH5qZwe
EEkJTDvArer2HKY81zagVvjdQZUVXeneMXGtfqksXMKwaVmhm64/ZwEKdQ6ugM51
49omJ+gbAPmNb6LmFUuCgc5ZLsIb7+NIeOxx8HJiPsbdxb2DRu76qCBH7shEwAtO
PAbQbZi7g7gQENHIrx/lO0Dyq2VZpgO1JGNlhk5MR8w7fkX103gjBZW3IxAhu6Bb
qncnCeEm8JqXCMy0hwbojHj/bh8IPlCrMPD2FhiLT+agIq8Ee+pC7NswxWfD+g6p
zdy/UXbsyCrhWrjW5KQopW+cY4rZ4MhqQ+gKjdJhCU1ZihCQmm1bbYLGC3rk4oAu
YjKSp58pr+ukFzVX8S9KSaGpmDQbJPh5QL5C7tCxFpFB4ibnGotMGomQXo9w9+MV
Td9FfuXTqf3ebA0wcEv3NqdzUqsTedxpzr8/3XQRDuThwKNM8R7zS0lHw4mOOPhd
C96uoIH2ANAfUCXTrgEwFGCDcOYaDQd1cYQI5/kC1w74N5UZOcWHW1Wl7zUVJdGl
rc44RA2NjnWp0NrmNRz3ag+qTUiQCQKgtxODhlz2I8/+uViosWkAnr+qMuTMq8RM
tdF47GA+Plf255cCorDRdYHcnfl8eaWMdvaB4NPX7ETVFiiBGYxH/QGWo9KKQkk5
4RMlzxU3JaPu9AaTBvey/YAYWSmRYtNNwTtCUWKOzcnfj9C79MLfVbDQhWhK6INH
6edOu2fGQjhxnka+3JyacrGEiMnSNjzvZ27hql0ihKxaohodAjXwp0wG8kMT5DeO
KwimajDIRgRbhVAQ1qNzYGbeuNPK4QQ5Bp/OBFtfzPK3z2aK6dj6zU/IeZhDJJiD
ruLc25Jlrbtt+vuh4zaFR/N8CizkCNrPpKtxdzsBpwO5w0T/1C+3DD2Fw8lj2Vxl
NUUzRuRKSuh/P0SmETkmjAeHScqFOEDMp1FR4akAvMTM81FMqHmH/KjXHdyIfY2P
W5ZOlMrh5g3OXKRmP1AyX2e7a7n6M/mEeKtT2RTOeBahl52H6v/xUFyxt0/7pUqO
thN6hP7NENtfpC4tYSJDU4buttN7al2OIcsXOb5k1Bmj0fgb4FiYYhC+mANNDlAb
64alydAckmzOfH/lu2E4ANhKLP1CclenuGiSKyX8g10KO+fYL9jicKdFYuoaDNnl
7DaUAFI+1oxSrC/XZl7QrGwKrmapuW5vKoPT0fc12p3hBDmw3Q4xMjtqnnlKs0Mz
jNMKbMerZBq6Uz1qCRbtoOqWyY2cdb65oR1/c2JRdDiHWizG/Vr2gZ7MKGhFtn3c
yMQeQbnsm46DOE6Zz9oJIGUCH42PgZxZv6U4AnRgqDQrdduG4i4r+ZQta/oOriRm
Pz5/XX08GHojySrawyLD6tDF5zGfa8JERxak4K8vRmGYEoELV4tJN7RN3U50L/7k
B+aUuCC7/2rYRvq3XI3V+s/RyerbMfG068MKvtbZVzjUAUxTePPVd715gVUknbIs
UjcDPayQyPfXN9TvbN2A3nRlKZMe3FNvLmRgyC1PDUfGdPnuEH8jTaq74W5+fjtj
gXvg7/lBRsMDRgyZ92NacQPF6jeAtf9FUdmM2kwIth/l7v36X8MQ9iMYNSh4gaC9
HT/yqV4S9Iz6Waz2GdpoR+iZEbRkXRfpSQz1D/o8VeoeEnT6X4rhsos2kAE9fkx2
IIOv+SApg94yajfmDWJuV/2hqZSybVArEDN8sZ6DjEf3EDFWLVqquruJpKPH7zyO
PO4ZUwwfgCenp7LqV75/6dib5J+buFroY5B+lmadDkQJf0U5Vo52/Wv5jJEgoA+T
p1zSLwldtKZ8Q6sPRyS7Gr0rIe3c7fOxIaH5GAVOEocPafcOzX076XIV6Ay0ZZIL
d7Lt/NSJoIdfI0VlQEGbOBz8HkQ6DRBN6Or/6VWXpLh5/k67NQV1c5rxhDUclLBA
15jkw+6KTDKJ+bJekExQYkfCmsF+jdJ0DxsLDSuZgo8a59jKEvAWYfm/3vEsBaSR
XnYvvOifwQrScXCtxGUUg8H+UOVHJuShzfQBrt9+5REzvDYJ/BZexu+0RWP7/jEf
IgP4vjI5hcCD4j9MFdV5Dtkp9lHdArdHN+FPtsNjrEFK/9zmuSIHLu4VxSfQPeyQ
uN+c7wH772yB0siO795qveVKBQb7lYDETSU+sn4qIim03SID9fjCQyrhpeIHmRO0
F2eMLWH1b0RRLy0xEX1qDY7bTMvMyfzUjWG5LPV2V6YP0XlG9WOpPVTiJ7qb+Jm2
c8MCtpI695+F7EtJmjY8OXlxn7P4VNGH4iU3R1PeRGQfmZoonVOgk0jorBmQvifw
3s13/Uz0O8FeJnJBBHBtEXmHgbtczXSaQ7PCnEQ6YGuZl95iuEa0BtgrbDelIIQX
7hmrt+v27kbEDHKu5gjetAcrQAFsGq8cj+lB7uzIgzbgbW/gpWkBJbAOS/BR49cW
DYaLnQvJwjrHXxSY5iU34q20ZkSXcOSzbvK0N0xhrnqZDEpDBI+MCjON+yV3coJY
YPWbaruhDBdHY7A7FeL0Su7rWt/80lLQKhlOIHVQh2fqLixN8uIhL4EtW/Om+4cp
7Ql4BmSzHOb3aQmd4V9kBawaqzUSk3+sBB6xV1bYP4P/lB/+QGwxZLU30imFaptg
/LCpyB5JV0lz4Ym5EOOLpXvVA1QHChqYsEovhkrA7uXXlZSVdK3ukq3VJNIKfPNw
RL3+xg/D3fs3hpKvJi4dfhJC1HkLNMzuZx9Kayd/D+K4Zuss0AqiEit3+piHrmHp
Xk31bbIwF8fDeVWGlCNwH8gOlVB15Rlh6TlmxszqOmo8Xgo5SJDGJ3HH6Cb8k20i
de1WCPMus6SyHkPXG+yeWwwpifKY6BV0of9TCXfuycHJe1Wwbl6HgtxFI08M4XA7
IIy3D+Vd3sGrg/Ls4YSN2Rkf/1de1dWy7MR9Ecxphxh69vUEdel7nmWBOCqgp73t
/vVxehW7ID675rzVzbTCPvBLXeMEgJKmSaMFObIuMigtyEBVxnUJLQMPDzuqZBLq
u9alyXyktm8/0IgV2UYZzedG/rnUisUFTMDsggVZruvKAdXBbP+JR8Dn0VbIGl48
u6kViJlhJXk5viYL1daE4ccPoT56ROIAzxuT9wD/UXiRz/DJDuAjPPCCiowrc//b
9ny9aaO29avwkHMgL/r3mrnTFzhFp9Dw8gYt/oW42PM5fBN4AjLvE04at6tmDod9
Fsnt8KON7iSoyDiMWTLrdM0XdzyMRUWBeZSHoYBWwJ2NzFEBbKWjDIaX2S/vn7Ge
644SbmrGkNeJdfGRYlMHlUUVwccWQ7hv6gp1p8qDDwC5/h3jMgU4q9cZKt3EhxTW
8RbIEyfCE2ZR0ORaO1Ojev9WzhkUKOVnzgoF6bqTbjiOgRINs6Fg9Vjlim/0hWDb
qEqwTg0/90cZ8Y1XUPwfK3K1JFft7psQ/GVZWy36qDrMYT1hMhHuKTrVHIBLvAHV
yHc+NNUjPByIx0ZmV8tlwZ1/IuCpZILUIE2JltkfYVP7dO9m2SvASsdidr3aOsiE
B3spef88Ez4tBVdeT0ydv8zc+3jA1DwKckcEXR9T/OFxnjOq6Mma+wCxi8wu3o/c
hZ9e6L4LIfnTGLN7yYlRsvsPjoiC9AXhIv+b7qp4JpF7x0C2d/Lp767asFEMLMjH
JalbFjOOrPifinTRqqEPVP57BZP+YEjbXjOGi97oLC4oJLq5scK71V09aAvd68zd
RWTouMamqghvam2IAsdy6jmErBYBVp4LeJDwsH5ccfASPmEq4I0xTiYCEx+VD9OX
9cqRlvnWJJqShcU86B/8dlBbNxsChtZ1V6G6uViIufEpoZXEYndqy/bUBFa4H2pG
IY3EMj+d7nRTHXIJ99/ItKgEPy8UUH1oFzHQNuwo1+1FU/smA7tg9iRl79DceZT6
h87K4UfIoHuTSLHzR/a1sGU+3E3d6YlK0JlEiDh/92Ir64rYcHH2cooiYnQaa4Ee
beggFE3t1FmKka0AvMOZgpJxoJoR5wK+4MyZwGkOnL4z1+/IcY6G5NmOPM0Nxecf
7ggseFAhVzqCzJ9nMIcDCzNJ73KNIJ3TOzIb1aAtM+WXz4vtvb5s9RL8a+YkDd+F
O4olYyGCe01ahA7jbJZkd5/7HKGVbE4elIIZA/mw6kFKDjcA3KNY13Rh/AuEtUY0
4wroLW+pZFqusjHIdtie7B4/DqUR9UheG6NanZnNftQkIOekbFrWAKXpWVzoxQAd
hQz7OzIwsfxa6KgEV4QbiS+Xpd0eHvvsuvZYgkxOpAwBjFp1jI8+Xb2FPgw7r2Jy
jufZ9UHsh4WIS1/EajUlKwzw0tMXx8DB4bmVrTDXgmug3euLJK9CdfgGvgsbTplX
bl4aDPuUi7APlof/jLh+vsSfJ3nBBoK2R3s709eewIAzOM6kLPCcWVJr37/rNf4x
UNK0HIiulsofahwGl2p/gQnfZ5KZAONuizsgVDfOHHIcLNc7zn5X6vXbYexjlb7Y
e4fEtguwcw8Scgm+uqdJaSUwGlgfNPeViws+I6MOwxExR+14b0hhSrMqk4E4EDuu
dec+fdYIt6u6N8LgZiktferfJbMhOzAPp0hM0ddr5DP1CkoUlwVWy6r4syOk0/CB
ax8yrFAw1H7sZfhgeaZsvZLTE1NqM00w1C2IsPNzmOyfVwsSWoBC7PXlmlwRVgno
TFBbIesUowOwoy/BpSSM+KVcFQDA7rHRs88DGiEan9FaFuhUbmJ8VvAkuTQxjHeP
Ksg5wm5CB31gYOeb4Xd199uKOrTaJ+Q6A/ljOi2b3ZePzXjewpLo4YCZ1y5iiOE5
FIHJArIAyy068UdhobxLLi7dV5KS0KL9btYbWcQJd0GNJdpZnUQ1cYYimgpFpITO
0VvDZUXVFnaJ3W6rFqQsaQCIRtat8hbu9I2WmdR7NBbyg/xYTGbBa61ItEBVy6a9
VvKWuFQpMEX4oOZgSX3VELcFeScez1VPxUQxRh5TFDD7ZxWRiCk894Nfsmoy92cl
iki2iWB07+MaeJDgsTdUlctdwCFBqrCwwU9MVr77VlVTMHwGjrPaMmrEW/YOo1on
2uUWQfEYk0TAfk3HKieTVQLxcdxhYP9vvTswLl6YNqvZaiTCB6SEk4I2Xh8AJ0HM
p5PPxd0sclEVEaYwL+sKBPUBIHUM370VAemFY1epp9MNUJR0ywDS9EnHmLdST8BP
8IHdRPHLVH/QZEtqDVZs3/6rQdmBPEj3abB4mMB2qIuUPhWrPcuKw8yaRlPaazOc
As1dUWcroxwGwnruGSY2jZI2d8n+LzjOBzNIR4yC1KmE8CmXno8V6N7P/sZKdVWg
tGLPQSTQ9WEho4frc04GCOL/7h1/H2/rxGycC/cRF9bOdK0Trb/PuNyYpDay5TWY
/cXpkgccFcBEukFlEoCUarXB2aJ2dThUmCk5Gn9ptdaZ1xxHDmZgVlPYOrjY4IOS
2Dy9EKKmP94J3RN3JJSxSCCjEWXWRcPsGesyag3in/XJUc89xCVmyqsahmqCQrmL
5yuFvBJs2k4pCAnwV1LQ561rPphdyojHzbKlDx3MdMN8TjpOLCYWGHV+pBgky+WR
eX57P4WzCOxQWBem+QGWMZKsnzko8MGGS1vxxAneZ+kJqv7AIhqADzHT2NyCQx+S
BiYCcZorrHHxwVsjYd3iHE37nlgTL9unsuCuCFKEl82lOfPGchpKxUH2DV9QGVXs
5RhCUUvr0rRCPnzCjIRWmCxQS1+DHiz+e6c0xxYERJtwflv0ExYjM1C0mr35yLez
jTI2UT20ECZPsdwy0mwIbUnB2CX23mB9fBZ4d9SmAPJvH1XDwMHLSRse/c0vEAqT
aIDDw4g/SoBk0NUjHlP7lCt0uA2gvQMdVJqM7WNMFnVTpn9bbaPlEeYZTe1A2Gtt
6dqhaX8uj+WywlJjm0fSDWS+OpgQov1H7gnVwvQ7UZKK2lRe7TnLiuqV+AjBkq/w
625u/10FvmuuRAaVIc2KRbrYRGbRGq4STtciPGdCyF72YTf2FSwPcJRgrb3ymy8d
P3GiJhKW1edgJRH44dc3rRTrQ+lbIKY0xWzpRKGXslB8X3FYlbwd960wMiM+Uglb
1YfiWxA7vq9P++kXJqRgvVozTp8HUjVylJUdie7lI3NDrr1LkYg9hzw80U2/VhCS
i9yU9erqWJ0L2HZbDORGlYdNOg3ox/84dl5AaamUQT+/C0eBBu7BDnChm4U844k3
djo/ZSQgaBBMgT//OR8rQpZrVmjnPTlAwoBwpdZfGueD6Xaa1mNQ8zuYDuHDusid
XUIWmZ76FRj8BV17veSiyKfQhocu1XB3pzLvZpyQG/fibWdcV5XS7ijhFJU0Kds8
EYpBHYdCpJ1G44f+VeIbjOc3phYU1qVBFIBWZMMnufT2DpIovnlwTgjiz0pOOZ6l
NU/4l05RsGoOdWa/ozzLIqveYykoH4mpNxSjTFxNM+mzOlUz/1dg2Ix/N5XaTUH2
9yMGHG6KzBWctx52FR9sBLVWt7fIvC+ui4+EBdd1yx9B0h7yg+pQKFMMo4MOeqF5
DXF0cxvH7l6fEKcwDyRzg7jse0ga5nO3uw1gJieT31ATAOoy/M/tN5EPym0kCubD
rnbzwOVg/YA1jZWwW6dHHGcMLEZHv+SfkYZjyVYaLUPWeCkPlErGe065vpSDy2+5
ACpZXUZkdVLcyaBjM0R8Y3ocnLxZ/3aCi+dO2VjKEZoy7YELnMNfR4ZOZUVUas2q
DpbEipk5iZQ0JpH6ghDBFRB8SG4f8r3pN0TFlvNrHBtSv5abQAHkr2ryBb4ZqyXB
YuFUwal4paghytnQ8i/qWgX8dxEbXk6zKB3gyEIhaRj02dUliuDJKUMvgoIe5vl9
HcCVjG8azuTR5y9zTY3OJThKqGTvng/DM/I9R2MRJDC0RaBZyrscV3099D+LsrOj
PHULHyhqPyrcRhitKIj3dnzrXJT/Q4hxiU3nd/EHWPE2dgHRBRpKU5AZYnG7Dpdo
6XrLpYW/iySEeD1oVDAMmT7khP8wEHUi7Y1CNXlGBE2nI+eEKq0yzvXZe7XU77F8
ZLqA8tEmLCrIwUqDM7xozKUcPk+QlmOfzlDw8VFCbRe1aGYVt+ca5an3KTLWEtOw
oLMopAQgY0hZkKlTMAg1Ve9tg5YHv9gdQ/iEXmOluiTSuIvc0gSj2gCIwPsTUiqj
+aRCvjK3HhaW4l2nxwZj0dR5nCj4eVE5NgQLCvuUzl2V+5Qgdks30l9blxW7jRiZ
LlYxbIqhmOV6yGEtcsmCr04c/Q9+leH4OKyePHts5aKUnFb4LGahW4JRV8pnHFe/
wJWNhzLa/v+oS+pPkrc2lwxX3aCcz3NzlLTuAlCOF/k1wCJUx4IonH8rvdKsmV4C
MHU/2+aFmMgcofZDE3bpFDHz8cHBlOJ4j7uzg86jEqbufdNI338zaYJ1hFx+RHu6
ObR2zEN3giZn1XtRp6UWo9zjHt7StoHS71U4kaG2Rq6UzvRafDteH4G1A8vSooT7
PYoOFifedd6IXOmNZWVN4bNhn+3i75EiuKsq9wsit7VB//TFRAETzQloe3YpV/0T
96CdUg+a+sTmoaUgi/L58WvjV0D4hblpwk349U8cbgpLDLts57lAui71yrWgzbJ1
CTBcqui9rpvo3AKYeP3QoQD7NiNbFA+W/U+ShcT24LeRVquCYZG/rLgPIeA6/92v
79kNXjZF3tFY3RCj+NUpLT0IVEX2F/1VadvOFQawRDj/3yvkEXIyQKMVIDJrvOlB
rlAmz0zY8pMaBYZEfrw+3cR0T4cf/T+1LWwFEM6bB8z4Xy3cZIRqJhg/xvrQ8Zeu
2tDrq/AX6XbH20hnUJH7sLdnToumnSHTYmd5cVYQpHW539DVTnAJUG/xwdwavj70
0eTMuwx9ZZIEZnckdbZ2ie+Gp2nl6B0apJLLiFzD5ccUjNHanMIs2403qo7c9M/E
WGkfSRIpmh9+82alRgmAEvI3A7B/VHELSkIcZ+mYChV3kdxURvig2gHDQUw661L1
ixMfoGzxxwRs9xOmXcK7Qj42fNzX7L/2b3EuWsIJ94Ic425Zd/1fFcERgb8gZRGs
3Ms6B4pq8tG0AwZ+VPgv/F4qmDjgK0MSTrNM2i9oK49aOxoExf18rgcNyRJyrruA
DU7tgc9/0r8ab4OS4F7lmTPxhDeTm43v/g5aN9chKNo0CimPkLedvQhoJKj9rRm/
cEBrqiEfPfi64P/k7nfD8fyp2binfhcQw/mM/V6dLNWhZn+/kJctkMFxH6scS8JU
BXWSZSwrguqKhEYxUIgyaar7DOyYf27e8dBNI4QNYQyBeHqpk9wmd4qtkt5WejNF
iLB2KBSG0Rw8z1E5BYybkDR7PaDu9zaABp2vs/y46ZUIdT7CXl+NYK+MUPixykAA
llePXEWC3eejdXvi39cJfp0JUBjcLll94qpKeNTHVFuhRmf7X80PcEuS1oF675Rq
FWQFor5HoQ2oezRbSggoR8ViHVRih8YySYp6PrMX2/DGt9APoQZGzAow7CgJN/vY
aabJ0ViFPDB6JF27ODy3liUuBol4g9zahoJtb5w9Is8Z77XYJpgJF0dSvfBQ/XH+
ySLPgYd2kB8TL2fcg9TNmUkpybwtNJHd0nXd4vpnRbljO6CQK1Q/Vax7EleBz8Vv
f9Crl1+l5T9In1tPzhdlRYba6s6KTxk+Utgvwsu31YfMoaiUxn2nQOhL2AKE8MgX
1j63a+WS+PWFnIdFRZ6YHh8V2ciPFScwp/WxKCVKLbqbnRTWNBphOko0v2SQeFVg
yAEHnpjJSWmTrkWf7Mkzq8H/nN/7eRa3VOzWzKCrreveadgTpe30mKdFl8Ic4nzW
022pj5iEgXzZ7Tm/Rn99d2H3sSC5IFPXqacHsiB5ag/lMfDiPOXMpHkbLi9xSf62
Hy5kbjobx40HXyVYoFdWRNy1ZumzbuoGeLJO20N0FjyGtQ3ej/vBSvtjBliJKbJk
veBRiXUYySbo5mfggg3YXIgd2hcDGOb38Wvrt5uszJBks7aCXs7ZA7TfXFxxye3e
TTwBPKxA4cJrwdx6G9fWseImFngGGKidmBKAlY1KAnQHipFOiiMc/iUo+suQF+mi
rcrprsArzuzP4qvXq0ny6QhWmHy9ZF5DqiKDeA+nxTOFc12vTh9iZNfjwiG3dMpm
b4n9HbjM59lhImMkcQLTWpkK5CBAusAg+sX3u6NT5xwtwKt79+sT25MFQk/VJ3l/
FtRQCR1TNZ3q5129XVL1T7cuY9kH16pDDF7FapWavtXrNvrEL3TW7IfdBypTlVI1
Ly7hx7PYJQdlt0PU9tXY/EEDJesZeSkp1e2GcCgDA9Lqws8ZYP9YhII4rHX15tX4
N4HKxAHJZv5nDiWlfUCLrnprVz3uHkOd3mncIG+0VPuucU3PwHV7NUOi4jvyR3L8
+vKvFCsRo5SJtWGpcD3Uw6Y79TC2fbrnJ0obDbhvCGZF0ZKeisw9Ut9YPnd1+9PI
DwrkB/jWv7hZCK7wSgL4l8qmH7BFv0ckdQt9nSr0M/LZhk7lyWhKMeNhYPpbn42Y
uHA48tgrpm+g30QbbSUzryarVQ+xrIkJJxfWKahge6QBTliuddeM0diriwKRQUxQ
uM/OpNEjAbmJ7G8F3siv6CLwa0voHufPVWMOzN2ZllOAYHWACqp+NiWzJo4ECpgp
Z0e76LGW8AzeWK5964BLIoN9R/IWV2cuJ1TftLCf4Za40WBosHREammMKzTOW2G+
462mzsZB6mN0iWjqB6V6Nfr9SoEwInu0F7Tb7jPWrZMGDRBYVJrdGrqlctIUiGJt
G+O3yzpZLjuhqLNsZoF1ZcvdF3iOBH3RQBarTcyjSbvOkA9gzQXt+P2GP2224ddj
hDfHbCEEJE31s5LLoSiauCszUL7Ks744x2OnyKO98ub8bj1YAfFIACsckSzOq9dz
KEDdLCmByPCZj1sWKsQAasLTvbLenJRynFZnL/631T8nEmcRaeSn0jSMFKyZEq3b
TS4fLyTcMiPA5qngd36i2pxkQnW9C7yT6eQljqkPA4CnT8K7vELnnNvIocEXLj+3
X/Et29lnP/R5DXDty4+JXQ6lVZqJz07dThFQikOw+MGEHwtmJ5OOUcudxJ3PCYbh
qSzW5Jhb3mW+qI8STBHQvHZ9Tr66g+A3/EDQB/Ntk5lEr194eb4d30CqAdjSs/Ls
/EOqvB263OFhFc+9A3hlrww8sEFB2rwUoTtJMhaD1K4PwzS6jt+DrVTzfyD8SUXJ
Drv9ZebgXyxnOqRvEvLHhWdf70UJQ/jat2s0M+QAlfODL1rIDGWcO13hqXovZbUG
cvfAPathNM9lMz5FHFLibp+eyQVNrnGgWA1+nC5l5A3k6GZHxlprnQ4ELtmQuser
XvZSvhxr7KL5gmHW0oI50IpqdgnIMKaZn2cz479sUTtfVAYz2RFAmZUVwrRuz70t
loEhkUgmpbJ77Ztqt9R4fbNsLrbOuCbbs7UGUfc+ZZlK+LNjoRlCHSUm7kZQIgXG
b3h3dKmB0gx0OLrdneX2MBpYX+8dNaTFOkWDeEC/E4MAEpktfzghoT5xXC9BfwjA
2UZPj4tw0bfEyUzzSmoXSJggxgb+I3kYoXWV79oVFYPlPufsCH9DF2kHTifrxb9B
6x2u2u1ks8RTXmsQxmOQw5ynQOVkT5wMQWw3GTjOJGk7azIlKNlHlf+UKCFFfTUs
FrUiCCtVMxxzqYq5YhGOpHmtxGH4Dgoydn+pjVxOlszsWHvudm7G0RjTXD6Uc1ET
1acHURgcsERFtCI+iQxB9D1HeLMEfZl6wXgdTs0hseAe3cvHzwyrCVZOYE+vOMBS
YLnZ/cvlXUfDQTMPFmitLd9vc7y6BT//zkLbyhzITuLsSph690P2SmdPOSikq8ip
mes2yDZdDllf0PlZTtvVHBDP97v3dPmCoBGSgVhuK64eGC+PLvXJ627h/0oGxmEv
RYaFKdm8hAsmhIWTkTXSIrDiHaVuu6Iu9FbaXAhSR2rVkZrEs3R/LUuzDTssxFrT
YhB0+wDzvfjZG9CmJ4+WF/SIHHzbiZv7ZzNTCGFAD65WjWe0GknUJegjopzQag3G
7jcnvgqw7MyGrNCukwX7MMe2Sk+eZUNXD6ILM+F4VA0y2wIkGheaxTjqk9736IgZ
yxKmDdPiC0tkoY11Q/YlpbtEVdAEl2XWn34GvpZTkUe8D8ZDhxiCsDNSeC7HEa+M
itq1sjIpEz/ucLtZJrcLszW46kW+Q/yQR+q2Y4WV0WuG000vWeZdkcV1SY/Fax+c
y3TNgZ53x5G+0nGDhvfXCgvExhXLuGDOu1EkNUqatZK8ID8Wkoh+GE0SOfJPvlJP
O3k64YXOn7lNc0lQ8Y38qpL4ceT1oCcTHxBRumbxydWpHo35j1cCEB9S3E3HSfw4
yP4sFYImJIurOq9HzGD1dCaliCEEHzRvjN5V1RQ5Bie498mgK6T6BWzOVc7Tefur
RzxH6Vfg/HgQBk8uYIc8USdAp0IWh1KvVACWe0AElE2/kQQ3MrlBFMSBp8IqoCWO
ksiuKKcpMMLO9ZKJFk5Bl7vCvE4KAeK4l9y8/V8h0lIXwO0+NyBmEkddIaGVlokO
UN0nRA0JuCWW1yewvZXKy0gl8EsGO8pSC0lYs2sY8p/hDINgJeLUaXjLnhS7NL8Z
4Su3HrfLhOArKOvlzLBIo78yRwbfiHQfH0Qbp8aTQautP20rbgcEbfQjCJNNdR+Y
TfPCvPjG/F8bZ1GqZT1sd6EBYB9JgfnzSvpkZb8O0AXL+ObXGxExiTdc42AfWPj8
ArrhMHn+Eiw7QJKO2t8O0kfDniWnxx5sec9Om+rSywaX3U0fhhQOUC/BFU5cwmYn
CRrrVdph0xagAdaolLDeVkHzzmxAIOQVsW4MWcUGO6Ov9gRODoHygkiVH8RbHEta
zakeE4u8avhUM/VeiuZO5MDuIMas3L4qjPFz5OF3zkz/XHH21cpYzH8Drc1uYONQ
lRK4DpV4zUYIbhP3hWvmHPmgRmqK4d7uJI4W4rIs2mlUuFGUNkPNkRpFY6TpRUOT
EsIJ090FtbuRT95KcLXE2sOZoXcTuX1brU82zqU+dXJ1gq0kjzyISQsUPzx6XOxz
gt06ul2m2IiS2/d/+94UlDZY0nmZnJCJss36je1mjxlnukCaARTRzCFwnR+D7JEp
LisHNvggzh4R82lj/O6H+zs3otYrz7SnR9A8t4FT0/2hlqSOLEDrBGCTd2619M1y
9jwNhveygmOLFgAcm5js7N5/VS0mL+VSPCbOIyClJAVMPq/zsG46crES+Xdw/TIY
vi01yOLRN5Eok3HfMemQJWE/QILOWrfOjzcajILKItZc+Z+sNYkzdDsoipOs1/U3
Nowb/iaAs0JUlbcy9RQsTH1jc0CykzldtcgSSMf1BEk3aXdWGRY+8UDDViZZarwK
uiMfFE5USNjAfISJ5rNOq0oLyTqZRhmZYE+QmddVSrM0Q63QqyNq9KxFgK5fRJVx
GWhogQSbN7SX/d6mX9PDuf+wrqRheI5gNOWwaET/iVWZt4qhBNNIuCHUps574uQ7
h5StBj74G/0d1obWUD/4smkp/b+YLbyl7xPHpyLIpx+lwIn3iEIfaSnoANlrz46O
eQur/A1mGYm/hD/HbZZNlZcww2RPie7zf59cg/FdnEb49rSFCNARuESTsdOPWRLh
lgMQIJ6pFCyeHM7AiwbGh743z0yW10TebcKJvrHY4QITRP96inQZenb9cXRPrnwM
LQKi3bOJsqRW5jlPg0jasgNTq2GzKFUlkeF+RCI371wx4D/qh7iPuQEHSgxXhAWj
YKqlqqTgvp5ddNaRqk7/7LUQ4ripuzT0AxDX3649NrzmxaCQ6aGRSzyqezCKWMIz
auddSrXm+iuNoGFUnPAHZ3pnqJFffEK6ZbT4jb1I3pM97ZveH/WJpteP2godlcYx
8UGsGj2pEnF8xF28cE10/WuKFSMnImXXWdn6xgCzPcBybuDb86PO8cIJcopu74Zw
7JuETGaPYkyCYcAUTdtEW5bULoSa1qX/OfocMGEC4oBX8Txx1zfHfqWqJbCP7guc
AzsvBwDIAeNd+NoKDtnkH4lYQhYxdfiKrgtfjVFWKvFP9SOm2CRbynQzvVC87XLa
xI4bMuCebiGEmhh2OLL4Pq7H7l+uQscihVdZIedpSnHRtbcEqIbe7Ewt8BtHLrKm
CjUeAz1avSSsLoTx4TJhaCmIEVghvYY0Kp03og7XCFgPCvktnFIucJz1jW+YGJ/p
3RjRJ04sh7XM/dutGz21rkZEttRopJcpwk+jp631cIg9ad7Yb4lYrnsAbLE6gAd0
wBAsrfaYoC3PJhJXqkAVYLNbjwbcr0CJ/wKla+cjK9g/fVbpPWElae0xlg8gZ1XG
7FEDDgns3W4vkf1+SJBkbQrNuqBc7u/K+JsdZVYUi3MEG2rypbkWHcdkmnIDTwnA
4jzbTFq6nlrPt0d6JEBzlD+km6l/ms4j9DRGbcItROdQWiMfRXXg1E3Uj8Gbsp7F
c9vMP+HfPBxKMXCAkoE0+sBE1BBmLnqhHTYH3CnOcJqK4bkbxjnK8cGM816DUIqH
1gt2WVYzub9OfXWqi0p/uLoeMz1fZCStvn01/MARkJVXB6QVEypmclGUJhJwqWo3
NLY0HIdZYRLGqtzV9KEAMLw87zEcUs5L7fx0kroiauCZMo38LW2Z0HBZCG0i6UJV
mLvtbWbPP+E3qlPP9GNJ9iMHdpUvWFGCJpuKCK7CXEQ0mF9KeiISLgkZGaiZkRw3
bPqmeFQjR0WC7E44F9t/gcTcyw5mymcYgc5JWkR1NoPzOtijbki8RjJXJox+tUTN
izsreN8GQ11UBVCI8hUBp7eDbS2TwUtNXOtxBY7TACn70hngavKxSrsGcJ1Ofxer
Op6QQqVkvmxj661yuWdAtfIoWVMWy1rHQUFkNwRsZnaIhGSpbYMoRAwYTS/DpAA5
yN7UNi0Q/lKqZrZcQtjSW7OofbSv4gwk73xzKUeYZlcWbMkrEoaSk63tXkQdyra/
RqnH8A25etTSrMEQJhiqpxLjXz4GDc9WChWPdvTzMw0XyNQiFN1t5laeYfm2fCue
b+bqdFHBKrZhAgAJNqBY7ZCsBDkwGiYfD77sPC0i9SM4Wjm14Sb1MOermtPkvWWt
u/lQoQYTiVSHxYtMzH1H3jR5V7cR7Ewv/58Ssw16TzDaE94eNO4hAWP/yyr1T4TF
LNeFXjwbTORBQpF88bktoPrLe5kxFyxaVqRQCgnQK0TppbD45wobA2D3AAdoddRp
/1BUbfI5KU6sdewWKQ/t5EI8Dz3KUOZIog+IYFCNwYbYyo4JuVblBhImIPheyGgI
IfybL0OlcecpDLiNm27v/0NdlZHALmBFZtJE3huX35pJLI+xaXLuVBxZDamzybPJ
AjzaZeygYdi32kjh2a2Ng8vxKCv5xjvjsH7hwS02YrALAx2xMbnHLZm9PYSgSAVK
O4l5Lm58KcO/nXjt52u4LtTXF74ouA1fwRzXWIubH6vtaV3swH0v/QutICkOQgHT
fZjhzhhPxQsAC2v2f0Z/DSGUpuJBwTBg5qYZoWnrWOdcGTFSjLYwUgAYIS5SXBiv
4WD/pu266NKcd985SWBPmcxTWEMdREc+fx6RFq8MMLYFQ/wz1r4TfLrgnzWkyM9X
3PuwdJAkv4pNolpHPWdP9/VWynF895WB0SKcBp67Ig0pJeUnFGG7oxT5sNTy8EqE
Tln5mMQ9XwqCVQ2Wsr61Iz8MMEsmTLDdhqKZQyCIt1qFQm2c+4I16wzKN+mTcboF
h17NmQSH1bLRqgCLP75Rto8QwE4bD64R8MfrF4T2HBy/BkszlzopQq1ZLjDYJahm
POfd/zK+JttQPnPxbBjKRGVOIy4GoZ+YMONpan2K2PzRN/wcQNP4ea1TKT8i7nkD
HM83yS7lXIvDcUaCF1cuVO+3EfeQqE0CjgPE0lq7FfnvYvCPAP8LZXsk9aJvspDt
yjceXIfmpJKHZNqp7TjvOSrPNZBTCS0RSudLaSsbZLK+JCIInYXs/RA52vmVXqYr
XY4KxMR8boPlpMUVO/0213FcrdcQh622LiuZbm+FRz+z++aq92xe3UBki1DPIR8c
dRmoodQqRKzFA+OjxPGHo/0n3yX6IytfeHaVLUY4MouGt/a1hg+lFxw3QIoTnVbr
I1YTSv9Tm0QmQM5gqlf3JL5kq52pdAGp/GQDQ9HaqT9ongO2K3/NJ433gRwgPWhh
tfDLZqLg8/yxnllhJATMgELGBnr4OW1BPERx/+KoJkPJxE+mx+lVyT+q9/TY/XEF
yCSE/xEExEvu0t2xX+vk4S3tY/AclA5xg3fKAZU67Oc7d+1XmKYmBOaM0/6LjmWw
MTsmlJdtPOz3oHuPNOi68ltPQ4C3XLEY11hru5f0putsthiYtTXDk6P1xq90lCHV
BAFeivULid6vcJN+lUjFjA/Mui4mtTAHawniQxz93+uG8Kdp6TxkL8B+juupl2JL
c6HhnPK2GvAteIFMFoFUYEhd8cBT1a+NJag6LZXE1qXq2YNpRZX9mYLjvUNrDZjc
4RNpcuKd2Y27gAvEP/TDQIYcslADcGPYKtN0bdqcoH08Pyg6R3dNbSJYRZi3snjc
qo+i8gX565ghybFUTJjjZ7AIE4bXhnDDqE2ZdfTKaEM1uDwtWuxUb17QCim71YXO
pEEx1HwGm6uPessYzXCGjrKkKXjizAdFM6TKp17FdbKVsa+kRaD1diAmIPJ2TfkK
FEvql5WVhvcQD2n/NGtSnMXzw2RyqS4KEFrPJWkvpJ3Un5+MN47Pp5btshdZ5zBt
iKvU5tybAOp9V+qD19BVun0EOykIiEQwkc1dysh6wRBrk3P22Gk5BNvmAq2gJtYj
XX2hXbKsNf9Sbahu/wg1mPpAxKyLUEoLiE7Uky4r/XJJx2N0U76KjcRa/cEWLLx/
l+V5vgFHc0A1HwC6klwbdfs+ac9gir5/+X8yqa1yhmT1nQxfB7LY9K2tC2oIoYMb
uNWXBOzm/TJxf5LkNt3Lys9zQly05uo25WG0Ez4vMfp19BCTZSDWqnVnfaN7Wk45
Z1CgKz5GmNgLd+s1/FaPZlazSimr3XXd1bNY+AbvZOJrBBIrnN+C5zSnv+VvTLS+
pbydll81fa3uueRbXA0MPEy0yfdHjh9/mwlOyOQHVZi6LjPPMk93NmXr1QLe26xw
WEBaKfIZgpDAfuShtPGkQUUslTwYEjkWjK9FGAEVb/puvPn1A6NtvBMhiWHP6y9n
fr3lkgBkt1YJmRCa9lMwSJA4l7HBr0yBDLRLejaFQPzGEohd56Vg+L90UUw57v15
W/u+EvBNBUI1Fo6zr4OtNiv05criMgvMCeGNoma4vWOV1Op83wDVrmTDY8zBIZql
gVgJc16ISik0IxNdDkZ7irE2PEMdrXxL2jjcKx29mKaFW2NpB9xE9dh/AAR7L0Gv
Ftcv+RU9WXcCPJuCArgtJnEwb7zqDVvlBVk0uNvQ3auL7a8KAy54X6VXOfcaKDdZ
8bTman21ZyoNw59d4GlswRTYCsOfZk4Y5B+3stHDjJoBr9A4cJOy1N7gs5SkEme6
oaUj4VMqUWDSV7MOqGz+GLjr2eucjKF9Kj3+7eodxHv3ZjkI80pHIlBnbgauDkG5
ehEUC7etePrK3ippehy/kLEQ5kN6ZcNDfpMUvWBweXo4L7zEY6SQA3cCPF4Fm/jl
v2CEvELcWWvQqGNZFZMKBnyJBAB0RFoY7ZmHsJTiy/J2z+U+1Htqp/aC2NjGauns
CP6qo/jCGK9DZ5RfVac1I0zv98xaDKVVCwGFlbw/Xm9vu6bK3jW0oaC7Kb0Rv8L/
Kxg/Ju2GEL3xKXxqg1IXhU9eu1A9JX4rqHdyvLtb1Iwt6sPaOFyk4MbZSXRG2Ubz
uz3jzF6I6V5+2Coj/F6eiHPysyVeATyjAseoqJ60P9h+Yl5nnV+e/p2NzDkrtHz3
wB1A1/3B1DfVriZA6SLlZbPCFcjknwI9ofC64JW4+Y1vb2g5tTE/5DCwaWCge68e
ZUe6Zf4KBEEObnsQebQNXzBU0XOzmN1VvVoIsIi1K2Vh18FM+0bAtX1sjlckFnHg
UIs4o/RUytEruZnCu7QWhVT1pRiuuEGHxGdZW3BFGJHugjyPHcWMuilkdjjdPlET
w4tmjWahAQ5DLAmqCz5fE4iuI8TONc7njVAqN0ltOOxia79l7ResRMLpZY9wGL8m
r5sL/jl9wZAkXQgM21XGPRv8Ild1rQJxNLu7AIzdlCG/teZdDmoeUg2GuVfpbWDV
ixNA2OMGLoMdZ9APvNmzkQVd5fWJ3frqx8jXK60Zx+YLXT4RObTKVJNjAk/hKJ7j
fILvuQaZ1yTnzG3TQeSjuSeX218dPyDc7RUS8JS0Lc0VWvf/2u5oMCGs1MNaIuxV
27WjlDX5iN4g5MJPV+iSQszLIO6cxWvy5poseyxDgcSDFhKUWT0NkEW31YyFGm5Z
7ZO+DIvB1SUF9bVbCfONJChjx46SIlWCr2iXDzJe9thyI6jRTQBLJG3L5f6YyXqe
7qOh6MZi1RWbJpCbRN4dEan5Lj+i64WoqITZ7eTfIZsn8h2abZ/K1t9eaA5D0N7t
lItEfJB8P36pvHFRRYO/uaMXJCI3e7Rmgs7dR5xwtmmPvVhNupyyD/9Gdi/KA6YF
oGNCy20KrhygXeStFe0RsdNCVjFAKhgXTXTYMlnI4eezyxRCyKWaWG24j1UR124U
cdTGdaKgxHlBs2yIzt+ZiSoV0utiKA1ODXEkj/HMe6aKIUBWLlTqaSFW5TOujsEQ
/q17bFtZHCwDhIKgmX2ZwbrLwFj9hFI++WPakFymgnL66Q+8nYipW1z1/D8r/UEK
ZLvX0X7++z8vKzZsB7fHRfhRt10YM1C2Xbq+l0Kvakz93N6UNkJT3k86i0eNPFz0
AA8s3Y++b6X0KXBMrGCDm+OEsnwAWtwjwK79479NahYXQ3Lu+H9lDUmUnxIWsmcw
nVAcCVgcQO1pwzbwRtyC1kJ8M2vMDChhof7SMy0pKdHqj6xg4Gnoau1JhyTKKJkt
1kcwizjOJbb9Ret/nbQQxI7sZhN0Yf/hIszsQU5jQ7k3zLlhZtFrUUwBQcI76ZG4
CqgJ4S6wm7PKKuOd1SlV0Wh1a4DNUDBnt0iA1FujdDD6wtXIAjCfTIOtdkDqfdiH
LTGxHtb0iAGbU+b1PCPbhkV04OMrXOrdY7r7O+9OjUeHHAU/vEKy17i+pLIyNsLO
qgjskHzohuP3kLtbxf19eqDWykQzBLv9C+drKbUe1bjd5IcZZCnw1QNT/8i4QCyb
h8V1C3jV0Oa+RPZ6/kSxXCEcb3QoCy7L8OSH6wFGx6qhJ3IQD7IMLStRcR2pwgio
V+Z3z08l+psDp42M4kLec0zfuiA02/3zZP08T4quTUWQfoO1MxLA/m0A2Xtb4Y6N
vph6HSyDGlUMfTPlloLZaatTpBGXzmYBVAmNb82rAIGjqz9iVbSNGx/2O12ZM9xR
MM8OI3hXUMYSFR5DZUpqlC68j99PHexZLwwE2DCLtL5vhfLIk/vblAcp5MEUiea3
rZUHr0Mf9hRAs4Nq0T2RKI7FLl9zzj5rtCmZXczg1bczAQvSViYfskA77U3tz11Y
9lvCiNvLwYTF7rkbvUruU9YJRZzaUDbQTRPsrotHce+4w3Wwl5cFWYuj5JDwUFXX
dBPB3iaPSx94BqVIR4WawKVL+OeDuocD6XCIqADY4UkMpz1/EwvXe2GuZtxEHDIz
5E3O8V/YaloEPKPTYXR0PMtlVtLmWBpGicgTZjB7xiaoh45nNLOqKSG0cZVmY9UY
kb2syYVPvaT4HMFLzATQ+LoankcKv2r1PJXvA9LEKX2ddC0InIRCPbuZhMOpjycn
uwM+WeBX0xXrLpeq3nFSAzUFP+k3TOfeMiOb21Nr2bwiMtmBwScDxeyzDqjWAS5Y
3kNKiIRDWuRD2agEMObaR97htJ2VylQBlVzpOMQFXx/SNp2QM5vANF5+YDqbIGmH
46AN++3lB4k1Y+4tWeyjbqRFfbs/SyJytzLdLViKNdD5IjRVupx3h+hKSUpEDmgR
O+LAnnLaW0EAOCYH/xldaFXY2l5dzoaFlc9nDanxPvfcAopbJS7WJZpjimWNCM3S
lJN965Cn5/3bjm0E9taMv3fvPIeT/QQPV7CNVP7lWWObqoCU3OChY/PNNgeUHwsX
kkzJPHTSiAboMadBu4hu7Dm7FVSw6w8lWMCqVxg4wSmAnCznqhXQEXUCx/HflXqd
5jA6EmoFaZWUCDCDCTo6TujPj9N/cGay42NMgEpR3AJ1vouu4azGUgCa2rMLcgJk
Vri/UhdznqRL1ThanLVJDTel5cF+ApKXF4BAqY8FU+OHzx7b5z/s5/Dw34IdeN4e
0AKM2gSz8QRdRvcE4KdvBI5j0bp8gv/uJnJiI6IGITtE3dvLRqqaVhAqtZqor1hu
XofmJNUEU9AIC9QrBjtRKQdKNF6Epb1QQnNCCeCNR2oCOdmeuZC9bum1JYZzKx65
N1/m1jqo0+/LJM1br6uNLeIXiXoqJhuxDa4OehU4jiPr9te1NTUINizkO26Xz70O
kEYdV67YtBvix1fzuqe6auu/Ep4kbtpTNXOSgT8qt47jrb8Zw7fyM/ZlvEIYieOD
Mn7IyU9N++rFBBBuws9GHIlWxiHKs0z70sH+FzboM0/s6NZF4lzGiHxv11j4kUrL
06l+F6aMpzccb24GdhYhE1zkDNoxgMLdMU2U7JLBCG5csly6Z40viglf6BfCgB8p
+7dY36nIrCozL37VMeGRx1ERES5y9W37FRITwEgZoMlkeSJLZ3bLmoH09gVy3b4L
VWrDZk9GtOmloXSKDFPQUJTBHafxTOJ0Bq/4o9fZrrDko/xrcm9B7sC39FAt/T8r
tsgwYzuIxVBMfd2p9TCvCiHkDoOb6NUF0xW/FL/RphaFP2OtWhh2wKscOlfNwoWH
100tpKiv1ZMKUVDS+Cy3+sKIVZP5RJ3yHPCuy8cjhWeGpfDX9zeWZ2gtZKnJsMat
ulAM+wzKuanyeDZTeIZMSXkiU+1a6lbxDKKiviZfe7jl2xmDwW+YoVfJR2jKUyP+
UIEOttu5IoInXFNQoiKfMrw8/a5Bu/WXu8KJR9pvMfUGmPmoHvwaXjwlsH4y/ySX
q7LeGXQP/FANDXCkboBQEQI7ESHXF68ylYMbNe9sOawIMfsvAeZBK9pApnxEisDd
5L/BUaPtXIqPhjJVIvxzdT3meVXfTw3swMejMOIWlx95jdxlOMk1t8Yw9Rq1SOG+
KYJoSgFfkNoDaW4OdEJarOd0YXB8wAnh2VdVfLGX7266aDeAvrgSOtqnDmVCDLkS
KToTcHcQis4QPI9Q6T73i+V9IrgHn/WdnbDHWvqm24ltalyN8oaSsGCYxjMYqQLi
WyD9iwZBXKtzx8UbZlwux503+9UxDTnT+t8tFQJDDpAdF9OMqfy7fsu6daguaEU+
kXXynz6KGjQFDKTf0G267Crl6qjGQ1GqyMXU0kYd0Negu6bbDJIhqFFLiIF3BbC0
nPURHJ9+DvLx45jSMcYV30jkaOdW87B0Kqpl2gcFORr9sGz6/HAojhKvG2JkP3e9
gh6/MI5/lFAX6QBqaxnsyiflp1Dq33aWwbjFWKnFbzzxAIUXXtRmssVyZY6wzJGP
uBDZcba6kOON0/nWqqlto1seuSaLZWpeMingoNOTDXbUSJ8zBq8i6Y27i68ZYV7Y
HnmiXyb1UcLsGPXog1kGFUAgi5lELbtV4PXtqhMxo+1uJ4M782iDMbezhl2F3qU4
MOoDc40xeHRuLHLntIOlO1SBwXkjhQsa7U8zgGuyTaG3wlrCBUK6aHWFjYv2QusO
Csoe4LLpv2C8/Ac8TTK+Mp1mbSgBnc7o1UtZhsXUiV/JgB189f0R8KsKq2NIS5Ym
jSoDP7YabBk6FPeIyDIo8rrgrxzHwWoBCAgzAHply4h7Hqt8dpMgANC7BTUMdDtd
lbwYCehqbrM03ZhVEWkTh1Mh3Li4X1TC/dyr98U02+mN/A4mTAEAab9qT/Ymiu7L
dapIupFBCU2+507gDwgje1KhCNmokAn1RkIzJ3Hpj1z+rCqJsgQzok2tkkLTNKeN
XR/qqucstzrjXzTm+tmwIZ07zrbnesfMUvKjnTKmivyUSTvcJRZYaG0boo+cqR8Y
x3AyjC99BY9n8USNic6kW/g/dfdvgLlLf/KyvV6G0Y9VgnGobDvywzKzACTIBFj0
c60+3Vne3yvj7xvKJBsvpHW52uYz/DDwU91q7LWdYmop8MSuPmw2yUBUVL1vzk2g
0Ez9AqoGtziUeg7+TiyCRzV4yBs7HAaGWtYdb9alHeNpwGLCHu1oLao0lACQV1gv
LCPY5LQpBDkKFcFXHk3M9tD6zxjwZlyLTV3p4cR61dXkyFgHiB4jmuqn7zMh7l6n
mDediIORoOttIUzOP9CCuLiCmbWwt1mt2Gu4E/hQLCzKjqR2Q05hb4OPyHcI/153
pIwt0pyvh7wZYKRq4vBl4fxd6MDxhWVqoKz0jMNz4bAxvgv/uRWYZl3hOilfQ1Pf
5iB7OUIfCk8YESDEQZYsxuandGdaOZQJGmwE/xv67bh47++YoNA5QPfNewDzKXnR
vUCR7Hphhu4MbT4u3HIqJ/DgvBrJKFf8GeBfsZZ2Hm/wA7gMejn5le2KkN/GxS3C
ekvczU7U8/5KtjuZ8ppmVcQ2L3oNAWDTwnubcDcJFZmB920M/kBdnANwPnPNHU02
ihbACdvvPgRB1ZXoaWX1hhXfq9fzwz5pFZBwa3vjn9bbjnCFzIvVDT3wvy2jidWP
cj3Ztsk7epF6bLSA0NBV0qUq72LPiQ27Ihz4GsXoBd3TPw4XszWIUIg6ISk6IYUF
cHTJHdbC9lu1xEJcK333BB5jXQc5oXYPLzUkSZGrIIQdHHSpk0gw5bQyNIe5YpQy
aF2o+vdQPWeBkubiBHKeKe9BWi9S70S6J5rbOGdpNdbWnp2DwdpwiCvny/2SGX6h
/Ct5pu7GIXaiya83mcuQqAB6XXBneaEmcNB4CbE2L/jNDgBmYTpf3wDWHDbVxNjm
CzJu0Jx2hxR3+EORqkyL88o0dtaRBWVZ/2dbwnbrtbsCXk8RjpEIarcCKbJwgT2D
QKHLYC+fofZSXuoK8Iv74hd1c9NVPc0f2gsZO50fuL3Kft8xJv5x+7yb3KwzN/r6
dgFWJZM6WdWxkE3J7WoxVacn9Dld22/PQ6+RRzbmHUvfVdZzdURvlWbPVFgATzUw
e+osrlZ4GhMBujrpAlVCj2jPIJecgokOq+wHT4QqbYcj+mjsK1D2ygfdP0fhwQWG
sjaKwo24iGieYwmRIB90jIyzwD/JZm5+6vpyZPILgLok/Ejp/tkwuhPoZUOSJilR
UlDIPGAsdVN9afv1sWQrWHKvPO+7N+5BcHIrbBnrtO1eWm/BJTi3cWO5JHgtbPmY
yhb1jGMjF+wUTE/ZdFjstkrFWy+L7Qv7lXeb+9U4mw1rP974b/qEiC6GODIuesuN
htPl0Ecc8ejOPXDGt4AyRd2YWu/yjGFmLa7f4bSq2VQuyXpOTXN9MRJOfRdHNNWJ
4J+l0tt620nkVGIvewTbvJ/Semw20dWDXgvRk/+XUOaY6ls3OqUFJLzyrSzbpUuO
eA8VZd2e+C0C+nIKYiCAgMmLVpFdCeK23/+uGNm5Z9ouzhB5b9/1BzhdG4JCogIK
w3zYvzG/EdhdegFkzheuWQOWZ/GvQS3qtrVYxjhOjieYHUs+u1CBHlvcadGaCiay
ueGKNeItRnNeVoAwxaOKeAQi7XFMDh2O2kuZNZTMJ7X4QCpXCuYALV9y/Z6TML51
H8tLa2ZQJeYcOuWE2azB82cnXTHxjvSpc5K1dfFyF6BGNlv3I0RgT04dsQGRSJEu
EP0ZIaVC5gZ7tPb3xzCXLi5tmXCIMHLK0Vw0RosylxhR+rujMHatjQUBQtylh/0K
p9yQGK88qzgF0HYC4cF23o4pkeROEAeuoEXbdOQaESW4cZc+E7B8Rv99PmM45yOw
oCjCHZ7tdfWBVwde6JZFk+lr53EN9vbGr1bhtvqmvvh+nZKpDTgTnH4BraYBBGK1
ixXMBfnRlez/mt7jkY4aNx3ladGhiF/UL+E0ukXGWkFTe1b4HQ8PGjPz22JY3f5a
AWdrAUMoLGZGjHlqjz9gplsI4toB6pMdq8l7OaFKXAGLxFpX+Fx+DMXv/GWmcVUu
syEdlU/0wkuVJXfJcEma1Z8qd7Pv+e0zEnjizTeG+ghLL9eyCZKatMQNkhKjBea7
RmLP9+jaXrG3/t/ZzvGLiwcDtc33S7hgIcdzSYOfSqkhTVpgfvE4ZR1eGifopfxO
3xje9gY1+QbqNK9JAI2M4RLqTjkePTPLN1EauebB7+tT/Nhuuji1L+2sla0p+W6L
grTv/TAVO1g3zhSslA/nhEU4cd6Tqqtgos4pxcdPpdoguajz7/OaI8/Z00uTEjEB
vle+RNFit7oREfIneqcjz80P7hkx2BPJNphRzu7OvMAjZvWeiWiFXMiyITSE+336
ERFjv3kVKVmL0lQkOPNUuoz4glnU/0SqgEZAomTwFPJovVCH/mVQxDga7GQSRbfi
xlfdiK7Na0a3I+2uq25kgjMO2YBCUdMgs3sXnYC2bQoEAPs59WYjyI4v5zyoBz3z
SfaGKtyeRGOzuGthAXckLg1oYfs0jI+yKMcDxfcSu7sRBlp4xpSbe04If30jz3l+
fNFh3YRdoIEw2DEbP/NB4rsqTH9jQ3UrjRgnBcBt0WZWDDnA26LcuoHXfo+xMxi5
O4RXE86AbiVsqYXpVlyjhH69OyqwcaQOZ4d0d8tfEZpGtxSwhBgb8DwXDXMKgCZA
Z9m+DFXnd5Zfz5HJ10ksfDYDx+3RJksmuwSeJL9VM9tQOsapJ8NWJ0I4o8bzlDOh
X043qS6LSoKpxBjXzOThohokj5dM41+Uz30ZkcJHBYJcV5srxqOjzQV1sfJXEExh
XRE/ehatl1TXFNmn3+55lzce0ioxoNLObEvXR6xu559mz8ffu6Y6JTdrYhst/Hb0
8WVZ/QTL7W0xUi4po1sEGK0iDMH0lVRTfnwFyMev8S+w4IcVPM/sPzPdBm1cFoGC
YsRcZgEkS5J+GPtD2Qhf1fKLBwmEj8ltNAekeoDaNYxx8AdoyZPKC51+KWgeErX+
D/czNnXLQxs9sBhOYjFUIn4YTdkLBsEpK/8w2TiNnVOYfc5e7PiSSjBxIhkKEsVj
f06uZWYivtJ/az05bDgpv18BYBHi6T64xVPntumRebJDEAECBQiDWZu2fJ9Gsj2r
iAWT8Mme6Nj/EIjIYROR1f2ldr/7oc+u+i1sA5HfVUNqvxDfICp7G+yVd9AmZSv3
dluUbeMmblC6Hb/YO+oyWDUw5mIeSCl9yxkD8iotfCcyGv0ot9FwAv3psCviW+MO
QWDGDPfS4WVrfepe8aeLI3ddHNoskH/GPdd8hC1p45JpPwP0b+sSF19EJ0qAeUzP
UPPCyIQSaZhTb6HmTViWKTRyS8b/pkFUwiKuj2Zm/XZfq6PtwWyVqotjk3mEkL1U
fgOokr/jiVVJlmKPluHOvSiG7vL4BNHmH/ErPOGg04cerCEL48qr7ELLItUdkFPK
U+F/0N4rOx8CEYwKWNnaJt5Y/OF7blKXhEuT6jOI8RkBKQgK134sKK5fV/R9UHY4
PGbQ1xJ74t9GrD5QdljaRrWhzxlCxGn/05ZR3asqll9TqrAGeCr1YYxPpnJxAUKh
8aBBraApJnPikEaAo2SfOe7bSoehKwdm5GWhd4Qu+B7SBQEO4YdwMf1r+2Ev2Km3
nPwLVDka74gs1Vy6gvqcqlUeIOSpnzsm+gZNl/e8DOew4yjZtixJNvMd10t7y5Wp
/WplapAPfNAWBtH8C+9+gCoVVHDrzAHXxTev+jbUpKAd7Xdvl8MYhSCbYx2Md6d7
8sAlLKSULXz8aK2a/7dXRyvealrqxQWIm+mRW4BfNm6bFuVsO4BU/nL2k57Ae8Vz
gz4zuoFU2AVyOhqJ//9N6qmovO5Rq6kjgwZZN9Nm99kOaCaECd0VKDgeNspjspui
C8H1sc4Ty1kkH7ge5V1Yg7nJb0UySOlkrio8Xpbf3kMtfvgbtf0vhhhTbrry+Qve
0k4ifnKSfiLhpoXhOiMbBCAx3wtSrg0w3ZSvufTKFi4Qg/CJXJOriO1ibHG3KKIh
ERxVQZ1CyAQ8NZFVWHs/BOiWPYLUSTg3kcaY6CYXbX0L2IVDWEYtx6IkP1Mk+FOR
InWRU0ejOVUxdFjTSGsM1Rin4rCde+KvlGUnhsiRftcVF/ZKCQclVI4Rx6GTzH0a
nznPcw2s7q+OSEp6KVRQ8ITvJLPhIiwW9zRYc1uTMjgu+LExJuJEKM4hhn6ONHr+
0O8uBCH+q2oPcJPZDdcPiHgdr7b2k7ncjG5YhlkIuTYnFWq92bPN1jkJqHZCw4HU
aAqB8k9K9/5rtqvRIFP1EGUl3RWslioXO4esEX5I6HjkbmmmmxzVP95tlwP2u0X6
k1IXTDmw35H0dnGn3vB1ymt9LLVdKPde1KtFSdjxM7TwTCZTn+o/bXPFvbiS3WTK
uvgY2gk5BFNz0Bbr3eSCToI7D4+g0lHb2jSa9Di3yYkKKbhyzoQ4LZy/wQ6kQRy9
R4UVX0bUsr4vkpLppwG+nH6q0P/DpQmPhV7TuGFNvymU9rlMMYQ8m8ytGl9O9Bp4
ZwQElekYiTNRqQu6AILOnF3vYXCldNobvEr3v+KRoPebbOKpVRwWzJN8u+ElsPe7
4G2K2JttDm6ycadR76Xyp4omrHFVJyWuuAv7rgh3mWd7/JzDtL4rzeVqXWuVh9nl
Flxuaj6lVoHxX5bvwnfrDgk/IWr0ucMR0qKvvEHcBoPUA3NDwiWZgM/Dh+bZ++Hr
Em2Uo4C6GAlR9BbIeAJbHJ1YPTuSUSEbuM0P8m0Flc6oqRo5EHBzIeUhbL8t+Uqo
gO9iRMjAoSSb48QicAHcigLHP4qIFgHskt5lDUXxyB1/oMwf7ldiWnTgxjTmL0HM
raPeslqedO7ChWTMzntAka0OKeFadOFLjgzfTDBvlzBVDKEyYQrVDc/ufLu9aeCR
EpAnSvy0B9wW3rZMDlJZLUT4l72fgFtzi0Iypt8rxAt4bgPWwXqSwnWkFmwL5UWL
QP4vGn9w3TAJpRVGrGMyxRHubjhLLFD49OY9dUr3UVpPNQnh+ZM4Tz8se3RCiqBk
A0jxobiZxH670+xuVJmOi3hN4KS/MYxtEqI8eOJ2MEBzgzKffM1SONZAEY+mvnNC
12IDj3QFN2jA1dccb6opeEGktzJEJyUrFae7iaP3WeC2AGJUUigFaCMaGzBcW026
3fomKQp9zora1TApwMPiS2l/Psp5+A0kyX+K0IockHLBC3EDA5FZxdYNLGBZRwrX
DO6GIEhooJxvEZBX20XVzFMcOu9Yol9OnQ3IZghmgl5JP0BGeYdW8w6+3SbmPlSu
1vfvLTLCD14j+08hVt/s9xtotBN6srsMPyN8f7KXaDjUNbYd/zR074laM4RplRcr
BESD7AEC35AnzPzidZC327r2RcrU2ahGPePRD19+DepGhdqu2ok2x1eZt6vCINWz
KBwvQ4/uSgPAy3xcnpM65AP/JqOLo+PGSfrctM9Qk62/szx6IrXiBLeQ6JBI7zIf
/ifgsP/0t+40oEVIMcWpJLv2Vz0iwfi3LrFX1UXVKW8CDfiJx55GqlidbBPvNQ9J
RiHtciDv9EPiDpknSKYaUEvSzHTUrNHnEL4jtTCQ+z8LhBCn56cjHeuYx150Z/Bl
AlB91MYw2cOhm9L795nPN2kY3Y/oruyhQiAHeMaThoVwKoYkvYXJLQ4XORiM4Yql
7p7upUDI7xYyCEPTRXDJpxw4HFn1M6Pv9QGbh3NmOs8JuiGQYbgXg3rWEpqaNTPv
gHjOhax5eFdWIx/P2kAprWyDXRueS52pwFEHppo4WAuAAmfGLhT8YqDIon0X30ZQ
NJ0dNpnep7PJggZKILB/sIdQCvfENiIEkxUqNSgUtkmwq+yVqnt+c9FjQh19wwO8
E1syDl/PLjnoW6FHXLCFKGsgUHA6xIDyI690EFeOeOpAxE++kPbwYrYVWg8wjxLx
UMl4Bn+idmjR3zq83mZizs7O9g6CuoRmNAj8UQO7DmyCTCUEcAlLCoke4uRxEYwf
rkc2RmfRhsS7zdh8nxjC0znSbPho1/nsRGpA1pGeHVWSb0LbYWtgPmnrTdVlipFM
cYjc2dRYATyIyd47CP3eXKPzziuJks0IegIRb+OEkNWt0ljC5Z0SNkujjZ4TaqSl
6YuemSz/7nL2iRRD8NQXz9trUFDaeAz9W0r861TTQqGSA/Btnbcuu2irpRHcwncv
q7urqqqYzsBO2kbOzQEq/tJd0XYmxfRLS/qGjWDU4i5fanCgiYrxyx3hQriF510C
2NSFrdnASYVug2myvq72tnlHMQC1/TDc7S3h+bO40i4UlB6giQwmxlnmTe37Wd7x
TGcJ0fxnazUHv14y3b9rSuV9LVfOcFVZdjBH7p9CiQsIe1IbkupaVXlr0rK36Mys
HlWXvLgxgM/dNe754So7pLaWTfDTPOfsdbvANcC6vGZmFR0ARQ3kyH+F2lE5bC6I
wNEHREygionAeo8SmvxwhJh25qE7nQa0rzcV82dpARHqJc5AkHyMJ9PBo8suNZk+
HM9tFQFJG8QU+PD+nB8kNmnuEFRdPRZ9hlW3/bJVopDoMjRkvn5JZ4fSSor1CN3Q
n8fMqGblL+5DXBOluUx8LwCZc3g+u0qmezLQVZj0AIsiG5XDKhattfUOOdoQ73md
f2kCsHmrDSW+VHrhdw47jCPvUmpOdQw37mP7Xlu+HOyzyg9/MX5pQSg7UFaraYJL
GWaL1Am8BnEYW7aMDgvNn1oo6qWpDHzhFbsilIIwi4aX7CF2S0aSE0xOhY2uDLg6
89LVT0eGs392n70DW5FQqwsKSutqh6bUokq02xdzCHpp/R5i0qLQ0Nm17FLPaIx9
j2nLdkzc9gd/RQLwoGVgmrUgVTbEtoBc/qSGYQxyJ4yGYw4kBQLIkNmCwtF/JjZE
SS5PCVEAuDEZuJc/lis48y9wJQD89WbsZje9p2+fVOHeggIBxo8ENLB8NamzAfwu
UKnHxhunGXixf3MDHhqSudAIyYNtbmoT5wrKkBx/n8CJhNC0yq4Mg21jK8zxeckh
Dl5d1ggcovmL0ODEiLJZdSMnQPGXH1eOr22tXiMnJw2Q95+mAS+khcuKYVjXeTOO
Q08f1h1gVxqx/5lwAJzfg9jExjV6n2b1TmMEKzVpz1FftIbvBqhpNrKFnkhyQ3M6
lk7VOW/cydvGFhIa5X+3NTBgdVhtImhDkVhnYRFI+THXnAw0+g+fuEaFob4ZUNnt
3nQ+hN+nFSwuVt0QzWyt6hXDex9aKsVBGOlGhctCkLv+w7wzmYGI2QxxC/v0EL9R
T49wucT0tX0C9BnR7fLoyZNtvZYGnxQw+V578TgjiSY4vs/HbthSdH+uQDOKN002
aVzcyF+Sz2a2UM66wbKqj48jaCA7QhYEmbaVwZQ9NvwCXojSoz1ILDQp9g0XZw3b
uh1uI4Yw1H+/YReFSvgS7BimehaOXgv9laVZj33gXlMF7cEJd6DsQIWxiUnw4op6
vZeQEg+nMrkt3S/kDn/YhW3CgHRkCoPHjntgv1y7nYHnUDyYj+smC4qwH6fMYPvi
Ty0WC8woi+m2URXD4iBsxJlyjNieUR9q925DeJagNcHHFkcQu/liW5kh0cjKX5wf
DBTWzxsKmBwj8a38lyQ0AUiCnw3nFF+yBiBjCzZ9KviC/d2qE1MYLEuFonGiM4Eu
UFGSSLZBlclFuhoDmqow2+YdAjmCGP34M5j7wzPXywLXppFvl1vsKWAcQ76RRLR/
0VdFxVzJzC+NeEFDEsQ+bEEwEhnd26n6Wzyz+G0ST+mSn4YGXXgYD559wBucaPBW
or3KdJL7qytTstR+CXUCzUWI2fuUXO5lNH+ZOQF9crzlZvOHtVFGpnqO0STxtz88
MQVD8YXJtVpqzN7JVlOPX5PlRKXkgn6wBSyWHed8r2KCthSF77pPPSspzjVPi0D1
wqrZBChUg9FO2Wh0ApsoF34JNXMBWW4HdVyAPT4njWToPWiQs5nM31j3vLHYGXsG
EJHUe9KIbObANhC4xw438oadS58NXUUJjKJWad0Eq4Uny401hvo00Uoa4hX7ChF2
de+sDOCATa06wuMJ4eRMbqP6GbPi4xm3HLbS4p2UbGdJamebD9VTFwIP2QdlfCpz
BrtrJ2gTpn2Eq5WeIBZef7x09DbX2cuNiLIwEFynf5H4lDRVi9l6suBmOQFxCCft
rIJAwRN6px9E7B5wSRRa/SQ1bR5VBktDTRLvLtPgmK7n3R7/xFvSILlgkCo+1jbO
8CZEzpguURQM/deh9Gqz7ryjN9oKto+dU13WJOOeNm6fWCNStSeWkpjeuIvGXo+u
kj0Xd/gen5QaKBjnKc80f8udvKgFcyf9GXeScSz2sqg3XVIQG62xsv8MXG4JEbVq
jqBnErvKEbTFEHwhQWZ6rnhISu1PblF8TuHO7FEmr45OJ6pdKAowPV0lgQoYKSJ4
CSg0fMv5l2giCZS2Lmaw6MU4dswugQ0kX1GJUZRkFGoR8pDMEEpDMGewozZ0ID1H
Q9Vjb2T7OLrGLkC+SfFZDatDSAXXwRXcFPg13CLYRSSqJKv3qZ9s+4EGsXwNIiCH
kj6dTcisnSntVvG+VrM2iCBOfaxhWz3rLnC+AQB06QoiuzLJ0syduc9ICULZprSk
gKcJRelW7YDZZSo0Xep8U20A99AzR47rwgRf/KEDgZ8bg9A/3Wm/bYDTbw4pZ3s5
LaICQMBiyIdQ46+D4CtbhuC6jLu947bcnZ4IJkmwqc7f7WjmcKc7+Ee9rEAocqTp
pnP/OOYvJjj0GdCwODVdtBp4EJCrKHDfPOp5q8Oi74xAMhN0181ms1ieQF7lR4qD
LB/e4nOyUpovK8GMpr7EFpU60jifWML9GltYmT71Fps9Rly8HOYpleVZaKMq4FRM
1e6NWPPeNvF1dwZiQCYa8pnAIIDzyy1n83H5jasNTwNZfkI6P5sRPJTr8oIquE6e
wo8hF8O0N2D/Lr+KhvysXAJvX5oBHQgwAiV8odcyPDcuaQDcMYEtqlCq1KYlbUqP
HoFbjh0k6k1qCsrv/DAcTV2jxQc7IEnHYynP3Q8XOjwhpr1KEXrofco34UtdgWzs
PV8lFYysmT7krc4MvGOtU8UugL3yyUs1RTpoy5QY44i1Owy83odz3sy4QRoZvTn/
kA6MrN7Kgr02jtEFT9BCy5Zi9sPhdm4yAJy+RhFaUoWG/KGG+iYvBEbAZBDFs8cF
pjkYzHGR9u1tA9VuIJWKp44qU8rECAN/3dCbFGcjldAhCF2JvlgJpjpqa0OFMt06
cKLPquc5Ci4+M7tFHJWyYxzyilsHyE3sDiE2BiSIKr4UIzUXLtxkJDEDYf18Rxca
jbQx4E9cXjsHRITQcqlOBTuNyHVB6vb+aG5nk0zyX6dTjE97CAIrxmw+p/zHHIvM
5kY3YqcTTxDd6Lj3oun/JGaIn2v5YFuSg6ZeOC1iEKVKBm3vdAKD7R2NkYVmNv3d
KC073spzTuR0N1xJ45vtc9NGgJBJkBUti3JSKh2WLBFtK7gEYxfcDjR5Y/KxpL1Q
aBwPbPTjB9VzqUJaaVujNTE3aiipJTQCE/i21fAfKKQMARW/S37XAxbvs7/G9NYl
9Pa7U6OrdJ/mW2UgJhfEq+4bGI3FV5S3w7dL8KwA94ETsCI2gb2oy2Yj64iIFPYw
0xLvflxiPf6OwgW97C1F9YzaN0pWRgJfZy+ghKwaoA0hYaPWOcZ07BjdbtZE6/si
RzkjctLDzDwj4AB0jpBZAXoqUxq35Kjpa6RxcaHfQYXJ19s2lhlqLBmT1XHxH2Zk
zS57eUiinjDpfJhXMRfYLxiDG9ihINDyYag2NqFTmZpVZgTa61MY8D8G2fjCYjjg
AhtNqhLVxweSrhJ/BPR6oHyjDFjtgvQnpJwNALlsohHIEsfNC/L4TViJn2Anzdpu
XnPxZO/VNQZlA6+wt/AAl5ebuGUgfXzh4o/TEPtlmOV028Xkj9ue7XaHlc1ZSUq4
M9gQEPd46bRfbUYa2Z7FUtL/wrAn+cSX7sEz8nmL5tK0mfrQy11OI3ykLNgEZw6k
kjPwAm316r3z6Nu6UvyahNxxseG09DZ30LZgDj9h9Cl70MPRX8RUff8NCAqCB/Tx
muJHn8lY2LfcngXqBinujkxf2x1DZTM+0c9KfC5TShbS0uW91w43KvkKBacjEK77
VA+8n8+QJX2X6we+eGCmWmg0P2BMDfEJfckJD43um8pfUVcugleY859xLRd7lukf
PhiGNCmId9aAxFwlDFS2uDl8qdUiCZFs3K8sjvcBnkLQORxnttiahcLajS/n3d8o
Ci/AjtTOO/wk4Yr0GPiqy+eNVmPb+09liyN7UArdnQ0BvJz7Y0I0mGip6srJQpYL
Mv0l5m8nK374Kso/8X3IZQsCbCUv7K81t43CyD7kYAPkoorQO2SPxqzB7IerENs3
AH1MVs0qJJ9wVoYYvPcEVOesp0xG3uW5exnYP7HFtiBeV0u+VVAzgVXrjD9ASQqj
wl46P9+TcoUbMa9y2LYAOs6Gw6b7u8cAQL3DG98QsMWEAjGTB0AgGjw+Wb78BJ5f
Zne4D+aZYPpYAHK+lvOm6RJPOZtpDtesDEeIvmpMfk7F2HUDSuZSFV9Jhop1o+wa
1SIMEMieCnhkRmkskdEs4L/Bgj5UCq863sBRzpM/ZZfTYhLsQV+LkXqQKCNiR3pL
kHhZ+T3gkv5OQwwgD9Y4j21m0P7YiGiP5sWymjfdubjLT7s5c03qBvxzSZBlS6UX
K84YO84aIj6M5G6WOS8HrUsgpBBYuaqSUIhxy0llGWs115M6kv1afx5JxUHuMA0V
NGU8e6LcwJsag57i1C5+BTRUsjl6CwatbTED4bgYXjQu/m+QGR2akgrjwTuAGqWQ
HwizFkk1f9qaGnF8kXdMVMWG0QXhVCgLKFAV042HfjZV9yEtJnBk+PDscTgwCxNs
oWE2OEulbtARqmsXrA9yjS28S/ZSgWWIb7uyfPHORKCDZlILLLVYjarpJPoiBTtL
BVUBtDjwKlxbwtHUgZhHr366tVnfef5fkmUIFfSwDZOo3rYtRqKBYPhJeBC0f3cK
OKOp6NdtG0+hwNApGov02wYPy4WQVnKSuq2rYlecFpK99s/lPy1nWkW5XsZOsG2v
6XGjHNQKVzaA1GATKQkghK8xMM0x8lJ6ZGSb26JWJlkrMgXCw6Ph8Zfd7ensEEOo
HZJnUce/C9yqxhRnc/e5PVue2MbHsMUE6jezuU6m8XxOgMtOZ5WwHFXIFqKH8h9U
JVWrIDSR/fQG/H6X2sh09Hmmkl/N+XHfPGqfcdwyhUpaz+Su2kX9jFinoOiONZhY
cV+QxqFqNp6OwhHvjx3ZPB9CWkE/fRD66iuSIa2pAbMHe2Qgt1xEP17WY+Rq/H3T
EdTht3rdfqtVKcNBGGHx6GuqCN8+cufYz4iv8NZ6y1PuO0aG9BdCz1topWSnSXyd
uNVuqN5xIRvjfoy9VxqNHhFXcu4A+Ukw3DXSHfdgz53IUkme8Xb8E8RdraWBTj0q
J+IDSsdfeRZ5SNx2pNTiofntmQdCGe72DmqVUTuTBBdaw8xvECfiHsgFsTfMzGnI
NkcmUKZLCL26PRbpguFAcg5xNQ+I2uEkQSeKzfAFIr7T0i1Q24nB0RWHFzI+cRWi
8jJh8FSG+E9GyuEj2I6cbNif4qopfmQw4JQfz/nfIvB+BiWzHLcS8BUenrgYa65c
i8JbslhZFPcclD+Op5kkPYSoYAWItXy7nEiynho5t8C6AfW9XpP2b8g4xLH3/Nvj
ix7RWmtOUSgcXYMoyzb0j5NGaeIJsX1qfWzS4sjG7xOdaI55e9KqrRhl1kM3v7tA
malymgoO1ngcW26fDjGQrDBDKlQNgjhirHlF7YLXlUGRWJpTQEATlUXWpGef3//p
RUdZkRiOQmO/KKSc7vrXnC5/pWsTXpwQoPsfAgJ5Bs+0vBIEIMff8kp/fTz/S1mj
QveFhjgV0cn/WlI3rycVcrqpoqZBXAK4UunJYgXnE6RNhUU5zYYc/iwV5AbcfvFH
5BJUpqcsbz2bDQZtMZ5aA0G+d0+LwzFgQu3dcx2tFPmU+zuAu/4I3RAl37mDD9s2
8PesaYyaRwuT4jLtr3Kq9wta+m8rx8xFmvBgUtQFBAJbTkFBn0UILSWt5B4OQgfz
OUwUqOkhlntuYHBAZX13QEW7SyikhSrExHhrkEsJ90b+IjY433w1S3WKb6BhHH0y
owg4dRKl6kyPPcMJdYIWIYw2J8FyBxT20VcE1Zb1f1R1tqU+sFScZZk02EcTN7q+
IlS3CMHkqHnUMs7IXRmvjlkMVZzOh/zmU1AvggxcorjqT0Pax1dI3qqNG7geggex
ocTWvF8oi97O3OztwPefaDlbBzpf/3k9UcG22LYMX2kybIigxSxBraTus70kuZlX
gcMvrIaA8Q3NzG0Dm8NM4OYXbRwsPycdzdb6huTRkJvWCDX0d+PJ74bMBmPhOd/g
X+SvrH28LJqJlNnE7DR1vXRCobqJsMJHy1dECYy+NK+fGYlVBybinDScCIF/bZep
lmwmTuSTBLvsxRahb3V5pwLInxhbmHquLHSUqxtliQ+3F0voJi1EGLBITGBTPWVL
LipAHZpTj6e1pnJSb/AlP4YFnheX7oLH7q12gOYTEAujg0knjkII2MlQMjGCs6OC
grPBWVLwn0xjuntM8Oz/hIxqJq8DMbHQYZU+rGM9imDC5Wvi+lzYltUYtSDnStxS
VF0qu6QFELp3bGazdHVEy4+JB/IZ0MSpDaBg4wrvZrrEQHHCZFD7RcOBIyMQ4ppH
P6Xb/3j21Ak8lkYiiRyQlVoUxSf9RugN9Yd1s8UetQxcSdRJ02LDoLb//wQkzmZA
5BV57CQsIj+0ikj5R4KDqbIke/6chBUdB/J2lzpC1zwyXq1kBbPrk+pW/Efubmq1
QcP3rfK1IDCJaaFwv2oFCAmoEYjG6TLB0hb19qTNd9Qitbrsqt7Vi7LYe16Ns3nA
MjqFiTynUxVHcUArSf+kGqy0+jYQ/O74SxbzSZ9d9ZoCmI5UKUm0VJa0qY0tizfJ
OO2juSbqEx/NDxzvFU10aQ9tQwzAaXJsYSYIaBRpADfEoHO6szsIOHvsJEQVhzNa
4bETxVGQE2htjDSD9p8WpdSSwCocInX/OR9dtzsamlF5XalGAcVYbzjJIc9WnCd9
yaY4vpUK6ARe5YfAPxoYaYjwjmKzcGz9O1KjhssOeMZofT2dAqCjMSmlnPuqio+O
NSW4u4IKVgnY4UBdnzpWiCA7uJWhhwavRfFxnnRUC/BYUmGMvChzvs+dufNMFQNg
fqXi44+3k5vihse4GT4VvgOGV/HqUOSVlzebFoqBcfFG60kIF3JZKPeFfXXK5NHW
f4WHumfly2h64QBz3My8t5SBbJxdJZS+8wRLDtMHANNoNnNv7hPce13lC54aUagO
+cdG480PFPbjjBwfC5zTNs+hxLxYFHJiyFyHbZGngUYrhkzLOTPXpUA6ICz3EORS
gnxBnsGE4jnEGNCPtedRUBROVxyg9Mhi1nWFOCtKQvJcK6ijG/Q/OPINssrZIWW3
thbvHHSnjTp502NwE8K9kF1qQ72IGMy026uBWfQzNIS9yt4jqgrjJJS67qyb30UL
WkHLatlbsV5BNizzDCj3EpysF7J8sorPak9DPpVDeJQwM2k9v/AWk76RaTykYp1s
WlWRoaZZxqAMuXvTRXuiFACk0cDODm06BnaG3sB0SiH1HHavhJc2IOCcOTZPp1Do
UKeOW4CjvUBTjBBaIuvI+Z9HZRarzqzO1pTpGscFVp91pyeHQ7WhAzfPHH2IJ9gB
dQDeqGab8pVeFPhLHXmwKpk4EGe4AyZJPghStEkCHAN4XbX+ozgoGrzhKRttzBuJ
14DBA0ertjIxcYZEYaqBGOgaPVm7GGEQH52kVdwKGHgqa/jAHOVYEOB6gLo0t7cr
dN8J2xahq4p/TtZmOehAFDsZC6wvw6Ns2rGABlHYSU6mgOe1n1yDDanQy+ClcUIf
/iGXNCmTScjQ5ugnetGv1GLbCq5XU1M33QlEfZR/158jL0jwAJX0eoPJfn5kpfjJ
tcQB0dPY/ML0HCT5oP5+OhQr+WdBo2XRUphhcY8JBM55jmws/As4eZGF9ddS7Dx8
nFkj9MTe2c3C4nt7T0zgzF6DOC3EEeZvcdmQjJTDWHOXhQedsbaq3w+YU0gGLNhG
jCGs86ESHbGS5CgkIRuypAoD8I8evwtCO4tPcD7YzxrYbMOdWW+ranuoIzf4+umV
2mF9QefLK4WygaJ3L1u53EJlzaxZqIdP9ZoJnnVwm/S2a8NrfSoUV7RBnSP07LGs
z/bJBiriIWjkG8xABuOZRmMNWzEStWeZOQ7XeV/x0C+AKYpIDDx75kBMKtqA5rpI
jkga16cdemir8newnZGHTxz38C/DVbctoQh1RdgS7Rz2q/ZQoavUMtyxSOZ6k+Zx
rxFszEuCh2GvQBRN0qyMYYOYDiujxuOQ6LPPxoUiE1+oeGlFV5ORTvW8RvcudXsg
TF4b85d9EWiv72VqKQ879YHtj4XYHCas8z5dbtfqkZWrvNYKPa8LJZlzW+LRT68T
jzMvcxAs9ZwvK7Q+UPDgOxVu4hCz/AxWZmMDJfBFPPl/pyD9srmfXb9DnenKvwQV
wpDb9l175DpNj8lCJqH3hcZxQeyBuLZbjhi70PS3r0a3RH66LWkI0MKk9hqdxs2s
fIYJihCh+ulX1YfprMvk7xNKb5WiUfgkloXrTdnUvqjytxm57ZU+Pvr578BW5XxX
e8TaGbV/AwZhGuBcDx0dISZBsupuLH55hnqVj4kFYndh7IFlQU7e7Bbe+zxEkM/h
/TQHnjZ13lFGfyLohU/ZvS+1V/kjK/Q6nt0oU3zgOr7C93TvshGgYSnRSDrkdoUJ
zSIsw8AXjitPTEhpX0Chpu7WbVQHaISfd0UEbdNnkD5OZ8t+PJTC1rLRjBEPH+X6
D7pWaMP8Miy8nwFkbq02Ppy/irEyH5S5IAJfhXeES+RV+8r02Nkj0kwnIDi0xca+
tulZ/dZvLVeiwa2dsPgldTUTNo4EByU1KlqgKeAipVeX4NFSoGAQ1nYiUIJ8o2qJ
CMeFAucfeqBC+Q0LnVZQGpW7asYyAG7nM0Bj/TzyW1S8+O51oXQGp1VyySQl9c2D
WEOhjcZ7g6S+1Xd4fxfNzO/87kEs/KZ1gG0o4zzlj65aDauY935GHmtQbUMIU0F0
2dIlvs07DzPQ5VwFVSLxg8G45I6t3rTrfZE/1nTVosG9werpUD3ra7FiwJwvr9H1
rWwHhmTGsT8J6s75l7smWSiHi0WDzWa/b7qcUN+eIjvfaC4csincACJ0NqRw3HXx
76i8Z0U3SoZURdpNjqDNTEGOvbcvZEmaeexsOcKxE+4nxRzIqpGiLLQ91naEkxnF
au8hNaSqrXnnbZM3o89yi9nWM6pdaFgESopXRSHCsyMnphxhMi+R2tQfwDZOWgau
c+Y6kiVWnT6VKCGip5rfU3UXqTqZNgXVfhn5ww0VtnaS3qoTiUFfnh4kj94GNerX
hLkIpAKt9gYMjTs2bwquhtssDWUQ0EJCfPbcYGBye7WOdW6+GP37LCv5otsGM1i4
J6vCFpjUF/7/D20OVYMas8yQKErjuY1R5/Y4avYc5Sh1rOEYHz4q9Bq5RcCNJZYG
d84ERlyWVh6SQO/ok3HBgufMkt//t9C53P9tDeLsioixkmSookGF2beQluk6fVr+
SRX2cSNqhpRwcSH6wQ21cYBGE42J1u42ctmEyhpO7rNScRS0ELUNPEsqX8obynQK
IVUOAqUT2dx8SmdWxz9IxNXvhXwuMgOGM1P3KoeyuKDqgMnGWBr6i1PI0mXAxVar
gqIq41Et9aoJn32PB9uH7S+nVCu3H+kLtA64aA+FdB1VzHdYH29sum3kdbjoHDea
+HtgaVPj3YB4McjMeGYr/IBOLdhSabf4llps2793ixK2gUEZPlWYwOk5XH8OL0IP
5uZ+wVptmp8H6cjYxkGi9LfDERpWc+flgNQwqP8dix5xZruYfgUrMHyDqas1ZL9C
JTKl5yS3i3LgaeFhH4m3be3j9/KaDvYQ8ziyMltKEH21U7DJXL1IwIslSTYB5wQZ
fiHM1sWB21uwrJE5TkGhalNseTsa2aa/UmbMZXg3nF041QDdDWPqX1lXGAwISg57
0b89KreEF2EX9CpjHnF4N8ec3PriCODdHmvwwUAd0UNPE9c3Yt8lR10BrcS6IJOx
4NnL8rhstXuHCi1SWGmxL4uSOgAupWu7jWYmhXrJXQyNKuQvpLMawV7F1Umd9pYq
C8KYPRFcW3qnzmPGqBwlNMCUQPYJc40u8q63TIqkTiDzKWIZURFBUELbktgMjdjK
WAY8kH1+bbCsT4G7Yn+SD/E4CcYa3bU1D5V88hqyyh3nkpe/HGkKkOYgdGbkbPJv
CTdxWi47McoTjLNGurWsgSswrsXvFW8kB2HArgeY9JOBXcVOu+o3hSO8OG5PeJi2
/F4zSTO4cXu4GJeoPXf/IeURnfWPV70Z8QisMilAvwwG1eszic3pCKf4TrW+eTo+
zgSdaYJniXBMw75M0UCpHdVibgx4zWue7uvSs2Cli100c1UQoDCvG59dT74fR9Rk
CEMnRKgkyRATzI5aXtiomQbGlVLvS31p0Hoa9fy0+VU636cUDsj7e9V+M6KGUcxJ
9Lnh5GYyF8iRboN+3Rldo1HMzHfb93TbytiOGayQaKKG1nSrAsaTdS4GLjk12KPu
Y3e2x8aPRF2pePzlgyvlOZ15orR/3mq3FFoDGRgl2p5MpdeJU9LXTcwTSmbHMsMh
JbkeGAAvDp90bg1OiAVD6CHfX5N8zBy4EqwrUrbqViMtaX9ZT9dlfs5FeSUqXeH4
s0dZ7CE7h6K4/IS3xO9pyHZXqY8xs9S52Iwzf6RePh1gkaDmg73j42BUEn4ticGs
LReuMpKr+WXYkWgmmlxh5cK3fVqmIjlNdZ/G/AXyQkU+/CsxLnJTdYnARO09PulQ
hUNqw3+Iq/10+LlSRfl4Qz1Ge74uYsleLZ3a61LwyoSPKSRO36pSmgcxTCT2X4mA
sodaLJ9b1N+uC3EHuehXLdgS2mFlw/FIgiZhyNLTuTi2+Q8AVuflAdSCFHpK1VBT
dEK2/PkWbL9WFBG1hJPOhTU3PWBEekl2Nw1d63OAE/1WSJOYvC0I6Ka2VdgrSsoh
EzoNLTDTvXkGaIUUAZVssNYA65zzxHsloCzoJ0ontNy7GZfJwwCzP2+xEcBOOE4s
TzBaj0SeHyIqzhVpAYoNMN3lFxJqg88wxWcodAhY6XpbPuFTkwG7w93ev1RNmOtt
4wKFTiH5AV3mtLrkMG+5dHMypeM6rEbzSSSRCc8d62ysH/jXGWcFk9d5/zRd6TPh
cbri8RbHfqLKQJFTFpbxAX0JCzuTyQyH+Ngoj1JqgwAJvUDAujFXp+ukxe57SIIu
k/ydaEaBLQGERKeUnJjTpZ3zymrcMUfVfjAoyHbAq8tqRNmNw2GzB+aYbCk2JxyI
e2M5/KQgpZkUs8kE8+q/QPspiqTeIK59vpFfOfMKnrm8SuV7SaoQd9W/anxSVa/O
QndIzj79cmFWgzJlB6o9kOW5NyVpzcm2Sgsl31v6DyiaomTntxP+NM9WtVAXNpTr
DLUxYN59OGaNOZVip8H9qRitYEngI2wZWncxGZVG54v4qJce48MB+zrfwf4L4hX8
7J7nru9UNr9IVWBfc8udgrhUwKxrfXKBby0dgzzFbcB1B2Q3j7famSW1v4Rvvlix
JVmUzW3Ol6Y+Z1ZKP/A+2p1XfNJHMbKc0uxD0pLds47xncJ30oY7S23BG3Jq02lK
vpL4K61AOZFOSjAUJfW2Ot8Vll5QrM0oW+okjcGo9wyS37PtTdosYXDDpJuiZLf7
eUZ0A9KMW3cdvLwpye5LeanxjsWn0f3fHbXIfV5OQslJWag3JwczjF6klB9cgjk9
KvTnvZhFUz3JgHsV6sMNQeIpKMin76klQyj1tjSe06GCnHhi9TL8zNXY+vRXjS4M
XbLH4V6G5kQ2cYEwuYgzmMRx2UNmxuVVoC9TA3W/nGojxNsC93gJeRSGrxznloeq
SSPBfwklno59i9dx7S5Dj9vq6p9ThEUl4+0xh9ydW6GKoesXV2zWhr5OE02shIwD
C2ssb5cDEps7ik9MOi84m3d76A6GFq20lIlvOwOck9frhvWoA1Tq61NF2dMrryrQ
SP6xVpQUQo55xSTy2TzaD4NAFyLGqdFEu0M09yzIXT/7f5cc+hJn6lwNHNmwwT36
oIEMJXXgLGLtR99Jm0Ud/ZFKzgZ89ObBn/gwgljLsUMwECDIEFkms0Pt69nDxYlu
9I4can/YkqukFtf3GG8z8HxrhDIVUw+evMTPJTPo603uEa8LBd1zMrYesJxtEvsU
WBvGUkXlpi78vsE51/PB48I1YX5kx6YBvKYvZ6F3by8IV7GGg7D6EoWtF9ryp1K4
rE4aLx3kSSfC4f5f23XRxXuC8+FxkPwvjFwv71D8K5WnbDFV0CMpQOVS65DXlFp4
01xNyZ+c7sSb/r2a+iR9AS3V97k4l/HtlpT0EOhP/2G5wqlIpaVBf7jLNmUefmql
W0T07mZF9f68H0AxH3jAZAhcyP7WauiDWvmlVT2uRzQDgVDDh+jubOBg1T+d1qnj
8EC43cSgTWvM6EU3M6hrNjtWatSbJXthknKuyWgLkbK276zpOxP0qPKd/0Sn382e
LvNaBBCLti9PMAxwlRWLTpOHEdqGtPbpSJL0uBpRLeCWd1LRNKlRx8k541uLxHfi
R8XRavR/eWOZF4LxgsDDyaod/KPdoxzuNNF8s4Nc0cGa5dCmoDxLQxgP/R85oKC8
7n8Q/9Ye1BRPShJZp9rBVHy+UitWIuxnpiVAuxSJwB1am91Zc0ruFz8N5x/AWrie
xAMREuRfyLmASKFQiv4i2NrSICgTcMAwIze0Sty7xXniRW+R/fZ97NOtGznDMM2a
UfShH+rIy91N66xhu8rZQSmSoWEIruhemhAsPLrk+wYokRUF7fK2ZgdnMEd5efWn
O/TSB+rJvEnoFKsbD8ZIXJIyqg81/Gz5k4gasqDQZGsCmv453RjHJKH1vo4m7Qe/
BhRJoK8MnMHMnUpnngRQRZ80tR38R/ZhN/XS/7nlg1R7+ICtx8dQXY04hEhtGYMb
V5g/NTCzaofbXoGBfRQxtZ5bCBcC5xKmsjIYees0tY64E9eKKVrsJwjLG1UYmeoH
pEtAPY8o1YSprbf3umP0ws+cITuRPsOUVfTE27EiAyyXRnzOY8QszbYHVsL3G69r
m99O/a7X+YC6qJ+S8B2D6VoAuIKVewzJCEmuZ5S9bBPEea1Rv7E5guU19wIEEAX5
JZjFEni4zuUfYzZo5Y+qvCqB9DA9/3VTVaN46MmaAcSLwXHv3DVjyGffvaSFlMFo
CJCwZeNeOybixChlPTEoFltvLWeTo+Lu6vDPZR2HcJ76k2PY5nPHTRuf4vWjNbhv
9pwy7rbtEkCVOKahw0p0osg1Wk3VNV/FfwK2UnMAsSBoVcJKNe+ZrdFHPOXC2h4z
UsVtin9qUqb3DWEc0WM5HrHM62zQvWayeAXPdnE6vKkdNBQw2IUi8j2aa79IVpj4
SKnQswLgOGKWmq+84pIpkpmDAhx3hufAYsR0bEUS4kmTioXt2veItH8PIGIQRpv/
68mhOXU2Bu2s5wUqsw7fFNMNg/lBP4/YKtgAasM3cpSZF36GrtiBVs3E7ga/yGYY
FnWY4jOQ+pxxxBdJPkvbsjS9kdcyWfY91Bu+AO//ZktnxFul4Lyusw+UOmmQVgtQ
KIV9Bi2tb1Rs3+Z7pxqPneqNQs/nKzsvKVjzwtocafuIjjoratIt1X5xMfucnZ7a
T9aUddYxCTvUAXkn+YQr2+rorkj+rTmfgaalUDrVIBZHFpKHvzoEjr9lJDyp/eAc
6ImlL0r8t/G9XPm4XbMxNa0W9bhCzPKC1VWrlTY46a3/yYyWgFhppUb8/DF4wEZd
FW0WAywW6LXenf7Y+0+keWtEz8Qx8tc5g2GeYW/+ZpgaP8t/u+HlMWu8xmZMT7An
bBnfZ2Kwk0HrDtwm53DQX7Lv6VyQzQAIefa7rufCuveUBGokpleT1fNIVDvtD9qB
rBlH4DHXkCLy9kUep0gnTCGCt7lNo3bFzmiCgaCXpXPWeKlJTg4g+qd9R2q5evFj
0EkVZFoXsorLznIVFR3TrkcwQuzNWyddtFdD6kQao/UKXSp0aKEnugq5GgpRnJfO
RrK215Y90h2vsBa77713rIKECN29x/PJgePaovdbBdmo1mFIwlyiveTNjlDhmI/s
+zd+ho1xmUW281CtQ8U/Quf8h9KQsvw5UljLctpSXZc4Vv4VMhfy6PZ2if/fzFFL
Cya9qGLCseWt4qD5vr1ce28ndwTZ7g8+pXyF3XEKZtSsy7x27IPMo5Bnci0GQeBa
iPyO7/adCG20EV/AHuJ3JeipeGorX+9AhO62z7/Id8+SNIGfIOYdAh+yAsVdyLwt
wLAbPxjMYMYhpvKx9f8/7NrxhJM9DU0Bvqk3O7WIxJBOMnYpnK8EipZWu8QxhSI1
SasZZ7KJPqYvm+4AUJbLtZWoKzz50vDaM23a/X3PYCSHxaSWK41RREd1aqWozGgo
Ey/KfSG/+Ru18ZNqOsau0KqiZNcbGAvGGdKtOs0UToGDmAqaF54YvGQf1I3ogbj0
7s4mPeSnNGb+WaAwQltnlWhM43/Xa9L5r9nlVxN3vf5xXp+5ATccr0pK3B79GJ8K
hpdpM2jJPYPqqY/8y2kFLo9OAVT40Kgxz3f9bXnX6+tsA2BjnstsZqfeqfrVbR+J
Zlhst+3qPqwq7PzDNC9U4/bRAT1fRo0fZFcvL1/rewFDXgHyHlH6b9rT8/pCJRyc
qny2T17p0u0CPuer1suKaC9dry5HSWHp4TWWB97fg2OKlo/txVM+hB0rtEQEN9Fu
14kjYgwqNZcwkUQB4kuYmjUsjY5ZOdWA45y3D/2B+jjNvJ5T4cFuplw6Bykg0We7
Z4G60PBZMGB1XBbbUrCDbZgfC91EpnjXfeObNEdyGWeHz1TcpKvgU5yuKnoHjI7Z
ClVvJz3qyBA/8PMOogUM0NL9184AaXOWNb6HFZ1W4gOZm9MPnDrcg3zdJz11G7c5
X854hKHCuOJ6IOvhYAiTimFgQpdYSuLWseaIHP0S/u6A4cv0pr2no0dtZ8SgBx4m
f7sH0NmsuKjOq8MrbY9jK2ucxMnAaz69ctv3Ms9L6TWaNua1rCNhyC5LV/yGumE/
nhQvRws499O6c9fLUzrI9in45QhQ/hdRvg7FGkhNNJ0HGWumfHhpKgv1bFVTuiGv
AUFADfS6xAEZT2SFDn15jC/hkL97TMuDArOeCPoLQpU3z7TEzxKMWjNu8rwyjH9S
yTE1e1IxZtTCFDp2Soci/GASepmuRfv2skzRgoKVmb8jyim8QI+oHnxT7h4BuQVg
ac4cUsHQu3Zudtaeqcih4YoY+4edty8B644PFNdYU2furkX+DcCa81r18u+UmbW+
Uc0ptcWYX4J07Jequw3NxRv3Gd+v3k8i3EPNIiMvm14yiIPkSoOB9l9AjGDwoNMY
+5NxJe0RzTv2BkFfnd8DKYS+U4NfvZSOkzBmpGUYW6K5Y69PDFvMqLuxajFPe8t+
+VU6tvyB2rI/3h9VlQNmzoD/cK9D+iVctPFYDC+Ix7Uss20ynH1TIxzPLS1Y64UZ
pvpQIjL69XaRgNhkmI8l84Q7aAGJcluY7IaKtkFwCVA9oywpIIIoUmZs9GswbsXw
aaEtZ3kATEmLTpjQWSYolcqpIiqCvc/DfN7iGebP679zIUIPvQmzq+/UOY5loB/V
PGUBuwuGRW5zi3O4u4ItY0PWtbyFueG8kYTXddMGubR0UfUO762SlgDtTu+bc4L1
NhrwCHGY6NpG638FhwzahByBOHwUkJkDpHiMNAPRl+pKD6df2L6WCKo3GPfB0UmV
NUfEQDNbQdNoEHXs9Im1/BmCfCoNDnZskmPcz1d1fXOesIsfV4mf6EVENrx1qdaB
/lwqWxPo3eZkkyq4PNOV66ub1pPjsc1PTB/RDy60q7ocy/ajSUDP7pFv0Gry+EbL
qCBSddriRIE1V+UBPxLA1i4EJ2k6P6XpTaTcFBIxGlj38jrtXuaTPNV9GYtICkLM
eouw2kjy9hXFM/goVgurDKai41HOOXYbCoTKwiqD6JagueCypm++Pl8x1P8YdVzO
O7ojZhDzzn4S3OONUsTOdsNM+hhGDTSMAu5mM+T/v7Huz+30jDJJCndwBQqMa9jm
Vu4VRVyzPkV/JyPSSozgDj2OsTH+U1cnAgKES+jMHhNGkwfKd4ntnmxCg+MYVhdz
MLQbDL120MxCh05mfRlJVX/ZQCe1bfZy8AecQnqRP38Ndf8Dv8ym8L2CMS1qH06P
KoPcgj+CMy3MNQzKQqPrBLDRYr7QT3t4nAngzftgh9NYvTq0l4gYZJjrbTRDaXbU
KybJOzDPV7nK32o/xTxod+GX/+HPHr7TWVzP6MyFkIuIbzMIh0WzQmwJf+KErV50
LCo4kwACBGbYsSnci1E/RHs/WlyhsKGHyHnIfwY5+UETfmSZB0qDbsdmBhjNZo01
uTB2JNmMW0Ywvg/AVtjsDV9jX9wYxvM1t9/ts3mZNVWuamNr60yn1GCEkV29p535
YxUkmtuSSct0SLZJrFrr+7LvecsQxUJ5GAxX0MN47EA+I0+P8TnnudJnAO6BVQEd
InnDwLFod1DXBkpXq8lKgPqEZS9p0bQsppjvV+HTJEsNlhYsYYT5h8fTAO4kqcdN
VJboxmvQ6z6lbcErDKZIWmSdueFxy3OH1niN89Fesk7fPEuzKecIcujPVj5xwffK
Dcnl6uFs+jN/SduYmlemfI18G2yGbxMn5RYSWAbHl30F0qALDH+X5ihHjEqEp21G
cVskFEGAdKBAmAlsvyDkauk2ud+1s/K2BG7a4XDXZ6SUzNzNYV7CdFt0tcECNj9e
uwxfH3o8v/ZIy5yKAz6h7YZYrnogIv0z3yZlMrP0dQ5vfL2kvqV4SC1cDakH3XWk
6FqY+MVx0bmRezR2p0CPFYvhp9JPOkwuNrtL9p6m5sYfceSgxlBb5adkosprcYYL
uzEou9sN6R/fDmFuZl8Cde4Nuy4GGeDXE42BG6LWMLAxKzYYJbO9nKvdegytazwN
7Wfqtbg427Qvg6BfJG8HZtxsVCc4v8gVHE1EMLgJBmBFRrxpmQwsJRxo3mJJMf0g
TVeAKnmHinFKPqCUKi+sQMSZOASKG7/BfKw9k/6QgYAl3jBfCWc0pcIzR0RhA9PQ
DpWKpVV9TutdXi942b+kQFeVBic0oKFCoAZvzsdPkpje0bvC1Ff6N4MJiN36K1eZ
r5DMwNEQYNNH7LZwO6ktr8UOhZoNuJtuEpM28dQxq4pvHUdVxP1dM8Ojar2vstG+
Xy4NotKPOi3kYsaH3tWqrld78fJ49erG42bIz2vsjYepzjdBAXin2fWzu1VwyHAJ
W064TWv/BdcDJzqqBZAW/HxYAAM9eDUqqQ/DMmFST3j2gQKxQ5sRc9lhuaoGHkiC
5qdnmi16kKkf1py7eVAH/upDhHzIwi0FRavVi+Pg7LrQ2+7DpLeXN1e+MchfdfEA
Yu+RMlBDAtdwoSaBwLfOctr2o1I9WZErBfThGfUILHj5GsKrjiQcTdfqVy08KlTH
LEfCX1y2kkR6YMssQHf0pRrmrTgvCv7PXEYDRZ1wK1XTAQXTWhGaebGv0hPnzgT/
xkrDN0M13OzsB2rqwyIVh8R651n74uaY22xuWyKvSxGWTzjzI9/kQBuqK92Uwh0x
slZHpgGzxebq0m4K2woM4ookC11PEfDOngw2jfFJjFvzA0pbQTbIrSJOMqE8jTW+
GJXyvWJemUKHYNfGQDHnx8s8UEhYywmXsYegEOUwqw8MkDK4kz3MQU+sLfv7Vty9
YchDxv3fvY2O0doJcgtFCi3HcvzhDAgZ3CPOXWEkZgbRjPzqKebaZshNPqC+7+/R
gHWgUfoYgIzGqm5svLmHGAItnYoLKxU7mAUv+b/fXfNH+ozSjVuhw7hpjG9iSQsh
2EAUWqqxKSt+JXKg6SH1LULZ705NWoA/0ADeDdVn1Msy+vBGYnfPEZKWni/WbOrw
DgoPFC1rG4jzZnybk42L/CE8T5sSb1f1KDOJPgcGapa1FBHaSSgBA2+/lL/li2lz
FsOyIDUkp1K30D4aQJZOFz8nGlG3y1b4ju5mJkZLEhvdwdE/0z/nuTilG0wLvep6
5uJZ3TJQiMibi9OcfnWr9PtJDU0e2kvYEtrIDR+UIzATGGfswyhv4ycHrK9AkV3k
v7OwoMYipNljgNmuLw8QJcWLsi2cHUigfEu0GHp8yk0DQJP0/9uxoHGgNSf8O8a2
Qg4tOwEqNY30NPxCTmcC3WWqdkGivNLXuzAe1hl4MFYdCmcXkMRyfc9haTztC1v7
JpjNriq0B8pUv34ucHQE4XNOhojK/Qh/M/7uEjfq4cse512mcU1Ozf0f5uMxQE4h
5pmJWhB5WrF9i+0mj8icLvsO8ZcTpGqt8ZbDd45ekyaydP9dYUgJsKkTEe8AXVkP
Uwlrir4jkuT/g9/fBWtIYi8q8DtEEyoeEz8J0hI9nMlens9owp45N9KSty9/2gJn
YUfK4CLrZEt+QeVMGGsa+dbRZ6WSjnHofIS/dqxYQrkAxDp4d6fLl9P+zcLZuFTD
KfKVdhVEC+NLexQJwzAkbJaRS7RbyJbrGiJWvataxodmVvSNMcfGuodJSs7xpGsb
eJh9/mbLMtVdsOVkFXBY7Ijkgl2TEkyZYkU40IlASaFpKG/r5qtx9XhuhWQq0yj8
/3s/5laFJr798lX8yM+QFH+y83uJqdq7c7bBnvCnk1K072edzh8BweQhsjxWiPsd
P93LJE2DZiC9L4xMD916pKK88krPpJuaACN4WrXTTlxug2UCbForZMqf4kOgfh3m
fGeSjLY2ocw9uEQ1xJkPR0K9jVXHElmMd95X1l7BexNtM6PMeXQyVo8bTaGC5X9K
PO135OYPeGmYtPqXpTAGveVsqkvPEuSwaON9BrUrTDiQhHZVmT8R/BKhwx50vWCI
yL4iLbOodSl+Q6RFO273SfRbaTc53NAcf3+TFjQb5QHLpU5DvBANQ+kZmmtDrI+H
yqIrpbOgnTQqrTu3+8vpzM0sd2/Plee//OzGuLLPh9C2CikfQXNSiT3BGH2V/JSp
yKfx5/AryrFvCMvSZ67StBWCnfMn200XcWwDS4MW4JAKLqijh9tWqsqgByEfI944
bNN92F9jVGJdMfz+3WfCqRPNiESKIYtCbYCjlKDQeo5rWVBE4laEmo2RQaMfnce0
wSegyXzDQ2HRjQCeHf0nDiKbDySWtp/JHVjh2pHLnf7Nymjgth5wPSh3ME/6crR5
M7hBWtbArtCGudMoCbFcsJQxSHhKV12T/JJKTsMnRPF8LV3O78MAPeizljPOARwr
ki8++5RKJ55Oi6/uv7wE4kL+EyRrQ0SB191OPWSXVZm2Iw4rbD4f0OzpdYz7jyn4
I4uadphTDMpF0EpeBrPdg5OEnwVibi2hXAycAg6y4Zot64xux/9g0dv0MBeRyZiM
S5Es5dkF/D9K5G9TCpeodiwEwxEwAuwIOuZfXte7aMnERLZAWC7W+boKGgAEgkxw
lIvG/MDPBU6ZRaC+OqnK2EeaeXDlfTOJEGOdLvCIlfio3EMnWr1kTknH0ijUTeXQ
5yeqMEsc1/CeDp6+65BHJ+RbaaweZWDIUa5Yi7fqqY/TaI6uGBZ+PZo6Fd2YKKdm
647jVOW7SZKR00JNvdNwg/UX8C/K2bHAPN3rqZQjKLISknHOE9JSl2JkLSMXJdc9
kFZxeCy0c04ur3X6DpCl0EmEZKDl0pgkQjj01yW17wbxr8bLAAMev27+lSZRohvn
H1lToAFwDAyds0XlvzQVEh3h5R3ZJ1g6FMlqYGGZH0kOcSqqPdaKmfXCAgOagiJx
540+vA8P0vuhuJ4DrXzdP4h/z7IZgxJoCz3R+DERG79TOsvPsOiWJceSvA5ECk/L
Ye59A/B19K0x1I0gEEpSyHSMzUgDVFNUM8DZ66iWFRA+NvhJ6MtK9uwrUv9oTW/i
zpLFA7txao3K+GnGezPR06Cw8JpgvE7t/aSNPjU3nv44zBMm5GPtdQaQtvSlOkkx
lSx1mN7E9Ck/OepxEv5tJKccdzwfxAmDhN6qADfdAz0VLZLE8/A7TsmK0D/JiDDD
qik7S4MjwzTaKRGaq+FD1rKNgHxmlP6R7ft8jUO7rXieC7nuA6HH4nneRfhmwjjh
t9re/PXhD7eKHX9q/bEzc9wx7f/QM7fgiNbvk3PWSdpKaIkJMWgA6Jyqd7XSd2yY
2pjc6N1hu2OJaU4RaEhu4JdHVOz9MCWE9BX5EQ1aOJ2npeoDRTZB7oxtje5r/RHi
htr9JXeFDtLwut0COFrITPXpZ5If8WCtxF791P2LsMC6OOBAEK/yR9faps5MsiFV
CDLX7LoUsXOgNwCawu97ugYQaWBgDKbVExAX9yXMKzleonaxFmqCe34ga4K1M6XC
o0RlDF/VaRAeJnMCIbrGSopvC2TI+0ukLUVoa4gLqFssA34tChRVgkWVn983vLIw
h4HvuO35Juq9Sd9ci3lki3tV8qrXTNKQYeYFcEMm7cd1difuIWhAvIvbNYv7KyZV
+3zG0yFR8lkQBqH/JRn28IU28fXmwd0PRPVUoGaUPPneVMHSL7XTY712rJ7+EQl2
hk1pHygRzyZd0T/sl5qhIaJStK+FiK2DhDWBG2eIuhcKPd8kheUCn1fFGVypbxaM
fYuC0r/+rGaRK5BshtyrxBcwOmOyIpkO/1w8vR2pGwmDQquK44vw9dpd3oWmfxHV
nXiJw24WRLsPgzQZwkzmHM+R0fZ6OYWu5kodaeLUvZpEV1h66DRQHjKEZmtDARrC
eDyRpVz2ris6bhskXFSBV+fE5JAF2laRvKIpwQitIuymenwqsH7aQ7D+KYKYR4xl
UzIlgfOUC8U7QVAs0TN3LISWWS1jVhU6ZG+PDe4AkbXPfxdH/+f0k7UKwp4V+L87
R0Q3totxHOxCY83lqG5WSLOelC6qpp0jWY1t+gciZkvX3l1FL0FhYzzs6Xn9K6bS
tfelz14KjzcEvDmBwxAczoeM4lsny1Ud+z0YaqlQi0nuVKnlbmG6Qsh5bDraj7oK
FairO7CpLYxTNJ51QhzEsL/tkDk+L+JAWg8BgGVmRzQ4buC0N228KJKOoApBC4zm
Pocvr6Q+XEz82lFxNGekVDrF1bp5Hcn7TaF73sZUxkIHPGdEa5Insh4J9EdO6Jh2
kS4x/clEUTD56AuPENs5TirkBEd/TxRcI7FZRylgx5gzMIzMZzJvyi2fMJCtoEO9
BwjBW1DuCvFRZa1fpeYHTcZIPOvUEh03gVT2jEWWlzCWGpzRvd6/RLfqaB9GUySX
02PHneoF5FNb3UpCUQcDSFyde5o/MrCiT7WvE8HUTq3Rg7DlDHzqBVBAZ00qAYLu
mIrak2WgSKpq+8FpnbJhyw/c3Nbj6K3DcUVJkDqbsQ+Lx7yVvGgVUz+CwT+TQs2p
FAzpxNEaK5VhL2Kv3xESwplzIjJkdEbmjG9zHEO9di5oBWpZf9MC41csA8E6OylL
S0uFUKzRBtihwXDdC7cU3W+J0B4uzIluveU45hkyvi2CThjgkhBZKaO/8DGEzv4D
2eJlcPUjQ/eXDEy0gxCDAP8xavJer3qBkF2dvDHZh/UliIC9UEODtzdu4vjiSjtP
ViEk6OrD/B4zeqGJv7yUfqzYZ/6J0pjT3dcxwvmKE/8Kd0Ze946zdBCmKYbljAkK
Cad4IHvhFpv3qo6C58Kb4LmV2KSWU+Aa/NXJFV5KUPggK8daEi3IAmASM7K3hKOR
qqZAMFxHmDcN2LhpdPZLK1lria/LOfXC1rZi+pJXRty0Wt+eCFxaLfi3YvZldWcb
GNKugsxSd56/ok0DhoaCPyp/DiAportS1K3V8lYBH1kX11h8264qxV0QRfbbWblH
PgePI74kBsc7/X6UA3l+v1bdUc0pcu5hID+aUCJb5M2Aae5Q5hget7yFA3ymnO01
yVZ2v20mZDTjw+uFvwOcixs1xpQJPYzOrLg/90919DXx/bw0J4XR9MZTYgtOBh1x
iEu1X6bDcpaBdimrzIEENaxCF9KfCvV8W8XGGgQj2qO9XLbTAo/XbPQOqxOhCEy7
SesLJZqSLYDxdzux0um/roUi1RyrWsC6oYNNebA60EA9Tq/hW7gHvwWsY/Njt1ue
OEZYIzajqvg24CPog6gbgRvhgI9cRSMgZUXaAXa90pNcpiOjJiQ6GMrpfvn5xm81
3EHEpvGRGAVWDAjUTrljdIJyw+NbBtZpWqDc/pbQ8bngwNfQxpLmWalgCv2MsMse
qRNtbh008o7Hvdc0VH8x0g8nivm6CyKth41RwrKKTKIhGvFmyg+ENZQ+RnuCKitG
g4dN/SpfTBISllZROo9d+VAb07ggCd8WudDrkfDNres3LXAaHuO8wlkAToU5eBB9
W4Z3WxrUecwJGIJQNDjs16SSRJeD5ErvqdzpuKU5vTJ6YcFTcik+nAuQ+X4Jd+Mt
NigV8EEXF2sUSqyL2BTDCD5UllruBM2EFz4LgU1FnPGeE/6m5ez1/ZDDcbptb3Gr
pGaHVZh5VO6ggeCoRVG9TGe7jBpKYEKt21bSJ5YTmf2FDub8+OZdIOY+Wixem669
jzhOchKfRnF30IUKtCWwHoCgBzG9yPYIy4D/H+ld6St2NBWgaVrVUlYSgx00VxWA
DfJ7ScOy332BjkCJFRGQkPD+KouiwuOQTNwtGFU8dpYoROVsrDPHKOnyXgLITnd+
viFjX5BPB3XXswxcMfGB9zDv5zSVt1FvYYz9dpKH8aUwZX1XVZY4Kk+/+kD5mVUS
5W0/qGDq9073gnJVjeoYwPorxv0ZDHX5xCdVfchDNqfqLY8u2aONjxDzh14/ODs8
mbptrTq/Awkiw5uTA1MYho9hYWD8nsQkSEAfnIy0IGZrJ3s1+p/TNwauGgiHYcG/
g7WxCqEVr48qZXmywyXN5yuJMX7Yi0Bq+gp/vZnYaIBVHoxFlqnhb3t5VDrATxw3
Fr1+U6TGRBUn2BmDEPr27aFycUr0eFYPdXPBjll8hU7PeSbFC7IxCy25fzcSvrpW
gqX9wfPrzq3/ZO2qOuY+6jnkRz6XlLmJTq4ejqBdNaHxI0YYL3j/nsP/CxNNMHgE
dM3EJpaAH9UVZwbpnFFfiokiaD24LNBp3QNLtagTnp1hLKO6E1pZxGih6rwo8NdC
4MomNzFosyvsWHk1Smyf3u0MGHSKSY1B9+udtcgw/RCbEBVsrsmhenxXnGNTgEmc
+e6CV8RSoohI1/dcmXWdQJyDSHnEAJErsE0hZqWBEYr2MeN2cLl7vKGgeFFoy5OH
Z7jNLXYpRlBh0ZchJ+Pn4KGEWFXDb/dzaEkEKM6yjQ/pZEVgCT6yd+9bnk6l/ZOg
jYVhtO/lJlzT9hXqOkOm7hfpkY+ANbr5/O8jvXSCQ4vugJIWKm4N1VSpTjWcnkKF
/ar7ItdUbEQCkCXV9+9EZOpmKvvhLkSp0WRTLpmy2RNWtHyCsnTj5cZJDPi9HgUq
9rtwSV4u4zpCXyP8XPPa2g+bDMRHMDG2OBL2oNNtU7nrpkXhrr0YVbfXNZmbPbU9
c2OapbieKQeNECHWOiN9njgbz2kvfUqagO3xaZHIzlE33PllRKS2yPzmJPApSc+/
vcV+ifzf0l6a97MOdaI/BbeAZ08MKfr8BUnEJ22sNofWJ0kGiE4TrjDvRnDCB+KV
G/R3WhAtPK4q6W1R32XBEXZqDLNEao5Fc44LAdz71leM4lt7E1cKsZ1CszpaYBsP
OS5oBGruYeKqy8mN/3CRjcZA92qAeEJeeibdW5t4CE2zbmDqlTvFPpzjj4V2S72b
07sm8Sb1RtApEjAtfnACgn0AJbLZ+TpXnj/aF9ISVEDQoO/bbb65OlRTRl5bY0+2
hNDrL4y/EoSvrJrlaPot3fnUXfgXZA6dvCn3cM/wrZboy8aMT+3de96k8u6F+Q6n
trJe8DrhJ4NQsiYvjkLtlHisco0+vcmNQnCsE3U7b4mbZyW/HtNtdq7YToGVX37M
qZfLoFYYkcZDxPDI7lWsL2NXcheeMgnvMNi/CkaA29W7qVALZMpYc0Qzpy9JNzuo
YQ5n5Ygi04On13EhVxDaxQS1BYNlrRFpTPu1pi7eJ05hbomSbUgipmOGM9KiEZbO
NxRzGAptKOUruUVdmp+0Pq1jhj6O9ltV0A8lc9l9r7pPleSL5NwQ/6U5fGHXXXRN
dLOHlzf/AD2wz9wOw4pNC5xhzkTjKFe8sB+3vbREvRMIl/Zn6F2+Y5oyuVC1vjYI
M2i4VDXNeenPIzmF5sOO/v0bOSTbmHGfbkbsFDJXdELVFLdUKsrOQfDCVCk1qs6U
75Q0JX9obdzLP7OSfKOgZ/kPzVnULY6jUigGIJR0ML7weEYKWg0JJJ1zZ8KUOZZK
6J4ezIt0XPde6QNjp2ZX5NOU2T2sdnVNuN6NFy2T3FLHDkFW3kh/dLJoEP5xHrtg
y7U7KvJVAyDiJyBHlh/pU72VoKnNH5IZ33nTv7Ql7ZkMpDAl/PxTQq8XWWTvQuaX
16kvIXCS31dwDKhi1Xql99fUAZ40C8n7jN4Jy6oUuDoU41JcC9Z9r/eVCaVZnEaZ
VsIxPx7VMULr0R/RGvARB6HJ5aF+Y/VQ5jbtlFJr0msHIXxK3L1nSqKD1bjNLoEW
04W3BtIgsp4XWzmZG/1PszyQ+oNf4LN5sjScT8Gh/CuLhXXLncjA6CCLqaCHPwSj
RKSb6rnLsn175+mK4t0vqJ2tGTMS9z38itZ69FtPODyDHIjMdEDJhFjHfntj7mGb
HaYk+MvKp6yaR9TTu/qHGmVhYc9gyzEGiPt7iL5taPo12pPigdDflF02itQbj2Ee
vFr7JOuGeW6I5aIvIZxnAe39wfYvXJe6F14QJNwLURaxx2oSE7+Qst7a9BBcmGrj
Uw/80kjYbqC4B/9jHkNtuQDzxNxA31ont5LhqVWdmklqm/BUAY14A+WulMlC0rDw
2lbchQZlTZGmL9KjM5pZUJpCXpnOWCAmjVJH9UR/hBTRJFcIzKLr3EndSNrE8w3G
0VOLO+29j71GMvkvl5z6bPQTazwnq29BRnKx7o6KifZucWskmHZXBv/P1SoWGZEZ
iYjRIHOv0LQMSQqoEg7C5LZ/zFtWRL2HqdnfPvbPbX9eUPAeWGvjsliRBq/qOY+M
w4ho+VBjqeWlsgrG28JRkconQtRHSvh5F1AaDxv+ZnkE/zBPw6tgnbVFe0tJcRo5
WtupmCZegAjgcUZnJNP7N0GT/hEXoeO2wMD09vprfHy2Z2NTY0wf2IKaao9rcfCT
W63yfWidJFgb/+T9WVfTOAtd3Obo7LsjYaOSBkoEu7XbU9+OVAQUEDiW2AIHMtNo
KWy73jOFkcutE64rOrFbo1ciLhm62DKcawf7oEqlbQod13rRtBqq45jwGRQg43+n
MTc8AmPpZY8mC8N4DgRkNejoaIHk+law5iKr0gTqL1rZCxMKg3jEaFfMsHrH/Z+7
wYIA1yFmL03+ZsDpjonnSXsLDwuLJdypLlFMJOJIk4UOLmEiwpc9CepjCwv2vkYJ
bXTeVAn52MUPJFMkm7CBkBZJ9SRH7xK1o11wzm8PSZuBr0/f2etgw77EX0xTfa0s
nFxIf2KcegWARS1tZNOSpqcq53eqco8wf1FP7APpm+v6iiDJ3SbB6IoUkQ7yqiDC
i34MJ54Zo//YwqUZNiC7I+u7aZAbXFp7OMydimv7V/ytQCX7kAmKmQmM81crjzlF
zCR4m74qAMABig42UhZ/s0G40w9zd0uGz33RHbUxyEm/JLMJz398Myc3FSYAyThe
wV+rVUzafRxpHs2BRvAor6+wYqy72InmhsRdoBpzcsDTCYgRFnZUc/wybMsTylD8
lQ28hQHeUloZW3o4dfmkUoFfxo3gamoLdypHQX2Jg0bJfbhFxWLiD+gbBCfRRnl/
Doey9DzyOXrkMY0jbG1WeE1oNo/6kWE1ovxx5jRsLs61LVRJXj3XgBpZZxyntfGi
w38bPCS6eBAFwb8cnszF0lMyq86jnuKQdg3F4VtAd25jHw+RRERfQc3gcg5/BOeJ
JY/OPAZaT4Nur6DX4w6o4SOPkOVbm0dH59QByxv7v3gtTP9vZN4n91OjeeEpRuzW
fw62Jm7BzeY5ljhq6hDa5K/1Tw2l9hlMc7kzi9KmYXIaHkyHrjyiT69/oKDwlJss
WBSmRtikO/vW7nEuJ5bMJ55hRVbdJJzYcO59kcgNzDa+wxkC2rf0+D3joUKzOD24
O7ayZ209cDE6hrJ93U3695CxZ6wpuYAGbedu93ip+Cdj+N3cQimHsqBqfeXv/C43
B0nJP436KxS22/skuw+L4q9ieIFSL2lwreOUqobThLTsS8jD9Yi5S33kiWWbDOTq
OVJqwwm6T7haXiUK38ZY8jBzLGMSd0HNow7OJ+Kp0hC2RgtOHyuonpkMUgIl15rU
44VUsZvD1RuTLMyC5EkoCEg07iU+iaeOGGYDTWkWztY5lOfWgr8+sWyMKlccPUNg
ufsTPTfg8QPkdbwivrp/Sn3KNAGb0KxTXnGVEqGMO6gs6rsjGD2ULTBF9El+dZwp
Z+BUGRb4s7AWysKIfxRtIHK0MQiYJj7HiFNapUKZyHRvhqyZH5Q+GdjB4I5OrWC+
Iv9ZQpVtDKNLnPL9XOthKeNvRjW/m1OKycgP+lO/cDGL8/OLQhEKt+Le8DFQZGgN
iW6eg2O+fGabFlLpeZkjNBDnxAWQ4djS6xcWERrPFwZ2+9ATL9E75t7JQbswUQYy
2I8NzF7/3en5TNOogpehSO4mJBbl+KoMFmEaaf48POEgHcXhYaCo4/ujiGcRhlIa
EAplyC7OjDe+OvKWJ4j8+tGRSXJt5V2qY1rlR3IcUSsglQ1ZmulgTWnkJ2BnPdc/
C58Nd3uXzCZnsszFA7utrZ+fnsBV7OESxeFNhcnKsePHpSHV9Fhk3BsbTGW6m0pw
ex8SsWB/olH4/NGmSBCWou3XPHHP4avKUrAv4+SNoOuQGG9buHlYF7oB3fFzicb3
RsGPWSINe+zq5/YCQb8KUmS+lMFLhoOf4p7PRTDctuaPTmmWFiGR+7OWJRv57m+b
0+/vD0gGjyeGQ/rENNMdli7WOv4U16Z5enzRWzVQ6gVEM2+XGmIEn8R7qe7wJVR5
9DNMwoeWdu9Shov6vzQgluUpQPrw8QuZrY6nRiH/e8wn7Zgtkh+W25vhf5HaUhIw
a/Wf2ATFsnfyxx1Qbx1oUIEY0SJL/Bg4afamRKlQRAGz0wM1PoLvewIRLIRTGsDn
KlKZDszg6EkQwyv5oaRcQB6g3RJd+ueTgeUfc8XTxYTVsVBWFtWzbT1aUNVJkKKo
j2OlFVTGHShO/01gC3zOOrn4cvBdSSAi45rFfwwOa55tTdineSyT8JcROsImyZ3n
Ry3WnednVCkKRiY2I+Gd4H8dvzWDfkCiDd7AGVjXgEkfTWLKS/RPJwflOjel17Zl
Q6avUOXN9z3Y44l5UA0wY541mHFY8arINihcvmxpkyBRvDm7NHUu5XiyC+62wabI
ztBmhf0k1lkXV3xbppF2Pw7LZ1Jfr1opZs/yEGZSTJ8mgx0AWIy1F4fsKrAaHH76
sZrLdZWrVlHcPwcynlV7OCy42sZJOMkwOhZEfAlGtuk1t6zrMMBCcSq3fZ+IV3D+
s+r2fs2Rc3bqM5v1cgrcIvdhFLdWOfH2kZ87cQ5CSYSCBPVcYRl0HpaKt7DRHvxW
CdzJgjSdgRW+Z3k/kRtNGCQZp/qv57cHGnSMT5JwZ5Ij2+MwER4Xa7TBPJlJk8mZ
W7qjUuRCX+os4lYQUgIex8dwBQMTHRbL4OubupvB+msyXPCQt3z84XRmcCwSURSj
3fa0FJYxNl4Zp8d/Qo3sVEWU2eIXMAFXzqK4RH2FIicRspwAAPGcxXJlmaOs5uEH
9Xl4Zz8nBUByXgFEfaY22TJvZZ7rtC4mGqRpNLfeah2HGe1ynxRr34tIvI7y+RIU
lFgJW9gNFnnox8D1srENrX4JKcRB744hIKnqBpauuZrR455j79kWe99J6JRI6K1q
G0ZibC+E+bO7mCfWjjqfGrGv93WS69iT8Z7Es9Om17AScs9GoZ+RywYDLOHPaReQ
k9dFa+an0VCY4M0i2UgHHfmlVmQvwWYjzV4AGvJEUkFfCGwsSy36HbzT95cAEjot
UuhWiyeSB00YNclB6maWM5HJe8N+8ilcPihmchgWRYi8S4lQv3d7aJkTzRzbbV0G
Y2HjRYiBf9lKy6tQYTQIWBQpLiXdVptub1itMjjsIpGbpZMaAZJzhToehrGIC6W4
MNRUWD68POLGS8QMELwcFIHvGEJWMlo+p4q0N2RR+AyhHl6z6PNMfJkwSxmSNUjJ
z8LHHQpgCds1Iu7Eekk0Uj3vkkn1d24Qq9NF9ZdZr/JHZtZRrhb0KHadmCdPU0zV
70CBH3g0q5JKukhEL/JSh4qqjGWJOjAc1gy6qov01ogZw1PhuGtbXYnvH4x83+5+
IjVnB0zddWZpY6yk573KWwlDS3CaVY1/5UelSK8fXJK7aGc7zg9gLeDdU6S82TVm
vY+kbIivObNvZfHpQsQIPRobAkKSziSU6jNDAnmxTbtnGoo3z9gFj02wO20qjm0D
Dz5nk8k5u3gdTSLJIKmf3dYV+sr8YJ9a7hVkHIpi4SJuJtSgryFZEgDOjBGv0xSI
ahf6RcnpDEALoFuhzn+2IOp/oBmSEdpuo+GMx4iP2kfnkBt2GiZE8LcD0fZFqTaB
yTT7kUI5DwwexQ9u4MnvUcSveWvpMye46rJsnJqeQPqKRioUI8aas9U901vsDtDD
dYJ2JS9KuigfIH63ThjCb9wqdIQGt71RIgn8VceoIOdqj1wVGIbM9ZpZIQLCVzzp
WPqzEue1LIc9R+diz/mC5CauUtpwu7voTjM9iVrAlBo1IxTNX2YGbAS++7OHe7v/
7LWGKczfAlvUSifav0r6ULdlMHWHJW5R8dzd9xs6iBUnwpUcUtNaI+L+9k1jh1n0
4hoDcj6pjJAA545RbvO/h9Wh32i/DyDZGWslR+kfT1i+cF79Lgy21VSXZBUvFE8B
RfD8uDYvK/vVeAYKp5QxW4JTz9FV4wDOGWsw9aGQHUNjjySRTPWgnzC2okoANi1/
CyI2cOqpersT2PAIVrJ8lDM5CmBoXWb9WK2DtQgqLIhU+yL8EIhH8KtPzg0q+BAU
pOLlzl2ZYPRLDcNYc0BlxAhSTSmZE0zX7RydcT24w6vNL5ryckUTZsKiYodLwZQy
VOx44mJXD3MiKcOmujouGbPH/dVo55Ko7dGK1teoQpE/OAJxY8wVfEcF5h9BXRgZ
7FsCyBhMdXFdThGt74Z1Q4NmM7RQY9zM32/5/uYIx0r9t3PB1IGkSl1ZW4Tb8x76
H1etDp3iNtTrsTaPE20MXVUvDYsZl8ZJ/xlskW4TWvbjtEaGBr3gnUdUsvMxrAal
Zdn8g3autdGu2EWrbm729jaXt3ghk5TTniLBFg6s7hI1wdemR1jrS+yMZoQ5Sekb
Ral+a8BuBKj9qMiGMmnJGoiYFZYFg4BrK6Zfp/yQa686oMBtgUaBgSRiso87mVJ7
UtY9wtfejDd1xT69JlP0chitdts4oHBWKLmFCy6bdSry4fustirELqgG6gDTTk2b
foMOBtoTlwaNtYm7IqJCLmIDQHriS0hJElfODh+HSYOk7KHBVuTJMmjzgJ8IvIOD
H0N/3qSC8ytUrboYti31EWKrp8+0nrRiaeHQXqjyQ9IFDhDR/0+Kt8yhesdDegl7
OQApLDH76YyEVVpH5Trotp+2OckGhWSurOw8yBWBdyr16FnwT8vGFfwkh2N5qF6N
bCWxsFnrJ7VVefSuWeRqX6qqpI2H/TiLx9te5mcDAcVvI5ZJDJ1dKbffdWCxt/PK
XpLl4g8r2pvCfW/lVH9TuC0BH9wo1HoPakHlVZoBZfDwlDz7vAsCUGDi0z8nI71B
aLotY6bpY90lolxMoagIEI/pfy+CjiDpSGi6xUDQyMIZgxEaEuNJabl3dUqQOtH2
+EFRsOvgacz/Mom2FIzeXyzCxExxI6vucgT5mBM8UfdH4alEKcKNnk1Ijt1mu7sh
9uGUPAC2YyRqkpusAGGQOj5ykffr8k0vLhJqx27SlfZR8FX5UytuyOnNjwx3ejCG
sJlkezfE8SWwGxudIoLXX1ivs396am3QNyfi9GpiTR9WftXIJ7zRcEqe+1u9dvFG
1EJs6DQQ6HgbEKuQgMHXN2Zw2imEy29KN/+nXaLDXD36U+JhYNCextSdePROgGJB
X5UG39yRxsedU9hLBVmuxOp6d3yhBhZO0VLBAJzVNdBzl9I0ZYq7HYeFcj0wLbOB
/E+9wsWjuBbGydEgE/4cYBzqFSAaOsaDPNOe7WTssBifhte7hgKh9ddIbDePcr4c
8s9t+ghgkBU3/Ifg4ixw6CREWGAMcfFMyviFOSuwYH3QQvon5eO3UYgLypSTHeXl
Qb1L/cmpJ9RICCTnvfF1JKKROh/+SgZTzOhY3ca5ux2gacTahAZSleyFLYkjHbBJ
HvRLAPu6cLNdJt53Mkp1xs0ji+4Ilj+uMJ5F0gP1UiPHzbmVbdkO5HZXWO0E1G70
SbHB7e1uL2bp2PtFFej1G0bN4/Erl/uKsNRroExvrcu7wCw8PfxlTWIGit4/BFba
QmTFrEQeeTeHO4KCg+/hdiCn6xR4GMp6DkFC2cZmXQlr+YN+dne4RX4CNDEHYVwo
slQnuUX7n1Uu3SXAe0y4q9EiXgFCLdrngrYs0kYdhRdZHWm4KVPl7Ymcz3r+kjxd
2PLv81JwBT8KVJT2txku3Ser5+XUJba4YxdTdqIrT5qZ40iAcMS0HpumWbO28M93
KcueZ93WJCEgUH7w1xAG8/Je7Gtm3vVwtnOUmSFsUvySxzOgB9saWQK4gdkpLaph
gUp9xqErW5Pt4DAScK3M9LrIIkDy253xWTLLhbEcQ9zfLx4DJnQNfpit7nY9r0ge
4htXZ4m7LGMelCa1AayJ5LkAjv/iC7bAAKgP8imzbcbZlsriT4FDieuRAHjBNyyH
iTNGUKRLzxtJvso9/3k6jB/6MvJbaPNcg3xH+DSXurbtUEXxtuDOBzHzZnv8ENXz
64xwso3zbWiwmqLJQoxUJvrEver0smjAoA95T2RNBxwpPIZURH0yZ/fj3/HUWhyH
fDwhxikKg4GCHkakj8jwI34d5VdKUXUHLeiG2cQL/XzMbhbacEVjvXUBzv/BGJT8
MLCXhv0dvH9a1326BNkwhw0Af63RCA3E2H9wMMUb96aXP/lzQKeDw+cnPCEZ0XGp
QTecTg3BTQFyP0+Z6UKJ7lpxnfdFTic/B6Q3HyLCxkX8MOvB1qq6l2UKYBwO3O/T
oheTk7bTQJ0zHf0FIEEjSnh20Uo3mkKVVP28Pb5s64ni/uGmtx5OOEnhenTRlf8F
HcNxh/eqUlnabwUoRAAi2R9D7w+/iXpuyRzagAUKLq7SKccKe8u9tqJtKW/UvsW/
Wn/MQr22iDmnY8hciqSqpQysHTKSXkLm8wX3MmYyODhq/6NtuV8tZHYxCEzT26c+
yKZQ0CYb3Zj/gxTn+uqz7nQd/zVUwjjrbZ6rMBJ7VnBlXao1UrH/xwtTb+cDdoVE
qvdvE/OYPGDbRIePhss1P4d3Bc/0us8NNelv7AAcLTFCSIoIV4JyPcqoWlKbfRjF
Iag7n7OMmi2O5yRkE/k7ng4OfQUcTqeY/bEeUlWXoECj6AxewQu36XIGdCn+HcU0
swpHgMlnintcr803Xu0lt1PyCennPKDWFicOnHCiftGnx+JDDTo3l+nPG8LVWkEg
3XMdumzMDxR/TyAQ1K1ljVGd1lAa3Zrj4VMWNtQBYG9flKF3lZvYyfsFMZu9o/rg
u3WFZiL9HMUPl0m5o6sv4xA6GasPgFI0IObSVni4OeMsd26k0vLDlxVUd0k8vQLl
xkZpE7motqtFcgj6RlFckvnoSMe6lnIcxGtu02i4VYpFWq+PXWZHOyJMoHoth+YZ
1y0ibMa8ioSYVvrcwPM0H9LlA7fzTKrfSiw/qL6ZlbbvEOKXJfBcKuq7rtHhLYUy
iU+mEmbq8G6BMjw2H3lcYyNGFgKypOo5NYF/ONEbtYQmlNMh7qc2FQfuqMmKeDG8
0XC/qQ7mxrYW3PRezirumBXUmZvHh4JiSkKX22xH69ATcJUNGs7ilnjKFUvcE2LQ
f6wOAz+i/NtCzivA+lgjyYDuzfTbPQERsdQOn8bBXxjb5AcZPuIFs41dqEm49l0y
iarT8N8cVELD3EfycU7hqfAy0MIWmA7sgobV4RJEC8JGb1NVVz++toc/kr7fAwsN
WnWJY+05M+im4xzrX5T7baKyBVWIGKA4WBMFDJfQLes0fcRILUFgKKhfHezan18t
RLpqO+Tn3irFDy4sAFZ9tYDaUhEUObdWn3hSxahvMo8f1stBAZQ7pKPVg7I6MkvL
QWSn4MiDSg8Frx4LBSc8wAGJ7241qLbETsKa6vMTywhs6eU9mxYF8JqQfNTXNLFF
jJBabXduxcs0WmD6UgQiHpvVg2lbBgRAZ9l9oQD4qkJtRxaokKzBY1nkPmX+6ruk
MxHLSgrY/LEc4kXZjAOGK1WSkfHYskeWnFid2e89lHJagjpBMt8BOAoRB5xbOx9g
MLfx9gpXbn8ZCuCsHDBmBEU5mhgDtEEmpROpxqVj1KcgeEZYuvsHQX48a+9aYoPi
AN3zwbOCAYMss/pO5HhzbAaWOeNXMgP8Bv7xO4f6vfadB5MWB7hsxOK7jajiSuXv
0rKUdI0eaMW9+RHC+tcrZkZDTenfzFXNXEWvlGFtN7i7hg8OlhDxX2MHsoNM/d7Q
7FCglOge/F0WdLKYOGA9ZLC5BsCNrvqVbhRn02FuGYmYbj42alXuxHIT+b8r+sHQ
0Vtp4Pi7quCeGIkYbW02cE+DbtxZG8OAG/Cl3bRFb+DoBLNwIDJYP/TZpFve82zE
05P//Nouj6GP9qRgDudv3v0kSWaQSYCCorrT9F8nt1/r4nR4RwwFRfcZ/PioGKlX
9XGb5CPz6JeEDHyKghUdEtvaTPMVT9uwOFoCQODApRq0CI21ovA3tNrf3GlXF6ev
LVP+qKhRpSTr82+wDPF9slMWTJtdM/RnRNEDrF7ZHXgtlNlBnfGNDIymKmuoD7dW
VlW/Xyxjc0wqeBreChL17i33HcERI6LTitq/w9Fm51Re5DxDV7hsovT0Iu2x//Ha
Px3OzO0H4IG0u0gHGmtls2N+5zZKPnOU512jiJieT0wKETg1tmPo7cy8zOJbeUk7
aZ5Aslc3FC3USVonvJU7xUdW5PLDzl84cwYQa1FSedN3PwVx1oeiAfjZjdV4AOyd
Dyt2sWdamKA+OQWf04XptSu2asAM8neEIYYhi+LmfwRwsMzPMTEFwhGuNG2dRGZr
WTXzrytrnQg6bjW5OA5/+PrdpYKCybJYmOW/c3GucWpG0nzJ3BM/ZgA16+jzOLtk
7sFNCl3e2or6lSnw5QhmPqgMQIw2MIwO5Axj4OTW2S/462fcbmm3VhzGwfk2F6MZ
XCiXZvF9rCj1JV4urRWpfxk2VqpyIk1ag0tf4B0mZjVhfOeL2Nou/++B5MdCTyI1
vOjZ4VSG3ZQ8PKFGNawCSej05I9grwcqd6JzNzBlZysEk86k14HA2zFn1i5vD++U
64lANiVKmzCc2gOce5mViwghYUeq6w2NPD7cR8jMDQCMP5GlUz5K0XcYPGyrxZ5h
4YOFQfX8wXsOfr33dmwxSd4lDFhfyY/5j3lw6ZXug1927cDnoPv1V1I43KOkVFrX
9S3k4vfPWmBriO4cRgceR8EHS3g4bGVM14bMrWAyreZjXVvSw3hSBL4pmYxztwFU
ma+vZTFVzKqn/WLJ8zX290Ei6bpUYhOzsOIYeRiEPylvDQRYbWZnRXvc+qME2A8H
p94Z+7E3kkWeGqv8ZLv6hMpovC1DIieO6MqdrqvYCMoFNkBFM5kiIVEhDvM6YtGg
3dkkt1S2gaeov5zuYLQHU81VWZkqdDKspTFiNdtHWm6j5r+nK+6RQtDUwN+pYQNw
i9z2cUBP96KtlKW0/19EP0+i3XZzsJ7S1aaZ3Sm86eQaHX7yP52b+E92mxfA88+k
gpLwwdiW50kkfLwtcZGdN2tbgwtLh9k18w7j6GiLPFCzoeWLecoc0IzIpI6b07Q1
jm75c7RMsGzGGFfvyxFUHqAmkbSGhR6QEpe+bcJ1UVlEVxo/1J8mnNnQbHxbJE9m
anhZZR7pIrn/a5N5pgfGsEbpUDop7XPQcNh8S/p4AOS7Ev1RbB5L1nB3PpPxJbMW
CrwTP6NXljg1/EjgQKL1UXlZu22NOLosQ+e43X/dDtnliniYG4evWwALRiM5GImf
8J+nAULC/UyqTp1bjUqIAALwsraQqYyc1DA1J9k8m3EQpAIQukwXq4OKvcZsf5ro
vBdz90PxhHVY2Fdtukoi/r0at5La+zPhf9daZW0wkIVpNjpFrmEP2X1fiLs0AWQf
WnB3nQvm8ZsWHgjW85/kBUZziWVfDoC2ZRQZi7jKFU1fbi90Lrwhbwd0MVDJ/yZN
PfbRbXJ0arYExR5nqQ/YaoNCD+bt2Lan7GNUTKm6JgpbzpNszr8foLrzjpK1bO/h
7HVrWHNxapHKsNgoSo2T7TTpA1Ec5MT7zNa8tTNZ2VFbDWlrhe7Q/bLBVEIKkRR+
9YlSiOtg74JLAP/7HRTOGILpMw0jEAA1a92l5wDkDCID63TSuefR+rRa/ouJgHV7
UJ4OJhZHrR8RChl7W+f2tFdr+N+Xy7XAWoqaiH2bTrmsGNvifFRKwJ/Xhe57Uufa
Jrc3fKRIh75M+rG96AAOrXR+dKgJGvedh6UeXlVeHfozJeAl7T/2gCGCYDwgh/5F
mS4arva8qgzfvDqCDMz8nAUhfFv57xyNcFFZEn8LXgc8UrJdII61vVgdAiXnQRFM
h85GAOohK3YPDB/PNSnPNnhSbBo+EOycsoPFtuTuVSJB7NgiGpyuQbdIyE1iM3pH
8ybDiW9vsFBOd+o69gi/rqb+k254z3Tu1EebssprZcaQT8+47wo/skgqXwqtRMbh
RHCxe1zbMhYyN43jIN4kan/gkGHf9hSiISTnJq08BjTZ8rajT0M2JLxja++ZfGZh
mL7jRK2Ogn8nxI5siC2jToqkFiU5xdGd/rzWkQqvxE/rsf3aNvKypVgRxjNE3Cy3
T6wPLyykKkaoIztLY9VyQ+mh6cuj2U4KVsuqyerz/v7lzD/RPXhis9gkGLdFW7cL
xhrOt1QB9QDft+pJASK8eYtKd/X/IHRKWvMlqALdTS7w33bapsWjpOESCra04UUy
56ijzpQYKY1CSJaB0AVgVhEa0eLpZ6CNQcGhlw48vrMpyfX+wlURr5vDyZwYRC0r
Ax+mbGgL3O1tKTqp3X1M9kfXnMjnhwlOCSZ7nvz/frDGAI1weZw8zm/VxvrL5mTl
clCG0AHaYjfg5wp+YG5riZ8/nt7/N0iQsH1FMZkaeh9as6jzzrNb8nnNOWP8AmES
K9vjLRXYZ6LPwyvaSrul0SWPHVggsilMl9RlmJm6fQEXcv7BcyO3yANADgcVCzz/
QXtR9YxQAsZJxJVf8yFNL29bxMQpCgsVqnLl4zhugCXPB6BDf1i7cboBULelmLeD
4pfP3qSi9QCfrv9X7NEXnTqVWxUmqc0V5OIwRHLTACQDge6irKHABbvpqQtTgx2r
w6b88ioHUyJPCT0PzskM0iuRtfdn5mrPCKd0R5N4afvcVU3T/pJPaA5Kwhcb9nL8
Fi+JNBqa+WTwzeY+1QGHbvx/6JJ1EolxbsDevifEKQsmr4Br1xsETpPUqbk20QB1
pc3fYJq1hwFcy72BZAtsdVAt7kmAQ/VfBwVMLRT7xIu85KcbTcKPfy+2DPjWQ5L/
ndnHjxaE23C+Upx68JCHPJHui94cApt6vjKG2wJ/t6hIuS3LSuON8aUgOG0aOCig
X5gdZHlgc9Y3s6IyWR4Qo4KVV6X7hdUKOMxOFnyx2XXWeEVdLolfI074rn/IaE/t
5JBN+fjxqhJtjDzOOnapziydUo16MBxs7lvBYVmTCFQx9ITYwatwgLyCrhMKOyRz
5DIsv9b9dXjJPY+wTx9ORNcAosynSU+orUUlwh/fTvAYbfke+cNB6qlsVCziEjR8
69cnOXVGxwcyDexRHAY20YgtoVKZ7AGW8H6u0yrQlmdCu/4/ebxaGAU4fZoUunYU
jG/+E8K4kQi7UBvTufm3Nd7AaB2J+AVGdTP2J7OPlS15wi55U1shdtp6faT3OTVS
swnmDLwSd57wm1k7ZX3F17HbHd7Z3gMcDIeTDlWt0ka/bJjD891G7o8X7DInD16V
za5wMmSlmG0bQ7+TPkl7kCgeoNe3BXc8IikmLbmr3Cl3r1qt47NMGcz0BkRtYgwg
bgr7i53Lz4Ss1Cq3LNiUz3DNow/nX8t9iKTJNxWEDoVu2iM4IskZEuwjCHm5albr
k67cVRhR/ZSCxNbqbzj17jD0STQdzD8usoSrlypgm4x/Zo39CNsiulSesMdhRwWi
ulCI5rYi1v/Gtbzj7CQ6zQhSNN2OwTrbVVWDB7mWjBnTRmVciNXzX3G7T2uWXWlC
alAnX/JpnjLDTg/C1+Eq2Rka7puYXdEx1Ai4OuZkYVHxtguN8z7xVz0WC0Q5XTwR
4Wa6BLEwZa72E0BQWzub8ixBB8zPp7pwuHyq+CIJoBJsmZLktMlyBSgkYnjPTF65
F7xICOiXDfmTdoIRmlETpdkQDzTJnUa+O3MepOTcdSVkvEslikSOj+o85Pa1iS02
rgM22Le1rcDPBUuhAQNtlH9skbueT7JIk+tSyQCaqSWwY0gE6yLDrSm4VCjzthkX
1XzhM6lnhdJgu2J9GTZ+EydDHTuVIXguYMi6QTG+R7xZijcbq96wP/Dnm5pcdvkB
ns8X6VafQCdDRJne35163a2unPMyh5GGea8nhABIfUbQq4UjTYfiWNp6JQuJiBk3
G8ZGG+BzwwQg7pSeOERAYAIhliQdMkTDJJKOqqLYc3A/9OLpeL8xOS1Lui2xCHTr
XpPKyXCbYsRAsbnlKEPg/ZQ4GIc81oGVm/n2p4dLI21hSBe8Q/RzwGvNOdduqOmu
5iPOyw+biN+Z2WxhFGgd/bGf6fwfxqSL051MSt636FXzTSGS6HKQigKJ9tyiHbON
TrEFiiQ1zMWaGcq1Va/Uo1zx5OmfJOtSmhcHYw/A1e7sLWj/65IUajE43bi9DFfY
FOKggvDcYVm2oLO45NhUXMPrX64QqTJx+lv2nzcItAB6LbO2tDItkkRuBXHD9RpI
1TN7NlbHQHO9SqOQ8oSBE5ZQAqJhR8SRzWM0H1QGZZawoHbebaSuHg5v5tNspb2w
C4ejVh9B0D7JYBwN2rxu+eW/1ixPWzn1C+jpTrdzeGWCjP4XiCQG9q6YeCeX1SO2
vjMdDpagCnPY8TjgKA5JeUelvi6OtZpN7evGnSrEpyVX5cq1MzdvJA3fjquRSvPH
EeMiG8pMldMIcEnWOpLMxRGMVkqRl3uq2AdUQ6ndTUgPP6Qqo8OP/jfVINsL+QKW
2IsPu8u/hucB6Z/sUoxjqdRlP/O35scX+ydvuQsVurg8Zg95Jquxh5I7u31KeDnX
a0Wy4u3ML6wtRRuLGbCQUbDYSrV1JmdHYtDqEMN4qeMxgj24Uv6AqbLe7yGGs2LX
GQFOPFnV6cMyGJWE77K0O792AjKES6yDiHxM8MddS/wg/14eLw5RNucof36cEDay
Zi5EjhHzbiVmN1JA7p1l98JLjqX4yJ9NQJErYlXNNhA2GM7rr/QQ1uyAB9TSt4VD
cEhHQhW1M+4A37NzV9CKz96v/SeGwdSVDXhOj6H3izHFLxY+NtAJhkOheLUQcMPZ
6U60zBiCBERVPVoqw43jNEEtQdauVbWiLi5VLyQRSbPDsx/m8buK4k2PHpDlrg7d
wHiZe48ASTQf2EiJu1m9M8NIR5T8j4T+SS52HqLpDYLzo7X6mV2dawAq+spVIkxB
+7l44uHHORKMkKcG50OA9hlVzEkJsi7XAWh9MD9sMTqReXc5ieSLDCNL1tWZ7Gwx
3yjGqs3N6HzPEj0MaK8t0+3Gpxu2HWCY927sm6pgyyuPVjgbu7qdPWMjwjkqSm5K
VT1IdOh2tq2rSZnlcY3JgPCppOdk3L5+ENFt+H077Roa3uWcDRd/QC+NP2aW3ihl
khAWsQqpteFC4N+nsFNFSjARk0mHcGrPjJeIIwp2oez4Rsb5BBmb1TfhjXQHtefI
toVj9J0K5cVHxDJe35hOXSzbblyNWiJ2QpIGX12OHsCVkvNQkh9XW0qiBUCpxzVX
WoRmcC8tx9NbBjyQkle75ZqBwsALrbgWcFeAw0GMO14Kxl/UoO+ojklT7rwYOWaF
gI89Yfk0qTu+fA0bOoNwDT8sYUSjkwXDvjEy/qrNsxEhEHeQo7q7tlmDwnGEx4C4
AV/514Wtw0cR7gZiieguOFJBrOToYdgxo5FPR7MIWlqd6/IuHQSOlP6f472/FmsB
Lv0lgGbZbbhQFScPtzzkKiNKiuuUyGVv8nxU2GXZMi4d1CpwodGAv2fbRxYt/xIr
G4J4Yqq8liXp2HMdE9ZtutlPIsCrsKlqUF1ptP/H841s5Dj3W3UbQByU8Hod5uDY
OLxtyo0IHYSw+0liI5gqWnkP07SBQe4dOfNaQJMKzvVULZUjTkh3TkKGHBfptkqh
cUz9iJd7HNuPLH7p+f6O1qsDSiHrV4IcAHK++/BBiOMW4+luFBvSGWcfKcvEM8mQ
ovJUwohB4pVWXKP5gRBaEqhlhCx3Xqr6rhdWLXRePGog6IatOlFQfsUormxGXdhI
22Fc9GccAx5BCTi6PHUf6EO/VHKoD9qvLZ5HW5JIi8fmndGuyV7K10zUQOWq1rDS
XGF86bIRcjRaahFP33LX7E10Z4qWLljFsL3mGeRfueYtIlF/MxK01OO+JjcZaLHM
2OvDd1MtdPBq0KHUQyhvwsr035+F8LGFZd44siJwO9VT9TpdDX9yOSitqrqTMYwQ
oP/FhAkKIqtCe84HVczHrPpJxmDbeJkwkdl9F6d7zgYrJKTRkhF+LOqUzTF4GsdZ
SUE8ho2clrfTYBThavt51YJi8UMVAfZWXrYdlwDy5A3Q2gPOBKfjB+f1vZAXPgU6
/PcBwgXK0rb72zFmcDXOOsLecypEQXA69x5SFh6cV0yyGjTit2caBysiLrbrMHeI
Dbiz/ixGDg/C1JwXenrLQlXAHREZkyntK1K/UyG87f0j6CNKz584xEkkCbpB3YEp
fSwLCKHocIN1AOD0QHkvygcEcsggBXZr4IkMJEuq86woZ9fq89pIqlS61rT6ivlz
8QZcE3G4UOAAMM6Z6pWMKrTYSuuXlkLkQ0I/MOqzBg/O07p1C3qzLNj51Z26fNcT
ZBoN58/jzh6G2zxvxESC0jmdH4sWH76NpRwvZdJLOa5NF7NGgDR8KcK9PAR+uqko
Gqy9pE5ZbcQb9092XT1/pqdFg0JozEl7xTR0SlgdzXmH3IoBphpZp3we/I+ZRAGX
oMlC5lp1sR2GeWaCdDEZS4GRdHAim4l+PzeU0QyfADbYleFx+D/cI6t9knmUb90q
9h/fLE0sGHycDrzuOvW3Wm1MOiy6BtpPWV4Gy3nqWxy+a+kw5RGBPNTPnyI0JBXZ
mt5CTuvNsqyx2yGfx0hGndgkJhJAc1TBUmt3Eg6OETuj9U62OCNAWopSG98Ok7EU
/pWBaNrMrVbjQCmjKjo81vveEz1Ed+UjLfrRSP3J9b3/1WxwbMIzrI8BofyQ3IIT
znn8yd6GKbYhJTkOQJ/bh8nfscWbiHZWByWVGpMqowYK7darcsVDt+Wqiewda7e+
ssttmwZI/a0Nu5cUxF+ynB2Ld0/1flhRJ+Mf0IaOyzyuQ0r8wNtroowopse/hRNl
ccxiyxNdRoSewJ9PvIxrl88BokI22L+IXjERLfb22XlILYkR+TauDOjrKxs5cDr3
DJNqr2dmLo06qRv3XQCkc7X9736ebJPOMaQTG0IQv2ONAcV4MIWbMtbV0E64NeM4
vBJObtxH147zCh7LCBerVflUsEgwo3rIsGRPUWC8yOPLC5T4ngwoeFzVB4+SDx46
RRCn8UC3H9mtPaZxKFFpB2YlGxpObTs6Z/oM8arFcS3LuBlpa6bjdnr2OXN4mtGR
HcKJ/rl56cjKoJS4Um+tjncU2Ian0Poo6vLyWLEV3jRMg2+gGRSq9qXMhn1L+dz7
cg7IEwFtdd85vzDDeSXRm0i8uFBY2oYd+3W21B2RS27TCi/XHHEMYL5mYdFhsgsS
+rT1YG319lVQf9eCLlJbS3ourt6rMaZJLdtPTQUwZ5cFOPnhofsDgtqQJ7bQAYI/
EmWjaUJqElZwSWewmQLpFlxC5iSSgBm48TDQS0eNpW+7nyPbx2oFVbKmOduPVNZC
Tsn3Vt+j6iJ6UIXthM3w8MzpbeQdLdutaiESARWJES63X2mmaHV9cjzKzs+yHvGy
9hO8+dAVUg4KIXj1SgIuM5KifK59E6B31+/11pSrksXcyFkmSCrH4PopVHTVF2zC
5uOOac3NaieBQ2N/cgrjiA6LLd3UAEAq2gkC9MWWNArNZkSXcno78Lmd2B88joON
km3za9CLik+BhFtOlHqib+1fytHMywRGtyfO5bQzUyhLznKASy4wix7kVFeubwED
tHjr5vMtgAJgW8fO8WMMOEnaefIQWek+c4c54WzIIHMASrAdaoyBHFqBgN32Oxgr
dk0NUMzly8dVK2IaScC3+7h5+oUSpRaUxeIoeMTZC8v2i0+qOMeQsgKLjss8gPpt
oNjpjNJUD3mg5ZjWDKv1z+Wfv+9R3flA0f2E/uFlsGRtdLfrlVkWhZz95Z/urOgo
ddEce033uUqJ4s6ZhATO3m9tTYviPE+MC0Jrh+cSNXsfpskHtHMvoQbVkns9kwld
Ki4myx3WmUlOPHFeUIYkJhSy73KrXEd6XP6ferROLBXArRlGOEY9trLD06uomDp3
iCXNo6UXNmxD9zBGsj7BHg/0UEH0zSiRF/hzf2/qQEk23O+k7XzjNjlSJNDV5x9k
7XOJFya4fMtK/mo1p272wyrcJJaeJFien7H9EL5GLM+o3nzT8q11ypOIYKq/iy1E
BPEOFdlTxtHpbSnVt24d3WVA8X/qCZv4ednYTmyZk9phsxnSYD/fuQIH3PJdVmzM
NstCNcFeCX/8Gyyr3waHtklg/vM7WkylrACz0Wrj0QxWDfBIH6T0AtcxPZslQVd8
Q5ozMW0TxIt46gWMxYkMU3Y+quOtzYYK2g6bGCOoCTIlGJ8j3qgLRQyPyEa0GxtM
ffTp7jxTybUKMW4dK+YtfqNh4tV5Z9hp690A3kfyM/lEOPF57aeLecCObA+FNEgF
LutKaTkmidsOVFd7LM4egSveoiWfpj/CXJV7Yxl3ZDzd5R2w49Qj9DOKoUkyXy/Z
jBzRscaxJdqlUNf57QPx4biCHNj5uVYDa/IrcZQ8H5XXlf2XnJtL/Swy+q8e+KXS
awxJCVQv46yRX4t1SUsLV9KJWfaNwhl1DFitVt7cY0rFcMGVbwsucSp7lDb3HDqJ
MkUXzAHHlUJNnxhgGn0Pl2KhUuiMF3oLLI43ISRl4WCXxp0DCfpSGX7R3leGZEqZ
N40qLgDRlCg52YmYP3q37c5bFLdPhfcJKDeSSr0aRl1kmTu25ifOPQkp50plHNvt
UccNZFWoeMtKO0ObF7FSxkmAFpNFzHsFZxn85ZQjohDghWjrqvMKPzlqYBtlR9kM
bzxIYvjrYgknyFAHuKv0taxDg8Yu0SOXvrMY+lfj+Ee0yp88C7ESjixvMi1XHQEn
TaQm7o2gsME9B7zAPRIG+CirQcZjfnXXGSYRazkzRF10v34GDnKzCF1RctuQ2Id4
Y2Co5RC8l0QVjQhX2m0GnBNHiPgyUJjbHEB3AApicjpgaH4WfEMqsB0eeEVsnymw
mxuQAaDd++JI66TiNQhgpi0VpCFxc0naGQxHS8Oo3sFTzKk0Uz5bqmH1siHOr+y5
yyHlbVR2ZEa4WcYk3bP3A3lfCOEuKDpC6Omxn634KTG/0tnVN9AaWKbWaSE/iyNc
8CdFxgB84QQTkjrTXJ4mvP2BxMvnE+RR7aSju3hvo6AKFMeQMWhknELaYPY6Stjx
qklDYA+59qXfwuSp39sry+zUXbD0Vk/ca/0CRfXMmvmCA1HyfPBOgeQC3iwKkzl3
Rwe5QWzv/ef5jwv7wxwttTvnUTdZEk2GwWT0Gw7qXxsVLtdCNDok5/QikDBaqRLV
GQy6dtQMsr3JDYMeNoM41FXhNRHXB1E7AJQ1rgocbWeYrAZScNZp9d1FiPC51aWn
tUFR1hvJaa3YDaFbpKSlSfYtwSRv05uvIFhtGg7I1cze0P+NVGtWtR3otjK3XBAM
HRIHzsQvYD2bSt4vljV0bijAdxxMl+weLuzvJ6+SsRYmr4AQDMbyTKTWuFzjgRsY
hRFsAPXBwJkfAMhb9S6nHIiRtxSLx+239TwYi/p13BkEWm1x2t8chcg72TCy3weO
nfcvEeE3HpW+4UexDom7L7DOuKl1z+pyd/pOB8plZQO9V6hLp0XJMLW38ZYDyaW/
mOF4TCy2waSukvzvIl1YWMX7OKPAh7tp15Lb2DhTaW2r4v3p/RvKae8LJFL9tMuI
XT1/g3hlqT/D/hSrl+l5wLjrncopvNu0F7hi71i1Cigk+sBuIndxXH8js9bCdS3i
ZVUNfohpa0nZriPWAyanggq6Ea/+/F0Ht9Aqdrl3lDG/78/HHDG0S8lBYL9jsUGg
WhXD0DI8vbo0DLi4jHPYvUVDCA++c3JP3nuDTqEs+RGqh/s5lPZyHgxh9861qymE
nzWMdKaqg1p8/vpC6yuPqwnYUi/7YL13eMYNuJMcZfCytaMPLPVE7v5mk80nsSFa
q9Lw1UMKEl6axtlucIEIFfzpcgDgx5zvJf/xMEhUiYv59j1fP66YQUkombmiKSKw
+5auob1pVkXrffSv+MOUbvPmboswJr+ZY2d8vqXIV4pk5UMPgRtuNDw8KoX/UP0k
eNhoQ3u0QTjKCRYU8a354jMsyHiBuzwYfTE7I7ubjInAlU6nV4bPUNiTHDAke/j2
4qxKx7VhN0eTQ3yrMc63LTwjDgCWDNx7gUChFc4NAexuYM8ZrcthHdoyBppPbXIu
V9pI0sOj3OWMwIaYSM50Pjg0v/zcj1/Geo08/3HWRvk2ZDBe65ibDPatrhcln1uJ
lDf5Dy3WWuKUNyaqg7yZBCDtc3/w8itiCJexFnX6s2aC/W8RV3nb506bdnVrlZvV
GVWfUDBZOwQqttTVFgigsVBQG0jzWs98KkTLt9bw8hnIlHka/8KZcuUjrYSvHSt7
7hI3vSRlBkcNt7Fbogi8MrBysbVaJlt2voMT16p8Hmu1feEffaeLFNicR+0ln/0L
FCSOzGNi2//5nm4m6nxj9i4H9xVetKuDQmufGQZrr58648k4qOdue2pGSBHFbV7E
3Gd3tkBiAhWgGlpU/LLAAD0QecJFCE3SKqybKvlxQn0MZc0ji3dREg0312U6PEHV
qArrWpa5dEFWeXf0oKxDhR9gA9ajrCUcrmpEsHI9JA9Womcmur8m7JyZgpqqE5W8
kmP1OWMg6XqLDba2DwQpV1aBh20fHyBZoF6xbPQt5kIP4sAwEJcnkAgnLX4OUD0N
lUZMPKZeYa44wnA9bluDoYUifr0vfegJG75I28nrFDsfy1TuLXqUPlmdEwo1riBw
WRfFkv6yNxwTdHremj07wZrTke8pfyChgcS+hG1EQirL9qdYMnnzsxCIW8AyfzpI
a/IUePFX9ZwBs9EpAdAygADS2kWxinq4PGvUhQU75hg7P6Dxn7Y81XaBJl8qnlEH
Xco6901FxbhyxgzI39ZTaBXFnCiDB4adUIT1d4ELuLzthpUL+M4gImsQQhTA3UWO
5b9jjCrI/vMLRMCrABOsk0piSM+EM9vVrUmm7nmuaD4Zq8P4hwH5GjS2UcMUe/z9
iaaNusJQUPhaGy7HxM3pBDH9SKodkDt8jmwnVgRT2a7guXjEc/+kpe0zgAIQ+Ic1
n/upM4wO4ArsRnrO2GxQLln8I0i33epSr7T8KMsA2tKY0XEngnRdvYuwm7+KSO3G
SzBCFpqmNCheY2Sh/UEDaYmWwlLTdz1zJowU8IQO+jIoXzilXBAOWFf/FDz9hMOj
apSFkkCVyvnrVJFguMNjOkkmnUGSC/V+NPYAHWU980D3n8MuaX1PuAHfznh439qg
DCV3f01uagozC+CAHelVmGy6HZA8GnEA0DLwSMdmRRW2T6NsbfnO2bZSJJjP4GoK
8t1cMotSUXHiWvYQlQWKDLi5ZXLoEi8yCMig6htLEx2CPjina/vpviVtKVHxSw55
jPm5f0nOcExd1zlVJ7MeYyftUkJEkXwBqrKIojbaYyIF9vQg7TezPSccLe5ylDyz
CQh0pi07FrVQh73s0oojIdxC9BWnitsh4k2G4c1LgWfh3/TeMJXkedEjsw3VHR4y
SaZ9vUWCY5YVcnSdhGrrT90OZ4bnrXydzupRx0SLD5DtkzHYD9Yl7PCirasGsntw
CZoCnhYJjail3qre1hpcjS37V3c7Rcgg9lTK0UOJDjICkN1C1rM3mGXNihLQW87K
QHuWwUUwLiwWUl8VbvkiD7UeIOQPUGve2LkrjWwBxhPAmghlXp2Csgen7k/A1gkL
YU38eR6U1PtHLK0s1mmDnglkrko4f4SdfMinRSSaF0dSP979Q/fsCP4dTFmyqWhY
2etiUayiE/ZsMJorFq3hCJPDJ6VvcrGlSZ8N8MAeYeAfKfcFT4ZQR9ULoK7XvErn
05cgF/ho4wcApI4kvifvTjjc1/bahjiyrkrHRwFEYJg7khzu72qS26sA+71OC39B
IHvqOBSV6YwSLSUGjZ86jECWcb4brjMislic2rPZ+RYu7W6/dZQWqEriOQiPlvfj
wzbS4TRAvugxEW/gaSvN+pKY1AyMd1kmckgCl1s20ieRBCqZARC/GJBwyYKoP9Qs
OGzopJMIluoGpks+iFtBHBlmjy3kvxgt/CwcjrRtasQhfyKAsFhuCFWjj2uTO5J4
Ryge0EmrUQ+VRuuiMiPsHlDAH7AJHvMrc7GR8caF9E/4RrjY8sKWDtnmLC7oPb8/
l0lGwRwMOL9UsJ/gVsgxFQWSnDe7NnC3TuPX/Yk+P7Y9JcZh0+cHU4GqB+fliGkH
bm1te1Kk3Ls6mkZ4ahqFLE02+zec6MP+dUertOVfYTDjpXX8VtFFkTiuEce+6VX0
QtFwY0QHqoA3zRQ9//IAZ2pH3IMTiQhVM0JN/Jp3y4xgrCik1AybV6JhADN+hOR+
k6U3BMoWSH7lWGJpuuCcLDre5kUGjweuHLd1EHeQxwUPzqCXi8N75qP25GhHwGX7
/SE8GWIoYsjV+tAULcgHrGtftwnU0TnJjCKQIccH5GkIG7jYGencufMJaw6qZJyT
F2clAUacniixdf+TwMqOPBL1pVMx394KirFtANYU2uB8vUQqMNkvmsnEv7W2lVxQ
i9gAQqgAIWM06ZQOKO9bDsVeIOZJjoY/e16B/N7ri45Qfyk1TxhWneznSpwjhJSU
fVMgsc5amYDQthHEa88IG42Z1td4mEHr1sY+TxUtNwE2mhlh7BDKRaJu9Jh3cl+j
YNIe5H3TTbnDKD3ulPHk02FwD5sMYnwcYuEYsB01tjK8JvpssZepM+NVhbOEwJhu
Gb6g2ihTRcZ32g+R37V7OToMu4W5qtvyHGGy/yMLSFTzrJrbac3lhSpRMz1hN5hD
6kqFGrquKWY+gX8GpcZeJ4oZUDeE5f9USk0tjFoUjR9PrOv6FZQ7A5oP8vlK/bij
7u8I3MIIUYZVNhXGNdlcxf7LXSJJlWoDF7gGjMCc6LAHtN0w9dORmJPUNCZNcXVh
hGFo668gxOw5IiszvObry1+yDMiJk/8YkhXkaXWesCl+3NCCLSbMP/NoGn8/K7Mc
7JvgjbgDbhypB7nkkEIBR2aWYWsacf6x0DOGGWkIzHSXj6yEVoeAPLD7SKOSBcFR
A1xbSTgzv6Jrh5WH/V6WjnBGIdoDRX+jaYjIVTWVu5iedH2EJS81UdqA5nWtsg3P
r5F8vuIY2VAG+JeTUccj7aMVWIJvCjlFOX0g7co9tvdABSHE+KhJc6wYQVgzACgV
Qy5DD8iLTwXYplOohD0p4UrHuAVw8K5zJWyYiL8CLcYbVol5xUSRicCSRgPJpnee
YkvXuGPTsG+2GBedtxz9yxeke93sJBJtLDWoe+Z4u94elmwI13RHo7AFJPZgCBy6
/D1t0Z16ULUjHm4UGd1gRg1MdQdakLKv7UsEWqfwdevR4oLdGS4oQ62tUNoCyIiY
DnP7HtIm3J7a9BKZHxIKrVtWNteXiBpmy30GO48VY9yYNGivgzByaGZaJSVBfh0N
y+EHMxeqqU9ILAZgaP3u/+05NDSG/6MiW52ni3zVNCMjwDLXfxpysmiDy14Zc3M0
AkWRRZrkzAiOlV5XFvJT7vDh6buIWyeargqQOgIJWExGByF9DjqFozdEddTsmRc/
yv0WoFWYhSfrTU2oOgDKHDpG9brUzaBwq8XFqIS4+0voPOXYwM9XlFDvJJF9EXoI
mH4zWKeHeTbFtq7Rn6IOQ+L4cnxiNfZlZloAxf3MEuO6uFRboHvkX0EqnJZRtX4a
143nKYZzPLYXV5wwF/iy7hl9o92lZB40WyOIQBrw1sB36DLNrAOTFWhLDuSxrJsR
p5DDkcimhfObNxR5xgk3W+v4SyJ4kVSUi9ljVJoEYopv2w9XwGYXuK1NvgWzcJ9u
g+NvZueBoe3uwM5be5lAQTbyp19PBxOYKw6aSzmuTOD1YZgtUuMY/R0fZd6jVT7X
egVnNtnZUP4/o/MDUU3eNKNHOx4eNGgTFgQop5W+tQXezJBNO6MGZdtUd9FVPeZb
A34SEGju5MJyNVn3j2y3p/a/daTC2jm+HzauiB6m/ytQuiqQJxBy1p8LdQEbqxsq
fA7nraj3CKes0A0YiR7NyGP8VXobnrVWwGYUDsjaVKLv/2h31/DJStHXyaHbKVrE
u5WN+lTqhTFu0HXunuTG12jsUqiOdE/YFJ9B80WwpvIxtDJDek43BXO5VcYu+1Qi
AwsMAIbeDzDNKt62/vdNlXxmLSxQBQNBxgLqy/uB0LR7UM8i4BX8behWNdpUE9AH
yhaZjord7WOisnGS7yXXS34y73owxixk2r5lqmdqoWmBgpjCO3Gm2XJ3YJ5yLMmf
mvHCga38/V0v9DnOBYJPBHNyfxyp28Cr1mIb3xLPxIKq0JMPPN36ubphcDTN2t9T
7HEwyDtgeIKOOhonquT8p7+n2i253v/n6HWfkIbys2BTirkll0ToVKfRMPfIWpmz
dnHcZ9zgqQeRZ8CpNvqIoVIB6+tZEbfH93iS30HQ3hXxSafvw6S1+4J73YsslmEH
HZeKdwmaZKo4CbIE+LKoS9RtYXoitf6lq2QiR8sLT1Ne20/1SUndIO4p1pIG49by
rppM9K5G+9fPFyJpYSofenlFGL2ETXNC/9xr+GmY7N2eoPUENsfJHE8x2zsBOsny
EgO2VBbV2c+jrx/naIkNT3MWCv4WpikGhfKH+v7utVXRndhNZ0153qZc/SUYeETg
Qll7x96qczCI5PJnx7on2lZ72EycZwDq+EN1mfvMSMX4pNyJ0VQlG1RzU4i4H8c/
iAfNXif6fVzr3Rc02r/2cffCu3dr6nOyPLPnJ1dm6rjR7hbFmDFiGIH9taggdXmm
i7yeQiQaWut0tQPgVdj+mBc45KniRVD7QEp2s+XsfZtMO3xqHFQe/WW0QlPW3pbq
CLxedWR5bqfq+0PVa4c4Y/Y9uSo1UGWuYhMtQsh/9FVKhPVabyt06ihl2umBI+El
TxqI2UOjw5KvtW+ZV9mTezF18g/vrlnb8zXUWdeo5Ddk/9oS3VgwwKw2ABKaUpQJ
aeRNhlqbGr2vPiwNxvJoXXcl3UcBF114OnG+/h4xB8RXSULQlDeWm4VVgRmXrWuA
z8iuKeh0+PDSWWA3tS9XNDaJ/lyRCqR/pUr8OK3kZbyAxf/11qF6UrqJOHcHzMSN
yNhlvnJBW1nsISDW8VqKtBk2/CK3klQqwUjMvut+rJ3BaGJuh4Gq+bkhTfh6tPK6
ocDb1Z9Zd5a2c4kUzcMnEJYIEiqT9NxwL4BM5M60RrRvhfaTABsZGljQpiELRmcx
TFMEs2GfGwsbe3KXkQ5ZIRQjZiaG8He0zul3Jh2E3mSYDqolnNWKKVnczR/hAYXS
LbPos2v0lk+8/ZqsD9BMbcFJ66+nMQXw0YHxJLgzwmYtIo/HIk7i5ScE+3JomuFt
7Cuqd8Ixbw3vhXNWUy4m32jp/nT2sqSqnTtkCBPB9VxQ5J4PHgjvNwrfrLIVzl2W
KyKS3sCfvl+M58UTap9ifz6j+f5T0MItpUNNpNsKHq3JX40k4mxGkBIuwoXf46Ot
jxHHNbqpOuCWg7953Z/ZdP603mMz1g0hO99eb/OJWK9Kb2Dcv+Edx4rE4RPuf9WM
Jz5bdyCdBkQpLTQU0eVVljs+Vzg6V8wgOghF3I5oDPExHKIi1Q8kl621MiDPDKUN
RsG/H3ui3EmXpOl/dXk/YKHisVvA1mgAJfBnFZPnXdlkfr0mjs0b1eVMjNnXPs7B
1eHQZ0C2laayNLi2+9LUIkX3U14z6vasDICFYnuX3ow5oHH0chZ06oqUnJ8okjEM
H5hPQiu0kOstmFlULDIK6MUpWs6u5LWevjaiRsRezcFPCBOt9SL8IygW3vP/z9bO
FacAXWltaJSukpDrzLLiQUB7I+ZXxCGqaB5ZpBRpXGhknlWCHWa46wac2rcS4icD
nSKGZc0b8ciqiQ24RkEMymBUSFlfttDFu/5UvACnrlAI7pbRoAxM8YOKY0/ZFiHr
S2Azd/bZdSOrSlY+hCiKvyN6WvOqIc74GYll4st0FSlXi5D3XlstWF9ocmE7l5l6
Q69y7xtzQLetsQeVnCzIfhbxJAoI6dlwPN4cU4UF9sDUFsOZ1xKWzBVaBdIMzvCN
OUQkfFlE5WxE6lxv8YjbXJ8Hr1PYcxlhHhgGDeQ4a2IXBFfJW2/yYGk2Da4rQnO3
9iOztzGHY2sjk1OEH0OvjRXdWGEtsyRYUDjrWMGRQ8ubXJ6LlwmS0FTUit/VQLzx
7jkCIm3sHWPxr+76G5xSnTvrdRv3nXfy+HlFMuZ8ojmTm814DXEwmo/pwwQF5tjG
mq711iXgkTa9ZlJjY7AOhyrVBOW0Un62nm2OBdRq0eSmT99u99cnqC3ra5Fj0DWU
f0ePBhoE3OJkvgAOOPTsOlnmPNS9eNMSMzOd5/2Y/XbZgjeYybNlbspVhxQW6fc9
9+vECMk0kSQ33Ft36S+fpesN/XueGAGvUrYUdFbK1EMwIlxkM+r5UVJv6xhxN58b
6Yyg7LanwHjw2LgqJou5fKvlerBa4Ha6qTlh6hoQjIWhlcTApzjTR7j3l49AqG9x
u4ZeJdOBEXYeRhbhskoSCcAzoTmq2XEy2wPv+8/5ptA4nFHBvRdKSat30eG5CSAf
4J5WOGnHi7m8c1bqNY8kMnQMRxTYJdnRAysCVwKQ3pMbGJktr15dHH+fnAQ8B1qq
zrrBr+J7fwdVs0caM9eFjvYW35FFVDQ66OdBl8bxpJnJTd4yvAFKndS03dnD0iU8
nlUiF+VDHCWQI+Et04p/5VwqY6Hnx6wJJqme+ZrgJ5IDWLrnc3SFf0Df0lbtgkY3
qZ2zSJpoO0WWdfOjBZOyrhUs+UFJPS+Z6o++QN9WIfalIPpfGYQGiC4xsPN5VWSY
Rgy1N7SgGd5yEDklAgmQjiRZUoXCcda+jyDFHrvOjQLdE1jDbwaG4BLZhsclWaW0
uy1Un5Zmz2t7gqKJKS6TLmzgDwkW59nTHHIHKH5x+XGkAirUh0WbNKW8FncbHSLf
3bDfl4uFPMId1j+qyHZB+OMXeTZuoBf88izlZ/ISf4dLSmczZ3HoRErrIbarum/C
W6Njpy+GBxm1pt0OjPikT+U49gYLGwDZIGpE2DPfPYJ3AcvHcpm6dX1TZ1iUFpef
piscq/caE08zafEgQVH537BpdbafRsUixAM57XNgrCaXZLNFGqwr7YMjo6Mgv9zM
g6ekEY+4A6rfs/7nEB1n++WkK5ErYIw4xonydq6ZvI1BlVDmT74J+86AXAOKdk6o
N/mmH1gRjmTr+wbiGnrKWGZKijpALwwNiy6HHO/X6bA+/EJalKfuuQABx3rolRBf
3mWndQqisdW5vkVBGbHEF+oBfhYTSwff4clcgctJZIeThnuVbd3aJajRDunA9FUd
AK1VzaadLKkXKY8W2+DylHZbM4+F2VD+aLJfKfF9rYfZpkrYNPLKYHBoxgZiLVDt
UETkgWnJW0vA1gwd/mUmWB5OtcVlnEgeKzo8oUamhKOga9+9qhJD0ocYeb9xKMK3
BPxUjVmN2r9zDLLdGGQOdEzYyD0S6tgxlZHUD33gGDY9qUBj9YZcaFjkgwnII3lW
S5HXpAXn5RtjmzxruYwSg5KGmX/xNesa8kFvPl1GvqEgS+KP4dAtkzDvFi2cUkN8
vh8qihJiNn7HEKUdoN6xEfQ+R/kJDMc14muGgZI3fsRqkrES4kZdkd9lR+sI+G/o
dksLwtA5QSC6BaovYVX6h76sQET8TiykaDH+8H8vaEOuQIplOHzif47KLUYftjlG
oOYHaKbJth51WrobJBgsxZeCWQGHEjLQ7m2n+HCX8WWpJSEqatzQdtr2dEEvyMQR
n54Z1r3uUR5JpGenfMuV8s39U3x15sEJOK6KXlnSAQHU5oufYq9GqEzGuZGOvBW1
toltYkSOnTIB3SLWNIn00KnCp1YALu32g97ffXfdRynE4y99Y1FniKKzgAm6/OQ/
Y4NpEuB0G0nmDXVR6NDDT4l3veqnOWOVhZBRVsQ3XmV/2aen514fyPGe+3s/g5Y6
eCmNLbXPG6Zp91MWasvjMOSGbl6soYfZdzWuMdIf3BiB9goAJ5CELpMUoteUtvdV
7Il27rprfchteCMqco79dxSFUkc37q2W2GtJXYAdKVlxzRHeawF73JltXUkyKQKW
Lz/BFaVD8n+qy0pDUKpgsoNAUvip4yTZ1mh/BEwbpSrnbDLCoEJkMYYCu7ZcPCJ+
WdzHzwIofaq9RKgtV0NvKRahTfSdbA5SqmrxQUgTUUSQIc5sjT4Ic+UzqEYRWUVM
v0Im3d20m/3kygw/O4RefdkE0Mk9mT84TElCBu9jo32Kz0FG/DGCMTPMKwA2Jvl8
+cevxBjYnjCp0vtQNzN6Xad9ZYyXS/lZBA3YYfsalCMaDF00UW1OhXpf55Bqeo6f
bAVJi6MWyG81tQ280e1RCHoLBSkjuWGYvyJA5vr9Nd1MDyz3U6DZec26QwpCaJXc
rVJR9sqKkleSiD9Q2Mzxp6x/LHLo8YcVsbq/Vmb9rzet2bdmB3u7jDOYOXTBdje9
t/aAhQ6Nf4mzFf2YTVrwfF50Fjs71JJjgMKcIVVV0wwyDCEjE4Fvtn48leLRlP6d
mkybaoV+3UEQPzdZnvTmbqOcVCsZDft3rMKtWuiDYSzkQlGDGEcPIlWkQEznDYyn
tJklpuFcHxDFzfnjbpIJDP4znSPrg3aoVIcAWL9k2MXbWAYgCCEutY3Dg8MmbVLH
rvf4W+E6zUaS4rHoalv95RW1LQIOO37Q5dWN+ZEpHEbe32Z/Z8VaHo2s8+7GMC8M
8jnfPV/+xF0z1DuQmWyI1ZjFxAxt/bKTu+Z1IZQ/11P7uJ7HqHgV1TXytEBQV1HG
XCrQfg6Z1OH/C6yu1NIZd6lMWSw9Wg2tLZZVKHaquLDeVu8yM8bLlgX9Xz6ta+iS
vL/9Qh7t/9Rj0eE50W9sfYjGw1jAdXvLnAnkqYdmXbj5y29oO2a0Q2pj1C58UeME
Cjmr4FzkTwaHHf4eZpjGSXe/HmojJGwzhb85Z88v7uP576Dux5gNp2og5ELZNcWY
AkPQhjloNwQtOpXLsN4tbCs/iihnPPyGQe5lhp5jCihd0TnBcSw8aTn2zwIDsUES
ruNjYOd18AuBnBnRUCVZH+odZx/ymrSkuXtrnn6Ogz6vEZyyLp9+rwgYH/yLzJ7t
h9tb0FzxjKAXMVXAbe0KNPEFsozsGCs531n3m2fhyV/ZKYpxlx7UFDm5AQwXzhZR
ICipb9BxLYcPSBngrg2T1yY4nSQnUi3jOGzwlku2UUzFXod5xSKkWRHT4XGhYkoH
rSXWL0xJOP/xaRql7a1T0IUuOgxDT6YtM0BcGek6aHCnsfjabZuTFKUMv+x7OJMT
IpUB60dV7YUkNDG0tCyGyRAs4LOrH5ev9la6XETwKIG1iw49W0kx84wR09NsKgmg
i3qWLfAxReAgwhUKec4yGlmAl2He1HOOpxyfCpevZFwpUECdW3oJHbb54ZK40FqW
NjPlN6qscLCVPol117k2a5cTJMeN3AsWd89g4tt9MrJKGaFqFMdRS3BW6LGyKXwc
U1BzaYZ276jkUF+nOafth7sfCjhiEPuXTdU6Q1wKpffSN6BcMbID9l+a6zgFsytJ
yYA9BaQQoRwg/27FDDd9M5RoQQbiQrscKFdIOMfEB42SVyocKTo+7QFnLkpIfcAN
Ooviwm8EqaF+cV6G4oy0EC6TM7giPqfZyEuxqQDbojUHQrnLHZn3IGkXNYGpLQ/y
NHvewxF9rhC5pB4QoV6ZlhQLT6eqOAp0EzdWq1z9xcwLC3zpMwVQoc6CPKFaU4QQ
Z519fQ3DrIYhRZqnMdBu5YOXXsIDFW9lIHuAodwPhXJ1VvFFrqjsCrJwBazf2ZK2
wvcDNiIYGoSyHN2eW9GURpsWVa6/6WhsKBtQ2byhNwMkZR3LiAJ+loKYYrhMwCNJ
YYSlOPHydsmFaHUdx4mBlXCbJ/4ka9pPLzhKhnpkJJKXgVEGygqbQ6P8OMyNY5IW
6D/Kn6Y43EWYFeStOlQl12QQywdxpmnbwD7Q+CRvCHHueNd1AzEyZbpoif1lStoO
gbl8yTVWxv7VdqQztJL8ah/nGy6b7GTQGJ7KB02HpVbReUZUIaV3eMKNsAULQXlt
akAvj69ULFmIloCHIw1R0BBTZqJPCDixLtX1iYxJSEHLQBdw25rWzEUgbr2/Jcgt
RFiUmrGL5njxzIvIHGRZvciaObZBNiz33vEa0jVsQwNu6zN81gjuS47Gs5zf08pI
euzU3hJrgWRtIimalIH54TPL7qhU98M1Q92Co1123BQLExDNkkXl3p7Ib5b+/jlO
QNa7nOrSi0Be6U/ayohQ7bTwXjsHQ/0cZ6MluHgqTwAEipk3qeP4IO1WbLz00qJ6
e/RXJXSQnkDE5RvuuaciBGzNdA2al/9yfvnDelBcAY1RL4rPKRMiF/9Foht9TRRb
/FtOfDUaRp4aS8/r2feyr+dErp/UlhYv32eOsAAAUABIpSxEBGRF9JeZcX+O4djk
4jqU0yogsiogKjVTAtcxakFeDnq0p5Zjw8WUw2EAtWb6GPVwCxNH1uJ+e1o5qcO3
D2eQ8hk0CUJP706c+ejeuHmfBpLOCfknbP8EUfEPetxok+oOUeL8RQ2d21CAC6+5
EwKpTak0XopXQAM+RK3fY8pyTNXig78TiPTLDqwWlphgmSOlyBFvyLmm+nXaAM+p
Eyaz82lfWi5TJbQzPLTUSFmv57RRlg1lOK5sRu5HKAYga2zXwGh8qwf0NgPNv1kP
cPclMeRJHGyo+uwzSmtGN6J8uzBBSUZXDmFIEyH8vr9F/pQ9cuFS2WbGCvqWWsGh
SuX3lCc75HIXuQdvJWvLBSy6n1deH6e8ROYrxGIJ3MwVSNK61S7IQ+k9B0FkamrG
+F7Rni9s7WCfa9BGvlpE2XrngDKuSfIuzS1DdjtD1OxVaws0l6AXAM6RHgwChAQc
30sYH8wJc56aOSjrTHI5NodOON1oi1m4XobGqGDu9gbwWH6JtqwV7km6XozXMnoS
urxP3PvHC8dZ5jkTq6RNcDUp9d1DyaEWmeMU8BgsygLnGiuz6QL6YrQOk/iF3EcP
qEAZHIzBnF2ffq5WrQmjmyAaVaaG6soKTI73IVTUWRl7wVuLUl6LiDkRf5TJhIjS
ekT8KpUw1QsupHxV1MLbVvzjoj+vMVZ3Kt5hJlg5qkwbfSAe8Y37gCr4sRdP/XxF
VhVOo27BlDyvGpkbBOUgT5i/iXo/20VKCU44H0lVmqCqc71Hk6JH6TTC9vE4LuWM
9teKO2KMPd8FIfPY9AxQMwR4U9dJ0MKMaLn5S8hNbaqtXKAQegT1if8M7Cv4mNOM
Z95bIeJzrfuDZfSsb0/9xX6Hewj5v8yWlS41hhKqVEWNTfcubswejdikus1oidje
gGHnCkE745OD9f46VnI+oqUF2R/AjKJOg01LNccbZC8CU/3WnVCpZwBhzeJxNQaX
tuw/vnx3/jWeyf3Pri79QIPKPFokaSaU0ZtssKHM+qKsX9wZKubb0ze02/NJ3Kvh
VB4jICDkVywoGiMwEpl48+MawoL8OP0VoxNwHYAz1V2tH7PKbVbE/vOohKvpV6/N
oz0svVopnp5c4hN3o/2kqQjTgsAkaT8E7PpXTX/IyKs11krZ4UJ5ZogZEziX5+4m
Iasm8PsX5FPCF1IV4IuYm4wOVWoko18zNehqqVaYtgDmk6eZ5G3eaBNa3KTtBwna
NymQFpHu2VUHaBBJul4a4AGxXlf6bg4N7mzbMOZP0eAeocfDbUl7/WSVXKsOpIg3
yuqOesQyWtRjY6q0gRVC3hy95yQIN3vwNr2Xg0NoKX4vyDTRe+U32DwwarikRMJy
3duKLBflPz1U9iTvsxz8M3k2KrnhtiMfE1c8WT9RSuuZOzacyzZ8Ib0uSRSqb6Dj
ZC4ESoaRV+5baXIVJYWWlQZPF6tFpJvsmYLadLMTlNO0QgpeRLldbJXuCE7xDIo3
vWTVklagAI6eA6MHt6d2UIED27USIaXpXwPSpbALUFZF7RXFmWx0boGQNFkAH87a
M+ktP+U8oEPfV+HILlr/UDv6z4MUbBwXJbvHngyYGxI4CXLwVkH3XX7fptWdXGvi
lqcu3Gg/C+GPdDhkZ5NKlDlPbRhSHl7b5BOifJYmES2g3ZIFm0eHmJpZh4pVMH99
iZsJGc12Rrbflp9ongSUCEhD+cLrCla3JUNd+CukyprK9ZVwetTkESDo+6DpBt8J
/qmk6UzKWLC8oL1N43lm6V4MF0NiaNWOJPgAJHvX1IYcVY/IHzE1FfW2NTj0rRvo
k3ff5OFWh0Q6oAOSx5idUoDbrDZTOeAZoOewcQ/X+TydqI9krzJDL6wresLpYiHe
BjiLuaFOli5oUwFT+uxu5mIpSfUO6qQLzBF6LuEoHgb3jwot9DqU/E7ffYKkOPS/
VRHX/2CvSlLYiHXQgvzPJf0gCSyNtJXJXkauKn/nZOilC7aeCGGOisHMe96KQWn+
e3u6hKz51i8akkbMLauEzbd2FX33uU/Jfa4WY2f/YmOM61h3QRgs8ow8dur8Iulp
iY4CvsUUTzlR5uH5qDpjI6LDP6N/9pBnW3OjsS+3TRKBMEgpcDsR3FBbkzsXdvXB
I9dJINPwBVxy7LGoSWSbXc7MlC+M6mFzK2CyNstD4OHCn1LPowmZtyjG9v86GxPM
/gRUUjP4S2BrxP9aVO5FugPYsZUPUcavgtrGvxP8XnelgRQoCNDAGadzlhCEPG02
1gIAjku+MXfEs17FCFAPMJ0y5NcAPAbo+9X37Nq9hzHEozrwgcdzqfevR8bLJIFJ
z6zrIfwjtyMNR643I0j2NivrfSZONGTHaXH8pieC/5Nqi0l+1aFIkyziX5RXhw4k
aGO6qZDNE8a4Ah4johZTvrRl0Kg0KV2NhR4v01B+gp5yigL97bnkcb/qNrrxxCNp
TObstOSn7L6F819CGZPDboGJOqv1weChUg4eAXnFsWwCIvSHuNBtqOynL149FTkr
+988RCcgasJgydh18kF2c/sqXAev/80SqZUr07tQRcFMSJmGOS0bc2+rSxK3wVee
qo+IknaOs31/BRyskVt9O/TFwI1EIJRtlYJqyhgbGdTD7miOHJDlV2wlHTLuVayb
iaA2QfB7bLq2cCkTshrPK0TfKD5C/Jn5MNbKj5G2wy5KpYq6Ze/l/naCBop9L4ku
B7OCyQo+CN4iSiEHecA0D0OG1mLgaNmla3Vj1y0tQRoQSN5z2JvJXihMc+TZoR0K
Zl13sMceucdLQkmGj/pmZyAr5ljgvBzx2+O9S9s38Zr3a/zkT2UegCAO20YZ/B3U
dIIIgszCoGwIzReTmWNIVKDDFvoATqoNGbwcLgbg3Pl1ZpRWTffGWlggH4+fO58b
O5WPvWFKi6VymVvvevITpfUTWLw2RLoKdukyN4qSVye59HsioUGOdrr7OeHc5Gh9
Sl5fV/T7aaBEkckKHwQ+is3hAoWDww7Dc+95WG5YJCHqCxk886FA715Z9aAv4URx
lu+kd37/vDZWYiK7oblyDu4iY4/c1AtBIFRsmuWPqmo6gk9mIspjvbIZtXc8g2aD
5PY4VH1/FhFxJKeWzOVEKEhrwa/6e3o+UNyfG9UUf8a/U60VRPcTEk2HVEtkdkun
+u9PbGQRwfrgiPXkLxnzCKNn3IYCDka/9hXUi/6NQuL27+l5WfyS1FQx79vms6/n
r0AqE6yfa41a+7jTOZEfOycQ/wxwN1AyxI416UMhq6581Zqydyz0wGFgmd6aG+YF
NnNYiF5BiMA6KfTrtpO+rN3KvmYGz1aXr2ePizr9Sx40MX/Ih+9gHapVogGLmFPI
zhTWl7NlzALNi9XWUEYByfuNqn0B3NFG5fHEjutjduy4w1ZWwAs4Pdu8pN8GVl/v
NtZABIY67JUxPFV6mZ/8qmgk3qVig5KoJuK3tkJil5VOdbbY1Yia4j+wP+HhtwaC
6jpuQXSsAWxNUzNB7Z9M8ZYQVbjai3I7VkdR0IvdlTFA1l7PXrs+KOoMzy2iNdtw
ifV7fwpzq6Zhpp0jaYMNB4xgP8C6j76dfALU8uwDOpk/rVolu3FcV4qEC6xZo8A4
NA/HSEdYY46w5kRauz3jx+kMxqDe0+wJLQMD/RsaAKHywhvb6rWhsV9OpUCqVOEv
cYeROJT4Ywno0zexZpe8nC1vwGZ4bQKSE/5aOimyB6j9vtHA5vsAdI4xlyRwbXmD
lX7f255nULIojCDN5PAH2UI7ew+fMdJXip3ugbEV7k9rqBZv+38Enm4jerfzGhZj
QV9pDiG8U63xghZWME7d0085zq2d+NFUmHuERk5bvlclK92dAurIBw/Bg5MlyGqd
vpbajwXzRhBZVewk1Gt3A5+kT79ucxPXIG/WYzkC1M9xk+bHbV29ouSYKmOxVFPd
at3cBJV+wsOvBzz4zoTvKHXWuK8gOM56hXECieDwUYXDzLMyToQudvLRTGuvscyn
ORVlwlWtrtvSAG0ojxJGiZkXA4jg9DfWvUhccAuXkXL7ByBqDLghLRD6N1isd7YS
Yj9HzyApBW6DqlVCIBqlnj4DoleixBn6xj5cnonMYrXGd8WANwfakfhKzfb3HW9s
O3UE4WJ+1RMiS5wUx3xVMqJRAZbIVvfKQg6DYbXTjiy7FoQn4HbRQUV4EbEQFJaJ
nRhwNojYSoHrBQ+9cVtak9bYf95D7xfxyzS0vDJAbFB3zZj7UhNlpnhi6yRLBOKX
D6hXVjZaI//A2d93gdwPNmh7WPhO/IFLEapCvPrRA0OxXA69IIASjIR3tKlA2qxn
ClUuQcxdof2awtCZArybNVDqCyFzaA9JEq4bUgzduaFbELxNAnRtNS6JIw+/aS9P
hXOTApv1DDH3NQfTYKoIwsyMpxy5LLtMFN7WVUWT2YqoSMUyy7UeM8v04khxlpcu
fW5+LHxxbrTyNdpIEsPZLO8LfhPbg6FnH26zR+xexNBoEf6R5rzoFekMa1yiCSvv
cMM001njnAZsh32tTAA5KF08pL2scus1omncOZzjgMLKCvZPE2iJFmCORVxkNz0z
/uYh3j5p7HBYb/yTpNLJGiPFpyCumQRd6YJDTSrPYAFByC9SHe7MIqrBI6VXpX1/
bwa/G3okvCsugmnbzg3cCnk4LusytKuhYA4/7xitPN0cXm7pd2DcK/uDhaGutWOp
YWr/zdw1DSt7nGSKT16uchPIl111iW7RWarG0ravKCbi9ZnBk0DbrtDfoIUr8LLq
ZA91y9X4vpPyhZGMRUjvxOMhqtesIulvreMYmJ5bS5FcU7vtVi97aBUx1rJ4wbKw
YHxRqs7/TQ2E4zELNQlKc7+vq3yvqfUYqHa/cJft7NCC7cIYC/AaPw4l26uOMFKD
oQX7QMdCtrBtXibydy1ODMi/oAA5T0m6MfS4EB5EH2qrlV/aG7fpxaM3S2Hpo2vl
pA54qccfPTnZO0k1c1Q12apJp0oyhEombeIAygP/1rLZKt8V8WjLTP5obokKfg3a
MUM3gI2rY159U1sH4jcdTEEXvOBRr9yX8pSoSUCQsau0K7NB7CTgwkVp08AO0tOv
kRoI0cHKfMuYg/26C7PX7yrcv4ePiL1EBQLDxQis4cI4Y4CfT0d+7VOU3RTaqUiX
WxUXYep41/7nzF3wBiB7Z77tYHqTyKfPtrSDzsuR5al5pu4BcadXw1OX2+Fr0ZHX
+nbgvIG6fx/LolNrNDgp9QzEc/eZ5kpTN91GiNmoP+uYVLQkhoc7aAg/jgTvDopN
qfGdKWlwFsyPBjEW1K6oQPuOBni76eB/H6hq7Ri/9zD7t2T2twC4S6shujb4YyPU
2ysciH5LlMc2Xy1hdXLC/pa5bXhocGBcXjamfbUyggDlIvn+gFhTnLW9+40GIBOC
IyGS4JhVluREpaDroH5hGucH1S2CnW+xyl2MPn4GC6csJmSYp0UzAIuZiDxSXksl
Yb30Mo6d5pIEeg/j7r+YdjAE96frNEigaYmC1y+hZl3/oPbhs1KYPs8Q/won0e2d
3FgKxSFd1OIyk3B8R47sj0vAM2VMg8weCuSrTrD9qV0bTCZwoZ63L9lK9iH2l0Oj
iCI1ghMfC6d2X0vRN7dyzZ4XECC9M46VLpIWuurIG1g8pEGomhj5iyCKDRSoiIer
P9A3xmkbjH/ky9jWEBq+OHJupoWhkD5YruwqFeewHZVhMgbB8zIv7gGRU70F8/Pc
aUERQ2g/Fda8LjQf5G4ksp4OBlYbSQmBEzmY2yHCUheuH/0ZEyYTcg1aO1pD6Xqn
P+hByDFGIZ2zPkqPr5dfwYaz8OBZz6xmjr6C3n9zyVq8Kz65hyuU9iZCz4FJd8CD
M5wRdDOWwfd3IMvZ6O1lIbzi+d1ImJUb5mtK7zugN1IIjoW2hB2x8VoYDnDt5Xol
ZEcfpcfC+QC4QYCFWH7arDweYzpbLTJjmepsve5Q7OxrtsbcMbDezSUqGpGIWWwQ
IpaGl1zja2ZiAJi/Mu7XRE3N+aIrKH07yGz/NB2gULP2Ar+TYGU7bIAAvFua8ak6
ENz1XbiyOzEtOTdMF/3CI+3HZg3WeQAU9T08LbOCBxzLoqskZ+gPpHg31AwyZ4qP
nWGjT/Ey7TOxM3pzP8DOwhZa4Was6co3nLEy4xbxAKqbCdLR1+dK2e1NJrNQnbwO
DdzXbRdydkf3c5n07KOoGo2gPFVCPkSrPCwU5eP9UFllyrDsJDbcVe5t2iTHMWwX
XsP7gqDFraOXVQvv1iOPtvYca/+JYAx4oSeYFHeShg6xAfv4yYImuCp3zxojro52
X5Qp4xSWprG+R1GTi6pFLMMUzOir4f+Vbp+Hl0HVmIcbZzE8WvMBksUKWRo0Wibd
KKSHmdTDRwZwe53JqV1RvkdWkv/Adc7772qQUl4dnItdaWfZfBA/wGYxCfKp834d
4+bP3m/24k9lmUdbcfkl9y9qRGoPCrOCRTODGOePkR0Gso1N6+oip7zzVwgFFuZ9
RMRKsOQ0dR+Y11oXWfIMU1W5pTMoB8Ix7BdH8nTXBqa263774o7vfx7W0HtxbBAp
9PMNeUTfuI1iiIToJtDKmDKvPmkMFVTbv+cFLyz1Pb4Df1ZJyG6sUnOO8/gnExG+
fe5VQWeXd/E0XA0A1OyU6cTUmdX/P5A1l7R3+aTm6fxoNGEpW4RK0n3XjuHHtZ3k
j8kcFISw010q7JgXqAzI+zlhDu1DvGq3lLtVb5HP1AFjkfjzG3ipDY0AE3lNtIpL
dqcSmQ3V4ZKLRVWJnjVacoIpLIS3YnUaeMo0VM/ygYX8cbnasVHwfy/U46EB15u8
YHx8PuRf+vuxLdBwEQ12S8h1lR5zrJ0x+5YX4sFci1izQazv0B6NR3dhL6Xu6Vgr
If8ZbHImJu9GseXujnJKBvBO/jd/xpeJ8S680oTlFkTsyk2fbEqf3A86dpjzvHW3
0PIrDHK7jHyjOnaoDrQLObofyLiT+aSe7NIK/oTbG6gPCAHgmvzpEgvWV7v+IS1k
QgipHeKmhcOqatLf1PsFUGehye86dbHSmiUOH5qwoL1s6RNeQdAduZWV38TbH4bx
1m4sUhrArCe6pvbMHSJAosey/9Th0ads8Y8xATpGaNU5sD6C5+/51o8o7JXmW/Bs
XhPBl7yP3qbwaPS+mIL4dwL8sfKPVHEJM2KrA2nbY5D/W9VnhYj96hGRncFMl++g
y9DB+hWxyUu7p+l10sfLca3AVRUlp+zmo7GSnHzL9HgX3uEUBOEUhYXHfPhuIYpf
B1d0WpoKRqJOKGbMH5J/ToMDSjAygJbArKQkNcZe6gs6AuJmQ0R3M6PJCNpMJsVo
5tdeHSnp63tExcqg4aGHSCpeqcz8fVpcmNb+OqnlywKyhTkDkfWlWySvFVZSgEWh
ErK08fHxHT2ZZuIW1f83GzxslhJC2PXR18ReLx1s4ka2f2TjJ/KrZQ4gmVU3QdqU
TxG9/BIk++x1bb2EYzI+X5AckQlbeql+kI6x57cF604hYS8mpw0XecdAQignUvM4
ywJq/A4DH7NYjKKwez1D0/WgYvdAMU6PiNL7nf/B1mx37A7Ei9+oSRbCWaPAhnDH
CHEQehLqK1D0Gg/S7Du0sbmxM6TvopZ/YT4/OrE60OkPDS8dr/kLw7PRCfXwFK7W
cNTtnVibpKU9w0N14vz8AZGvJmPz9ieDSdkPsX92fpYTOoM6AHiJ6rDLJd2exUrO
Qi14M7qS9O2Fd2MI2D3HJq9ZYSNZYzvMgSA1Z5otxsfLh0iZHLvbmKorP8Z8/O01
NzXf0ke4jA+rW6ZmesBb8Gg9v1bJB4i44y6wjBe0UUdyxUN7Z7eMkGOXSmet3TL7
eyHT7h8adhFRaJt6RGlkw96QsELuMJ+jaZh82ySyAvneg8VWkubB6iCGnZGff+ld
LLjCL2sp1dm8p1v5bnX5rbpH8gFrH2oD3YaG7vS/n4PHpUSqpBHXwInYNtIN/ZTY
/4TScvwjANv8c2obQf3iwqAxaLmw6HHN4VN+gvRAAE5c5wtblMvhWQLHoLTYBl6H
yI+qSmT7mFmMIy7SDkr3HQQrQdi5N4h3GuSGVp4W9WLWIl/E1OPfh1wVKVM8QjR/
aiVuHeAcTxwFT+nv6T8d+yhObtt+J9w5wHcx4DoFqlDSGK/2QeAW85OP93UTBRoT
Zz/ezda1g/f1X6rUhhi4tWSyhxUz3ftGWjYFEOrY2Yrw34t6sj7vxaPBzexNOTYj
HsomO6+cDJwxG3GsMVfxOezFoTUk2S0xlJF849jLXNCMZXGxRPgUGZi44tgIysPV
HHkrJkDIfwpxCoE+owIXUqiqUrnQfAVqxmJi8meA9yfgoqVUDdjDma+ZvWva8tSs
NumaSXkg99TbzBtyR1nYQw0LoH6voi3t8OiEknYlmqp04wIxpYAJt8gUxgsSjzG8
LMmIdrhlJCxZ4ixlqh8EqLBuuB1uwDY60M2ycfnakkBcIVlY48Yejxrm0T3YWWsK
L+5kxtFUhw02ENkMlJgZACiMSj079869DdbPyWbR1PIQpuSObRY8AmBQxhAaVr3P
EcFcQO7xm05aWB604lkp5HI/M7YU2kndNmEy2IhgT+6mdxWiqc9BZCUIdDSH2ahX
2AOuDbJ4rahVbGuucmzLxa2H16swGv8W94lrjzu1FXzXtEPvSq+47lXgIQ3ZDSgh
nfio3M0QybLDjW5t3IOxM82zxXGl0+ZN0m5oJ5oti2mUxcx4YCGcLgCblJvci5i1
2HJKdVOyj5HIawQ7wSwe0NR3w0xZEQwyhwtWRF5d23tHHEHZ9q6AioBG4MJKZLQG
tTLFmm7fP9Johwtzmo5aUmXCUlCSk8ME341KMEFw+1srYBg9QBMAEThClK958y5L
aSOBH+e0BtT2e91fsfWG0RKN7qacYGGICLhIwuc7EaWMU/yNf6mGyEHzSlWNe3wj
SEeH32NA0JnC/S1m/Okstj7vxI5dPSfK6597CiSDz3KDJ+umTtCEtn9PNYSGDNUY
LYtf9gvJ/glA49tzckyxATCwBJSEirVTC5Zl8ahkyxmjsmufoJlGHMa3i2SO4U0x
qqjs7oz8ADkwF5HIuhc8qjJK0/b5YTzJSnQde3D1zqh9csTx7Qmoyvgi2GAHROzH
s+6mGYThDHWuZ+DDpz+P/qD0jf2j5HaEHVJl84GD9o7Gk/QJjrlihYnWM4TFbqjH
x1qTdyE683g7D6juCfPpBVr8LVbIsYsG5z8oZtuX+eVLgGVhLKcjAYo1C3RzijnY
SrZy8WUFzqxOlUVvk/Bvw+5y6rKws5ozy8hIJcWRM6QAKCExgW9ApX1T3MstJHKj
na0JNpM3/On4KmSgjz6iPIuI7MFitZDaV4lLFCxhHky8eNdhzWdTYN6bo7iV2OlH
Q848xltorFX+OvZ4g56Lia28zukcug6yxkjB0LqxAAtrG6rX1pqBVvpUBLNDtkbX
mck0HAhfx6MK9R6po8jr1P90YP8i8sPt+Vb4JO7sjI7WTF8+g4ZMj3otxDA4DCDh
Iab05pI3X5JpDz4Mj70VE7guure9R/wP325BBOuxIkfEI6qHKqMBZZl1U2HBVrDB
3CMouMFd/7pP/rvJdNYq+HObL0luHKf5irIQX18xueYGtGZYGx+Mo6BXrNH/oPQ2
a/xbqnKXoDPGb1KgguRBQPpyMGBssS6jzRtH9IyNg0aFZ+RoyBqeOniqUZ+pn3fn
7PFaX3PoXAVw4RbTOTN7uv56NN5UFOo8fVL5OcZyCrTnl/xEmKz1J5u/0xsJqDJq
CWtqJji5/mmRGykW15fgoPrYCGmivUdTz1uygE7Mp+opbWy1bXZkFsEWLBw043JZ
SVaxXvxF4dBBYEuQTCk4emBhEG0GlyGO55icwAeSinHSoBIE2gVawmiO6eyyynAp
1LiSkyLpUF9h3g29g8+b1JZuzgDPTXqJVMg9b8PL8jYAeG5y1lQcpaOVQ6Fvbf4n
TYNpN1xy+X+IZzuC4RIgFpxANp4fji05XzTafoy8UMjIP6OS9b+2eNjcPMRLYLDm
N4FjOetDNirYmcXHdQEe3bll84mZOXYMfpgsOWZIRzS+SkpDfWJliHGQ2x35i98j
Jx2m7k8RGIS1eT2kDL3ZWUX4IL9ETXxAg5t6X4HgIvFVWqDYVYriMzgV9sUPhbaI
RiCwwOkgeZW9t/WR5mI4gOIv1p+to0xBTexjnJoGON/7di6PnerZnOvf33m8JmRK
TlnSX/EmC18R/pios5H5aGiJBXxClD+8IKJd3m6ZjBpCC3Pp7IXcTO1zmNcGQr54
xvHDjU8wuRfogSqDPWFwkIYV8rXDeR5HUgKRNY8PxnXweP4hLvMSFIW7bnHD2cy1
q9VeBlm1vPevOW5xqx1r5H/xEmI63P2x6r4QyTYqa551IyW1DJG8S47OkwpZ0fIv
u1x/ACgnPwEAHM0ME3/FVF2AovFgbJzaH4iQq7kvWSIo2Dv+AiO7j1LwhJMDNyA/
f6RZkJBTzlXXj74MWtc8riErjQoEcp4YpO3umJC4MlOMi7X8J0725wIR3X+2l/ON
WL5ZFaGQ9zMzc3gLW7l+USvW8fp92RbbOadgLSTvCQaQuTYtFKyr0BRg+y1dlHCz
Gb/zfrgHBXReesnKyvY+Sfr7lxDPRIS+iDYjinnv3eFL7x6z2/wMLKYacxG1lfMb
t2aioPszKCbYEMgBgj3Mpv7G7HZQwuRhlZuj7Pv3fnk2ppgwLozGU/OIxagHeVHG
pe8iZ7eJ1P3KxNAhNhfsZ156xFjXNJrRtlNKjC/+zSLl4C0kkTpq+gY9AEYS15Z2
UlCHG++vNlcprOYlXSBxhJW+IbjOchl2lq1MssEKdGtQYkBHgWZKcbJ/TiOfiTR4
nN1jUy19j7O7bf9mdOqKZyQqgxq8k70cqnB+QLskvNL/Y3i7iaTRxM53Sv/G9xxN
xM3cB2vaeBM7FoUgMei8Zj13e7hRY8jmCwYz9GY0RuM7DSFJvXr0o3eDwReuD4DA
Sh+WQ1eCbudRDesaKuZAheM6//H6sB+GybUeL6TardN+mUruzeInKkSRNwqca7dj
3HjYDJMes74y2r+mshDmKSqV/iBcOAL5vlgMUZCk56Br7bHz6UHzborvBW2l87ix
uEgA8ZzXpBSruKMtDa4waUvF1o1RCQiG3REbQUksxrILhTjahShNxweH1K9Rirbi
5eJmwsIk2UrqNqc2Wqppc7VfWqu2ElPRcfp/0Vzwj9rq+stVyABMFvRGddV0ImPn
aWPN6Fz45eGH6tS11z4X69U9xhVx5Z6L/QNNVpJomqwlrNwQMsYzO11cTyOk/1cS
rdnuMeQVHEN292oAfPcuxqYF1PaU4q6Sy6vijJbI5bs0VlxxbzV16268vIyKvT1X
zCKYwfOgbT55go9JD//bC+lmUetCsEJHqREAlShNU09CVLrY3hSEu3rHUkp/Lgrk
O6mXY/jkUO9Jv6a7MU8L1innMUOxGYjn2BA6khyYuNNcWaioeLEmKjfIxMlAfIy0
IwPg5w+M4hNxiaBrPj23vW0ctMEjmaHWc/k5jw5yxexUyR/Ne5Fi30ggKf4jMbqZ
K2FfNg+qm1saLouX0reGex4p0SfKAAPhA+WbTthi/HpDgoewwCbBUMH3Kt8BKvq2
B8TXdt5sm/NFmksB7HfyPM7to0sV1Nxeado0TqIKPeoKStzo8hkVchCDxo3cgqOG
863mzrwjJhV1w40WALkGnDlxTWJiDkB8Vdj4oO2Z0x9f71vW2zrkQkXOg7Mm8sBW
0mor2yWHkJpGkXJQwZpiy7yEm/YdxUGXcXHxTHrydDwcul3cW5vKK3ARswaFwwTe
0Nw2pndIWt0NQpN1iRit4LkYig1XECrlBGssCSAPooFWkY8iXBghObWFzL8FzQUy
RKilsz/VEf2we2TrrmAkONcNvJUBR4YgTLOkNPJY38bUPtdsPSq+vHlv4mJL19dz
CS58B1Ght+2lzhfuskrVVqczPnF83KPQmS3eLH4o5bQlZ+UgAW8ZYroYJ6lYARH4
lhl7eI+vKXlcn3MMeDMFIdTGbRBOsrZCWPVJ6AIGvkSCb9+DBN3m4D6sWEqKzS0H
ibVlz3fiWXkeUrAb83a16+qt3gRE7ORXmClVPfsEMS6i1rIdy2AJRenIuhYZOLAU
k7qnCdymxiMsHpwwo8M3QuHHWk4lYH9MzNIlD0rrPnNMxj7ja67bIbMwT6J+l3bA
QUvPseZ0i609LN88ZdwbG1FsIHNxjkALB9CNTKWeiAwmmZldv3IB6IwNhXtxiLxB
xO01n/i6MFRuesLNWBscXri4ZWiIWxwhoYqSEl3iwDjXXKOu8pvZDZ98doQ3NQKj
xu5Jsqj2jwqimtKKEvQsNNVF4jKRWlZTcEhCGnPVEpE7m3fTpKsNXyZKblhmmLy+
I5yE1PbHXtE4hcmwMHs6qFPDKlWlL1PCS+q8zRvmDM6zS69LguVTgR6ybKR2wp7Y
Fl/FFEqMmjiSjNSM1TuJK00daAJ/3R07rQdZ52OhEuWpefTZarZe+FLNTWo3GiQ1
USRbNB6fDBznmh5Ax6Ti9+AVEmcyL6alcV/01KnrdnVYznwemU4jAVhPieaUc/oI
4vfkHpno7a5+FpDRy27mTGfgVpZ6gHJdEvSfudqom1euvn/nRkedMQ+0/vU+fjeR
0OKyp+t2WtOb/jtEp+GU1jFCuh7XMMY35n3giGUY2vY51PjcIodlYDX2AqI6YnmS
adx0tHjEIq6wlDY9FZuadMrNdQJMeofiMl4tooLuGJLaKGfF+npJuPRJi/r4NbRu
pYP9IOFeeK4bfPtINWtnxGeXWC/F10jYFiUqL6V26riCRGAAFCgT7YAIz6WUhx1n
2FkMluuxazL5/7hC8R/r8yRo1U6d1Ez5qEeHE/4q+tLQlmSw9M4ihUfXVrp4WJwm
HCtFilfZ8a7QiTWJJaHTeeGEc4P8Suixiqxv5qzx8h+tfNmmcM+KWBjhwSSH4d+b
ztSkR11QtFQVFwgJDacWXDdFx1U4ldNiT5hdSvkE/jt7sA2WVjxNAKTgGR1TqF48
SGWQy8iZN3xJl+6fZh+lUP0HFJZEI3kQUzZTIypgZ+r8VC9313zviuDrSvic1hrQ
ZB6q6kysRhjA1txwYRYhRU0yyPSMxMVW0V6OR4s4ssmYr/7hnRvpQmV/UKajSqKp
bowhttuiaMhK6223p5fNRp1P+Idap8mTnAjuHzvKZRTf5+8vyyu0Hfjidj+kJHNB
osUb51JYQKJFaEnp91zUkQI37BwkF/ZPsPj+G8slvdDR6mHxAFfx/f/v3Tp1d1PQ
ZEo4el8T0MmxsggzThkU7W0T1SDzzlIGy5cijw5F8TqVNLxRA75TicH142Bsukg2
l0Xst4bFE/MryyA2ru6WccpgZJTrkNcX/8KnN6xkSGxx+NLUtrOCQd8tG+JFJC8c
UsQPDDkDWDbNWhz2OZ2ZLJrneaxG6IF4VOWPnB/XnE3biPUk7bDpL2liNEyOVpBw
j2kprFvhxnDjh6/QI4f+YRiQ6lfqBYi77GVDz/vbDvP+bH8q00KzhRT+1X3aijQe
Vq4jl+2dtY8K52pbUy76YZDRgl1L/IU9/P8kJ4APTFCiBw8YTNWey7TcOpZ7EtoX
letGV5fPJFy2IylQyHuiW6lb7ckBnWh1kijq2jy963+97A9IZyyaGrDJmB6U+VQo
+RKdEPGJkdzJf7HujpMfmdyvng58FJrbuIfbtOyaAPXqgPVtOb25ynB/e5llFE6o
pSkwyZ/OVisEz0Ar4Lv0joeKyHl+zSUFlt/1ENDmQDzV87/Y0rY4y5wwiibqg3KJ
lVWNzODw0RUX8MjfrtHIgKwFSQJ8EbtxSQw61xS6UT4TFpldlayimNSvNonajoP2
9tXKTV5lyK8rzpd+XE5F2+/uE0G1jwbP6iuHQSIXXL8iS/r21P1gUW5IKkgJ2BZf
UEDdpV4Z0/Leba0NCPnQoBtDKBRUmrSUnojIsESuCL3mxOBE22FB8DWIA3S5QXxq
nltWAuq+prfyTVwP3dqKeDhpvuiGzUS9hIHPgpgX1TF5WtWE/pHFgF/zblM7SkSz
De65m80M84ZeoaaUSCEiqhxtIVCG+3/XgEzcstIZMBnkUEXFKFu76+JyNZPTCKzF
Z/gi5Btx9YgJ5Ni2rE+DcVUvWcHzvbcU+Na1Cyv0j0KgGHTWPrJQxgrI74TkfJe8
KuvM/flleqGagk7ETDkYpBErpRRnwo8FYdwGITf099dQzrL6lpPBPykffZLZfjRp
zsqAySzrbyBbYjD43Cl3CSgdb/RIFZ3yRKtVJ7iVl/64GNWFQ/fdILaYpJncnQ9I
YXMbez1kz+J3euxJFUciFr8p2ZKn9IH2nF4XWGO+gAKHF4UWNi9Z17wLXjMfPh+1
zvDhFo291nRwerhUX0br/dMbuYOtMkVjm1wVvT17DYzivCCLhl8ARBtXlW52lxrl
0U0chfRQuC0bxCmy5J381Y1LX0XzcAZ7po9h5j8VDXkNEFgeImVspCxkeqsStjLC
1NWev6uc6Uokq8q4ZWYzbBOO5m8rzlLknHqLErHRW9T0S/u5kt8Iv2KBLUhlQdoM
FhFKVNLVz/WWFjCYp3ueztOpXL9L8ehxDVuV9nYgI+Uzxf0/i6p7AGWlw1uDUW9l
qYjdesCtCbCi9cGyynhaBBqRZ2SKQtXu3qf4GauDJ0tQ7zddrDFYd8J4qwwN/N6w
+SQWbh7ZBC7TkClqXwjIaFuVsxGWA87Sqk/VQN1XRxqDiQQjPZHjLegonowu62Pt
4SxQoboA+4DkZCX9ZL87OgdU7mQXeLDksZnkWLkJY1WcUsqLgAFU2nhSbmbNeVNu
F65S17ZyJDaZAl4A1RclL9DQ/ivLOEEuIlQuxf9O9vAeNcDRN3+YheNJxZCs5ooW
5rU/G6L2dEfRZlEP1FhGJEKiOEnym9oDGUj+8kt3+CGnXzsPPQfOWHtx7szZ2EU1
v64yu4itV8GT+WUcbXg/hdg0rkkWcT11ba2n+cBz2HD+Fmo00BGXAhf34aLdJSgl
1ZAinhYBnYUnGla6DqB04UKiGXtbypFZ7r81etewDHDxd0SXh0duhnyhHGDHCZuJ
2tjf7KIFpwU+FWsbdT5DPbiHPIogsKObp7eeJA1fQI6QZhN6YGu9jv049R9a8y5K
RIpbBpbcGqKJecN7DzUb7ci4bYdXG2pltINka9NVoTRXho3iAFmhBD4xKzbedunX
PCsFCnF/BvgaS5QJTRgSMC/ifS0Hzu2BwDTEpVQYdpEo6o5pUtzsCVHz2UpE26zH
HCE5xofTnPFnmvP/u8l67ZVqiiulAKvDhS/q4v/4YS8tfMYmVaLdxm/fCs29Jufw
mVB98GQUTQtGzNfqG6i/L0rE22vQjt8qldI9cw5OJnUsqy7Xa0X2M/VkNdeFr9NL
6/NsWZRhjxNHamuAlmT3aFcwBah2uQRnSMGbLYUZHUtUxEKP6ThTZy55Ghqq+GUr
EuYNzOjHM0cw0KcgJVReMJGR8GZiZFyAbg1gZeljQ5npTBSssVS9Mrmh5d9+xYu0
8BKVNGOELdZbcvCW1pgqE9P/1lP7ixmRAT+LCHPEI4bW9z2kA1gQJhyQLxbPzkhT
Q8wD5R9gbv0zJxVjGgIKuSjwBzlMK6rZOKMLupcynIm5vRui4zf8NOP4VX5hA7TN
joBQnL53E3l/LQU40nuw2PNG8t+Sq14/Y9L2x12Jjd/XuHwBNSXxLOKVZ/iFdPGS
tZVqkX2FIT5RAKOFm33NcAl0n+ALvurH4n8zVflDx7JY/HylmRzq3gfVcdQgNZaE
aZq822f34doAXJYSUSYr3sJQsSA2U1JXt88/+vN5aHChnEBoI3m1HwE76mrs+L20
vKKi4ya1Qtsk8hlzO4u7dawnoeQBgJQ578qCHuhGVnFsLbxY51e19KI+7vKECsLT
YPE9djLiNN9IogL3+j6RoYCPOcNxszBZJlpLdQTPpdzf9I8EWZYxfAKhVyiCX1zt
7gnf+mMPD8ryYP5fNY6CCPePB9b42K6Y8IS2oihJnPgf8nGYwDXGRQetjMoUU6B/
iJ1ZIwWtIQ2NFsb3dgad7V2eZ7UFzUGambcaJFU4IDEEPskxeLsjpNK4hidw0Qhh
WQb7WU9osgwCGnAriRFYtKOAVGCEXpTHjVK/pYmjh2Y4i7PCkwV0V/sk0KwcZ6a5
3WKjWoLwWcVZPOK3C8Ms1HwEq6MLVQEwLDTNEV3sxBTEv/926zj4qwLPLpYCpqHn
DxBDeoA+NtW1l95f1YhE/ejDbNx+q7uTZtLk9DpyNGYAZ/wGhNKpvt8KX482V6nr
KENn+Z69oD88krlsqwPtX7uZWMUWF6lu8xROU0qqbx27QvOn9KqhsB8hBHjkkKjv
hSY68ytgLIukPUZliCsQyAlmybWbAXMGe3FeJeNrdGG2AHmxJ9ccnfqql614O2Pc
g1kabBMKDcbAv+dB3DUKsCjmr/i7pKmg+uGD2JIbQMbCYLAuV7XAht7BaexR2IzJ
mmzSyFoP3ptPyWCbusKbr92v6LTcO/ceO7Yi3q35XKnuC3zFZuUwi42Za+5A0jr6
VMtOaWSD1sOU3Pki8hQeAYhLVi3lm8ndxlez8W4t60BPz1KmxxU5+v7KsGRiHIR7
wKLm5x8Oj6UeseGDYa5t8zmwYWMs6zna/6Fxm+CdOQbP8eyqC6VWGxYijXSgpcRX
+SYTXmZgXx6HqW6wRBUZ8DpWCEc2tmEyoUR+/YHy4y3bQRJyxzv8buQla9mgcMrx
SPP9v+6sfOlD9bw80AqnyYvttUZzdfv/WZaDqswA5Tdqyc3L8sE9aJhAw66weLu+
3vX+pgiYPRtM+fLU26tZb+zwRj2TRP2MLbAeFUcusod21Tcg7baWlmIF/qX971bj
Gst1MF9/CMLS/pT7KLnPRcMF8RP5QxXTJ2JgXDt/yHKabLiCjPR8ppuCTNyAoEqo
1bmkA26b+G/NzFjGjMRbNu5ZPyBTzOIoNRgZbh2vRcS0pnkl4Cs0Tg8e74Glc6m3
bbHfejJPVSz/UpXJ7LVyRs2jTOSt+ReEmGM70HAROZ745OGDstnq9xras22+miiY
Aj8Hfr2z86BfOwiivXstrRHRrkl6kI2aH8WS3lOlMW7Y5mjRGJqIonrqcCTnGunQ
VPvENaw/5/MzH+hTq4gyLeF+BFQli41kHb7RDgA4tmITVNpE0DM6WrUnfJ+uO4QV
FaK9ApHCcMCIOtWGDkbb/Th56r25ZuStxbf+ddJol1a+VZ4bfaPtZmlMOd+fTy6+
OdzMBFH4PKDHDxGtcDcCQaosaP8JZ3XlDHJ5iu31uP5dTtegCka/Tw5o7sxs9962
5xUEJt/Fh8xr1PlFf8CdJl2ubVwTolKBZj5Vg6NZnNANuhu+2OIpcxlMlRkvZ+c6
C7aV4KddMR6RbVr+Snj0aUKnLOvKWJgmn1vAZVt9w7dqrcJBbYcZASTcdmUplsyZ
V4RpgnNhzeLnfEIZpp5CBGdZPf73G+FPeRoNZkoevO0coBJdmhFi2l0G6/9YysGj
4Fq2MRQVItlGPN2xZVE+s1sC+xtM3nhVNQIaDf20QscOiEPAkJMICpR8B3g4gET9
6jI7fPb3sXK3P7Utp75b30swI23K7HeDYnSlT1hVr876zVBAy2CoRy9dnQ4+vfMA
rmfdnjc35MR9gCcvSnvuDRSdeUYeLnuxklucK2UTx5s8fLmhVtbxFH+avKoAYie7
9tjjPYZpUwJE6hob8xvIlsYjyCQnViBVkiM3mxvDj8VkMF4u4zMqyVH+huFgx4PY
CXoVK90kc31lcWPOkIvPzb2XmluH8wJNjMhhlSExV9SW+/mydoR9w4pBdgbZivSX
zHKqyHj4IaCHIONO5b6rhVcZUDlIzlpOFfBTUDPghoxH2ye7Nz1bl3ZtVRjNZCKf
xJKjvXrIhk6QRoclaRUUi1Oeqp2NOf89CkkzSj5chgEBDHOpeFO9za7CMTopZ0M9
KdfzpIE/gm+b4dJpTi2XRbQZq+dEZ9wyrwIvwI+qr00tTPYOEJBnIaD2Gxt/6FNq
51Ovf51qVY3pRNh9bqzIFnEpwfi46ag2NLll1pfqqD9Cc7C0vRU8aVwB39lSgi/r
SS6i9AiIHr41wE5s6shADTo/DTTq8+YUZda/hxqsUaJwXAp4AFneJlxmjHuhhhji
8hC9o6bDMmNrAKatg6qXI9+KdsaxjZRg4MJkB1zzmME78NPb3+/AUESHpzy6P8hS
8dPvkiAVgDr+swavwUc9y9lcIpjd4Rk90zebxcbWYzpJ/9+tTsVp0V45oIHX2M/E
N0ss2sZOi48Oy+VtBVFL2vOEQJhUAaUtFQ2m5Ixzfur+6hnCUCzxlXTLtGMz5NpJ
qrfcpITVZr10UaQwhCfomY4Gz7++ALspHFvCJadqSujNHyR8o22ew2UEKXDXjWK0
3W2BRFlZyWaYjadQcGzfYPAet7Rptf34C4WcEt8YlcUS82j9CCz1eJ4TfANFp67e
wEQ31BbCCZOPhFT134imGh/6BVvzuCVGj3XRisBpMamhSYTX0+zTsQH+zSwjnGvt
Ni1LtoYlLXMFv17X7EYpI/YMCT9zoGcqH4GVSFxt3P/RSq/nYz6X5//pIq1ds8eh
iXrX7atoW5g+hvHc2knCWQcPcHIEt7ZPmPkqERhOCtcQQnXWpwPExdJ33hFO8sWM
6B5b5ggM7ok7fp/812Olm3puB4I/BGCyqqpZGDeFsHO1TlaIdaPPZ+TQkuaG1rw3
1GpTsh1BSoIiveLuJ9qhBz1kawXNaTRRYmDJQ4MSPc4rZX+FTmzADBIG3aWFQvNG
oKiWRl/2mTC+lpYNnj5Vkyg2vj5Su8j7a+RFmEjtphMjazdNBA/hsreUScHX7mcp
sWeJB4aQXhJ+CI6nfxFnzU4aw5Ix6VlGClFDTH3UKWQp/w+VXmIz1dN8MtUkv42u
4efQ3J+Q8BD/FgkD/0k/S0KIkSxPYasP3bdVCjqU7cvPV0ecdpJE3sXAeBtqxnHK
eimUrZpl4tYMqRzbXDdm2dL3EZBfbtUPeW0CxhaaBrXDMkMAfBoJWOUiSkkAycIl
bsvWky4NJLMR692Ve33NUmvMRW48HxY2CtkTasJMb++xx7Mw+M4/0ZIQQK+mQnzF
O9ZaWLzornLfZQLLEiHu65iSd6ZgzXpuQl6mVpwhKLNJZNF+K0pgmZ+P1gTkbaze
f8gU5C19NwY1i7ftkGIHujiDjScSW10kD5uJlEOA07azY/Yi8WdrzgZ83z7GOlw4
sz+Zw28OyNrq2xtCK2UK9x4Hu7xIHyfRBqsafM4k7J4y7k9y3xKDmypIpxUSAlw8
QfDWbnEL4+mGj+DS5vzeYad9ti2pWmR/TJcgU7u4onPdCciaWtRFoaKI0nNos7bj
bVcQgRon+BRP0othvGQSJDINpPWkiKvVhKOs8MYW6VY4fPRCmmrfV/NIc1cx7Czj
x/2LCH32rDCWA9KvaYe2bEWeoJq4yACZAGDMpaa3zKd6rOHnnch6M6AjCYDXIdOK
Kq3NgyyK2c1K1A52h7FqlQowmT/hTw0QbyO7pRwmQZLKhGkTyQ7ZEtDZzlsXGNpg
082xBITMQZN2ibkULG8cIB35hfS0xdY7fJfScJRvzg5qZBM0B4G738uKVvJNwV2w
fpNca3KUoHp0l+I82xGPTRivFmHBSFoYIyvi4Vl45SC7WWqzyP6P6XYSUhNqHVSX
AYmicOteN4nCzJGxO4HXyxXFFoNhDqqX9TILATjjesk0iF75E0X+/UVKe7O3WNVT
sMEpTRq8Xq+dyA47PaB/T5i3l3J5qKCXibzM4KVG/v2hWiDYX3VoTa5zKypN5ucG
bDMQo6ImbQkcqGzFdbS5tkzo6oFUOnz9Pf3IjOwoftl633zqfsuzR9jwT09GeGHJ
Ly+hV22EOLRjIeYONQXZJb4Iy4Fr6FhjMudY6jVzBVDIaScqLTI9x8bU+a8axDM7
CxxgXDytuWCtaKhTnKjwTKYJsEchTHv9ZOtknW1SImnpBc51RnRXZECiyGv6hDro
JUIv8/5jBAk3uyapdJQVKPktUWEI8/u0PGcGqGJ0j3eio0nROjij5ErqiV5z0XDb
1T/9GlWWOgDxRk27c8Abe/GmswNs59c22j8A7ONysLmyxrxdeWPdPyU5T/kwJeS/
b8+fLxaN6gMOvjZ1I4QTZo9xzVnV3ud8yamJ0mkrCG+4ZEBHjbqGSDwBQ87o7fqI
t2md5AjZ9EcTL7hfGNCdZAXzpBzN6IIbb4IRa0qlEUmhMcico/0xmo9Np3ejI9yd
sVpQns6Y1RQBUdXCflI53SUVfhL/Fgv474ovc6ljB2KtS1JVJmsC/1CkN3dfzmLV
9ogMKB5QXsV+seOAfV3uRpS86yR+9lrkNG92xSpDKT2vHtyApJWTDodis6oWUI//
eQDZ7nVsNcyr6ojLLpyNyww+4XoE8AJ3xKMKBxS3PP268wyNpMi9NQd7v7SAJ02W
m34qFUSG4Pncgwgtun+kcWUKV8f1oy62oH62mes+++KuNVWBitnBBuhbeX/E9X03
TmL4l37DX2PcbSGDG2zo4+C+UAYI08oeoWjXvTNC/lqFMeaXp6a92+hGroC6jV46
mU9RivM6hQ2++SG/dRBxG9KIn7nxkCN+QCt4qMb5erQpHNXG0gs3MlUQ0BP98nnK
lhfr3SBpgRBbtibMFAfQdlgxCp8HBR5JJRlsRuM4szIB2ulffGq4oQlp/NPZNVfe
5+PH3iN2J/v0usT9C3hc0V6PfRVHw1xvaxeXCU8A4dWEBtDSnKxrHpRJuv77zCuX
YjezLEMt9ms22vzbcJK9ym7L6Ce2SE52RGiNii4EOguhg26hgBbdchzY1stxDWx+
XCaaP/BChTeU0IYaMBRV3AWFZlSAtOGpnf7oF8C0/R9TJvCfNB+rCNDm+1zriy7G
0AuMOowGBM0/YXb4rB8tcVw4cyH/eYSktGaUr6kRolgoVLvgFiRZFLfcjuy5atMj
h1+lCA2F7GqmJuLCRpOA6XQSrwnCkm8ugGO0Cd8bKqF3hZGFErs8IzhwQvN8vfHB
EhSuReAFUtaUsgw6yZ4+525oUqhDMFyer1H418IOubu6fzQ+eIGjNbi+PCmuKC4d
61POvz8u1mj18RGs9pNcXM1bSdIheJ1dM4Wqxoo51jZ672wVVepMCx1jaNcJXCUh
1sgwZfgB7HPIQAJ+xECo9qp/1JmoAAIjZbICKAKN5OQ4Xi5f7mBele8xvC9WdgJX
HEaGlXmnGuaQpBoEczaSjTnWio1gTFWuc4dInAFHMtcNRP0VnCLgnFGjhxFcCNRS
B+IoRiDzwM+DMXnb5j622fU0e/PgrJBKK4fdS29/KSEjY33TLl0H+7CIyNUrzuAq
V7aWCCwNdNDLMJWqbGW2suqbNH1S5DQu7CN1QgNRE/V1iJqEv+vt/olJq2oSuTQN
vXJC3n7KK0GnZNpHnrJrZN7iwWVufkJtcinm3F+H4ASUDBwLFlJ8afOj3WN+8KR9
GQW7HUB+z5xE5W6zhZIUr0cIB18XvQ1hXll7swLQLyQyRYTRKHoHODcWFozqfzGW
rcWXV4SyvwlpSUELn4KgIDw/KzR224dwBDTV6Tb+zE5Ce7WoQVnFdhRLeOL6Jn/g
pbSGyWAxmshrLgu708yO8Zk3ZuI7lEsmskaGtFZW05cOyIeraOEsz1rLJAiH1VNW
/Ci+Ba2UtMfhvW4q3t0qNNwCltVp9dPfEyUGT+pxn8kmSDZle0i6W00vxvo8kFa3
Ip9mj4smKQYg1rpPMmxaCdjxzqXTBfSxPOPNcc6DzI5J5w71lFiFRhIGay2PQhyi
JRk5ALc1o80BFkxY9sbKuvR6eXfF6p0jk8FOg+QLDKy1VRxvYeNt3r4oBfOInWf3
i/DOIIISBCiGJulOyfTA/uGF8DzmrXtM+c8pkEGYwEkPt/cIg1kfijmDtxpLvSyI
9WH5vjvZrvwIHVOEc8eZYH/YpDO5xKHLfQZ8xjr9oMuHb2Hggg37lScNHVg865vZ
FsLxvxQmfMk+LUEWYdPq0cFFRpaAn+gssh26z3gfiXBcuW4/wnLljLGt5zWxvWed
GmMWki2ZbkSQ8gEf0Rf5iYYVfgqMwRgz0jX4SmgoWaMDqmdc736f71G+I23W7lwx
UpwOZxcCVOSgT/o2KXxI74IZ+fJU7THmfAifq4TXp0qHAk2BVenCJK4L/yc+CEqt
ilVUvxkiAl7SeZvUKxPygokFcWE3U+bwByPvwbkLzq6h5ka8F/6QvUoomptwuY6x
cLoIp/Pg5bKEQwvNM3QI8UOmTZmtjYI619zXssjRZEtnurshZl4MJZMalrVFFr31
LfgYOM+mYKegOBNQTyyUYXDyCWpkS2AdZcgrUMO50b/z72+g5aMNCOAbhppJOVtY
LXiKA2C948SJcyxNpxD85SxyonyhzXlR160kj0J7Csi2UeG3YuuaOq0A39r5CYEB
W+6sGindK9EQJrY05OdifieiU8O4Ab7y41j7ea7h6xqlM5+M/U5eQJkJycPezxI4
meQM+/EqQPUwYFqLF00huqV4eenrcAgEu+1jwXkvkp2vdCMbEz9kHoVak5P+H17P
w1mplyrrY9ktpv/LEGeS+HDj+QkY0Y9FNUfMZY5SDLONn7PsICdercqlK0j+LT3y
Qzcf5MnKPfB9AJH10rIC02ZSjXCA+BNDSRm3V/+q1fbmFkGmsEvXpLnnBgyPML34
LmMdVS9+sqJZFyBg0iwKN57SKYpev+iAIGiDImLJ+8oRLsr3bTicL9CUvfx4sypa
LqBZLgoJG+VfG/aA8vUwEDjant8B0Gpa42oWm/uTiIPtqnj46044RDOdVJ+gbmty
fK7OEBpCmSJcr9vbHqcmNqq4qJTgAsgDzR9hOeEVGScfx9RBWi98WjWxAbKcnL+c
X+xoYac+foNnLsBcenN/n/7Prk+fNJmKor3hshzMuCuZ22iVADSts80Bp8QB07Ur
w1hzhFuHHS4ayv/Vi5HUvfDH0jLssISyE502oQtVJ+I++1kp7zWhb0ZsY+Xg2ARC
l/ZVmHXWOItHGV6gxOiLBQh2b4CZyqZD84i0baw91NKoqFtSHuICm+A/xedyMHt7
ZmQ7xvyhEtkTd/UW0ietv5Hjh2fMSZb9z2x4Rht2K9RD5r07I4hnb0Z5I8X0ahVl
BIQDIvKqbHlAiyNt+BBibfOvmcJnr5XPkFfrON95y/vuN4amtFOg8VCLCrA+E9em
rsw3BiyWkqS7TupdzoXHOkPfM49XgWVuD2qHGKz4CM1LHIuO+qe9ZZCSEHOMaT8u
nHNbxEMdOrVzT5RQkTUFobzS93qDwfL+SqEt0DeUaO5jKQws8d8oe30PxVYJ5syV
a2PQ3FjaRTkUrW0lUxmr2FRjSWg20JToJZje+yBuUYwn5LK6z00BHKZkfPNoVm2w
0exW6r1g/aH1yvy0KgBQwatg/VEqooMHOnCptZ7AwOkw/Q/DZuFEANVuj+oOc5F8
MTOZ+6a6hsMd+ZPdaP6lpJgY4HQFKZnE9nAipem49GkvmD9jjBgrXYftOwahkxHG
cdGqe8UOzuiTr15A/8mM/vQ8uFjwP1jnW/DGfRD4Tt1+6H7bg9HWL2c7yVZJZ2It
+ZXbVD4Bl2FN9v+z63Z+U37asriLoWi0NVN/0zXtgWHQz8obsa0pXOkFK+DZz49j
d03tLQvK8DmPCoE0dDQ00YrZXmAfwzahwIoKQO2QxQhLcq+GS3+Hh/oyEjOD90rH
YgPu/gzgxv8sNzHIkhGDJNmLdoM357/urt94xNkz4g40DqaUTF/qSA/KSyWFCoJJ
/EDsRY3luaXptNPkXE9L2V/FTdZWZ38vTh72dlumBh25ArBzBg2t5xTIuMMurTdr
n/mD51WGjLL4sVjjYhPFG7zqggNRJm0gBHkskz7Id4BTedUw6vRhbdhJgflHBFQv
ylKOgWmczJnFr7O4VCzQg4iNOUBlGU3l2qZ6mIu+a3mrmq9okL38B/ISmU04GYdj
2V3x/9lBrrlUTKz1IG0SEJdSxuZXcpBuSjvfg9w4/x6GfhqyPgz8vhRSCmCBXw1P
ytZCFSHXeTuXkZc52EAHBWoDn/k5o5HvPOQzem9GuDB24TwH+G/GIkX1CYlLZOnb
6SdIVrumBCPaoiPW3ueirY0PyqFNpj8Km2ooLcDkB7f9vo3QDd4WSg0TDYJEmmBo
AnBJHR30kb2zDQ807OKUSrXjk1zd7jxhwBfigibrci5W2syOtQehfarOvRN0/aW0
vl6LdtlFA3a0804HsmcU5Mbs253SROea269b8Xa8QTeOous8dqaJtvFaN3gP9WgF
jhUoOunYcRQUK8TCF3RIiLokITTa3ro5uodpZN6drBZoO9DdMEx8QWSp2kPXQPUO
AQRaAqiGpXH/PpeyIq4rcq9113qiwiMOEu0dxs24XBAJuKmUi27scfNdcrJfI232
lcuH0lX/GgBifm1LUB6Gn89yUr9+TMBAbKPkubZTfH2omep5lqRfpZj657oKY1wW
Bs8hju2Ud0P9DQ4C6zekv1rMJZwjiXX3fExtwly7lyN0N2tDscwJIpAr0s5di5bL
HQ0x0tSeGxK9A1/hQPSLP3PcHwA2ZmV+05/umS0H5/GLoLCroU4zH9GoSUj8hp+Q
m7RYq+5boMebCWWBZcKkv8OX7kURUf8LbS98RDavw4EojJi2Yqx0CfxWja6fP6JG
tzNhF/hOT6lVpEfTl+IDZC2FSLqvEnA7+oHfDUpV5Lh3E6pCvBQCp3zivpoi1nmE
fwrro6lahWoR08Qbw0Lc8fPIkmItnUwUWaU80/+192uHRa+ItBx+VfGlIlEYWbWc
nFrzeQ8ui2BuErugZlcbEPxfjEWcrfw0JNA30dno/8SKXnKxeWn7Tr3KTXQRnafd
ix3DTIoC9YZArzKgqpmcFDP0gRcX/KdWfl27ctaUFtYdYHdFkAlnwog11qhzzng7
TitdhW7W/nM4KOG/bw7/i8ydd2dCgS9Jy9EOFLq3+2bTcnC8vKsCKyMeGICDTHsk
9r5fKRa0+3akBxL+DEvtBbKhKmQ3GqPFz6dxqBAmA9fd9b4MdtyI9TZJaWj7C8Xn
V1ITjRBdTyWPVik80IiBSpGBCox7BcSkS4p4Z3yWN9Dlst5VHrBA7IIPCxhG4o/u
0BbgXkKgiW3TUtyZRJrp/54plaLbqNinJ6GP721vYpcmQODV+NMyiQZ6qZG8QWNd
hsbe1nhXYqM7yFl46XD4pw4KRyD+MRkCFBhFnokbEvZC4AnbgAsJrK8G8jZ1tUVE
2AjsaAXtoynM/KifrE/J8odfqNRy8C4O9BvPCXSFoSJU0B7Z1AAeuHbKtbU27rHT
bUeH+yEhfasfGL7DlwbW4uzGk4nlqLLnqmJ/exCC/YNG1174Adukf33lPMF27AeP
iyFG29OhGnt+oWDZOpe4gGVvky18su6E4HOXEIvDh3uL6sIhllUQ8W0VxiVbWY06
QFuRcppRDBz8Tsohssh9FR045Ih18TzWFUHxj6nYkSltw7LEjgixqyepxE31FFbe
uebaGuzRmNAk36FpcQq2AO/MmxuGMYa6sUI3RpbnsVr1xVMV1zZSTHy2QlMemOnT
ZhhUvJYRT5ODj5Cs54oVCrYcIEq/6yxqGZspt9yG2q0M0M0xZfKznobwkflXwxl1
IWeDOMESwpDSR18UrbntPEuJq5wjX28XvxNlsY3FxB3jqR53uMwU7Gu6zRxne//z
mPBGHpDqtObPdTK494H/xJ6aByDGUQNdztrdhbIaz0GF6IZDBFXr/8llUHb1Vt7W
Za9jpZYKEpaPEIuydRU8klOG+50cpBWIM8JCp+Jk6T94FMm3LzvuFfKcaXdC/G37
aVCYjHDGMJxexo12BRLD9szA6DoZSjjvZVJ5oa5LNBp33BPh9zXAkEZlKjM/ImAj
WPc2++aRf5x1ZnaOwY20dG1r7tRFFQNfA377ta3fGdfr9AUi60i08DBjRwmyW+Ek
If3XOO8d7+TdSpBWhjuB+TuSIheJAJM9TdbRgGINq5645CIaUGOZlRy9yBUx7EdQ
ENUsUBB7XKrA0FAYJzuL4QGzzYH9csONkKZZdyB4PdNSHVDaf5BJI3ttzZQh3Tld
kmX4lV9vAW2jTwCEYXT7HsplVb6iNGzf+hrL3/csO/NuSJTxOMRx+XLtN4Fze9Mn
ws2sF0U7siwZlqY9EK/brK/MPgQHA8OY/X1nv+6myQ4cf2CTqJfw43rutw41ZQD5
CgJpRJEmEEmTujkWPEwk0uAFpmnaUxwVWbJlzJPdWDSPwL1mB8BqMhObPLRvU9Vg
UM8rdIcWPTK94JxjDaUvvqAqLDKQ0St42EhOrqHMuNMbJPGDG8ABTeqm7T8WOMvn
1OUpzOQemmSNXtYVipnDuVC9UzwrC6/aTUnYqr9YGeEhbMILPH09WDuXPx+FoqF7
NjpwKC9dMA5nza0tUpxIrCG8AEXRYQL9PhemKbKe70ORz3wUPJt9bksOXyyvspyK
iVpDi5hxWsFK5bKfkLBtKKdl4dT5QDg0kw6LkJZKialOiloPu/2wGsEDezaHkJiR
QuHXB+e1QJoYnsd/dC/o0Ld31uP2gy1AAznqbbzhElxk6zb1gbu2TVtSoFxLzDLy
HwImJANS7FdeEr3LRnlOqrbNdF9px1ufbxt64u5FNEtDefLXKjMW7YfBSibT6Tij
LeP2epc6R7IxC3W9MJnCR9GyZ0wo1NuZm+jbBUB4CUrxIO47l7Q0ZLTnHWqlI7yr
uZ/pSBfRYrADXIudOK/iHcoS+n1B3NguiN+pqxDwCohOulwBWyKDTD9grgBxRms/
vFKugTHtDEHSW4IHybxRRU6oncjOoTmsblTLodQF3mlaw/ubd05wO73Nm7ozk4bz
c0UUmVofNM4/ReQXiROtIE7Tw6kM4mL3sDjC0XQbhTv3NRL9lq9WRgqlpCf0emst
QVLDdMUph76u3pHSD+JCYNJNl4F3Y5iQvrD6/Z0Yy18aLVCdm0JzwiTW0S+BI2Ki
vv0xf4gD03Bwp2Uh6k7PsuSqzjhQdTbjei8RGGfGgH/C4JD/hdb9/LjxIWeHXbZz
9i+8CBLbejhN7YE4SahzCMgOI4o7KCiteEGyCrkmHNcxtg5UzfR+kOxTu0K/OrHQ
cZyhnkmP9TuAxd3YWWh+MdV8XfbRG46xlUiW/s0NouQnE2ReffcM1HTI99sa5n55
k5D2IdexNLl1Ri3of1c6wE86iYNk8OD9hs2qaZOVYcR/dIJ9vqgX087B9M6RAVPw
/9HqpfqncQsQLlszbQu/ecGJe6sj+vnvhUek5zFvqag0YyVuJhRsno4Mzj98XPQL
bxcglxIYJ4kmc0tf9ZxWfUjsf2A3nfuWHB8RE8vJMuXD2iFKNHmwya/00jToYTqV
k87tkoj4L/YJlZNff3vYqAE936r/ypGbp0x+U7CPDcOmTAMyb1cAccmPqo96OQx4
ZLpf/UVNNX112JbxQU0gEkxh+2BsHrG1PFBtd9QvLfPCOvK1slcQekolDHHfVsNH
h2spWG99TYwbF+HBKmGgNEhb1BfYTIq3mmtXLk5gihEGrnHYFNFNBNUO2W/ffgU2
wjLrSU6QkWKEz/ov759kN9t5FnRjtZc5CaTxy9BrGr3VYlBPGR2fy3yFodHMcqyW
2WoRtGGV5LvBKXrUbImgfSx1Vpsw0GGcJDOegpTrwopXB+2/VyDx0GzhUx0kMTHz
lDUfuE8fW+4wllaMPzdcmJ8hcQ7s5OTlxr4/tWw57mC7EoO667KWQ04mMlsQ70JE
Xhi8ZqJ+kwkVAuUh4UzSPFNkT5qiTt7p2RSnNtNfqMZUg/hSZRXcDhPnsU+LCWgI
AEeZmYIdizt5rNxno1V8uqjmzMndR7aqdur1Ykog376/2BeNIQs7Cz8Ti4AkDCZk
lRHNWllNn0i1RbjuVVt1ArLnijg396FyI6jRSy666wFlAPtBHwIN4kGgZvrfRxeL
Mo7rVaPIoZN0DlHwzLu2+QbFmkvlH6+exQIMqFq3wKk8ofLPwf5Jl7kugphAUn/0
I/L0ULOvi5DVJIasGynDq1/cLFuRcsnQTlkvo8TXAsJaD+VWpg+kZSbJCeMk0TXq
ofbeK8SyIn9Kq4tNT0xOXsnu27QQLaFZtv+zZzrCI8Ee2sd0SwIckhh83a/F89X8
0R6Tj0NTxHvUWdsV3DGnnQ0MdelVfe6z4Q2iaBrfXQu6O7D80HIUdxHaO5Cpu81D
NoeVteEqS+D2xCXwDVL0kazi5qVzDOi4WnFMdDm/g2wvLVbS2wKDtgDQpRcLDfCl
y5IBj71hHqafp5i2m39MaEPumuh6JpJwFNkDoH/uxPCuvI7QDIqktDGZ+dSONT5Q
5eyULQCYRzGC9se8SOGPvaDYENoBUCnpjgTRHJx5sJMvt/fCSotfm8/k+3lYDwFT
5Gsk3ftUOTlhf9jfUlr4CHHTBAmHRGTUkZr2UYcMPaXNgKylalOKvpadLKgJsrOm
Q9bTe2UdkuZJWsFQZ4AC3sMvrchSotKwrphu+Gun5gy6IOKtRGbecCQ+HEXFWgin
F6vhYKENYtn5jqvfhVKKxRbCtTWkyb/dGJ0F3kuJCaCjdfH+4b5nLkaGZGLBRXQz
NsLSBUzcNATxfmz73DLdmlNPkP7+pH0CawRbP6oOAwM9QDp8vbvHI1C3PJOywEn1
3Dcbv9nZhsRmNBnCQNWdxbBR5732WY69yp5Y3K4gFNffXChm/qZcQQOmtS1MCxsQ
7vJyLw9tbQdUlf/qroIus6LmmbtYWXD+tBEMRtUcn3tG43aQfPQrES0xBDK8wMlZ
ib2aZEEopvfm/AJ1n3L40EZXTJhnwPC5b7Y6HSRIlHobeRKviYmb3vTCHrFQRaM3
GRy3xa5JdtWT+3t3eyfmwR0s3Emu6K6ZPUlAScBxEEKjW9EdpnjYXJqqRAln5XOm
ARCOwlt3mRu8TySsXHAc/7dQwYA7XaY/Dmjjc4fdDaNTQUG3m4X5t+OPWlpdko9I
uGQLSbGI5PT/H74O4w4Iie+sL1XBucFJB/Shwmbd9cd3zOxD2TecSG0YBd1bGoui
fMYzRZInKRyAM88Hs4tIKBlOVLeXm3QVWu07V5klwj3KfNxWHSUiHaq5CjUkYY14
AVn5Fa9EO7LaruyH8XM5+G/EoTYsEywrq/DPFNvTQ9Lhk4T+L77JGP7FaRKJSUeg
TxhKcG+E98KFy5UxKZjLRsVGRJVlpcLdxjgZrgNBP5s7USj3wHhK6k5DYsozEWYQ
nR2eTfBdpSa1pFxmOEjJG1vLguRg++A65mU3KsqI2E/i4Z17sJu2w2aYaHX1W2Lc
jIp739AnH1RDq3NvQfwWF0CA9HnRg+mDXqbdKcupKbph6uAa+RM6igkMPuOOzzQo
zNKZzwFJeDMFSogiaQoAc6Kdfyx+8lQogCONPkC07gZppN5B0Hr5BWtyHuM3lQ50
qHATvvUqyfoQpY/FHDmwKXvp/R57nul1rdO9xhEaFJWJzR31ckrCVW183YKfHKVj
bBmudU/tuE1oULsCszflloVN76+0sN/cYeiddEa2MzOMAuEip3XFfS5jQck5j2d8
0xRl5qvKhB/A7jKGrIAhtOWP2mQv+gujZT0h3W69IgTGxVT/rb8GX1aebgS7ELEC
+frSPWU5WltwQ+IgMjsbx2lJNDaW9KrBoFal7PfFZQhenyGhCp3szx2dEPKmCk26
OpOPXoEK0hqELl/C8R2vEt8n3jBVJ3XuuH2NVUQUhmSiAFIW9zyzDsq8/gj1Ss0H
OfGO6XWSLfUaDRql5h0gDj5HqDUq3goJAUpaPFVP7Llw2i2l0HRKR1bQRpJr1aQE
rAOQsSEORmJWe4LwBIJmpqjSMjIq+EOLVaysnF2B9XYaLuMRkTCWGyzXIIMO2aS6
kumFzPi8auKi1GzMzoP0GagnVD8CAcB06a32k+hulAF4mHtUl8u5/N/JfyIVe5zj
X3Ee4uw585vxoOr+G+pek9b8pD1uTgyL0NxdrSD45oYEekG45q89EEYU3g/20Vnp
ZkFKxwpds28EzuZFqn2SBo6xNZmzMrde7+3pCqvbi7bSQGdnEOkTsKC12smqy8uL
YExyuAF8JJazmH2x5OCn9xqaLGq6DTBnVgcRaFKJo1otT+8r6l5LKOwPGKGPXC9w
d4Sm3viMFWVMtWv9r5bHpibPYahAt/4lSmn3GWz8hqfRsDrxvyX6dgX7z7RYmgsU
PG8JIjsg0EprjqphaVlbu+OXCFThCh/fumeIASEUq9Y5ROJolSPRcftCevL6qK+E
9WB+KkR3Xh8g9kWmmiNNwGQtiijZSkLPcv3eLEiM+yhdjrqwofqd32i/TKOrsR46
I60lUsqkBcA/36EEOKtcxy/Et0DKdMob7sKfsVqK4U+Fu1m5Srl4LPZwueyE2l0A
2yR+4dod47OvgIh/lK6mT9Ti1sTHG2dwOrJJe49nDsiG0IC7zly2QC0FkbNGt4zq
D/zUYscOywuJcbvVkCaTimnRkG9hpYN/DDqSC7FFTDMqFFb+nKVTu2waKuaADXOs
XPW7Y30Ep3zgLrSY/WHqmhRtSGyUI4fL/WBOmeDZnWqjjgZ3syXF4ndmBNQvsDCZ
stBsxpLT1Y/k4qK2VG7Vv59Lrhb2XaJWFEA2PJEMbtC2Tj2k1cMOvRNB9WEjbYs/
hinzfxZud0f1leaz82+6+JMN9gu82AB/ShfhaAWXEJCcg3B78btcxVIEqQaBjEJu
YWY+gjiFEpR9uOkQ/amI9F8bxJ6w/+bSNatzo1omSLKLuka+oPEfJ9BxuZpStFMu
PyfjByOas0b6Ps6nMEoMbZdR518RqmUU7ZHOus7W+Zc5CDXXXCKBfFZOuTP1cf67
cQzA9apMfzGB12EH39R8uJWgqwOTzRD+LGAStez4/HMaFR6ilo6gJ475W0dO2eIr
//8ZgewDU88JOE8cmXj6eXM1w7T1bPnI5RnXhxpr9uUS/P1S+4eINyHu4U1Vv3Ka
Y2xggZDwUfSwla4u7ExA8WhMPDuE3S/pWwCGUDuLuwF7RM11/Yt+UHhqXYNKutOL
gLR/OrhNjJmJqlIVfiUwmRUOg3WZnvzfREkG0U31aSRC04dA5suDkyIY+/tju/Gp
xoBrM7KVipAAedEcXYuy3Y7BNJgoy29il6UvHGhg/20yrp8WWybd37mBAJ1qO38M
2bnuA8LhQvwbqCfZq6I7oWeWaZCJeXvK2s/lSuHaEJ1Qq655hRBgOTtU/7ZB4MzS
BR0vRJc0e/npcsXNZTf78jurUrhR9Zamwuay+5VbNyy3MAEvtFwycLtPNbEhhnUt
FGpD1Of3/Ond0JOn+BDMH6treCfiomFnBXFWyUTMZ9cijUIozYTTp0wVtCsl5j3I
9kpOIWDYewnHZBppYOiJ9RW0W7LE6EP0hlhBXNs+nMUZsmPU7s74F02hQWTRkwGw
miRs1/vZ9nmtugNtwQcCW/DXN+/zTzT2LHItsWaHtccOCPNg58btQB9TiaTEYagL
4dFxqteQ2ZDVcvyMWRijoJAak5u/ZzvvO9WlaWPnBlIM2YuR4sPxdLi//K8U2And
2p3femjRxcTSzG5DlPj5LhZsUCkyAyuB7EULbYHEi87w8zaUq6AQiwq+U/seDYf4
E6TNp3bKQUqIg9kIJyar3bkl5P1zOuZwPrhqWtEbQlXSbC6ppTN+ChRzZq+C4gLB
DEAAIZ5Fzf0D7xVXolLSJh36qdAHzVn4oav5LvFmk+YyCmL1hqMZP0GAET5bTbLV
Y95Ut+W4iEfn5jI/KuaKCZcb1ZIOvQnNbGno13QEwc/2/JfuP5w7xklx8yM4LA0z
rW+Ng9rZPZ1OWlA0wSqi69wehou4NmcrFy/h+L1VkarzVEcNLV1aHByXJgDTAyjA
8LV4emxPpAeN4vbh/X702f5DTQ5q01zeTESxmaEO2VSOct4ElBPA5nGNBWXpS5cK
ELpkbkwlW1OKbUfVAhGRepz8vGja0mR4tueyDf/GLjAXHE9XvdbaScJKo/2vxV9T
EnW4tqvEld0ZNDRGG1WnEJ1XW/Ps3Q9Q3lvImdKBQVju9fiSZkaEBFOrdSOc+tU+
Otcxtud+vR0gVs7GeNxKVovL4OGfacySNKwzOQTinfuOKQSmZGfkjYmthxCt8xlf
7SC9uMPjP6IkXb6XD3ZZIzcvBRmeAh8CzcRjULakjtchRI4Pr7+EniXbW2X0Dpdc
kbM9MLwpHs5a4YOy6yvKrJ7raRNvqi5BpvIxI5MiVpi/CSeB/Q9ZMoJcRwjjLtHe
yMivF0EEwED/j2JwQi9FQ0xbc2zQNGyaw3EpfJl9wY9ZQPv8X6xzAtlDIF1KlpBn
q8/YEwpGwsa/Mqj0hM23VmR8+htm0eOS5xV7hEgqRNXdtibpZDUSvbofZetDog+H
bn1bcV2duHjVeum7+U1xI4mINC52DwhX8E4oMV5r+cSpZ7R5IskdIAx/HR586w+C
gg1h2OqNCmtzp+Rl+AS0Pyfrc5kktDKC0QssVinEgAQJLg5V3AGPrlp6lphn3Fke
jVIT2bTH6d9bxVPY2ppMmcuZM+TO24SMuaTPiUTj9JY0622/9IKc8rzJY/Ql+RBQ
h6BKcV7KWk7ecZ8W3ale1ULAdMUlVOYJ/RiP1KaXtSMVKIYMIsxKzOmBHqkH06Dr
cnbcAOqzLzucg6PUcxRhQL2gRwW5OKqU/PFNMh2HCSF4YyLHXNpn25I8oAWA/Rzs
WfEIx0r0/qdXw5CRf9hPI+hxkLasIqa1PyyPGCZX01/v8qMsL3saTOFRjfA4sOaa
wmqgWUrXPnYeu2sfWCCysLh6Wt9Q7icbmxrIQf6dDxINlpe3njP6Q9ttbHx32rOY
4A88/5xfeljYfXBzi8Fh1KS2jhpxTfMfdvXC17MrhjRuUHKfKYooVPgVRTN/tpJ6
LTuVkAaCoHVRfnj5QZrfjj7akL4Ut+IqW4a2vPl2t+IQgrUISbPkroy4dQGambIJ
plLyMEhInJjj6ntPYmh+dCWi0fDRhHOLAb/RKSd/vPtHoFAfBEHdcJOEka2ng1P0
ZcnKHLlrrxBbqoto/MS8VJCgJfu9x1EKsonw88xcK7lhOH/jMZdtFncicz/FI6IM
hVb929kSfn7GUlHLRTXngpQ5qUqtfuJV634Wa1fHr83OUeAlhB/jBvnUo8JwuDmL
LFHBf8uHWiEvXXGyfGSSiDG7FwSPjt8KgNkmy8dyrHtc7WODDG8P8iOJecGVzFSe
nSiM961Uwv892KP+Y988zR4AEgkmCY0shnBPQAsPXyUnpKg2bhVCjShjEFJ/iu8t
pwLPHco9E0P/MKj9LkHMbJyFhC7UBvBOIFPgs7EqnXcJTUAwZNUTJ62Pq4DAq1BY
SNY9JUO0OfFqsuGFDVQ/cPO01909+ZNffCf7baKFP5+/U+/N30cyeGvKtBfI+oUq
NbjUV1dGffblFkr9UtqqsOGXzjsXk1KnndNzeHoVqHAS0tug5iaCxJCO66rUz0Zj
RZLOyjYyoPmEMiky6Aq4B5lhnTVC5VqWFaQnu7U66g/GaqMfzYob7o9XSakQdbyT
jYs03tn0JoLm1SHpc3WRsBM18TZ19tPe/0LyJldVzEMnLa5NiH07ytoHtDGE67Oi
xbGXfD1Cc3R/JvErUXH3rwt8WkltjbLN7hL3ocCEzGVZP1kDUWz7gLSL6jeewdfE
axJPBw6BYiYNmdTPIVnmNiiFIlSlg3ohtwxUvQrF6RuH1V7TF1MvpZ4RC4KXu85Z
lW0VTdmJ8JtmPSMV4SwRx03F+j/kZY5zXUrEOLgMGl8qVPc6TOwRC1DuJFxQdMB8
YSGXGjFaivhyjSb8TEAHoSLesFmuhmC+1pV+NbFzS9y8itR8vPJH5u6fp98IPBa3
uh0WwiMr0Ai+Y1e0VEKS0pRtD/ZhmsABQO8DQssCM5fYATUBxzM1IwW9EoQ4QQEd
KR4CJu/UaX7NLZYIRRY1RaVUXHEEEGw5EBLH+adCm6V1WfbgZjTXnP2nrQSrXie9
MxkHJUJgoZsiXX7aQkNQB0kZ6NWEKtDIDdMC9Wn0mp2OGy2rj00JM3cuhkLajO02
S2aTzYsd9Q/D7FC7h08h289QSkwz/pv70+oK9JZCUkNIWJeKUYTUdKLlPOl9nlQv
SHAYkn6EaQJlpJGgnQGpmzg/SoYPdbjR72IkpBlIZdBqWtk6tNT1Nqx0oejkKE3g
bIGDfqrHylr3bfqswp2FdIic5QVyYAP4kOPFL247fV8jI/HxqjaPL21LhDXg/9XR
LAqpNg3rdmL0d6nar2NHZXc16vZa80rdrOItqbJ/isZWkR/2OXn7kuS8mGwGUtKa
bYP3SZqctkSoveKYSkRPmkemksD12/IrNC0XSdQFaW56VEEG/OoGWEH8o8K07eji
jIbxq9IykVWgS84Si+lYqYozt8zZMiY15v1Ssu1PD1jV6IEWJ2Mvi1kGe638Gpii
rXW2jwPNjdxOP7EMa12duzlOCRjvO1+LSZzO2exCnmZqE1Dhh2nJMI7D0oxB/VSA
yFJFcmc9RvXYm/O9olGbppuxtXGBWjVNYQ1ksFwiquXdoiENN3LcMrHD/dNt3jLv
oU6/6jrJ6/JQ5KO++bEqpr3SU40yloZfl+auQPQCjrEZ+0eQUB+EWgR3GcRVPmhl
snCJE9gv4kD+EiobFaFK6hezxy+xsQIk3TK6XJJSoRxuci3vi7OBzUQg1JVqK6Ec
UygNGL+bfcgrXIPDzLvokPNO6oh+u5cDlb9/MHI0LTmHWrNxX0u/tTbGlPy4LRFo
QNctY3xJA7aiKHgPyor33gGEtCDJjexwaouwanNEq1ZwfSApRWQAjYU321tr3+GZ
zhxdtMpGhuVsXfa7LzkEKSCm1lnnsp/5bXVQlDa+G74BLSAXoU86U7frMK8SmBGy
nYtkgUNv3nNx5Y1xBqaA38QtZhrQsdeRIqRkeZ4bgp2iTvGsSpG44lSDihfEK7oJ
Ou/Pse71zio4xDOuagY2jtV6CBDOvGWQv0Gb7zR47Vert1d4ZHmt3Cp9V5uylFG7
N4wukpfV7a8D9nXrgD1ZY0ech11BDAsFzjDCUPHxBB2aI6sHQ0mOuM8diuzadIt1
3dT7v13Il+2h03Q8HkIMxehYXv4f8Q5bAuFr/x3jsHMn8wz7XZ1Apt6E/8BOibIA
AQUWq9oj7tuwWlv3NbNj7jpdpgsLKefvabhBit6ieQaBoMsu+mHdSjWvIeXqEJHe
ZF+CrY5GGMrfw18sgPPIEMXATi3C3g9NvqR2U27ECee1c9PSLqA4eInsOj9vlYTT
ZFEwqJ7GyaprUhXcWa0bjURPS+/shRX2kc2+OE05uxlHeip9nZ99vLfX+xVIN3d9
1FTvLn+0/WiMkIMBC+73SAwmc6M79wElNNx4fy3u3zKjOTHM8Og6oKj4NRiYyKdN
E1TSp6tfa1t/FG6vWEX6XgYIv32nQ2ew70jM7FfsVd4y+XOHZ3GcSyfiHjwvxKiz
sX79GJOD8BvVpsD3GgFCWrMqKKmWqsiBoTVvvvS7sqE=
`pragma protect end_protected
