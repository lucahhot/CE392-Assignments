// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
p/luyj0mqcl4ythlbExUlmV8w+ZH0R6JBM1ndNjY7/77HX21bwJzEnfLXAJ4dy8uwoXNj+/m9Em/
K/qc4b8OPjgkrLDON60D4VmJU8SIncVRL4P7aHVqQiCUvE2jNZ3Mzx7vF8yppUClRw80HVpwl5Mx
Bddj3lK+2WrVLuaB3BLRrl1mq5JrQH3cVxgogPl3pqiX/XuWUh7HHN88t7Dq3hskcLm2gWNyNfmC
zQAt4tLe4MFc+Brsj2nbnziSQjA+Z6a+rdOpfO312bhaa+4BvoUw+C3A5ac1+uKgocJwlmpNkZIK
yhEsOZaHbtvtZ2LvqyfUlKt48XowEZsEXfcJDA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 91344)
ZGQDpUHn0k+sJlG6iVPsNScxIDpMo8meSvrFnq4kUKwE3FRwpPWZOP5SnGXUhbql09P5xaS1L0vD
T1XCEf6wS37mtwJZTnKMCXGFYwh2vTOuzj695MkM8QJ57c0GdCB1i7PWxzB5E++F4gie5fgAFNTt
uD8fLZjbx5YPpbXJnISUMtmkAHsD9AA5yNe83CE/chFDpS9hpeCkBaaLz57AZyNKl9mUUkgBtigZ
5bpVrkYIQcEU1PUZ1U86Tx9gsnkMwLCg04+tdgo94fyH1fWLzSRhze+msUl1p0LnNvAJF5JbwlsY
99V7H427Qfm5KKJYmqSJpOwmK13UKrlW7M+SxgtDOkGXsZJkWcwLnykm8yutrHEjKHPTO5HeoS9r
lF0X2Tmk3d7UMNh14HBGkz55WpjJ+rN+a01MzWIgwcNCOJCs4l3tpdQFqhM3fF1gFcgCHaO+dDIi
oNHjZkNJQuMI5P/809849q1ZBP9z6awU1bOPehxsW0XXYKNEOMXrX3jNpJQzAN7zSTIugW0xag87
a+cB1Udhvx68UHME0e02NSzJVZxfQOP4Sc7zhQT+qbrEGoZBw4/Pn1mc9e8TYU9Qa3quQ0IkOTzW
XGv+qDivbCDxLML7FIg3mJKJSNmgR1QePT86p0bgRDupdgZ8qt/abpqPJMxEh/YTh5wbWrNaMKhe
p9dmYhp/7wj0RIx3NGlOO48FX6SiEgt/L7ewXf6gzPx/uO7O0KxlEMJpfqXA2ZbAK0XYg/I094YX
aHWvsxHC9bG8KYlAfRuwZ/Kdyq65Kfp+7/Dk1jQJ8RLD5ElMeGYrE3n195Xqs0do7VLru3hpipk4
oD6CjfXz4B7KwDK+O3hlt9SYkXa1PRfZzGHp+Cu3uNRkscFMfKbsBmbEQSIG+8KnGnTIQeSe566l
EmxJhASPmhFzAUVLRugWFpC5fpO7ftQ7gpnLjtuP9cJYhL9YO6Rza0QOmBsDVxHV6PpE9D2H7D7A
29H2Q3CYG54UQiuqgCSNUjenV7urXBTNlwdw9Xo2Qopw2SxlrbUHtlWMflDvWdfJhUoC2VENl4t1
9swRcWzEZd9r37Ace5mPyRo4KykJ5Fk3Nn5wux0urm/ndulAPlP8a+euxIdvgMbiuGH7rcNfUDZN
M6qhjZflJLCy//6wdlKlgri/b/Tj+0A26KpvvbE9+VQk3W25rtLoMRjoB1IHd7x5FTlvZpzKIs9B
WPAqbfrZb+YOzVZNgb+waPlkzM+V7MEwF/R6kYqA0eRgPapyoxW0vqzbxRajoIjjmgXaNSRI2Bpp
orK1wLWl+LgOYA9DYzKEOdAEHr+LLM8OMeOYF7MkJNL/MiKxOCivrRDkjT+lVGFg0gtYz5TGvzII
KbBAZsK+6wi7fhkFnRD7qC5A/tcKsQNSK0LynXdgttszgzxt6+CI2ZjK019MKcLmvh6FPnLSxgfv
5f0qsxjgqP7xd2kVTF7VrI5jsewzdLFySthyxJ2YugusRzmAI6N489e57rlj2SWVvUvyyYQoaKP+
P0TfK5YQAgsuiIsyzP+Qa7/QP8gv9IUQ/OPQscfXxcXLtZ1B8D7RAd0j2ZcRfxXl+eozD9XaM9u7
LyXq8FW9P+pLM4AaG+6INv5zYQ9oFY0TvoyJ7QNPZIxXHIbCT3TT0FhMM6/b87K8p4lPWzRMq1BF
AYTvLtqPUOcHeuVU6/b68KC6APENX1IR6NBK+6l7EZiZacYFvZzcnM62dUmrd8I0A/sPFjbgWYCT
ddvKvw68IM7KRBoKGok8Eh6ERQpGMp9CZe7w6EOJx9LxboG4e0krkdI5GOB+XVaoYNISYqh7TVDd
cO1R5ULRYZzYCSQf92lCV668+wjyv7xHUAdB+3v6TVmLU+dmmk0YtcJ/WMhO55qbTE5EQlEelcmW
mSWDY3q0JgJvQH5/3D4otkbU+uDhJdn/oc2mPWTDfva9uclLTMhFCSgU62ri3f327HqApCyd07wk
rexCbWA/hctBW9eokeQV8JQ/0nHYMzlbI9SFzsyHN41ebsyGxH4k2ruTu2DMOLIIj7L1ftcLUzVv
s3gfUfT+wJt3lslT2JoaRByuyzTsKaJ/8EX+V8V0ut3qMMITAIjovA4pUlOr9otsKDqlmw2Q5GCb
EQ/xdao6izTrFV0c43yMHmSqZb3omjMUSrPjgogcelMSdqHLkdErP7Q5tH8DpEAhw+GO27pQUB9Y
dfKGs+OLwphwUebRdjVBROOOtNESWaQbDJgVII/VzrnvOZIcvchR6H/4vFA3z0OXdwEj4kWHQ40z
hcWdB3BEMNX4rJ9jO+y3PwXpJC1KzkVBqic97nw/9LREYjUJR3mzV3s6CdxMZ5S80bWbMWFfCUJ3
scKVG0L7p6AXMBrGvOT34q62CUiW7oA8Xx05r2jmhGQbvehK8KbrqsQx0mA/uqtn726mL9LoAFZA
2dL2/NpJCb7ao7dq0/NQFKu/HXv740IZH5invcuN1lNJK/yVXBDhv3pa3Jt7ea8XD5KCZLFQTG5G
uIjENd387qBaoyo7cgRD8ItzLCEpx5oKwKWizIMqccXpKVC/U0yMyhvTsPPemHkE6LXaLkSE8tcz
FfYBmqJdWqgxB+MwtgalDYhd1rmlofj+38OefxxRq3AUo2mY0W6TQlUTr1OqWSG4yRU+kaPvnheK
QeZIQB+o5aqXtCYDO3wCZInY6cXdZB0JlMznsMsRdN6CTxV9WinuloGdyhKYQ9qh47A9wX2OvW/g
HwmV48KtUMZt+ieBx97ivKd20AUDfI1fwZY7mq+Yfj5M+YgEfn2xmdhG8u/a4n0/BrfPg7YRJ1Kq
z0puRSuCcJA8OjycXv+z26DBtWVFYg/1PPuCdWSbwhQYRhU/EdxvK1DyrkuMqR6d8AVqeRelInBS
1PlljjFRYjFfw4Em6XnYsUfb1niRIUkPJb0WQ+a7OalYhcFLlQDVlotXh0m5AFRNm9+N5wF8uZO4
UXwpqi9imxe4KT3q2HWsOVDAd2XYlnDWxlG2BJwanNK9yfr8vjKM/FT6GuVz+LEjnj/mg27Fcwz5
hxNKLLTu1bvZtBVOXaA13vO10k8Ud58UrMVN9SqyRhEoqBxxuzijzcqcJWcNo8ykaQeqY/uZppDl
7PQOfXS+Lx73Xx29B4pWTm8eEzoiw7wvvh6W1jfQA1dP0uT0cvzklJP8YbVMKvbi0qwrltVWlG58
+fSNnoPn1BOLmrcvqDF/KtjXuqBJ+DsVKzjgE42gnUIgnTijGAFCqRA6Wunkxy8T4/R7Mf0uFDP5
pEvtOCfQsJ/F1a3G0PwCXWNQSlEagupG31KYjFq47wK/+fcCjlvOGbFaGnE32ouxpE2Zj8gi6kxD
cNphnEh7EbPHcKLU5fEiCf21swtmzuAVvWap3GIBlJoQBqCw2xFMThEuLpuFHiHpsnSx1/AWqxQU
AefLTRY1eROilgiaDrRZsqPBBhCZImJeSUJp47+QopjYtLIXtROu0E+duEuPJfuwoPQTd09yuLqF
5TKvqSxFwigVpGDvvjc8WdGDXAZBD2svpG4Ac6K+9D3Mlls82KdGdgMIVEM5KGSBRlTjh6f3/cQU
FpiZui+GqYLNdvTbnhCCdffHDp1RQr3PkcAmgf0xXWSYT2T12DwBP27AppvXEZqt0ZpQ2xzrF0J1
WyMXkojduKweHW3ilMfWI4j5cEdTsMRcs5I8JM/ixlzjyjTRK/Azv/R9Y21FbD0KaUR1ZkmKD5wo
m1PYb/kfyHjcIps61Olx31b0bnE8gvhjEpt3IppukBNWc7snUBgiejzUvQ57yU2xOgUt7ZW7GUoq
WF+o4ciS8Cov+oTFyO2pimk6pakRVSvcJ6xY4ghyOSBQ4SlqTPPbRvuGyYOgSZR24402RQVcWBau
1hY6wuggrC4yhjyRrqcKNV6qTIeCj8PcC/jXYqPppdMt1H5o1cytA7HpWKKmUiWVAqWulaOoVWzy
tkl/VU36tUlWQpCzCYRG6d9V8qjM/FaxJPxC+Utn6V1LNk9fk3pNgTXzJqR4Z9dthBRkzcdiZN9B
ahbBkgjLztPHfZKx7vtusVYkjalbEAzGJuU2EglQdwadsNEW+hNhVrow9mrBFBxmvc0++rGANmLU
qhA0kiTgTkQvifhqtehWdBrTPmLSMwDvLwXicONrjS2Tr3vYnOqSgK8nRk/Sg8ZcvFNCMsCGWsGD
ozLJsB9ggmNYuYAYvZwxb9LYsb17n9I9obUn+wjxmU/op6eHEJgLp94fXrr+GSYu0ktSDrKWoSL+
0WqTUWmlJty85s/E8BLlc0XW/YUS/5HIkR4upzdW51VwTQ0Msa/1QEgGUtRRmKfGu9BXp8lGO7zS
rsiTXGqEDLkGY6NdF259FWn6XSllyurjmhEWSOTyQmqXjnMRnADFlXciVSdUe6Ag5Gs1i2EI29Dp
+HHzfQCNVQ9wv+5w/DAbHRv797sjlJeWnWQ+2SGT4sAfhRsSUi/NUT3blAsRgOzYVeGQVu+YJeGu
AlAc/N7Uj57KxLpxTS0++d7JxQd57gTx1O6go+FzMoQO1B7B7pnnrt5zvvE0q6epF3kAWF+PP/bl
Tu6ckn4R6LYbOu8xHm0STqmuSS/kad5aOVQx+6UG97aw7Gi7TBZbFqJk6a9HFYv7m7Nf2AfsZCLj
JSMj+KJKDixPB9DhdEN+XBKVR1/ZM89otdXLmCAA/4KOFVAugs/mMGUCHBaoRfWoGK6W67VPT3bA
twTOaqySP2hQbXHtsrwVNnq5H7z+1a6/Bkl8Xk6MgPnIKP0U5AXPvgBEHsA/khFKJ1EXPGzAxEP7
if0ePfiDEOPW3vJqA6Wb/AnE9GB3HW6yow4f21WxRTVqLAEYLnaNyj1ptG9o8U+iWDMi6/dxNevu
0vxLEJ9HIarWntlwSHx3OmkzR5lAiZpwfzn8EBfYDhp4zUynpvfV9UoeHZI5TzfcTbbALtUdiO9B
Lj1EXNkyLfrLRkCoFOLFh+05/IGDGccg7Pz5yEp6WJip4rXYUrCndVyqZJLN3MHKcOhuEF8z5wxg
5eDSt9Bu71hKl85D1MyGR7wlpx68dX91cD1NEfyskaURU0Gg01iF+jA6uE29f5KrKkyHc7ZVdO8W
wJ81pCtXXCsc2nlUiP9VXz+BpFJRLzyfzjpT60setqIIIX0D/iu90PUwaGi2js9Hf0pa8OKHXMCV
/Gqj7Oil7p0rGwQKcxVmldS8/yV+dqezaFIqi5vAaduFcBxsfhRl0YVzXktr0U2mPHXsUTr9MKym
CCnGZlc2YMXz/RSp8gaGgsgzooLpWqCE1PgY6EzGbkw6fJz1yYr2kAdAKz1oHzg75Q6ntTC2/pBa
ppGvcUMYyqaRVA729QzEDiMyXGUduMJGfPy7T/xd8kYrcOKS8r/1KFL3IvDlbfRkXJgPPQOS0TLq
wwSVgeA1xem/iOgIaSjfcBDcLR+Kl8Z8dgfatTMaDv19KRzmFOPXk/6adTpYInSXRAM8SYyLD02o
AFHV3afbF3VdFxAo6mFU/mGTkaoeu0mpEcYeKXShy2TeM5p64uXs8sUaobncq20qt3OpWY6TjAVH
+Ja1G4i/7vyMZwKyakCbGqnJnFW8o4d46DIQOnYwE7rP9OO0oQYFGNqps+LEmAHIC36z85C6brHy
vnVkms/p5MG8CpL16KCL6wAY5GVs2ZjIpVzsp/9XUXJ6JvBG0WHNOGS/K2bKnpxSlU4qtUgiRB8Q
4VsE7KQ0OcpGGaFGtLHmU9KlFcqIvyzhVC/7414joGa0ahHO9dG1UqKjku0jYXbR6vcTHuF8xZS2
TGVF4ihuQQ0KiuUZMvQ30CgAHAsH26NrxRRSPlxgr6d52Jnc6Wl4mg+oA9Qa86RDPBARWeNpo0gi
DCLTZIsRw+WZEg5k3wKIDEMh01QMJq5tUyqAFDubi2shFF5Ac2CE6VNXw2Uxpn2bLys/p4CLWFRA
7sp+y02Bdy2TcMJPfNJ6B9d7948LOETM9UgJU3tmEjp1W6jiU9vAlVyY3qQMptoPXZCriDgkp4cA
tFgJWsXqjRNh/v5rPf7WSVRnvvLn8pt0UjjFwIPZQ98ffWCfsIYvmGduFx2PRBrJJNLNdRub/xi5
Jic5kBjVcOpgHZwQrYZP5lvm9wZvNHhKgFofKXjCwuKrZxW1gHPSBStvkRMw/KGjUNJ1r/5rVlEV
D98/5NydNUKNnLy6Q5w0UobC3y/kkV75SnS54l8wEr/+JaZtW6KkrBPYghpsqUbbVMtj4h7NGgUw
iMWJEEW/gyaayjLp3y4vV3x+HWvbqdAVhmMhn5p22Fob+VBG/wtTm33KdOS8Np2OG+2VO+5s8rBO
/+KwuW950bWn1KwcrL6kQhlrmR39kG+JiIt4uVlLrRucaOq2Zu+D/ykrv3lfqhWON0fBld/IogC/
D1Hr5pkHCSJdHS7lIFAioF/E9TpSIIO6migxW8zrcfrnXXCpNXTSW2QayJSsxL7yS+LOR8AZt/nW
CmCLaNWv3AGVUQyY5eBT3kRxdnhFRGRThhVUr6HBpdLcWhKYuf47/Kusw4PgBP/qH1G+RRKD3uhU
O0ZwZQmC9vIaYE6TVbfQlVTk52h3Tgy9cphUaEOIo/yDgEs62xsuIhNK016gShm3P5nHHBxNbv10
k02yrJVueFH8+e4QNdWVrfq2RQVj/BtQNpqkukvE0Myixx4scKm3OwcJKnrAzZifrDpHLmMb/Oy4
PD0sYjAJ1rcsde8y9MKQHIhVLXL0NyN4WGB/Ci5wEixJJOGGudvqUUxyQYX8uwqWO2KW2l0BuLE4
YGj/44ogkuw7D+7c4kfXjrs9B2LQChvAUlE60qytpLKynnlzGm84xMBaTpZOFuih9BWd0RIrIq3C
sBvkDp/Hf2NQRa1MUSfVrdrPPLHcjQlsZL2yD89UbzkWuJ9tU+tKba+U/wZ0qsq2TJA2kEFhUuwa
xM0FLQJyvnQhI3V3szFk2Y5wd1kr2f4svoBbDwDZisBs79hLRDmZNirtLjSMxEceJQiZIXjSyZIJ
Si0Y9ERHLpqZsFvuXf6NCCK0RPPHf8VxvYa8krLh23FN1KFaVkL4GOiJ1Mrbf61Y16/5fWt4+tIH
uy3wdQ8WexXHr5eMvp5IHQ5uP8kK72mP8HzDrY5aHb/SclBq82iw2dYwKTuCRWcuUSOs1GSMN2AR
8/At5f3o/nNoElm1Ql8m72S1/LEd7hhQyu4IdW5uWCi/kKRf8uR3UA8D+HHogRaWA+56dVYX8/jG
D4drj8BLwYCmIlOsRIpMU9ee7it5LguTjOrSwjcjtsQvr4BYlZMEnlLRjWI/f0qC+p+4fn0mTCiY
3xTV6qVbVaueaSisuDUpesKlGlGh+KkciwOx1fuiY1BrzmcL8g5eFCm+Or8LODVB1f2cL3a02p+L
pkdvwe9GAkivfnd3AdRa+Oyc6uEX8sd5Rf2eoRPz37eCjU046TNFPA1h9VWf4I64afTqpg9atVQE
F6ueKwM3nfeVT0pnn3aWPAa3iPbKVsJhcLB0IrPioptK4tPSdhDEJIAMF92BIeo7FEPACtV9GjJM
3hAuyGyQ1WAKvPbPtFjrIGqTpEZdHRL2Jl0ASK8v3ePo1At1KcAmE3/v4EQe/N3daTwX/q7SFawP
DCl/DMPokWUhimelLnLvjY6cMGDCQduBuTVMUyISl4wyMAfB68ofLr+q4pKqyZ7JkBqzVLl7pxQP
smfBr9nOjsU8Q6FDRvet/hLCK6SfRhnqVPf3pLw7wJ9Z5GdU1LPdB99v7bgnO1WO4T8NYMEbiw0/
fKYm5YG1EgcRO80Yf7O538ZSogs8lvcaCNZJX7Bx1KTr2Z5B9LlSl+w0NIt30iSoUzREalOetJEM
6IgsggDB+Kot7ypCPPDFKCO7cZuYO+0h2QoQqi5OHZI67vTFTHNO2jOlsF5EaPKdKLYt0BE4BHGh
M1aZxyH+xsxxq1x1Powz8qcZIJMwJRjBMT1fijukTS87tJMt3hu4drRIRqV2wFOAo5kwM2Xb0lfc
xS629+MH0ckuMB/M7E1O72Ak6y2v3KZxrpCYGWrcQB7sSZNaRGyVh6gB5WSjD15xQxuO471GfBuK
tbyP3qAJjJ6nyBefp3nPJi2sXKmerZSt462goPmQn8QPWoc8YSqZN5Ii1zkI2yWyoucXbeXE6ggH
goRWnNQO++MhiW3QFy7FyQlHTYprqGPpH7W/NMwGtjAISwM8tyhgYyHXRzcnIbBQGoYWbYlMv78v
b14MIoDMMWHnqLeg7zT21RdIpFMKOyuS9bTmVaWnfidYONeXLvAYt/EUzrOd3hN0zm0iNKuxbbDf
1yqTp1VYkgCGcyIDQm94+nyqfisB9ZOn17QebaONrVsucQB1eTCil/gLfTvfllHJTxph+XUAgORN
ZeJxIG6RwG5EBbGPJ1z2iySt6BmamyyR5MVysG35bmmpNGOphy4q+q3czEedqMVs1KlhC2e0BrUj
hoA8cDdYrXqUanZBEcTqyyRUyQByGdtC8Wt/cB4TdrQkTdEpug6swfur3BPIny1r9MTP+JF4J+iA
o8xTLg+4nS5Q+gzUKL+7MbprnirscIck7QUG+WftiXRq3EGTvTtLuVg5RDEWxybRIe1UG9PBNj5q
7mMLkm7EhuAVGzp6Xlhp8LkyVm1OxaCHvYhkhtUJAs/slqXqFzLpd95qjWjdtfcAbt/K14ZL9oGJ
VgbB8Q5iqvupVGO/flk4y+r0q2XXXNTnD9G+z+TM/sn7HEVON8EfwZegyDU6VCoRNDVbh+cSL4ew
JMSR4rk65Bgr3IgzJt9E8FghLU/YUak6+FpTwFUNVXoaYJ8EmcOQ1iGlSTcuJcoo7GGrhZ73zhN8
TJl3FFlTR1AUqWp1iuhAz7VmMyMYD6T2iqUSIeusPoKpGYCmbTsfZ1blsFiNN6cehreoif8w+nx5
YBqsG7e4V28Krt2cLk0st9KC2YV4GS/wN0vXIS7J49RDrcYcKw/vcodF8E2guH9hKfsjMeJMH67g
gf2/KjUrasoNYjuZdmoAFX/YXMU8c2xzcCPlXhNtBL+j2iV4i9NXNA+SZu7zd/J8YonejYG7By9V
U6rpzYjDgwVuv0AixpNpxaZ87UZgAyIrFLA063awHsVUp2id84SEk+Bg7jwoKrfsficzLROEfkmb
hhuyaNxcaQWs1E8BfHEejAnLslCWghINJbKFX2LW35u59aOMPOeZHlXSbUfMUOX/n1zN6zBNjZyA
MpzUj7+pKyo8qHpugSLnOwa14zqJGho27m/evbBPxOogMZuOYjPcdnEtJjErkCUOEKpt/QKnQZP0
HwILkH9JwYtxZjZH85srnJAXCDo91cVJES53p5VapgJNWDbH1wMEVa276NYH00kwlqofS05PKx9R
mMhv0PcPDCVLpf3xS52csH5bY/qYqVqrKddm16UDpqInE3Msmjk00ehegSSYXrlWFzKKOD5zrNMk
cEuF18FHbNCrM2/T3CLc1fXA0ITH+ukspbl9VhggDn1QZlUJf1Y1T79RutzvkAaQE2md7F/HrkUf
GRHlT3Mm7OhKaIgL5gMSjMpxIeVbKQVcvy/uS2+J8R3XzNg/VKUyiGvRD32/wpJI61+eG6vit6ua
f7njSKz3eOF/FGp0PXSrl26xoaUXcR/ILYM5ZVWD0h7YjbYzvwVJn4rz1hDdbwKAbRbpDkVjOVKl
76bEtA9C5h0Zp/TYAN+SygmRRJZSqzt3KF5eBY6mcMRlP5IXMpBAlyGCOGDFv4/k/bNCBkzmoZbO
vqHPbRq3PdSGdVQooSYtJOCOMxupXdd5i+QJIO/GKYaaxHgD0prr67j+QPDmdXBjfPasaxKPrVtH
q3Z+QH8ljMbg8Zw9MeVi3zP7h9Rcgef7JVxVnmJxUJIzkhWKqWNHJc2NJiKoImK+TdFuO7dvsk1G
bWh9y/kDgxNNOXZhbmeUUZNg3Bz+x/teKGJdV9G9Ri9+UFXvY4ErX83AwnGb6l7Y/G8bOsG/SNNX
qj+xS+nrHd0a08rtbfED1gSDAlerM42G9ByijW/EUppLFGps8gHNx5D/KhXARUtAM0dfRZj6/SuA
SuwP+/oHDrTZyIONBBNHAZ9rIeb9Q6KIp+ZOWtLm2EThfD0XiLM52mfn6qcbYdcAiWO65T5XtWmF
Tq6cxF2bfH6nJNZQH1kp4Y+dP0ADq3ngiAQjnhrj7iCpTZBF9Z7UH8ew5RY09rsk9Q1u6vb4269H
QEU3E/mkMDHA3xGfUvhQiCyilBHuIHADjLiPPUAmkAMG1Ru0H+cTw2USHzizn9j7DLAdKysbwrkY
EntS/DHeWSuABRxzDgxOYzi223J9tel1IpjG5NDdOi0rHBLDbjjF0GWA21fOkkRKxeu0HOdvx9Bm
0gq/sGucMDYF0lcjOAwfYgNBf1thGzw01KW9zml0ryJUmksmlI60AnDxAodsAVosF24QuvgssZHI
dt46FAzN6VshM+Msx6ntiVqR6TvBhJtSOhGr9fLOKeW9haJaZrpJa9fWByYs6NbYIe0FeAh/j4LM
HCHUe9LuwbysU80ROueddtJqk5NRxjbrcc8yXTvmrybMo0vspDwpZ+J2XG7Or7DuHRgsMYnMIktj
ZgdZPixyvnDlfytQR0HZqMCN0T1nKqCVBOjzLmxctDcDCToltotmHiKblwsBaonSxkkHE0+dNnfI
L/uJN1EBR+h9qWwIgTBFi0233SyLH/a9+jLHXyWeA8Uei7epaLaDWzR5uVoJ6IPMszpKwL9BHnco
iH7eN2B36L2fzQrJjhR7iTd2fu60vtJ0HRQzxgEY2F4LwpKIFL0jCFxHmtOYNM1lTQrCyk+9qeDA
R9WKwGkuA77VnzTRxC6rye+mBGGCzAPcJLQ/em3gnPSCM92y/3bIZWacc15UgA+5LMdoO4FTDwdm
DLhH+Vid/ruzPrB6hHUL0j3RHqwQH9c/EQPpImq54nS3DjgaCa9x2rVfgxTwqsfCfblboJkFSzog
BjWM4O4KREwZwzCzYjE7pNJyB0uxDFTt0Gm17LBfconxkwMNdXhWQPI1CxxbBVbToSjZJrOdjtCz
6L91+bI8/RKOzDSuiEkUahZDTS9WGQJKN0MNDejYe3MjvGHByAAa1AfmoAlciGE2AdRxp0XwR69X
aHA2W30Yhw0uEYRhHfl71+yeXZZdKMI+pn3lo3ZKvUb2el9CqMrvwFTPlgYiqpYPrgffXCNYKyUI
3AxcmEWjL5+XtZ4YbCaxUFx+4ie7eetfUMeHNVgQh5TqOXK9ePT0Ubs+SIfHvr2JOrTMx9+AvZjY
zFw/ZDcXuSJMjVCt3jpHdecxTaRMfsaxSaupRQBAN/Ki/EPuGnaOYGbc6kcyM6dHMRkWtuA2m6WS
p0scTzi+SVcgkLUinprbMpOesT4GdSbY/VffgZmazHfg4Vmzx+ZJCvsNMKwlp8igWRsyjod1wrHn
PTGkC7P2w7aIu21LZTbriSv/HnFyTVDbrMu1l0evMMqh58SmDwximUklvUvsv1yi0Kq5uIVwSPNd
fZzB899vC6dTL+bzyTbDV6DDUUGr9w22ZormoJ75YfIIhRM4k4Rn0nSeRZtmX2wCKQGqbr1NNr8G
BAHQimx2BGqrsEwRfbxZKrxxlW2uHFaT4FxLXPzG8/SDVXweiadyeyBNzhMbyYSp4+YPfD40UK/z
sH6xi7ypYkadGA4iGa35yyAMffZ0L2Bwzc+lD1PcMUpogzagrOS/qwPqCf0s3XbOImJ11feGW86R
pm+2hTXtPXv3PljrUz6tOOfLxziPIAuYa27CazGPDyAy1B8SrE3o4SQQlDEKwBhpP0Xx3ZZ5KhRY
ih9naTRJCmnCQ4V9nk5hUTuM/Qju8em7y9+bK5snYqVCZTiM6+hAGQwjRiTLaLul9RQGwGo+TAWP
iy5PhtTa58KEhq7enTY5JKEnkzaMhWlQ1n5x3vytezQtSBY2DgoXKAtLA0zA2AH5jmuDW3yVG7nf
S6e/dtCSZZdRa+Wmp4kC4T/FxfWOb/8mGejWAXSxsp0fvbpyeikjWTV9WLNK+fF5nDDi+ODdR8Fz
d4klaRI0rpBwk8M8OLFJXYXSveU8E6lFTHk5piAIdG/DbKDvBHX1n9cV4cP7I6A2U/PJsX/yzm9o
G7Uf9+952HZ36KxRRlUhr6mcTc7f453wfju6j0xyypCMelGLpAd4yGMnKBx4DSBGGJViU5s1cD/l
xoT6yRRNsC+9zP39+hlZMkCqyoWshTMl8fCYqRa0dfZFP4smAg7y311Nl/MzYu5aeJjnj3CdTHUb
1Km0eQIo91RTtNa8vU/8aHJEftLbbBtgaUk1ORPZQWpYmhqCnu4Vq0ZOVWmGwKzG0HFUnvNUpIQC
t4wPWpf3efwpIpy1dRGw8P6/w5qmOvXhQf3BtzstdbQmdmCmpFqyLyXK8T9IxRwrXBLsX695ef3B
9s6r7oRwW5H+usc9LLub0/14oGu6g7L2oqubuvSo8re259rh+lXSsqMHWUb5irjdCPHphRPw61vy
W1OPG24GNCB4YMHg0HPSrys++dEL9Z98LHLNGs9kbiYFWOVD8x+BeRvwPD70+dslgA8WD7J4Nzax
w480Jt/apg22KbpN2iLX6piwsUd5wMy0efIRfBnQCSanartM15OFbJ+N8CZI0Zwu/6+vC4CYU+c0
eXeQsF4hB6n8qUWb9QaccDqOjCUAjRqyiV6y2JggjC2k+4Fj/pF/CPpIqJXNh7fOvvCR00l4vFB4
H48/6zULa+7uJxU9Kfo/s/nBczqo9MlOuQfVl7l5o8mWMn1PfkOzORCVbaIsX7SBPvak/Yu6VyDa
2VszN6/0gk5w1PdLDG+Ff9IoUjxRwLsN1X2B7MSjtm8tDL8cNrTp2GEgGG61wLL0tjKNoaGcTONc
lX7YR6tvJWwVUCa1Jqpy2CU7O31ih3EpG2fAQc3nlO2DvsbmB0wlmrXCEkRExWNEuiWtRp+zuWEp
ffQFnOHMAZ5jnj9nCjY6pHona3Pf5X5N+1myTLzKwoJU0rslxrvPD9m9Fx6JdJ/mpgmwMXDS4HMu
cwCfLpH88EtWpkR4/JP42vY9u4MruYKwZw8wi2Zdg2Kps2dD2hrX7PvTU7nmx39Ug/Fd59CY/alY
9Iziuiy7ZBgUhD5/Ix+3PdFWiYnDdxqj90sj/xv0T+d5Ccl9S4oJWhjd5tXmqAaj4HHYnOzVpXrf
xo6aiLBrjqPXP9lL6OhWuFRJI6RttxPgj6xWRyZQXoJ2R0iLh/0TKWu5jYwnXcxKX1wk8ZscpIxo
or60EFEXtfgAXSz9Bo/9PMQaSw33EzlU+u1SNzxMUvE7GGICK1fsenNhv4ICQRDjSwwM3QuFjLuf
Fx/bEaPXCpyB9D648g9RW8fOK2PuX9zGD33NScCz1p0qI1d3ASJSkwzf/QqBl3TeXkllA61NySl2
4kgwPt3Ce9375iB6ePDNuml9nf41VUkYNZUoDsixn0RdOqYuUlbZ3Z4yAbkCjgxP+yIwgm3hjMzc
kundRd07uW5IgipRYlkjzKvHjo2c5YvVh/6/RoiPxWY/gWXRGFY8NjwxGLuLeXuIA9mrLbjnXmJf
fr5ProJ9B1fBdqfm3/yznTlHlcLScFIoVT5exCc2nTz5gH9+WspcOdFp96FcUAxkCbPo2U4blRzB
XlLEZWkgRH5bbfQvG53j355cOCVP0Ss0Y9ZmbZ6FuZ0k0duiE1eZKLbu1/bjK4IPT+NmYO93PTUw
4+7uXP4QGglX0pbo0SfLlS4H6bIMJTM3NlrK9SBiCBSttbtU3MH1hdGjZbAMOSFa+pUS2dJQyXJv
soY7Aqret/82tLi+m43096V86+tnahkaRhzlL879/6QonUDoGyFaxkw9lEOoeRaHZAMYMm4LkPq1
hB/2XiMhriThZ8YNzjzqnP6eemc7qlIi4w07/YhLPf53JzjXWbun6bWdxvEGTyEwc7i9nUEqDGGK
N7QJKbrLKEwsKDF4X5p0h5ocsH40z6JZdEoW1Hu0hGgZHHpyXM4J62G+efNpXWkv8nKz1tr1kTqk
iOTt8VZpjCvEGPLLi4fJ3f+l0UMZEPhVidzXFWZ9MuK4mwUYScZa9g2QmLFF9hKGYtlzy1RsxaP8
vnIqu0QzUy8fUj1FdLfqso524EJHey1Q4vJFbSb9sLFwi+SRO0md3xEbh+GARGFPepS2knxYlex0
mPHPenYO0rHjSQc8lYubOklJjIatXPFTgr4STFgbAtxIwJJNcX1MbtCz1Nm65x5jSm8yWRbAVnXy
be1kaaotYe5zIoyTvp/pD2VH8z3d2nV9PeEyFeOoTK/2d5Am0lA3KNC+RiEfmem8g1VeUPHq5ley
2rKV8/RdLaL7tpI8CvmT7QKPnk2n5QspmOoDpvtllB7/lN9OYApaWcn23wP80pvXXvV2NqK3pfpT
8vQFF5ctI2yWf1fOLQz4A2lnh2/wk7RlWLw9GpAfX9lsXq4xiOLE5X/0JPncpu7GAcYunsPFcH8C
7Au0BPvADnIf2shejWSjGx/yb2eOKnHvYW5kEaX3ETQY7/QPhegp3M0djEGWyCpxWoN6byrI06Zj
hDtoJ+mApj4I6xYq/kKAF5iC0q85/yZhJjhItHPOgn9LlLYZ26dPZtc8gOUHJ5xd4AwY7rJ8UFdZ
wdB1CtTVotVkNf/nNiSiDTuRKeSyeIW2BV8qfFXeYcfo8k3TY1xlCSvT+KYyz1joxM4NVUqHsflm
+YMVB6/M6HvQ3lb3ha2jy3SQhn02FkHc2MzU6Elnhw4tP0ZAK7y4BhpnuZa+K+Ag0YkIRrTJSrVI
2U1wgpHf53ZsT+ahrePLQKev2IAV2ZpQ1VMwRUWfeK7bJ8jys6R3qt5tNwNqdZWsD7dUeiAetmES
vl0MkRZ9WGcZiA18x/uw6EeOkEpKMnUD4bK72/sHOwq2rCjF7Ta81J6CKD0oYeXP3UeNOyY/2X8C
YH2tgbJymwJYj7/J9vhu0RXQip9qqKamE4AEUZQkfhr4Ei3j5FL+YEHbSG7L22JTk/YQAl9iOfuw
nL3vZaCJz6Za+t70NclvXnsQdkLA39L5SAplBoWgtdwe6tEh1fhtim+fgB2GoQxbKF+lqaFuMe8P
LsYhdcWG5ZDTUxwBUVy4mlRl+XGUAxBEjajI55pu5qEkVh+4auzBkQxxRDpi6SmwsK/Co5S4idu2
g/fXh8SQrUw/m6wC92QOw+Y9iMAcYV+9VE2FHO2pYcRlF4qpcREqQysX2D+N3HUaWwNbR4AydoAR
bSXVkz78ARVroinU3Dqx50QaSZVcUr+lpqYaNjBs+d+p9xohefMk421Zl26mgYzX+I9GeX1GdvG1
moQhAzv/IA0XS5Pl8x8aM4oRavJgl71zXWGZR1yIhOElMSwu1MP6Tld7k6QHTTftot/oLksAtJ3T
pm2y1TYdQJhlDY3Mq/LBF4a1TonVbGYqaL0gxdCrNdG3S45EgUDaJrVhINkErjNKxULHhgN+HLHG
wa6pZBemZN1XOSC4r17mXutpN0A4GXtDyWZzijPHKm2Hixs8LKKO27BcuMswWv5JsPUWT7Hi0vQy
POOZA80LvPXLyY10HyRXeZc6AyA7CnDWX7FDrIab1XBumu0YS/8a0DIcjZ+cxoKhJ03xPfH4qcsT
fIXgY6cF0YW65MzekqpDRO54qPSo/I47fVVEpKTsScNB4h+jkrjNatZzQmkPfDjXitTiVqYZM+X+
8R1ov9kljb1fdFDe5Df036RLlJfEOWWb7V/PiJb2OGrzdQ8ZK6Ft63XTDTF1lp6a6/no4sCGoXQ/
zw9K4P5AnPR563jtOyOg5RIng8J7X1vAUXrGzJfPXfE3xJM9+aduUBQF27DjXGP6v+z6HdFky8kb
OicRqGs5rJUNMAR8yAdRQnxTaqoKoxbucgOU1u1illEA295hPEa/AqR5+sVmJvVCUpjA2KGbS5b3
1uYesq/BFkzOmfvbeY/RbBgnGtWIkVlglYGv1JTtMi99yz19iaxxU0fGB74Pif9x1cbC8WorhErz
qGbkhJNIAMN2S/WCKN2ISwfDKejJJHs2+5cIgs2KhQOt8k4NzKW0y0XXEI8xIxck0EovFO9cRodx
5G2oxGAbDmV6iw6WMpvDKXXF++CuryzA4YCoXRWCXgY02EWwqX7bEhRpxjP6Sygtjnr75O525Owk
efQIy/U9EjQdF2FjkyexCIz/b3TSnSfKhg1Mo2SGgikfdKudLk4JJoPBd6E/hT7SxNwTnSxc95m6
+NssnViZ2R3tf8Cy/5MU9NyYQ6ezxgtbPTVOtwyv2SuBooAylriRL0sEUsHt27gRku7Y7GYmYcvj
ogDIN5BGhIhVjBCLXx4/rDrp8XcZ4ryc/D4prLgRcNBBGE/rzAETqJh1OpxOnql00hM+hWMoDtVm
o9Vbt5vTTkheApBmwme02lasOFwdVTfGrUMHCaYcsCIuQe1MQAJL9xwmuLMtwsKnJKXSxVj2Jham
aO5rSsZeciwsSHO9iBEAoAKI/gnBTBepp+Kz/PvWB+klpiCpgf+BqcCOWnMYE7FGudoJ8tbiu1uB
QAmApitLm67VJDnXB9zxAzUIsE2MfB6Ks0lUIkJbpI+IIO/bYfGyqe8mj6q2U8OD9YvGEp43qSRP
OXG/ZYT3PIHg42cdEwM/23wlW2XJ6Imm38dm8KOZt5IHSNdShlNiZFlTaiWaylVg93A1GPwwU47X
HJgCaf28qk5f5fjUEFbDM1h1Wui8XqRdvKAB2/Z8BahzkBrEJ1B0w2bCF5Gp2UknNlQ/nwFDmEOc
ddYagOqeNziqW3FfxAu2pwSbz5wMYxS4d87/Em8zpGzLJEMgi6raBRFH3dN0DD0HLKjTU9pA/aeZ
spvuCRx+RU/iLT0U700R3poNU6CwaR7dz4gzdzStqGO8lAOrCEtJOMO8TWdb3N1BGnCvJyuDKGnA
4J9vtqAzDmv64H3gQo00OXvwr7u6YQHzsYKqXNZsQs4HbnyCZIGoZdLP+T9K+ttqG4KmaAmjwoGx
sr9zBhMUyTKearm5ZTXcm0P7/KZtxnAMFBWRLlZhfZUO8BY9CVdyTQ7dTEH2cbgUlSJIOmunkf0S
WoWHnEURVquNN0OQSosshy1BxUOqKKB/jDo7bcfbfEIZ5BtBIs/K9RYs/j/sgx9kYY4WRY/lSkBj
g1LXehi25Cmn3rZzBTGnnzeGQVxNHT2A6hIF5CKqeMViyqbY7nl32dSIOvRcxaIA2hx0jOa/iAwp
092coNEmnFUz3BRdZiiv3o5fLcgy/ecBHwvh9XRZyGD+YGLMG4qlDZ2CE/MHYlbGfNp4iEB9wSc1
PjZocfppW/XpkzuoUgkSNgcv7ccVUBh+dyHC4PtkL0F9WnSfpyXiSe2SSkQQolVfhvbqvYGZHx1u
d3Dx1EjR0NZpTfpdXd/Rh43Hs8cmOp7xmu7s4pS0RzWUvr+w9FJPUidZUPmg1oKM+ucVY0/FLY2b
R9Hz/Lxl9GjDfF7v9AoMTs7c0NJGxU86N6aOt8AsXtFgzqL+oZqG7oa6hy8w07bNWf/YzfwfQqZr
CMpYdk7PCEqk+ui2Hntsz/XfeuS90h1xXAAWEyxbcehql+ciWJzN3HmRVUk+A/g0moHMWOQQ5dor
I+tkFnKUuRZBNlapOpZIooP7iCHrBaIQmptuX3XjVyP0St6OtuaFgHj3gUk/W0nCDopeLH14G5yU
cGB8SBjaXiQi2lrEXLgOrNw7/EcF1ye4CfyDdQ4ML8mJMTuM8cVRZIStF7L8gvW0Kf9zshV67Hf5
ne8XIYpLMPz1l/huKBfSZEarZZG/b+YP2inygE//D5NJFV54FSG2bw8lN8pdjNMyUAyqU1xwemfr
YSHMOr/4Ca21dC/7WuULdt8L6ck4e7TpLnYZwmNJZ167STg8YaIsEnqzTIP9ny7QTlLOLiqmzEUi
2AVTxs2rky5dYU3N7pk9rUoJniB/Wdzd04THVL5sN1amMTA4RndP0OoyVr74AYoS4T/evDljxKob
Kp24YkeLEAkRWHxk1BY/JkmRtgZqe6EMlOO7M47JsEpo13KSfRfcjJcjFNzqKnApkkpEUuZ83um/
rB4G04krNS0nyRZXiRaj5ytMnghnb85fvgUiCP2jkG5m1fRUTEqcEJ6i83qxRfzVkdF5plzg22N4
GhkleUr2LP1wkD3DUU3jXCexmoz3vf/K55mwXRFHv6FeaaPZCyvmYJTopZzr+W6EQPK1xTHVzsmF
UYdXj8PH9PYkIeI9nSddnMm4pWAXzkwQOFuSfykiNWXQc3RUMT/F1gSSXkTzcY5Sq/AeeLK1PWkY
bY/dBCm0Abw+zqb24HwRci8sbpPc0bGJpknY7YK2r9fZp6sLqKH7jNT1yt6pkyNspyZZqToInLB9
ZFibeKx2mXP7g1GZyoQpUKEkjR5XhVhLq0KkZmxGw/cx8e6W8TuQ3aMUIo6B4BVpw4DpiNVAcmUm
A+BZuW62fFt8Nj7uj7R56iMWIFcXw5zuoD6p44K4UHM2ZYk73tJebd3uB2q/3DyaMC6ciHFrqOZJ
nzsJxX+bS9tTuoSq4Xu2vfUXJICHt7+CaCk2pBCBLCZEDajWxSeqEflz+ACbZeoTnbp9R694Incj
QAq7a8jYXCrXh6ytNEGM7IuU4wRGBPTMjytO8WpGt+3pDUTSrQq/DpEjIDHCPYqdtPMGrY7vahR4
rETB5SgV0Rbs6ekIc/kU2AcSuZ2Ht5XaMuAz4q+OpvQyJcTAyEX3hchF9ndaTDT/df6ECtjxa9R+
wbu32/sUqjlcGt9eF6f1aYkzsQHaiFTG+a5JiFIAirhF48JEuQoD6wri6pzwRRx8NilALnXpnhcz
NC4TAgxB3VcQ9mV4Z7CLUZ/WNrp0v2kf2DAypnap7uOOKPfNRi1GWVNrmSqXSLDambckFePnfhZ9
hzF6j1IzL64IrcX9BI4Rs4AY50/Ji2Ms45ZGITnf1jbdynxZNy1hVypdSb33JK9dYde7/fmjT02d
IS5FggFaaG4H7XMKMx90Cko7ty3Tm+mCNopCe6byS7y/FcDZO/TwN212WG/i5rfOLbapIiT9kJ3h
ZcjARw9ZeH06go1tezhFXvZOiTIyEvh8/V/9aSHCGyzQ4RtaJqmG7NAfOGJLxZF11ujOzXPF/07v
l9z9n6DAMQtHZoKrtmZSktjlXfP4dDqhYG5gFiRSctxtAKaybVxqjDbbE+PHLSPLQN/q6HXRmOAN
Ply5m4ruiFypB8ZyMgkP0P4MASUIiynwg5QNcQtkl3Hrfv9EhV55yfXXYGUO8ikGnzNWforNb3Fs
ffMxu4LS5EdSF9J9B/mKqqn3NywIoqCjeuyf9aNx6QZaNSLcaJHCaf7GB0ZWgbopgyB+3K2O6+V/
qLzyyJmksj1PZmAvl+szr7fuLoaFVYH0Z8zheswrmIm7RPsH86ntKbNaRPD5xscr+BZLdgKCH4D2
BANwi/UQyWKNSRaYJMCBUaiTV29/UZm5CLNBcZ1MFtyY5G1oGVMcXNoqmf18vzKzMcCD5L5Q6Cbv
GWWVu5rveGapiTGSuySgSlmm6LU/aYjei3ZJm0fSRCWeqRmHnkpGzxpNn4mZpT2OiV873xvc84qQ
+SdYOBBUduDJi2bO3DD15DMy2c3ghkSNqPp2+6ySrVYp0Gt+gtbrYl1Z5G3Bfsg7pfXTdXJnwNPI
S+Z10i15xQcsOgMrMeSqdc2qcUJWRU9Jig0YOfKtXrT3AiwLmQO2bp0+gsLrcQt2vZZoYRQ5SvRS
fhTWpoIQZd8uSXjDX6E/xaZpdGYq/Q1JB1pTmysUxC9kaVbsJ1vlZ9cx6UOlUSiLa0w3WLNMH+YZ
Hxa8xbS0yOUKXFZQsm6+F0nrjcqTIY1iKQbTmD1GPFC1gFY1sSLfpGdFsQMJWRm4DlDALojGBb9p
U+PDQDYFu6hf+UyPbSla5IHe/pL0KPNTickRAQhYBr6K/wU2LQYgdM7nS+EoVY9tJQYxUft1gkaw
XqpB90rAkgGmm6yd7BfwESAcXVdEJHONioP7idi5Qoa9Rag118M47nRCah2KTwH7ud0TfboVmHpX
q/VdWZGdDfl7kvfs9geuQnCjmFLIbU9Cc9EfCTUi+8mtIGKbaIkLMxKpyJeaFJnDp+zPHQN9M6Op
h8jnoFk/4TpD8aBpKqlsLsG+DIQQQNpp9ZnzrQ0vhm8eojcNTJl6EnPdPS3J9aMArhvxhuC7XDrg
8mkB5d+HMHU1LEjm9KTsmbwnuYVUIRubGFAuSvFftoBaiz4IDdCVCeVQu6j6RvhUWy8dKJxp9IOv
krw4BdwSrOTiZyKjE3gV6dvmYHxWjC1DIdHs1Pzj0UUS4hWWD9fVhLjYGQtY3JLWXH18wDpzvQVw
D88iFqAbqW4/R20v3SYUqDEc9mYvn5j3zXpl0cUquu4kYYjZAXfrDVSVShooQTAN9mBr0r1XwKOc
EKHTvtolEAa6Gx73w60d5JbJYfIeF6ZtlwJL3ucY1uxrPhN4pIVctksoBVEud9M2+HWM8p0D26ZB
BkxWrkSrlFpO5LH660M3YIU21bqHhpI376eKGkccyjnqap4rVF2kuDyTH/LOLbB5I1rPjkLIZA70
ZAjC/tt5YH1v3v8HyuDFZI9hvaOhMoBIzcsyWMNMlJjE+RL6JE3xTFLhbm+79aS3kY2F2YZlFQeT
vCZP58Ac6QRXG8awnk/RZOFjkmmgnqh0kivCwHMxktHbHtxTFvEKbDoyd4YLoHd3i9Q5rlTQVrgv
GSiLvL55ZH7+wijDPRD2C5uP5A0QoBRDXvhFA9jVLQ7woLkigWjh4ir0RjQuSNtbuYjb46bdpBFE
GdQqx671ZWqLyEsjoWTDMKTojT4ZaCaJL9LrR3FX/f2ExgsPjg4Cwmi1HyFKAgEWJP7SlPstwHyQ
DWnBGRNWltvzQADjgi8FMLfvYGHbnUvYNrj9D1m0w3uuSiCgkXeztZ1uDhUFufrRQqL77NDDjGxs
VmAYDkLl+SkL3COhGZZL3RtqtHXjFhC90MU5oo9zHzd8a1onUJvn5fQSKTnCanaTYObGec2yEU3N
zadRg9AJTemGb1mxC5vjFC69EsXh2WWwTkw+NrSFaR/NpEZW8esWRDoiiUJmXkhdFLLlulVZGA7V
T+2uGJIroiln2TFxk58KgUqTWw1nF9E5RYhyntVICJjCUMSutIEL76ChyCc6XqGaTaxVdzGis1vn
WT951v7mBYPKKXDLqDS2WXzoBV1TwB1+hIP3Bxj41pTjWpAOEzztOEPp5MBK97h/6CZ8or6mWzfA
MOMvlz5n68D/dyjb/ence5jgKiiBdg7vxaT5XYHqbxH1DFzkRCOVljEp0fHcWBYJOKrdPFI9fKYm
HZFIzHvnqNVE+xwTa6gqcq1ydTdj06/fjmmJvxZW/k3izJhZhOoqPLq6Jxd40rmV7ztyG/wsegfz
c3EBjF0nC1k3WGB76CbsESxVIOGx9LH2PuTXLB5ZdSoaefvNhv+X7WetgwF4vrAeAVBdtK3WDDPR
kbFVF8cz+rLxbKO8uusPUGND96fkBdH/VJa5Z2aif0MS4CxEpqtz2eQB8rZahy3SXJbe8+8nmXf1
PL5MpF0zkTxn28cBsloq5s6kYfeIgYHGhgqZy7pWHUEyPn8WnfU1ePRJ8OeQPh1y5NH55jCAxiVz
U4sT81ngmSkP591ddv0vviEkEBqQMSNwSDKuLmIfMARm4wSKaEJuHub7fuBQZXlFeR2JSLV8PTdm
jue+q5axpXhwH7t+U+Bg2+3IPy+kiatPW9io9LL2kTizFmdmWs5Ras3RPPT/5ac/y7tJg+Qkqg/Q
ARcwMmu+dY36Bg+gsT2JNwkN+wmvkOPYiX3edc5GG13uXHvRcMXbxt9t5ijw5p9LCR3PBgWxfeak
U92tu9LJS1lD+7opY1YVVRFKO0FSjd4PL24iaECXuK6EcdVwCD5GkpzybnVdTtS+B5290Gi2VOdQ
c/uDzqJF6E9cyUkqqUNigYWkGAjoz1rpLAepUw2ZN+WGGb2bUblAe/ejZ6D1lkF8Zs/nx4hrpBA7
UI/+diUBM7vAdEVVtlAlTu/P7fb9pLh8LGix8jtYkd2zKLZWWlLrUOccydFw+838G9N1JuAzNs8X
s5vFATJNMv536y77JRLcUaIuxkbsFjzUgjEFM+soMHnLzXYYwniBC7YeqVIOYpJhWk04mhWYY7LQ
6AHmRl+bdXyp/6eJsJtvVS2YychVJRZyigfsIycas+dlTCOa3go3UBCtuWb5lJQeT1jGXQVu4D4D
/hIon/qlkU/HtfEbJvQz9IxWv0nTCTXkPkN/wG68OfwF3F2lc5kfXXpmKDDui6s5gCfykmjhVZOj
mq/Z5jSjq9LwoTi3bZq0GdGBkySdSQ/j5e0SciOR3gnmp02ItoxxNLfYZjZVhuN4U5m5j17Dqi4P
9Qkb2CTaFSadqpqCaF4dApZmWZT/FlH8BBNDK5TNJEbFAIcCZ+3DVcRYfprZoJx67yGYX522htif
ZYcCCMLj+uHlcsQBQZS8OTsUobjFqlPHen0Y7jQd/AaMIBJT/vvWllt69GDF5nYDhSpET3M8xqN9
5N0ujOYlmgeinG19ENKEin29hWrOa5hlIPu7kJIahsMMAlXwsz9paKBfB2rd1L4BnHQdZNKGLnrE
guorfFjrtnxg5g6xuccQXVKr9tejGTCZZNAoKjEktl0etmCO7d1z9SQ85fOFSygnPy4KzNw6jy+6
+dOhtHXA+UA2GSKGKBsxS3tOW9FKB+Toc4klOj4YFpzp0lX3p5cYX2limNG1oqAYDQAhw72BXurB
OqpiLor5TVoy8pXsVV2kTfSrlKzbOaR4r+JVSrKmb8ugV6z0SXA5Ue544j3tEMuS6gvtO27rEWGO
7zUKMXJ61fWUcbWIf4J4Yto8eMp4J/gIKJJrTu3dn3uUw6rr3XfC1uTqkkMheltFH4lOXzjERxa+
iZ7z9Mkc77TqS4BYnu/tllxNatIMNVOOfTvU/R8l+AfZSCPxdcNFqnj9eYLKCp0YwPTMuf4Yk0gF
sntijxNsCIfnOloPo53lxnN4TNfzkdgPxxrNGrXlcT9iQExc8AiES6L7uFH3fpiePUrdMtttWAS/
g2Le06j4+Yc4EDQFIyfGCS90c2iaumYxTm9quP5VYYAYuMSpJZNbBIOXtXhyqKgIND/S0Va+Oa53
nDvoptHLq9lQ6wMrOIh+xk34viQRlVD5iq/WRV34PvckrWxTjJJ/zTbOxn1OO8oShsyuJq5wmDB9
LhsZYK/CvKZBFo1UfxexsJhLu7YSugmCKKvNMQBiSRYwqiG7BnQlQIO8lBQQ7V0qRahD1CwHxELT
wIaj+DZQQ2Saxm+JRj+CRH5VPDGZY9v0mkaNSpHM6i7x2vB1kSm8hd1KRcUUfKwN7h58/+90Ovd6
UZvlcRtcXGmaxSrTTuPHsWk85z1uzyvJtvzblvp8Vn2evnz9vscZfu9FhVaKVHpL0u7mjvdDvcZP
k3qMllT8wYry8CjDCzBujG3iTqqc3dlXzDvSA1LAOABduKGOQt2d1MYR3Xs6evZ/LnE9K8umqVit
nfCu9aGGiWP5fZHmDDzh1ZFJcY6GD7Tc7W1gqvz/JS656cIgdaocD+NGR+SyC0yv1B49bwj02o19
pULnkgp5P9LAonvomCJQ1SKN18wfMWNnQ+JmQK0X/mh9nyMj7XeDe/tvI6mdBD/oDore40PwAG/A
233aSRNBvw035hIVbHEL59xUv0BaWKwORfSl3Ezs+2mL9g5xdg5ue6R6S/fxyMJcfInQ4LfkSR5u
0tlcJmMSVNDQjGoCD+H/q665fdSQcTMIbUyKKplYy1ZLfc4BpvWTqSDYhZt4qOnyE5P2/Efxcw3T
XZ1SdLKwAt1L73xk4ZE7Ht+j7sekbNFojVr/QqS+qch4NwwJ1ZFxxsdDeemYgTCacD/ChpcScJs/
ZqT2ncSQlTKrnpPzvjeHmB3c3icXEm+omWGOLF+OyIHQaCJIfwYw6dZfVQY1S8rMP9AvqtjOA1cu
0alKD+8K0rjqGgkFZfYCmo+G4qpnaPBrZHYGVZuUzD1l7+CU6DX1B5oV5U+UgVcUT7dmbXrTvERf
KpcdcxlF4r5ooaaYQWfk36i+NEweFFnGEhxFdgtPHJMJsgcdDOUN1W4fxzA8KdJN0smZVOKaE79r
lfhZSZj8FsK064kLEEazcrkZXve7mu7h1YLFinmimTOwx8X+faDsuZfYPvptcyAZj6bc0TxXA/I7
c70XB37uwTVNq+DIkwFIU/zd1xsQglK3xP8MrEcIULLKgGeBaofUXQH0lfR63dgTD9xpENv/EkM/
AJEK3CnjhMfUlp+xatNoavyC8jtDdiyDP4xybO2rsuA5NribrUaJfAYTfdp5D7BAIeCifpQq8WAZ
KH3dLXEMmoZQBj0wfqrwjQX4ECdzJH3c+Co8s/ETDM/NErhISspClgGp9MHXg65EVZ76pfvHiQgl
jT5XiflUkOd7GcHG/iz0o3cPfzVc/6nX4Pg/CHXclEq+FnACNsAgODiidVkQ8MjcEpTLkSYTuLp7
3BLdd/wNQhBg0caPj8G2W7ocjA8xytSXrdKpLuUHbIVwYHi3nTrU7EaGOTP1v+NK34CnLAhUV4bp
Xq7n+cY7OKgbLADes3cnN37D3ohRH9Fk9jRioH9UQjqPr7yks93cGXzzj2NJOcBdgvqNCk9oUeEY
vOhP8wYshR1WMSbTOmC4Dk3MxYdrp6v9goN40CkCMJmPMdLFqGjwEzAd9NAdl63XwrnLqQ8/Sc42
JnmNJHYaIWB31JkAb46kwtIKn9GawRXaICy4q/0e1HLX25cvzGXCOVb29B9gIySsZyf4TPdOnsdp
n0qys9FxTKk4g5Lo2D9x2xRMCaQURv+VW/NPm7moUhaaSPArLmhlcLwtoY9kR5/HwwvKgX7zudf2
+47AhjzVm9z1bYEqkFlaokZOD3wouFEUMQXdmWsJgDdl5HUC7AkJNwYLlRSErut8kzCehQHf9M6A
7Gyrg2J/S0vcz8bz7a1HlVGdZ/WgdC154yTq4l4jAbYD4Ii/mTyjODTzjwaK85u8UP9zlxsAgQut
g0sxmqDRmIT3vmAmepo0lq8ov5ygOSokvOA2vk/IhEgLocvdQuM4BagIhQC6/WY3GutZ0so8HIIx
NUHY+46plVcLPKs9nIQ7jEdAyPO8iW1jpwLECQ8ImqCN35eVnU+4j58XjiKyZMXn3tHWvJYG0dqw
X/Hy53mOTCrgHpIFGCiVSugjHKT2v+xvNE3jjQOjB7XmvwuF6fMFlmsVvGc2UodrHDcIdx3GKHKA
Iz9kb5BzAuKtzAtCRDXRdoTFqr5YvM+I8+81u4ibsBekIa5UED0R7l1xxJVRWbnofurevQWqSbA+
BwLIUmRLTQ0CN1d3nQILqBPen5dTdWWTISTWNPO8ww/mVotO7TgYndPNckSYZkX/2G2HUh25HJNn
+q9ne6sn1QgA8yjOY3PpwMCM8y/E137eSa1xgYbq/E+90vVijk6jFLMLVvKhJBrAW0/ZIIgXWv0M
B39DrWWjWCQ7ZQ0mFUcb4VDAqY9cENmXad9hX1Ooah3A9H6zPQVH5fu8xjD78kmgdlQvvmZ7L4fx
EnedAQ0ZNIJTT0DlLRQxafVJTqLcrmFLjO19Yc9rPAUnwi0HWDcevSdPCZKvvDUA8cH/7JU62SWc
m2+qvRdennoXNBnpJj3miNa3wvrqoZDQjQ5ptMJrNaEXAlNymTexNsoGAniA4FDrgojsMRxZh6YZ
0B4GKgNMB+Zpx20oK48F24GBWhZUJpS35fRgoHA+BIlgG87aAQs5y2ZllLqoysOaSLaNrUFrpOqo
tXmLYHUh/eFX2c6MYpWkitOVxsIQC3w4TKuaWqFq0wzUaBE4ifsYj3ATgRhWHwr6JDpSr4MCYstq
NitlSoU6oeZPOzYJNgDgQ09dPcLH8pfHB31KdhP2xW7meCHMSIon7Tc8P2lGdmjgWWsTb8xS2wYU
vPCEmRnsM9IGWdPslGHbdLABtx9HEjmIA6+p5dbn45H24I6zu55cz/3fRI0VwqAONym8wdJKKxle
7hPD750ypQZNLKD9l0i3kZaWJsRi2YiqCBNg+i4a55IAo2HXIgKlMjPBsr+zYFGKgJDXTm7KMsV2
FK26Y4Mmudz/Is+F1YIRcy5XrjXIV9aAOSUkxCnsF5nxpAWutuZoiBOP6mdbJllb3wXJObTuXEiu
HrZCrcqfPA2ZR+9TkchFTXrl0bY4Bj7lwYxgnU6ByJpbrKNudFZmPb1FtBBvj7o7EQeqkdypHc+9
y2brDS14QUCrUdABIyptwh/XJ1Tkyx4K3VWx5/lYxMJt86D1wiKczVlgXUG4ZyCEs4tTJGYC3QAg
9UvW8qL/+pjH0J7blJndLNY0dxCx3XsdHQta+1345XdzdHvpkspsbeESDvR3wfnEvbGhLiD7H286
zR5cEX6jICw0lR2D9I3+4qzmt8p0Q/5/myMkNPATHUiNUp38JhjuR4G4CX70uiQmx23KbL9DiCHs
uAMNr5C4heVwVnjf0n8zrOZOo9LZf5yhp5fCXzfyKhNFJIL2VaSp7UTKmESOvIVpNwKW48AHqE3h
vMtpfdxUa4rZAFR5CKpni6QY2fZnJrAaK6rnGGZrTxE9MVSTo1ZaQPlJwnNkRQzFRr8azJA72y8d
OxEF4a6gEDrMDDHzFSrtwFlp8ra8+H92GLU0cwIppyyu5nZwYJfiLafeDqQ8rMBvZwhB5tWePAgT
8CNpmqedNZ3LZF9nUXyPtZ0VCv205d0rOsK1eO7RAMI+oU52BZej32vt8yp9cJYFaEs3UVluFGGB
H5jfvLcorRlPgR5I3LomoqSBg9e4AyDFIKZwPIqmfMJQyU+AjMtpe/rsY+DKH0ll8yN8aZjxBqHo
zNJ+g5jyqZKvNminhHlcigdXZs9yh8yttG8hzLDvjy3FQdmcLREp5KO/mXMvW26ZsjOzSn7vqI7Q
XLW6jOF7scZx4qwebVahwLoBDCe5CLmktlZQbizMr9o1XS6GZ0XaeUkT2zDuuMdqi19mr02XbH7E
rkf+Cv2cqdOiF4zI3ySr7+ldB7m5S2YhohZpLiCS/T0/Ms+cmMYK7pfl3zupD5cO+kfxAbk+OYkZ
e9+HYzZB2LuID1RYlRHnAlwpWBBAtUVHnHtvVsBfMBV6ghe/rI2P0oDCqCYAO7WXjH5XpMrq7GQw
KvEx4ofR4hiZCEMPqYpkz7uqO41N7lJdlaA2ShLtLAAbOZgPEgTDnRFzg3LWe73YDGT7kJWv6TaP
PMOVWShPbadGNjDsdivLiXWYdWtm8hu17BjHAT42nK2Fy4jaK9iYJr1/t5mLeJFYUkEEElTqYWEf
4B7v6o3uquCXzpbloQn5mkWDVNkuDA9mYatzEcQTgBNGzFPRZxwFOAXy3+1CIEzRV+2bMXGh25xQ
2J8Oj3CbtYBKpFL4hhBkCcLtSmr2GL3ozb5ZFlPuq4+zes/Pg4+hnObPOGAMetyPJh8P68RbWAWo
jUCFODAGe/N213e23zeuVwEf3jDrXTqC0UfYIIcanC/Al0uCQ6u1zdtZMs005OYkbXZZyUPcwRCD
iZukZ/JbeMB0E9AgK3z1h8xVmaTASzFRxqGkaXY74r6Mi31CH5h18JLwuphuBwcikyf392cK9Y2r
i3niCvD/10zy71P+mJsxVvVxtjnOdYAIicMatDZybNBHyUXIf4po3i7MQOncmE7Wa9vG70ctS6oL
hW3ghliO2bG/3HOEQHtYU0fRcAHxm7Bhnd1JVVovOqBKCgbPzEMwSerZLwHXxslgBMNs5D2W0baK
4r4D0mwPlWj4qQ4DAQvzCOjooIkKm1kC2EfWIEbXS99tyG6pmOGqWkN2UOr17N85iL3zTuHX6ZXA
hdkew3E/qpuK5JivAUaKuLxglyiaRJvpLY5bb4a1CyJlzhlAEAGJRqlfQCMfxW9j7obYY1Ac48WW
gTJDNjddLWGTXOjLwPWC6SRiRXvJaooDXMlfKxGv+gQgqugvkoKrdcftonvOZEpj0E64EdCgYnmt
LJUpFWOiIo4bv8qZJfSjKf37wR7HOOJCTBQ1WxKtIgJX4s7g221l1WxiEUvq8GULerqszLMxGjD/
hj+rFEcB1t7210CkIgjcH1fOWYaGOtXMMwcxZoPqEX62EQFWGPIjoQCBcBRngAsdT8j3qxft0YH5
0cYZBlWaJitbCZB9dsxzN8xGVjEOLREKjC98r37TrHHUEy9W25qYKSogEkej5YkBgfi8KKNGxXqR
or9Oiynzox5dxpXT5GzlFnnS7Gp1lSKCUiQThaoM+Mxltl4kif3aR6WL3UHCjh+h/FQ1UT1Ul8fC
zBlX2/34HsSdT4P7JmnL1il0W2wsG/k+53wXKXV/7pzlw3nSmgssUWKEK6azp0arvsB5oQ0KnaOT
SxR4iIYCu4XW/C7KUYhlYzR5xtZQXK1nOnxQkciYXHroDBdIbWJ6rEbytx2IGwCFQyZbcNZi5wWH
EKYcK3xiHkWJn1k9ba0UA3EZmEZu2vwG+CL3zMQFrlSsctnZhnccwEdP7wFl2bnEc41ax6EK6OcT
8vjWJy+FXzmAesAg097sCZ2wchhSjYefudNb17J1QatSXv0aXgCQhB9s25HTLAy6xlc1K5Fntp7T
Z1316kFi+3l+kqAkFb0mxyOCLSR4su0KXqLKgx+diBVqswNK6niV4MIZ1wtqrSvfnIu4EGXQblEV
dNQG2rszftHU/nz4kUJEPyLv8GGD9BjSSHs9liXM9VeTV35nhy/wUa5+bHBZA0OZlMYHoBP0a8FS
KJ1ER6TDTZhMJYUETEbXI4RSb/3Zobi2F1oyNVRxG1NcclFsJdI/84DCCIJuKY3wz71uSasM4xnf
bIx+8ybp+r407OYa7OAjuIIm9KTNYkFPchY8IYDNwOu109dtWD/OkcQ6KijBHqScKEhhwN6iwvNz
6GsQ+N/60exj/FKEa7mky/ooikZV2kbJ0zwpRMio8z2/1Ddiap0lPW4vntOesyuFcf6mh0tDlSgd
rSpIZTa5/D0Kx48A1Iv164+b/veQ4dIQA+nE4ZnvnPvRl8Sbih9oiBbJd0CeDYyox8JOQD7JIL/G
RVr4Bt/OXHPpMnYxnYNnLNf2oYR5wgLQP0Dfe538AyJuwXbLq4B1xX9bepIItK2CqeovnAKDG/Gb
s4BIeRFAtxj7wM6me+glxnGHJwgH5+QAv6Pz1FIF7Da5y0yKIHR24INs28APdK0ZxoTqO88SpBqo
kruggYTNHDw/yEGORWCNfKKBjBZG/t+1nY/nJECnQayKkldGI6EwO+Rf5LyMUynqY0ilVATqs9M3
93UhtNP7TSuaSKmNooB2U75CsuaWEr3J39+ojmoQNnZmhMN1GTivWkNsAzxx+WFewg0wMRdw/wyx
IWPfEXGmnopckvJqINs87I/TO9H4o4uNFDl4riSNxQqUX3UXak5aPkilMu0H2ZuicBto+MLT/CfY
0eAlKNasSLEnXaHTzlmDuhK7YXf3zR3ytr6Sk+eUJViJ70GC7pWLeVDVZ5goHoZgenmMqk/LpyZr
WuuZZNO9Z9XyYAqq/xmDoFkZwtfCVyBU5UxMDb6LESu2odbdQP0dNhRBOax+Wm0bY7VBg5K7to6Q
ftV9I6Wz79/hg8+2wx05KR9RP9Zh2KEneqlwrZqdty+AEYPBMqJOIv5TxJ2U39IzAXpsVSnzIJGK
u3zyyWsOudSd3iKeh36n/HH7e5Ytbv7d1oH99oI54EX9wwxceDR7Vjckqsk3OPvsAyyZMgXd0pC1
dRP3Sxw065yHjUGYSU1xXCjLoqKJmAC+GhlZo20RO7hc01jCSDSo3FhAiBpADHu6HmLkiO+TSwpC
Srj71plpLnjSL/QCMSSSuWmVr2LLW/VAn7gj9gWQEgt6VZ9q6t9Guc8zKu1B+Oq4gsMpba8zuEMg
96h1+lY/f1j5NKltix8H9rVel4jAfvVi9wQyRNCCLtRrtE3yN/vl+n7T6ZayRXOokMVWLXaBAuBe
JheO1vj19YlSdrJB9XiKLlNqVN9qXMHiNa/L+Q0SIDlIfrl5P9qbBiMxfYFNDzCjfoycyXcp9XiW
p6lOryA6NM9i45hUD4OnhCiG76lsExhZu9PGeGem3ujqUx0ZPeKsmsZB0R+5ctzHJC2AQ0EP4B9t
/Y3NL8twnQO4RVrhcQo9hqafneny+6GNkMlEhP23/4WCR04sI/JDWMOrF715t656dG8RJA2MRijU
hK/pct1wGQHK+YCALLQS2o5rCIeYNN71aZ6I67CojjsC9LVfxnHMV8Vi/fjNwuE+6pVEkyNcFhtg
EJXelXmAyILHPKUSro5Lk8jNzs+1bla1Zr92XgInq7TIx0b2feixUbEWWH00pOE9pxBkhpqMPalX
COhUPCON6Y4MEFpdwI1nwGkE3rTtXYi/xQ98chepi2zCi22jD9vT7Pkb1SyzRCckxtqfXLsXy6yQ
5iCA86tBExmQaitXfzwit9tzlFbNeLhAD4Alle4OjYNTU880EVwKHLpZ7MvYXQdoTjK6ZSBqzOs2
J8K2u9nvhmeOghA7w/pPAEKbnFV+A9Zj8d5FU2SMa8By7L6bAEGUT+jGx3BpKUhF8nnPCaGW2usG
wtGXMRodKJHCZ3p+Qo8uxOR8YS7db+RchizR/kpjfbCqHeYgn1CxL1l9i37XJ+c9DYGOh+rKR5bF
uuuuCvSk3Op0U9cKi/mxK43a+MhohRNy+jsEGWm7DwKZuJwkvRTPr59yqI4O5WFJwddGo862GNTw
r85NulOujcAisc3ZRY4knBeN+zCIuXujK6oDpQwJR5/ciL7EjBZXFAMuokqbvusBLo3sF6pSLyol
YvZcws3A3j85wRc5MGAo1p1zJRdy7lr1LVYfSMDMk5IKuLlzAR+By+/Y6yn4oBhEkKYw7kOslXl8
OV2wPHwnEnw1hDOr7hrFm0MMCdjRgp4m4gO+MRPSeb3GkjcdIAWdgPwSo+cD5GUNecOh+1NbrF4v
XxqYXpY19NQMgwj3AjSwMtaE/+GPEZf9J4np2ENPmElG0dgnRZ+AoOg+X6tBaYg+A2ROCDbE24P1
jgVAqm9tqKs+QQ4oD7LHWyLaKSEbp5INhz1RfuZvc5aS99LGrnn0SopCuJlMNtMtZnFCYO/dFTEy
2lLP/xeCQutsY9bgta48CS9n7J32tFYk4b0r2kl41q5OA7H6cThC5uI7QAzYupUlXqB9yaM8jLJQ
+qvZ8TSppS99SJVS81aezobKHIryZhnidIni52sm5pUit4ViTKgFgdlTq5/6jSxIkTVnkk5UX5lO
coWhLmk5gBzEWJANzVTk/LYfnUDMn3hv8CoMBks0OOABS9DeqT96kkiWhtVnMGsvNpASDwXpAl6T
vk/NDs4O37n/nK5UVVVCV0MGhiTPsrNDKxy6DkkMpfLQIC5lZu3Z0TWf1PT4Jb0hDXVVq1KzbtHz
PFDK+uaTiTdjRKpyrVvF+uXVoYuMBTKLufKLQe84tYEyrouxrWUoClOQAwd3zlKqWLZ37jU7w7CI
a0mc1NOInBC47DCWLRgPDwTmHGG7YgFdH59BGZS9Bwm0p8bpbobjiRuHt+yKnRR0z4UNIT26y3jr
OkQYv7iactVeCQiVQlMzbB1wXTkpK5UriJQP1gfJISLodcRjSM8eztO1jGFPw2puRhQed87Dg3JJ
Of7ZvU7k7TVTllHchwHr/+Sd3W/u40bI0bIynoi14Okpq1+UMXLy5AySDDVD/RSCi1k2UlY8gtsQ
4T2Yao6+9j9lP7OWWlHWoSkDUvjHw+DyXcqo9LELUiPDMUaHbTj9X/VFFAlXg1tY6h0Jcd2deGPW
rHPE9zVaMRFdaHQNhghTuMj/SZkN/z5x6iehqS+s+q4Gn6iWdi6mEZiXZohlY0MVJbAtJW95WwW7
VPJIck/BTs0avcOHfZUOBK5dcP3cWclcPpT522uK5MCInopvES3Z0WfqFH5rXQYl/uf4oINsx9xO
IUrG0OZbvWtbbr70SVdnffRxTRcX+OdQWWfJEa894CrBL+oHJ8cpERJqn7Uqe0+OnsE+A5GmwJuB
W8GwaLxHYVo2Cp6P6Khk51yLAYyYUGeCjv2OWLuUZJYtSyYRFMa0dvY7CfzJk0lqflquMod9t3bq
FCa/uddmGiXkUTgUMp/y1z3MnLV2d/EnuvZpTSdj34cXOH9hjdoX9DCMskindUR5wza+dQgSFMOi
VUl+7ClEcWhfL97O+bSk8HNx44rYPHEURqejE+U40SHvhsXMCuxYVCYVHZ4B74t8rLjN1RvBSYoZ
yqWmuBQ+6ka4nX3yUyCAis5GK3oG7qgJT9KJ/8+/4cH4hvmXyqs5+mgR7d+F/rfRmnzpbtK5o1MH
Doi5r4Hl/EZINy/t69Ah3NIYfiZlsflT3MwbFrACu61Zf8ejN5Icw3wS5T9sVxVkS1FpX2VlCa89
8nlOiCsJVocJEKKz5rJdGQDP9kEn8HKktDdbkiBdswaVAs3njjF3i8mIblf3LJ0b3HwmNsUmYdoF
VZw2GWXiowiL1TPyWnthDYv1E5U6jKlz7LnTWYo5G/swUIRtys2EPbJ3upobtaTee///S/MLfF2n
ZvkFRR9zO1ttSLgxh75pvaibPrDsDdZ8I1vgtpsglNVy0PpPTf4G7E9NpTNKhI6eis408GspKntA
9l+BkF7VwIuDUL/N2Pd0m6tskjuQixGeRZFYuwPsiar6kslQNVhdbcE4DZzusYQV5o3lR7KEn5Z+
8LlU+mgrSlWJTDUDLjcwqIeZgIzvZUZChVeFoNj8Lb/vbkW+58e4LCyQHUtO61OQ7EOexCrHhwet
68oun8azPHMx6qVeoJUUFyj8skcuVcEX50EAkd0agjJ71ahXQo/q5Zlu6jrBImeHvMHYoaHAZq0w
8gHMvAYGlBmNbbKPBI3p7ic3LAday0guyL21yvcApUNLQLE/dSOOPaRXrllvPxArlhpyTQQ2lU5u
naA0i+4F46ZGP4/p+oQiRpVkucfM2j+NX/zHu67nYAahPhpmTQEbZHG2j31R1MFwvxUeuZxHVO1E
gVM1RRMqdEm9KJ9zaaucPDPkbSc53rmF+AzLzRWJiAJTyGofGsm+usM7rk/plwTXPhDCPYFFA4Gy
4+5RZ6JC+If8oD8xfv1HiR7x5dvWnruiS7zYyA4GDuL0cTLD1KhHn4J4A4oBh3g2UCdxQZjz+0Pe
mBQLRwwZNXyQI/vYxqD2D89XqNQEQVk7ygqr/wnSBbj89QX4kVFBIOEjVcYsm1vQC82MgivGRCkk
x7z0RpkGpqaRxyE93RJhLgMO7yL/soAQJ5j4k1K+zRpZP6j8diTkr5EhISDujPGMF080wK/WrxDw
Yc/ZFkYwzOlZr5MuSFd8LsHmQtxfQOMfIUAPPfhoIjbbPX62prrwFZCOWv/wkSOQhdKLuTdFx9q/
8iS4/svVOsy5Q6gX7ImlOyoH7pK1VzPEQTg1179wI+6Y6IxeBevVIQP9hkVfiu4hzCh+9IOcG4O8
08l8ggzqhTwar5zT7vJAlhCVjyZGFPJCerBy+xGZxcQstD+s8xK64jb8TzKdS238K0BTaz3o3h6c
PjCOUgx6nLnbd1d+L8umpuDYDHszOK2UOl31aKkl9wnye2mrtDWDTpN6uZciFe4exaH3ud8/KqbZ
wdteWLqbObZGc3m+lIzwTvnqVReSlm4+8ilXD72eVtS9laOJ2c46QqE4FsKgx0kiPgBBHOeQV8rB
x+N4fSxz/5E087feAyQzT9YmCd9IkK1T/WinSaEp5bhBxcaw48V7ARqghIyc5XOp35ioP8zNy2Du
fAl8W5lkuj2YS2XQTW2YMqh2VGEmvdlCh3U5og0dYRrjfw/OMuvXTOqZ2+O5E30L3jqQ9LnEaCUY
iKpwQlPkP7ZSuMyVVtyrZ5YOpnZOFcMoxtBmDsts5hMDTtLSp5/Nklgwoa3jhGhWqfJgIkqNLLGN
0Oi/FktgSTY/W52ZUAUokGMslZFqhCvay++C+aT5q4/HzEkTL7LfLuxjqZYn+xsWzOvchdmz4atG
3fRRafvyWI64B0cboEnELpv4bNGg+VuFxo8aOtQF6EBHBALIcqkHFdUyQ7S0Qct9gawQQ4F9OJeM
R3xkQ/m/9pxeSk/SQmC2rl28d5MCk0sNLK1LeAmJm7CmNNB8Z3ZBQUebLuoCcq8RLO639gXj0B5Y
V7NtidSHYoYql7sxskYfs3QyfOhvMIpZV69opFN9lniES53NZQAvXA0t9Nfaqzp77gzCb+OkfkA5
zqS60xAE29O3WoU90L1y1qvyWdFzfywBCsPRBLf/1g8u6pp+xQrEvUtlP2DX0Dj3iZw2S1igDYOh
uFtqGFK6fBVjw/EzXfzw5ako41RBoymqcQ8hhhoUYj8AdUB4QZlikQtDGw0ahiuwIGnG0LC1AAKw
3kC9eDwZeRMc2/Y2HDXJuZG3flB2vbLS5nnScdoui4bEoTK3bj7LW8nxcA0Iyqv786BVyt9q7Noz
hpbpJP2B5J8fTHUa3bP4JtMLKjado5Ozddge7voA4GxV4S5uhQ2gMtDAml8k/yyKjlPnpJs+PlKv
48fO4+REO6G4MdMfdtGUVgAMaOrNIKTfw6wdQqzBhufGPzYdsUXfT/USz2tPW8jBkbydsHkKhm1U
reoB/+3/aMp0sJ5JUcL8qOTEnn5EgDSjxjrdcSGvkl3w4uAB7yh8hUfK8qBBHoIxDjnbobHWbxKo
sowdt6KC6PkYorshBfqk4v4XrzVRazeE45eq431rvvfpNwGcZd+QZgSIebhbccu7vd4T+tpswI26
3nfrMUGOgmyUsh8XgFPdMnVx0K7/z+NYyETz5H5qJR8Zq2S3XE+KmZG2oKgIWCASsCmC5syqb8KS
GbuU03vIMTJyIYNcngt9vDvgSc6PBB3VcmY5dGt+qQY2Dy0ka8hEqXhhCKCCQ3AVrYgwkZCYHb2+
bxVQse7ZGoBBTgoQ1wBHebmQ/sPaahH6kagHbCz5yLfb0/nryepRlVw/buVfK1XKQaKwnZNyN6wK
KVf4tPdfPwnFVGr5qyXraFNyY38V1bDQlnYwsV3a6/HmHONgfDU7AXE7dh6vDrVtp9g5U3RPQKNn
I2cfwMIJ3aYUr0wnKSdABlrYuR5XCaq6e8xzz/RxLPuL0410SytDA3Q571H+PCnbMfKWqFSO1AvO
ArSsfsBIGOzUTQQarZ+/Q9uxnNkfe0xFwotIdhAVoU7qHGRk1RdmDCww3uk3LpuJ/GtgNK4zjLIC
7/Ke7mmtau8sMSKu6PEEWazkjmIQTSSNUWoCQM6oCauTc4idKqiccGbj1b1essTQNo/42Mtq6nTp
zevjIWihPzC9acetDMa6D9sTgZG0M836Py08GQzBCpjdfaynx1hy1t6lgYLDyQo9Rk6PuFkU3Tmu
L3ejVTnKf7rOTdNAb63vGxE+hgw8+hWtsIVtzz+/+PMn7U6ZKW9aBiWx0v1BaCKjtSDurVWibdDO
AmjqPqKIZqo1z885eYX0pUubeGa3k3UO2ow5c8jKuUFHbz3OWByvYg/5UaJECiaA2wP6qnKkG5IH
va2bjclcBVEdiEh9DfJ9c/cQTRcrD5pk9bDbzbw3XCIgOWcdS9PZ3wl6Or/Mzsl1IjeBTt+h3UeW
T3wCXE9jbIkDr9kJHPDmKcT+arOXeCWrAP/4ZylUb4FscNYLsRiN1H81QMZlpfTvG2nfLbDIN3qU
FFRSKRo4/ji3ECRPi7p+TPUH3oESYfcOpLa3uo3JO3ehpasr4fw17FsDnfrKMGM6FNqdKY9pmjSc
sVg5ZqjqeRF4RPn628Juh1EPX0mYB9cnP/c67rY+cYGbSVAaQ1jtyzFO9/4jei1MQnBmHbp7BUA4
y9ZBN8mSOPFGDug3PLtS3n1xiuWKfwf9i7r6OLJKeodY0tADyAl3NLvMiBCcuo3XkvYjNDyd2rXW
pQoTCFPnvMwgivJS4Z9uItK5WHTSgvh8urVH9JYVRLGC3hKiOPBVnV/HHUHUgewnYvF/hdj1RLT6
VpXbufhug+Gxfzw0wf2TvK270n8szfEhKF2SVmo6jKWDFRhbqlX3NbFF9EbSQtFKbS/fvSI8hwLT
j/erwX9fYFpNycmY7h9AoYBLJPLzWsVrYy553JajZmfvaLziQDUgGR6ZA0v7ajx3DrGquoBU24LZ
nkt2aBTp31YN4WszwUjpaVnk52V7WQyYcj6UH6ol5uxKe2ha26VPCb0J5YR1gbeEpO6mpBi/eSdh
SgPUIKY/++d4jrPHlG9srgUE4+v3g0s+uRngOQQl+pmLpsiP54+gqmmBzQrcNs5U8x0h9dip1aC3
4t6Ndj/axzT/JtfhO0hrqhZIygay5tooytLPEjT7xwDPAlrlO4GKxIlLrDtGbWmm58CfgF9p4OJJ
vpCqn6XLKs5dK40qVWiVphKXDVuwa8ZY9wJFYBi2GEstt4pA4IHNrByVWYCQW4NwZUkXNGNd29tt
OPGdcPOKLzRJjbtuwsQkke3rIp/vCQ8RdNkF9FlI/XOH98HVOWjfLz7zkYGcv7/s3w81OvZoFHVY
vMXZCf1dtBtdyxHQHERba+hqgSL33ode1bsPinKW2se+WIAi4denLIUksI5BNYLAuI9vUMewGkgO
+yGMG6M2Ay2qZKFk9W4SHS3Ro9wx15qLs9vaztQv2Iz0aqQRpTiuN9il9LB4OxJxLBmcjl6F4M+A
DF3VSzdcFteEg8L1QY82nkhoD/XHxbDaRwVGvt5U2OiKAMQgONbn84wTA75m5Yk6WizbWFC9GdmH
K/gUQj7/wPR+PlytI7P98+SOJJh7THlgdf0Wu1/vdNOMFdSZ6JlJcrVD9RrZVx0ORtsk6dQ2sdbA
6/+UtNPqQ3cDKz9CmWhqSLY0hgFmk3hA8YkyZNKWyjTziQsIws/5plRUd7NfKoK8F2P1oFQI3D0T
wNegR8GHzxEOVJdEE9jFaMkfbRSOphCJ/nb3/UIz16hGN2mDRpH1Sdu1jjdoICs3SMC8K90LHm71
6swJ12ZipzQ6B7TRzmWzBmnxwKF3UejleADuS0Vxl8BTw/uuABW30/yrFPAYSpPMfalQ+kbB9u4d
vZiWv9ZOO8kEUe60S4aHxIgQe1QWWD3ENYhdEhelM1/9rAELhbzVMHu0rVNtkafw83a1wU24+4T5
SqAyPhsiW84HO1rzWwZ8+JgAgheqTIxJyr7idHsQLSJbV5Ayk9lx6jyUAxWIpTJhMasd0ERVbhJD
kgUgKF9LJYHgcHM+uWmvO98MLgdd11403OZtKDglrkbc84HM5BLxPI7JYW6Ys8T0AOx/qMvOxrDc
dERP8edAaTIRJeAmDHqNNij4i6So6fQ7JDRaN7uZKIcK1kXKS+EgwcCmxbNcOTOYUYUUQ+jAnGRN
hIZUOIJkm9ohXb0+z198Dkp7i8cVIMqOILTC1LMBd08D6CEN6ZnDOiwUKPGOBScZkCSaCzIz3D5M
0UE9xbgDAsehx//HCF5fffpeifVyl5/gkKiC8ii3dNt1U5fvLKBv9JW7Kdv5B+yXSgU9nV7vspIE
pBOdvcKLEONDIW5V3WOWpRKmyf5WK0oXc8BNHYTl9MAC8X3bf9CfVZ48QYn/duCGIREoUKOPGxdR
dWAIH1/Ey76SJiFa0GJMm08tWr85b+ftoIi8/xGYvnlng7lMXEY/cnNB9Z9phsreiVG9iX6Dx2ew
1WTHNfEq6BfSEAucechRAxmAhAnf6umIB23L1os4JHtAKOi9SAGQKYiy8RJvmuNeMeST6L5TK8MN
itFBQQDXuw/6mXAOVJTtzktYSDAO+u3qHJQl0ROjnOLXmiKmbNX+kf8mCx9CBeRNLcNwOUJaRdZS
ggHbtEfYeWO3YH+G946UdVQ9y6aGMjKedecKov/TJx5Ob7ZisuT2Jr0Ts1PjsZxhWyDPTbN4lAcf
a/xzLnQrPgf1iFb7ESqut05vEDBfjXM38tbUMu/UKxz3sZc7EwClO2l2cF4d9UquMGCZ0vQsaFaF
Io/JHXdmcJMbnFwNM+NtQocLzpQjJqOQlW5VQPCEO/fsCDg5U5IuTAMnhqulEAjFd3I4apE3SMtn
E0lRZwdikRB2dTwGNtb5mk1dM7HqBGXQ7LE406pHYSV+Y0Vn0pOLX7namyYPHedacgGUIoVJuumv
UK0+wOec17ALcIfWkXQeYUL3LK484cFxXj3ngMdVgX1rvP5SHRjaDG4jMnQpjVa8VgQrXmgRJLK2
1ZKP+9FPhMjXT2zpsmdB4Z61ynkQ7RSob4EBA58kMWDsSrCsK9gi4N6g6z0Eoui8kKifgFY+qrVl
vGFdAzfVGsMg740ak6FgvT4JPJfx4OtDUAZICbAcccWpGvRzFRzKXvIdftr0otSiRxjV0sVwiL0S
Hsiipi3ohh4nxeJZoqMzjaEHTUcwBRS3Qj4WVrCpV+z2HJLvBZOBEP0miU/LLPzaV4dDEYCHBTWO
QxbwerlmCdFKu5YRliMgnohC8BC7tx6SXCXpfXtpWN8wkHl1kfS6M2TFH3GL6wd3iZDqXICYA6qt
pRXckucQ/tg7GxsAg1CKsYTsaTueP2fSRI9+sInLsTT8jrfVFsXxQZxz6NfgX+ANLVbdGKhOCsCS
++Gz2UBD+ahUu00L7XdI/c2pR6ll7n2j3eBllkVfbMq4qaCy9vmtkVA1yVZTMVs1M6PVO43RhOZO
HE1UvHwY7Za7ljNec9yO9UKg0Pgd+RXsiXhGl72hfCr0lUxZM6EDzjrWgmYvu2x5AepoRyPoqfER
Mm0erOM1yFDQ31xtA/fFpdKGsMJXLzDXi4Acb4igpQtGwDvqywBsW2XtGa5kdQDpt9tijiskgBQT
6wnUbZHaYEYlQhpHx0YuOBywSsklrEqp+DnGvI92YCq4KfvrtB0meArwJkeT+x/gJGEOnMKwouoB
qb0tTJIq2Lq651t2t2QqQRXdXGgo0ZfHIWfUUN8MWx1XhBDMZtlukRnEUTATSFOch2uXuAEwBJ5G
/PvHeM3kLfJzmGQInzm61tBzx6b1K4CexoFzsu9U1siGGSjt7Lf1yngTj+UprG82KzX2SzF0uxHh
W8zvpVtTpykedihliUoEEPhLJnVoq2xNt0hMila+ErbZ3+PAgf0qtFb+tsjIFfAfs03J95jtHP08
f/bR+Tl2GHWiTgdt2gyX5OxjgL+0HDBC+2J+tdCs+EP4gWiyi6R1mBQrcoPqwg8iB3AeceRBGIcz
nfOsmoJVCg6jtxu9Tk+qSb+v4S5Lekc2He0IFWmR6g/nfy7UhcJhi+5mVeTMRCSskuq028riqKQO
kP52crgkHX76wOAuxuIoMoW5010eP3JzbSJfAL/JC3sxjYnJrQHPDu1aFOYRBZAHs0mrQvo4viez
leAn0bKLJcjbEP3PIWSvYtEfdeJznFdOzBGCXN7wfHmsZgkXA6LZmYk/bhCjdnet0rvJPhak7IO1
YP4N19wiN+TSc2v8X8gLFUdJit0jy4LEUQJSGg5FvJ2jkgRY5bRGwWZWtrbndoKN6/2Xsrq2hL5J
Wer3fgWyCuyXOBNGwZ3Mu+a4JGJI7T51wnUe2CDXKneNS1ovoWdau6zg5AzWUqfmIYa5w7jBSSs9
Fgv1oYgVJ+vf/Bc9m59woWd2AhOoZf2GfeowFsMZTqFabT5VbOjGc7oZhAd1J0eq8wZaPyueGkon
vuxxDeQZAm3P8A/EHajUO4WlN8kpY7iTqK9iPVsMF/XI0JWjkNI/GjhukmFFpVVN+L1ezUf1cPcQ
4B8Lle742XhLcOTsn+kcfhrKMD2im20yKHJJWHtb39tGjLbVD/TZRaTOAV3jBFQVHizuzPeewtIv
fkvzLO/7W097iTRVkMyLwLPa1SaD1h7EH7/Q8ZOyKI05Mxy6eZAnr2FEsvH9Hs09MLQfT8jtAAJn
SxA/c5TmAL6izJON3EUJrtNpG7eOWrljp6xRFpntoMF3SeQsj0q49FeR2NriB3WQuT0Fah/hsLff
4HfQ1ZwVZ1YRUBn/EcfRYArUWKQkp42o12pnXsK7Y54MFuQ1c4WdGiBLAhNOXCXAa27mUTtcXq9L
LYTAXAb2i3fgAUadG+Bgqw70jLro3M1z4tr2gY+fyrtfAVl/0PmngWU6F1zScsy//ZU7EI6dXJyK
YMcUV06ch5Ql3M1Exz4T16TBDVrWU1+/hNPIryqz1I+PBCASBvsdpVzWRIE+tbeChzhB3U+HL+tj
ZibQf5ZRndRotBjJERqFMuJ+AN87f2NhskrWA1CeeQTrsQuQQ449JnWQz4qu7hvS4Ws6ZXYYnusC
XZJB0aODwrx5vStEkgso3sLbV7nginHeAHwSfQkWuZITHTsjl9FX7KH891grffOt2KRewDXaEv95
T0vp6hLGs1l37CHeq3R1DKLtAiOVkJ0AG4E/5QiuWNl2vPQqKi684vwk5kQXyaXgkvkZlcuUBzLT
dxGCubY03013i1zNjr/8Pc7qNwpnC77SeWCi/+2MzlSThBJglwyIPBft6yH/KK4GHujnXxTkxl07
XSA9EkaiCAWZDQzmg25hA4Nd930uosMocfvL6qq6ScRFgsgpO5YXBGoZwSDL8qwmfUHOLoN6T2GT
0tpoeaU/dmouF7ZiJzTK8gFoUXku+kobfZNsUaMFH43lVq5F+3tXzkqG9N5Yd/0o0VY+blOZ+F5g
tsO31ywL0WTgTZzYonDXyJQTNe9AhcNDydwu3bhKsvThH58EypvlX0mluGoRvHACxJgGHO1ObGl7
gBqzzNedVr6u5v7uYrJrQB7+yUx11xv+2zLZ+GAeHN0UjdQeS8ZzmvZP5+3a770FwpvavtkAH8QG
LxqZzR+d3gP1V6MqlZYy92+dwCFjDVI0CfGbhCe6CbRVdTZrXCURx8YiMaxTNFa3+efrHF8Y7fD2
JcCiIUAvUxPyLGgNVOPHiAbyqF7L/kS9YLT806YXmFkMbCuVT3QkC4E1mfAw7mbWKnNUpAdXVr0L
IjRzUb0HefyieMbZucbHA7MOfj7G428r4rKsBAdVAeV7xG9+wUL1o03rjqghW8NueJ0HqDosWEUz
DP1QiXla2+8yR325YcyvvW3gGGfr344NC7On+zysIJAUAeRxZsjw9ErWursrVgMRGCACbLPiFfcL
A9TprTa6PLWexHl5ZmTeALAqkQosNYEUv9YjyaXkIM0R5B1pZbV+02jRLPNYjc/lXH4ghp7djz8l
n/fTzCw2tBizeM+9QtKsjFnfe2Qef3FvYQFPwt3psk/9kqpUPIniNkxApZ0YnOcrgBJ2DlzSA/da
KE1zUdd4dD9P2RO39iDbMWE6m5sdp2GbiefRVhBAxceIRgWXZEuenxe1dxtlmriAD1YeBkpmGhgE
UdZWm2Yy6bJGHdfLfvonJFs4P5tsftx+tQJ39jsR3c9oChjmYJrM79MaDZN0CHPfoeksEFjhm6r/
+Mn5wkR1jmr+RC+kaUrmB0jeBKNaiMzXLWlSmoG5HsSBSGdb4eoW9hJhUTlSyzBz+ghuETYfp2o/
HOEz/6T/IksPAZCiWsWqd3Wv1ldulyDJfzZCBtNB4e0Ko/aVH7pr320fk/vZlWi3mHYiav+YS7MD
HvAP/bc4J0HmCZZCik4uwREZaZckjP9BwN2Oe0//UBexAEdmkHmMShL0G5WHhxUgmwwZrIc3xb4C
UcvOkuHhazv/9DV8E81/QU0qjybZMLb5N5xTgbEv9z6HLuJZ97yfM4XrIRWf2gYofGirq7c/xM60
jme+k+W6blhVkylFbYaMnAllrjIwEu+x7a06EvvMb7cidyy1MkZkTUHblm6jj6M1RaO9dMrCI14B
EnCDHvhocxrNqM71v8yibADdZtvcKgcUtS2BwQVmENLvvIdfN8zPJbLuskrA3qf6lbVsHiz5vwGl
Jr3fjjbnKa+zbl/W2d9GbCRb9Jla0UeFNfF2vmoKSeSqKhM8D6+aUuyj32UPUC63X0n4PyQHRiSl
fiCfdEjQZ+Mj5OoYBPFjitr3+pRaCeYRvtVs9Lpxhzz/jwL8JMNVI+bpOTJFf+X6iAtSwK4dEfgI
DvU73x9BKJrKAw55+uZHcn9P3zWJvi3ajBe5unGtDUlbX1C/bCE1Qz+kYjqHPJRIA4od0tKgttDd
XZeFDgj/a48555uIVQ/DoFYoDVSnDKI4AMgANJlp81M52tuBoNlGssMiIGDp/65Ay0qFloezw/eu
QcqYL8OWI0QrF6W4nCPFljoGi+vqvrWNkCVnoRFsNhsMaVbFeDBpcVs2JjLdWQlG8iMX7nwPMyT7
GcFO0gdDZEyiqzBvlvufBA+bjv/A1OVmG5Y0INPmunRnj6U9WfSs21M2ot6FPp5q9kMFL6OJcvkM
7feZcJpuQNuZ/mt45haoPZQnXa4X0fmgWrsFIhVlm0YpcR/c6VXbTKFCnR0eszUt9t6Kb71j1QpT
3QTUUvUh60cT4iQxjXSjRJgDGKpxOgmuXbinjo0OYlKMIAWl1IKIO10EmnnUh9SY6SJFOYaU5UaK
t01R8Xx52ae2muRQWqflhgfJloMmosLINULyU4tbNzS7Ch8vqMAhkc5nLZNlvRdRQFNu57WTK9tK
6woUHByBx0xrMTFNgiEphTEtIlfk9Xl4X6atDQq67Wi+KKZClFKIpaHjbNhp/VzrwxEJLbR0IAwf
bkWpRBRC2f5XdtpduznVvQRQMCf8pOI5dyPVf+Y/HcoVBPOhwcPtnJgcJjrrayS1GzaeW10vwpKS
hweE5htW5buMoM0WbEXMhWxEWKfM1TBgYfFntU7Ek/xRb92CuQ7OKEZqVKbWTD6zpPqAMSB6Jn3Q
GfUvzEgxj/LxMfT1jvCeC5G3rBCtbg1XRtTotgRSr31kdWuDkhA/LmYw4bdyFXIQiJpiAmj9GyoR
Hfx2oiGRk4NrajUBbiJB6XZkhDEVKKzvEs8LJsDWl5/hdu+EiIvzHmcBCMRrjQoSuONjqxRMQaDa
LEv7Is9nHnIq/zom9wvGoeZY3FNp7rm0vxGSHzEzfzCEeubpHOLFEtKPsk2ibyq5uM7u7dJtVjBP
eeMYatdictqBwoeQDF8A2V/uDIRMCqSjiMhyQDftcL8PWO5TQCIXNDp/K6Agjt/Je5wrm7Bd0o3w
0fxGDEeTyW4fu+lfE6MD62OCusB0AT9wIdzSu/UE+0CYefP6Rxwf1tfgKWClx8pwj4w6JwAcJpbm
AXtGdr3ZaVnwHFlSu0wbtnR3SJO9SusN0aaZGY3mSkmdVFqhWT5JiPqLFnn/8TL08g8f8iI9+Hlq
GCGIh4xJiNiObDXScujpfQguBTQTQWvffSzpRyyJxZOn4mPck0SkpYwhjTEjhaWGzpSf9y9tmv+2
Mizpxjw/i49iKBTN9aif45AKlgb8h0Ach+nKPJ0wl9V2uLlBcAvwiTPwff/jXZO9Zxn0vSgQujLa
wEtjDUK+922lF6P4JdiiKYI/n3bKMNJ/3diL3wpEg7bc3kVHUTYkNzGqGSjZP6KdHVa9i5NHo3v3
8+2McDOIuty/ZRsyLaFgqLl+asb7cHdMFWuuyiJ/2rr+xKd6hMgDfjzlex+pSvPB9zfSIHkWvZ91
cG1nqfUtkh1w2BKnjzF2HVtw0NLbUDbhfgwOJJo38XXknPKDa0KH2WGWyDKoiu2y03l5HiPf4GMF
r/y24wTRoRWfVrqn55GHS2H/K+L6v5drOrAXU0TXBCQkuwKa/YyJvdP3JpVQZlsnoJSbVBed5r+M
CN4mb2Aj7rYxqQXwRvagOD89VAINNdSP/0zKPOhtRk/sEkO4kJdTYc/eq0mlH+l8CUi7Vcn3cPKD
C/kiLlDMOT2TrSRwDh1cSneZf1bvNLh4YuhOTifbefDcUDImKRXAZym7DVk99vUM4ZpPfcqc22es
PUDfgXsoakwrsZLl/RJoYCOPGKaBh6bXMRkBGTgZn0cRrWBDWcRJaH84/NDuW85kNdcPNNtl8Xjf
79kFdst781MSZrW1vY1pf8RzzujQwQMw+XyHuZTFICP46/ogE4RjSu97IgUxrqDWsyS/lPKA/y+L
2VE8oxHiJGMw5AR/kIalvCO3OIo2LsRXB88fgTZ486fE9aqcUSXbf+4mjZkV6VP7oflSdOC3uBzh
DNBHL892rZnlM9XPj0HgsboQ8CybZg7+xBAIoC/695A+8I9APZQaPyyH6HBrVuw0QqsR8vqwbC4B
ArySAjC8q+cPYzQEX2zy6NO+cp5m2HM2BPepTSEUSe5Zb0EXF4q9UZSx4oNBL/f2x/86aaqReawo
yjT+RWRHNVvpfQKKMgKhPawZJNL6gbbWpzQmrd5yrWFZDP0XVFPi6fJWYo/ipb9pavewrdIaBHsz
TBorNTrsIKyL/5WA+365kp7RLLgZGnAYOBQySU78YBM7wvEPOQHBZrNPYBfbXVZliuIQNypLAUOm
ca+UR4FgG8xS2QJ8KLDndcKJo3awdsZKydk/bXu7ti+n10sNuE2rgZy6NGH0TK3Ic4+Leh3NvlBz
qPjZtjY2TxHhgwxrZM2FdUnjhAFF2aV1+JFOaPNbSrB1aUQkPSF9CU3R+QkBCFvmDNofXCWAKd+P
R9DdyZq86sbWwOIVTTLXjuLx2X4oRbWhzunRTKe93qEODmxXCGvg6Iel1c8n6SQTr/mIQJaZXIde
hQAvdH9NnGYtwO6nXCubHFyV2XWPs7CMpke1WJnm5kzUR+V2gh0qKBlirRsJ6aqAIlnCe963ZQnQ
SH8AYAVu+ZSaqyhgUFSmZ3XmJ+ddS4Pa96klj1cdwTZIs16KSwyiyMve7iR9PEf2RZU/PUzzdunb
MS8ASBFjt2Pf5CXVMhZNNBQa1g5O963Q3Fgtp81jKga56rL46gGkxaX7cpzkOvPj8Qz3EKyGhd8x
QbFEF+fWh88EXXL4litdN3eLuVvUJPCxl7Y2iyio2OWuzUL6wO31nsE58HI8bLkUxQ7bq4eQdifT
pli2sv39cdX/Ew5p1dRTv97FFKdIcTXzeAnjT47sBseVpwckUNLenkCg6DE4eNnjVGc9QgU8T1Ml
ljUIvjVo1imISHdG7/WXTHy/Mq2WSofj2m61yhGXt1Nch4/apQ+agRRtxY2wxnRB0GSbYCCJSUXc
qX+tFvhHbGarqr1mVQ7wPr9bYdbKesAmTlrWZH0CtFKFTKe4mXPnZEgqN0GOTEkWWluA4ej3/BmV
ZfS6zi9NZOw9GQvgHk2XFgAY95V7TNc0nyfIQLiMM40BIaSr5hcY681JQXbRa6c38DEMhTLT6YjC
JXDZhuiOvJVmdUqc2it51SXLr9AL0AyAmzKhktffVdv1YZcGVSc1aQqxf+P4mc/TU2AEW0Hj3sy1
YH78+f/pwolwbx4aZVxtvYGzVdwtu1wwLJIL3+FID45K/mhr4kIwO02zuSBfR34Y1EwHyaqd8ICm
vCoY4IuojhDywPzBfwxmvIheuyq8Vcr+0g0VoP3ESEyI3ICDy/UBbNl1cGrduw+qpNCatB/2KSsh
6oZk5s6x7tVGsVBJjwI5GRjrz0EMRLyVyRJTazB4LCxrRa0FVkdzGzYuNmCZtQbcZMZpJHc0/bai
6BAvaJxO/vMgVA7lHwVyBBv4G7vxRBSdThk4VIfaq/VIGRD836I1pIXHA7+4IrF3dSpznrrfTgtu
w9mYi5NSRlr3ezvVHV3l0gLX31cUXWR50aCflkEDLAldzg/cU8yPwt/M+i5BgoaUdwZ+XURTKeJz
xN+32OlZptBV2LRCqqvz05dU3MeWoTbERcfdWSFzxU95I+cnRGEjz/hL5Wkb+biVhJTXAwKOJIVO
9xMsaZGJyS8NWk3JIII2QwWHMEIbvSAXoy6wMjiqJVW9fPZDGbt+vgB4MmS7HzOMhgkbD6XpOpr3
oOTb1nkcTcUuYorXxAlKqwYjfn75MiM/oly/+G/hzKTvCqek61T5J6+wtYKYzBS3JNzFx2iU82O2
dBWbe/FMPYtF9o0GSvAhIKMu7e/vgJOaSzwjxCRmM/oRPQqrXhPhNLVRX6hq2jmoxOzpDL2GcSUB
Wfu9LXVFVHOOKwZ69Fwoj2mEDaHK7sYsP0YpzPyh+dyzlEqgWqmN4IEPaqe0Dm5K5NNf5rpH0Blx
xV8y98SywGTGH10smCt7s7dBRF6F9OMXYFXsH7Doa19zYg+7WRooxte3xcpxZnEsSJkZlmhzNr9Z
XPU8iKMhUwhsnLizJxqBCpXSTygpy5KPDp47q0o8G2MmxrkJ6CG/z3+0Tsp+nHVOCCKJ9NICqVpv
v5BpDRJFhFQ56zOMQaTyB9Hij1CSW9dxsUjWfrKpFSMEzFH7uOQW8TGHa7/KEoh7tzAn5Q/u33SH
11KymfFbCh7DzTp5/ZC7OzADRay3vsRAXk88fDdGrQDEfuAkE7bdQbfSW7IRlsSjTaLbLTGTwvfF
1uBWGeAO7xDTfSA20UWGM5iaNaM/BFgptrRPB1tzWVEsGGO5jVAJWmdzkOy+gAh1WlkC8dZ2faQm
IAaoo64Fwh4mVJ1wlE6aUmqEHz606AT369P+Nvmzq9l94ij9XTk3EHR9xmlzOQAzMCr3NKWt//vn
p3cVT8e2gSVFb8SU0JCbfOMsc0wBL/z+ApLzIUQyxyHyF/wxvbmhvvNwk1IoEFqKxz5hvXt1SjkO
LBiccJXdS+fs5JAzWYFXqhqKKW3A5N+BWAXz/Sc9uqRdT/DtUUNPdRTR4SGPPJdz1ahDgPKm5kRz
MG+U/tPqNVm8n2kARJkyRNteb7r3WcQla7QMIZc2IiVSfaDiZCSoqa3c455FrEzKXGz3AiOH8yKR
c0HxagKBwjUJ/wGd9Rt58pLFc7HPyoGT7zN3MQDhalqInDM+7Jaow1SYToN2DC5K2kvAox5RSmF2
vR9zAeJC2fn/q5vTCrvFqRg35Bnfjxldbu5AJJoW5BkdJEUgEjd4Z9NTt1Rb10Wc9E8VFNfojpwA
n5BreAj4DiJtTxslQsX6n5ZGsk7UTbT0Jl1lCag6qmaNzbwpNsHXu2ynwprXvbDb0woS/2OBFbqg
4KMX5AmfQlvRaCj7zW0D3hZKxnP7SqAcMuaXy8VwUGMpvB7c5yZRQB3KrG6MHDbbp7gLl62uKHLj
JX2plnOsjpwUfLYS4cKTJWiWmwuUnrWrcLhD9Ri+eayx9YoaeNkRU2Quq6kpbUw8RWmIwGM1gSgo
pLnUmz502Hv2s8oqBjQcvUUki6JIPKyCfJ5Kf59nZgJ2RTB4Cp9agUWQfA2tu6P6wY4TCuaPkMZ7
iJwYLt/ckw+fmeIvESw0P4598K0yclY3x8BTllnNsCAZs/Aua7fC7S1hvCvv/vthRQ/V3+vBMjAP
n6aguhpIPBejc8xsv7WdmEIXW9GHaK3beywDO4URwGfBkSUKueIyE67odWwq0LvZTfBZccJ/0WOt
kCd/CUNb/BPh51ZWgawDikmqJe9SBYUdumLuL9gT8RSf9Klz4TjjcRJOpCDuOWPHl9mNiOsCR1SG
rU3LofR5FKHolQv2tmFIlS0oMjrk1iZvcZf5aX51k5mSp1SePuAJAZOf89AI3B04E8XI6MWy/1f1
k31X4PVkleOU8CiX4ptKubv6aezBTR9xi9/OdhY6Vv5Jqn+ucOgv0HEZKEpKmDxffRbiJImkUakU
Thg23CegbWNf6RZbQturJpOXbPM+NRTnKZIpx7+AqOt7LeMw6wxD+kjZqL5x7uoSUSyFeEqIMiHN
S0Egrw4nwYaNU9LWqkdqYWmtYMLQrq5S0Lmsg775oZRyRc66lywmO4Zdw2hkmlTareiggTMbDtC1
B/diwtpBCryxyRikr6bmY4hHF2GjNqWEdmBItqICBhcJLiH6Czs2tu81CfdE7Yth1H0Tdg/KfnuE
vSHP+Yyva/G1Stwsqmb9c3zuunhHQIxQlmCUTbX8KoW4psHnxws97O/TXuGxygwOxs7kupC+jb7a
8JoYrD4HT2S1Aw5rNObQtuApGLYs9SdIK1WNG8wsIwvLQfW0ZGBFhT0eP8p5L4wkeBgzcsuiJpff
e/D9T8JXw5LRo+ccC0L3My2uUCxEFkZx1329wo0VxQwYRoSm5JTjajgxP/0KbHkNZq3XMVBXjQDZ
ri/Ax0ZBT8uZYFgBoHpNXX450YvocFL6UYkxvTqGOkKq4OXwdfYYKhvw93afoBy1uqYqGeLAdWCC
xuIbxSe4gmm3vIMLqu/84/6HzzsKzn31vKEJFlBbOCXlNUf3jI5sB1klcZEiUbugxLU9s3prWKOx
9zCOcToe/6VghUpdNn/9aYOsDVudPUgTFg4g29nZulxFyWTiq39pOkpJJsmGAKnZKC0yE1TOydFc
AS9F80JCnqPUfD736CYdLIjH4tagbni0aS3y6wsLoeYhEyN2ysVfdG00vIcNDdHxHQunMi3lDW5t
uUdizSN7Ra7vr+O+sdnaUzTqsdD9G5Wlbp/zAcF1Syr4J0fymke/QYBO+A3ZYaAu47zObsMDzC97
4tcv6MkSDmrymCKQ5HRAp2WAi6ifeFt4uYZ5Af+TKUbi8aXflV9khjkqTpmPAR17tPJEwFotKS1O
Fs+JsO/wG1f/cA7GB/q4fl+2f5S4gfLSut2QndjuKY0twLEYWgX80seTQeZbhs5IZm+QQNCEKLYw
A7FmgzE6LLzb8nj/lHE0uc4SMaI2WEaz3Vm1mCxYuanM3z9GQFMZsfxDz4jdcKVsOThbNVzbRPbt
9x+gwFw66a4spmRi7Ez/fZEeOCKpyNRLNqPSgphsWU5Sw96I3t4f2gitZYs5zN8LU/IePq0Hw2Gp
WRiWqa1Ngg4Ug3CAlaS3tZvDmCDQ61sAj2XyHv0KkJbHN4dHqyxeIEkWLSTTzDYmjBCFJkLOUUMx
CkOjxUwHcQfIkc/yphFyOetfuaIwOT2JyxQwnoeJi0WWzVQDR5VctYqYUCKHPb55Rw3pD+7l6zWq
6YZOkXq5aufC5nJQT+GtF8cHz65LkiFYsihFtwyB3qSPE8n6EVIgxHElbHqMf3QcykuE15ce6+Vw
UDd7ngAs50ClQt3o2AEcN1yLQUAGidiLKk9pbfpe74E1oOpdu+e8Jg9+59//j/60aSq0XwaBkb88
KQSkYGP813aOSoP/C5oe6uQU0N1CkFth5tqItb48Miax8PXDKbDHBpEg1BQaD/beKNZBwv+QxUQD
8CAMPJ4apgiZDICueuZGBO/DnC3ytAeiRW7duJLHnMzyQeprJ+Ndn3Xvgl29XFeo6KXpRYOIvaCR
M0mKwcJl5VV0EWByNk+YOCxZ+tt4rL2np/HDCI1F5vEh2n8GiMS9rnBdljplPwlCQ7U2UuZAVNEJ
eJ1+AYOv1vaXr+lV8KJC1hjAIH9yXcGcq+8WBlCpA/kJd8MHIWj7eTzEs8WWYvFt0DOOqVoWs0od
ow3jxBGNsGk1XMiTRnyN5+vIWqeNOD/qHpEz6nmRpnUnLiYb+Ty3DLDjdklvkPBlE8Pg9bd6yrPn
AXjy/lcyaiMCs/7yv/Cp6mPxze2deFueFHJu/RhZ+fyS3XwfuCSCvDSJIWEMQVozLYWFF/EB4ngR
8gojaoUltG52pdsbs064Nnro7mEn0tR2J58E0pp54/O6qalYc75NKfJeknBTFOqipFECklGWrPVK
B9e/Oi8JLB8iHtxM55DW0WHPHf1p9+gXJ7DdMF99g+XyTP6orEKaN6bN9LLvhdSB43QkUnsNqLk9
zqItM2YJgoefH5RTRZ4ZMONF0mU0oowN35goOxTT+mRjSM0de8wK4wfDDcTdLPR2pst53+E6nUPu
nIu0YqTgGpMfStaBaYLhmFtxPOELwyFXn3oja2w/T0rkwydRBX8PnPDVUnHpvE0aT4L9DLaX+uf9
pU6nft4cmsHKl9VZyNJ0HALNgS/SQnm2Njl60kojTG+2OhueosvznLbK50Zw/dVuB8XEA2Pfa3ZM
krvqb86srIt9Zf6NhgeYkRgaqBoOU6hGeqUXNAeKYoNR6BzqYQRVkMXWFt2Bjy4xyM3IP9LvdBO7
18uWRXoPISmvrb4D7MU43I+kGJX2wMohRsmDgcfRm18f4kqUxLccmcRmkQoi3KXRYYghi7jER0Sj
hHy38a127RJIBx8TEUtvuRZDWf7O6w/kxeyP4FrkGK8Em0zmiiHJiVWlF/RklSZOwoWwbITDN3gw
lpbmhEdlfZ8bMwvYUYJyznnSnteeo+wqMkn5y3/9+ydxB3YTJLhXAaYe7Vyky7ZCnCdXSWHxoFpA
TgRH2Aox0K6Cnb9AXTd9ic+ejxN9kioPwIEGxkXPQO6mdWkW6tjhNdxFHk7+8kOkQxWTsqyGubLc
X02CQF31lEY0DGx+rJkjNcN+nIKJ0qRf7dHfLrWc8DlsoEd5cxKDdetTvacNSr8gWBNyWOOYW0ID
5D0w6Zuxzh8myvloM7qGotykycSpbrY/8O+7UnphySsBS0E9KNOpgI4iEB3vInVm7Pq3pbTfdbF4
geJ839vts75XzwjAit47w5o3p25xLUKNCR1ngcfq5fNbIZG4AzGt60M5Yulnk39pqAB0Yy8xCJ1+
qKgw1NewX33gG19Ck/55XHvUUshpTVBf0z4DLza9zP5L5IxtgVT2R+HHzVyJqBj6DWIY+yahbcDx
KV92xk9sBKVL/6QSTQcsCrem8zP1mgLGfIwE1wsqgk87iVm65lcuEWxCIKAV8VYJoiHumRCwoDz4
BIm4XD+zdBZvBrO8KMTWRs9ahdSeWFAxHdl2aBirJKSnFx2kG9riaF1D0f6vi59cWy40CfF48hvK
qG6ChTnAUo2zsKDy50QCXuJzbAu20W0Lw2ZwqzgKP6gYe9O+DL9vey4pJUaleHo/ndCadRitXc9C
0UxUTzKHD7+VbSVBlvCUwyIaFb+KKeiLImvo2+S6EqzCQaOjD6iKi06AllsSsMOEOfmU4eSRI3ce
5nojlvpUuMRHXq2Cd38zdrmEHviBtQQkyRqCeLBPqsciTz84SUkZzikIDHRVSmM6JkKF3q4BUFnH
QtktXNgd3XtSBrkVYbCzd426xBtrEwUtu/2HlgyyJCvIFWfdwzJmCsZJkssjEjp7Be4X4xVpjFig
3uUXNlmvP3wQjrbxdY7BOPZTRB4BP1uGzAVMIfd5/0E0hacBFntz51+3S73IbAfjpcg3VTNavgxp
UHMJM8mhd0HSb2+E5j+fzE3I10N9/5oj5BVYmTsIN4rvAylngsQY2dF5Nt4cs4OXEyV5ewYSHQ9x
oobG+HYG00qlJ6+nFaOAAz41PlgLUVC3d6CGthl+4UL8bQr1Kxmkrh6EEaaj/g5h7pToQLv3gVmE
VcK7PRbMXwKSCKjPgXvDHibYDwmJX1H+mYujaCTQmsa/lY7N/2AkL3HkjwTkgOD4fgBfhAQ9jJ+E
+0Ag+PEp93ObUPVdWE/VIY6orI210llH8rA1hr3BalgAHu+IIeR60JJ0iHA3IIaqX6SCF9GXc5CW
BUGzPjLiCnGohPQcfcZVh+C2VBVF2pLEogGufTE9h9seOvFDoF8/CJljlDjXyDLzaQbrj3wxQ+tK
3wIB/qQ0t6JKFjtudGrzLUIN5ytHNW5JJTv3QfsYSa2vornuhLhxmRQBRiUWxsB5txRuG/5NPW8J
hNr+rL/axheZV7jDDKHA2pQAWasGqP7a/T+CMgbt+Hs0DrsfXeovK1J/+mTGjGjcwK9NqYfA9GCD
WfTjpCK7FafaIMQ61AWrmu4KgvrOvtZUqrX0THvlSYsqoxcmEp6VHyWlqaFi44CYfoqSP+kXsLb0
qy8U6+nUgKT8JHQSKGpXQdUJY1ebrDB/IT8TYGSk/0u5L/hp4pNHAeUrdNXG7Ww2HH8iTX6sBE/g
IKeXOs7psEz24uIB65m6TyknDB745NwcB2vWZDeyCiXCTSgG3fuQ4e873NDFV4CStSJ0uVqRELqG
s5R8nLbkwoU4nOxQO5PHjVi+6fTBw6EPjxJhpodnTrYqWIYWE1S6ISSNoewVjlSknRxXWemXOJsS
uW1qejrQIy0lQJG8PhKV065GrUaAk961hlQH2QgNOl0ApAcWEcGHXB6/2tK2/OKAfaY4MCR5WPOs
I8MXzEJ6nh7LK15hhgeU1br+tCpB7tMgAFRTsch3PK+eAUYabLhV84O+HLdzqNLOuJVY4CkqX7Vf
elGxdjlyFzzTljLUTitJVolU/SCMAcrq9mQZRN2iE/N8IbrMVT9+50gUWeuQsbTAAewbOjlP7KsX
emjU5hlJ9QizlellIJDqImz13X94XY0jWlI5vNj83PoFvTMz1kckmF3jkfNJRy7hdwnMauPmD+e4
M6J6lh/K0Ac62helTp7+2uc4PQoRqD1VHnWbPC+Tq4aRtj20F9tJqNocRWlTfyMU+qTpm4k2wJhM
r+nJ0bPJ5Z6gl1U2groMOgtcCT4NMWGsOQU1QTiOD6R2+KFfy8j/W2EUuLlP0teAcobAorshx/G5
sObrxkFznEcWnGhMJnywcXS15soW4A/DJbha3df4CNaTuivtTNeZ0ochFsQEgR9rVXv0r4NmxYFL
N0VSP9sNnUWOV4d9fBI3ba72mmtuUHUsirv2USoDUbc4W7584yyvHdQ/zii0PqhtBuntAxma6HgV
27JpEpDoLbRIiOwEWyP77RMNzkx1TBwtxd6NsNGDBS5toYPsZkb4n143vyuiyF9mG+c+AxahaIkC
8AxJn1mS7ER0+OyVvJrvjkT4UdM6a/sWL/b0xHoX+34Lo7VRdre/HkJmYiFXZxVtEh0eey0H4k2e
w9JcCbyR+A/x+EEXWTBXKzEf6H9v9WHfzVXMlJdwCvDM09u8BxC93pesqYrp5RjC64RRpO+0yM2S
2Z8+Z2vBe5+1u56Uq9nitjOEVOmt7Z4EUQa79dBAEtedgBrFas53+uSuieQqeWgKzWw7IULXRu3O
y141oBb/c2jbEzCUJpHnHPpNO5BcatetdMV1ozAxkeUh1JsSJtxxu6NsNu/r7Mrblw+OefoayIpK
X2GB6eRHKuG5zKkcoMCvJCq0f1Kn1gEs1Z5Mr2xlgCKboF7CBQuGEAMXxHgxFyBpgpfv6FtlWmYL
nxl048uFK/HIpyoQrAXvuzXiRtXJ6aGIPkoO/oJ8Q3K3QAwvdDWkIN/J6G4ip7Xho98lC8AVgxm2
LZ+Sc9v69OMA0FD2MTjSiFFylA2L+WV2e9R9JoEiw9xR0AQng8gVB9Ge+MvHAYepJ9KoY5KV22nF
eD4jkyVeouwS1au0JeuYXBXjPGpD37Aha8VDXoq3anJIgvfd84t7ckbZf8P8TXYFGUjvcqV+Q8eu
pU7LSd6zkXHhy8J6LBMX8MEpFGaV+a9Bf/FOILs1gnqJ1/D96ad9PuBOZHdmSn9Jb4Agjq7mL5dg
+mrQVAdAQwaXArDKcFEVEE2VsIxn8zMN8ivLbH+BDSwFPSHna8o2AF39z9mE+yb9mrANH2QDVzkV
gXcPrnKzdXKAoiGtkBIZgM53MLFQtAbvmEqqAU5o5z3cMTAJuhYftvUa7ke091VqMfFt4OGWGV8W
6+mOb6l/22jnb6dbokovluScxeKPNg5ZhPDisoizXVnmQLOjz5ix6jLd1FfaOzY46G6c3qS0YFSd
U4/0JYm8pIR7+LxJYXYOwID/5XeNW32/VsKxQHgTEgMZnOIHgqEQmJihQSCEZzNBcyFPLvsfM0Ls
6gVnqsGOCgJ4tZLTtQYMbLct9FE79kp34SgXZ4yrbQ4h9lc5LxOYmFe8K29FSh5B5rhB3rCFOs0i
NFhnrC2O6lwdV/Ha6gX9/x06OB580StfzSr48E+xI9Tq8XuYZAqjzXanYxGTLDyfPWefG4FU9532
DdtxgHQoBjhEAVxZaqp5FFm5GcaLCD8e3ONoILPJq4LM8YZMDDnXkFXFPIgdb2NYp2c+X/kSEapA
P27cCBwwH7tI3QKcVJWrww177gfJSaQcTMbGPe4moYDr3EDDp7dw4IWAkh5FsNrO/+CBLPOePNyR
b3K1X4CBH2EJOHuJcLY7t5u9UzXGGTMqkkVTYXx0wcv5l9bG1mAObLvF+JAYpnx5iLvQ+keJKryt
otGXXYQl7sVFvwjzUd6J8HO//Ni18HFlgQeETmsQJ2UkoBeQKCIrNll4N2t9suTkBDLj2ppl3W2T
xOfEXgRlVPz6HpPnDEyM2Wh6J3Y0M7zE2NXLBTNr7h9pRUTrCzgEUYW+Ryvtvg90a9H9mZV0kTeC
n7CANLwToq85krizWbNyUk3kPWBjIJwC6ImLdcv9h9bWyTxVm0SW0QBhb3rED4oSLn3Y4Oy1C4tv
6KzZVDsNpm+1AFncMBW3PETUzirbol2chEtF6qbk3BsZKrhi0Mmzpcf+fAbJInLwIb9HjGG3dZpk
qInubhGvwDSxX9D4gjS4au6RrPuf3Fu76iI07TNHCqJashtVkzx1e3FDR9S7L86V5Qxp57yIcr2k
DcC9CX1ik1ViVmFU26HO3tJvpPZBcWTR4g1Je1jLWF/efbmciRVtvXCXAJdXtcXkJsefUFSFqsA9
GHIdgK/Mly1POvvsVPkJ7VRAPzAW9K3zW8fgGRk4jFg4P2ThjZaP4L0HPt4sNTmN0N/++N9885y6
gZ3nSnHugHOhPfHX32gN0xXQ08aH3XO6ezKKELTfPke9e1TUtEPixfBTrDz84/FENMi9+G9CJrCr
HKg0VAG3+JTzlL+8EslhPfkZBcnv7tevPTOBoupF6lsFJsymgJJL3LMarJueEua/Zgu2PArBOH/i
tR8P4T5dVNaqvm0j5MFn5NsGrg1ywT6EK7BpCV6NCyNXxaTF1ZmC3YZ7SI8PHA39dECPkVBeAWQ5
qknG64T0fBbpul6ADWoe0nGjc2TTQ+PRTYvQLVYVqYviCbJx5mbcieGXTGWVU4cVH0MnXwYh3Tu9
qlZxx4SPvGsBjtlZXpqPA8Df1XX72UmwYI7dola1zAbWWBUYBbCyJ4lHWbPD8+MnQarDoBD5v/1P
ItDAWMupKZr+7OnRlGdSJlDSG5mzcHFxU7aV6GN7ie9a6QAlDMbnzQwNTjTNO53cReoH+7itjriR
h36dzISvf5qwsUPiJfk3EI2erkH/zKLfovrdc5/gUWqXsnJlofMWX87SwMvwTjInqHWMN82TGRwg
9A4M5glR/rPmgAN0BA8qgx2RWFMu7faOGxhUMfyJj067ywz54bKOvcldZJfKEYr+/CKPOzReuArh
K1cHv1pLri2+c10FGN2Bm3KGjO1niDZFeSvr9KQL1NjsDoqx2zZ9yCDf/jaKLtGPZwciBV3k/msA
9dkn7BZ4yRatehoA1744RicliUsSURqe1/qortxKuhB18AjXyt1O9TcXfMmLN1zcHsMNwinTzR4D
juRtlYR/l7eM3qinyNfRNGR4GfcXD2WQ2VWzqWyjiVH61reLI4i/g5opwMelylJZ3kcJPsvg4lZf
lc64Uu+cc1h35rALloR5pjSRF4zCOTaj2g8WlOUYSrctActeFvvmkCRnCNiVVFPTz7bbtsReHmVb
QjrUU213YQWgrUBtrtG/YEMcL0M+CTjFmhiEDUlWtEgvus51L8y19jnBewre+ld2G5Pi8lETdEfk
dWskSxEU6oP0sODpdPX0fCZk47CXKYLUX3Zjjrqbl4iezjWwduWONH2REG5+o+sIohozHq+WUmDy
dLqzpeXQSQkIVyh0AhfO9gQJ5/eke5Co+0tgSZPsO2rXyWMoSNlAiDyIyhGDAqIWNFGYncuJ//6R
fgaXDxVezUT3Gi4D5TCQGwyEoPbiPfnt/qy6qxoK0YTONLIHpbdeSGiZ2I3Jfo5mGGuL12T5LN9q
qv4XcR9/X5+Vs4IRlYHFoE6kBKTjVdy2WieEo+0mdBQUN4TpkqMJdmu/GX6Ql1OTIyKHvP7CnTpl
x2Rs1FsDzWUDNYWd2TUzDslU0CQ7jwNpG1Dn+umdtW1Skz1Eg63M9bEycpYDBUZFvXr/JYlyipaM
OplQhom/IiexPxr9HKq5n6UqMfVaeVXeLmmhGfxXyfQRT+uNhe0yuImEGm3uDeJPSUJ66cwify8o
yj0/Ibv/mjtlJ1Rsstj8liRBX3wU1MA+534D9lEBB7d3mIyl7DzsStB+qOyloW1LjcFlN9fbyFo1
qrosQIFxfCvBVeg3ookhhzrl48cnH2JALIm0WxmHjbR81izloH9S7BtoOCRQ/x5RKuc7lQH34TdJ
w7Y7kJ3t+Dzu4nKtFoWdHgF/UW88BKHEkca8TvHvwzT3q/cNbI5EKnTdafXPOYbMA3DptShoO1cG
kJZIMUrLEr/k6Jz2GF+gAypWfKiGQUvc3xcAYEobKiRCGIYRPFfx6UHCGlC6qIM01BZq8fZVNTaQ
A/3iJC3x5OMAVAPFRVE/qLIbOgWIfBPyJG0x6/phovyb66/3XQlHJFZ5nU6mJer3XaKWdum2kTT9
PLjxKKBZ7MX18Bm5MOr2tuJtJIP4piy3AuSg+zHUgZLyPyosGF7B/MAO2R+tT1g/KI/bcJUkf2Ga
pthlA/2HgATlx4I69yF8XxTYc/9OWk3aY9TSuPKHxWUIuZ9wwtFPvlQsqTvT6RuHAh36Sn93wR3l
7l8m7UjaOTRLJWONxliupn4w0t8vlZtPqnz5GsNpersLHD/MBx+0dg14mTYAq7Plm9CcxmzOnqMC
V8VR9eRar3HoKWtwPgtww17EsqbPJfzdMMZ7+9rELAFNGu2DaFk0kEG3WT/ArNXhhkRH2NZurota
lz4Vi+MTt4IEjYZFUmfE+ArFZ5LUlNl5auFt142/BtNouqJEfYnhuioDc3rnLNgoid7wJOafA0Ax
iCPbzMjpdrZr9sgZzBFE7ARc3wcLBHDVfCrbefAE8fIUk08CC1ogR0X1wzn8Cj+fwt0o8v9rkfDU
Tj9NHkzanL8nz/l9njZRNhxpEkEvGcsfCM9038dEJy+x3j1s2qjnCYsoYruk5zL63q2fgVV5jeMG
dZ5GYvs4nN2cd1PrBRPbb+cEdeVhir/auSlEuf6ruVac1NISEbsIG42uN7J0x3JAqp4C4tC8Viya
SPyh1nu+Zxvns8tAs/4nlPGdTdGP7BX5WMTwh1UUJt1jSREU+VrsLzWjfiDEeHA+kQTnhb3/Q2jP
rurTdPp8RrL4wQU6LgWBE3JIfCJmL7XoB8vuyay3q1zUfspDRdXZ+NXszp/Dp10+OnxiB2jRh6Tu
Bztelx11Bsu11jRQZDn1VfEANbJlEPv2jTtwdcObbCDOtk4e761lusgD7EIHGGikTa934GUxC3t/
gjHWViAcyIcfP8MwV2saGD5yjMQeKo+M0VY7NWo5jqF95ffL8Hnhsh0c0fTXWoex1ZKut4pET6iv
l06gadSfecFLGlQRgj1Hr9GuhZCbsZAxP31E3XyaMgxAMsd1p/PfoioYiaqMjFAe6hq0H27RqTm1
BMpwYVyjVWtYLrFaAt8b5H530dZj/Pusoqv+uROXxyqn/NgbcAPgJHneCUKF54eRO7vuPSRkIRyq
3ral0PaWmbzhFZsprd+0N07jUQP/OuoALZixkT42l/xBswzbZ1JvJLGTIMnZV2+hgsLFXP3onLWq
nR90bFjFQZX7PaJLzndCkcFvp4d9N/5z1oc8RuyQYN+AQmY3HYP9G5SnrU/5Fh1bNOdvDv/duA7l
GjcB4rRvZmVrX60h7GnPfea57EmLXv7+odtbQhbotYsPbDeiRC8VNOJFl3RLnlM3T3tV6EXRGwCX
9LzKJRnx7Xd9ecUSguevwYIpnwg2cBGLG3SDeFt2aNgi/Tu4jMwFuaE3hxy8XG+LSE5UtNIAWry2
PZ/DMfjSV9mco0WEYhPDJYQ4KH5KCFOdINGgaThslV6HZC6fae/pYhiwKgbWjc0h3qEl7imWMqem
cqBSk7+jVsSs0c02GmSD0xLCvfT3JvGjb2k/u9PibxNfZK1ivBprNWoFXp9vdpsNtpEhbO6YQElx
5E0ZFAmkCdMU/Yud6lz/KLUC/ioaRxOMbjDaXfLzOFS4ebqCDCZX0ccT5TUy+nhJrMKCKqDm5YiG
0wBHkNfoPOjg8dnceUgRPpPvmCB+LglIaNzGM+hV+eTYO0Ylddrdr8hDpXZK2kDNXuijoVHNdeJr
oHY7VqTcdf/sGBsxW8+Ne4GdouXxEkpzbgN8ZRnQpu6g3pDD2QrYxDdaKwLN8uAmJVIS1gAZqMDm
kxpTJM/HLIht/nJNNY9j8ts78nX+Vqs2J437wrYWOqP7j6dfBBxUq/uD1kxvn19UnioN1bd5AHmt
cjJMm3sPpCuVoJHbajCqFVjHkQVQWF5H1bJhvOT9QAzBU8S4VTdq4XqI8oRn3FqztZpzNMQ8Q+cF
vO5XPEhveP4dzxKn5+PUypKbpeIrPB65K8IZddkNogE8tjmmWZ4DTFspHTOOEGuaz/4dkHPJV+b6
eC8Oplz+YVoolHeYPYN8L2XFGQVKm+ZOP0ZSKcxZbpuyLqAd0xhQ3Hew026YHRSBE9ADrNgFCfI5
JOGlxBW+EA+GCkjLdnxV0VQ/aduoCjS3LZp0aD6CClixh8kRrdEBCFNHsm2kLqZOP/fhRMoQEVYV
aJ31OUEOem7Zl0fKg3Nryabn3LqZCr/1NAQ+Ku1hxKKEfD+pSfSphY2yBxujOnZjUTWZ9wCroDqE
mmNk5gxedHPU7QxNBlyIuBbqx2lsQcf+rpiAV2OC053m98nCWH1J7JnD40aN1NdylQW1xicNK3vm
Zumsc5Jky6laFFy3/cKSdIthknDHMIG87FFfJ1WzeF1SdQjixAKGlla6b6pm9HJd8c64puqIkgVZ
uWmF1LIE2JhGUX+WVBYllw2ayXmmEA97CmOFyJ9xZq0ol/2g3EvXrsGXHnJm6aroHBarxiQ48nJy
IiQzXasve2iqDc6JFLYM/gNw10IdIOBUnPvjElTcq0WgCrmHPpvJHHikdT3uUEKjVbAnGEyj+URD
2QgD8T91uiietUYWI3eZ/Kr3g7UhQCh41vApkWL/uEnB7JL3ndErYMmvNRDYI2Au1Tcp3U5ruX+P
GcM8Efbp0s9t42RBcPLtIvfPwx9tk23ehjm+1pGeFsKmnzxgvsAVJLUiVbcHejHAt9UIpONaepUG
zcWoCJGoO26S9ZorxdO1EvIFy5qca4u5z19PQOovQx08bAvyIpFJI8CF7WGRJK4T2Kz4Z19lDQe3
kipgjyaDXkEM9dYdVDwZpEn0ufxcgJpK9FFZfpXFIS76w50YjQ4Zd0qDLIhlhEGqwGm/VUDI6fpD
i6+iWW7N+47UoZk7rZldMeWg+lWJJDVeVX0HugmuFp2xiJi3qb8nWXBq2Pks4apkhMJQnLv/oqJh
u/+TRbgzSdGT8FHSjuCWLcjfcqUVwDg7ghRpIsz0X3//RJyBCuxlEI0rT1y98KkzEtxsR3mC0Urn
SPH0Pnu3fWqVzTslCCJ+U0EHJzpu5pX/vSZ4PzIEWvIF8oQO7tmPG+JqZLPfnZBvJGT2PG4ZLh1I
5rs92VLU57sUN00AAHzlh5w5Oscg2AN4HVhukq9Rk8jbpWcRDbIHCjM6UX/7wx+tnUZhxGo3syev
hxO2+T5Exu+AUk+5o0TyK3jT33aTGyHe/7pnw6NKsiEEyhJreqZ+Ad/u9ekYmaJXM0mxEbJM0pZX
Blgn4RUFHZoDZNODeDFwOFaHdcB+pVyXSOPa1UZ+/v8w+LPj+oknLZrJU06Cc5hofRj9nwcONMsg
IZLSeVsnV5FMeWAbt2FFoBfMD0QWWkKJQSYuuIzLiyyyLYLC1kLWUxK6kzhyYmC+hYne7ulCnvV6
xZinOnPZuJtZ39GjF3HE5+lsvPWbG76/6L9l1wrAWGaRLPU3Or6qmZT5eOgtlGeB0Ab6Wrs2cVES
o7aGARm8Opq0/j8jpJlMPgwFrYLwsiDl5qfYMyIizVIrlirfJoU2Wz7sb4jwmvCVh7gGIJAjT+AG
01Ww25GyWzjhls39oYOTmmrm8tpZaWHMxFNwO2LDcqxrqbR0Xzao0Wv9q2XmENuLcgJ96YwIfwd3
rSak0+vXk3ztz49kOMfy8Q5+DW+iOsWgvGAKmFJvoggAhhjP8SMvclWNBSrg1v3A9dOeWZwURkVx
zfT/hdfQtyctENdxAHisx+JeL2wZHEzQaM+gMKzka6Ww8UkODrfQxHUkBrhDDLoNJx3SmYxR/DBy
lFMUEQtpdG0DsPL0MBwJG/qJn2pNu7cgoVKWYAoxIJGX348GaDpeX1dNXHnFIvvKhrtUuekrZ6m6
H11K90DeuwWFNl5GBMTgNuVbHHQtlVF1upksoVeaSJtnZRp4aeAn2s/jmBkTiYEMxZATKhS8H2NK
JHb1qg0R0r/SikhZdI2pGIEE1t64S6lp8ueIijOmM6ZOs2fFY3JloG6HQ26K5JvJFekzhKP7EJWm
nGQopbBRd+YkCkwFRRDl0lkoasFIsIKgNSPXBKCTZ6AMNk0OSAC8STA1QgvXwZX5/ZTFP/bvzbcX
QuNZYBAeQYJq+A9KjydZuwTdqDZyEk9LoeQqyj8QFrGRM3BGZfOhz7lMhHX4PDGzcxKuCXIOou/x
7ynKg1e8m6NruSGbaMNj6FfDuZlmV3tQY0UMcuQRAcANcSC4eDFHVjOkwX3+UgthWGTzONONnhpc
mtO6RvH6FM3q+n4cXQgSz8vSzddIK+Ij2eY4rmVJi/q2tKktcT/zDjEVBiuFygaHl81CRNJsyUWr
Lp7rS635bspehhk2lHIazH6YKrRxof6Q2dyI/jg+CH2OqZTOwg83S2kCOs0geiwqImPQkULBSapt
bnipJt3XG60gwqqH+ZJnUjy3I11FQTVkwbD4baVnL4mZ4/rW1+kpC0akhDAEDMqG9y3OIhBcm7rN
isH6AtOnGB4Fy4znfrW3QXbDKnSeFuT7ir5iZmUrq3LtrpuK53C45K4Dv7HuVN3HD7Hjvworq/t9
3Z1fRsFpJ5G8IWbXy1YEeLrCI5mSwzYlzxE7SqXebBq1RVTBiRRrxFtXts1HlS/45f7dOs3eBhgP
foVS93dwlHEqQgiT54acezd0JWDnKj37GmQLyybAmcFF5rKxeB0I/Hp8wMW9ZkmVw3wh8SextsZA
/kWX3u9/V5h3cse+wYIaPO+uFHEm4atEQcV3bgZS70CdPmN/73hKQEmLHbV2v8dTNJ61eyrRX9sg
17xvZDdj3xUZ+9itaRv5Yiwsr4NgqMMaYgZ8CiFO6D4IxaJu+LJuOhfkWNCcecyuSzCPzorPpeTY
IRi9tFtgD2ms47grUtEgbv3ljSMC3AdUY2rdfyEygJ4s20xK0KyyC96I+l7YHMxciNklHH1tBgX3
Ke+pnemcRT6/P/UL042yb/fbFBR3pE+lhrlPSnVM3fy6JaU6Yg8TRiMDOxCs1RGncg880KkiA+DF
oM48XFYcIMWaiQAdHNpyA43WEZS8XzeMF0z+iTsLi8BtuoHA1dtaNvbrEP9eFEQNA9JxgKqdAIAv
LVkz4EyWjx430XuoSlTBxXPOEDcg+f7DwqtfVmmwaGlBp9L+2k+05ABBER0OvnYMH4SzAB+HPwRy
B1o0aA5rimpUsLUpX2Ydx6FLHCjXN7Plr1IKul/uWT/4/JSObHA5s99vxC/nmi0cE3zczBmH+HYB
kPQN87yGkC/GbXHctfptH8qaIGC3lN1Ei1ff8fGTG43qSeUmxHSbF2bnrO7c/A+lnTcRYjXoYNzq
q9hdfljS16h2IulpLceh9taz6U7Pk8a7bMDeuO1JzhkU/CS8U0JX73XnxO2QftXo/tx67XMNMK5l
skGZGApAZ53i+51szbOZAuiw1dZe1G7dX4xiMI1L3FwtO/V99yigSGPE4aDWIzQbMgseCn4kjbn5
Wgj+QqJMiL0TYTap9rMt7milJOwYumZi9cVnQIM997GSHsVzELjYpK+8m9hipMJRsjanloj6yvrm
nMnRPdJ3ZSrueg02lW/mer2zZnR0YSZuQTlY/l5AzifItmWIOfeZNE9kDKFSXeWMYjEejqWyiMSy
l4cjc1y1cuDW+1baifNCNOfocFaXTlXqMFvosrw0yKuHQRa0DxbHlBjznUbNnf1cTd3N6KjA9fxn
dX1qqDIh8i+YiuWBTJuBx82QgB/ziIhiz9I0RBPsPqFT61yz0T+eBV0s4Lxoj/Ep+PgNfhkvk9+2
jMzAti+d/I2adGQgyrWddwUmkjgHrwezAvPY5e7DOvlqClvh1o9BWqnp2InI1io0Icn6mTJGvLXx
3AwBKqOiGUlegfnyypiF4cTXomYcgTs0JTH2pSq1TNwTrqD5/AwbRvSxt7RXTIqPs0H+0ln4bukw
emHWhqXYmx2lLaxD/LV/6cA02ZdjAefYorz4AHKB89qy23ams6owxdu7XWFX5ayQ6HdpX0vCbBEt
iZ0vVQxzYxDwTfvnfIbiI0AYOIhiNgrgUwXm7jQFUv5PQhn9wZhehrYFe9LdKh54zndZl/DPVs7c
0Rm5D9P33/ekyyuFSe/MxWD5OjDYE3MHnXrtMgo8CHywp1HsDz++Eb7M4k7Bzr5DPtdOzZmynCTp
oMvM+qKX3BgoGGMI7teldXUEoS7Zh32OolV+mcAo/9KAyxGnw+FkQefK4h8jOZVYshRazirVslwy
dMC0J1D9ZZ2h1JLBFsTRa7A8qk/6CwlYZqOmPHzFepi+H7/Qu/oCzCY3tO1vDKLIiiOyTGTlWip4
Y+pcWSqsE97Dch7miercZJmSj9TtjZLEGXrfsIGT62SixBgDuORYeMosqI3U36K3UkO+k+XzSIJV
rrvoRiKSlDaaRfPUOMwdo8mkohNqeQCzRwpABtl8TFobcsBMP6zDqdeZK9pmF8aqtVL8HihJB2vO
rz8ryweE9liSwgXboXolFN2eFkblP1WcTy2mQPmAryxpPc4NYj35KeyrduGLdszEZaWU2YmZK22j
lPQXuQz8d9kyLmWYdcmRG+yPzVbjyAsU+xqB5/Oa/RI8Tv4E6hQFj20RcN7e0DMZhOeOwmoJEWHS
SpxM/3V/1qkOvbv0VGqV6t3arUmBtoBL7WgPFLBjg72w6eFOUa+UdHDwkYJvPP6Ion/oOyUGZjIk
6XqcBuTJtZ5t1QrKtQ0figy4mxp2XOdzs8yITUYE++IIifFa9FU+JVoBOp3DqTy3ZLnNSIcrcGTv
GmZCsPxuNSd4lk5IuS+AkYP4XPGiAFIlge9WsB3avPCeGICtAHIG01nF/S9HgV+cN3pPxBnd12o1
eWT1cHfrKoudZEjYqQjY7j1589yrx1dU7dam6A88Hi98SpiKmbMHQcfwEv23zwl9Da5ADP775O9L
LboISffXsvrgp9RHPg5dXrF26n9tevr7/lLyggOm5FDN2iSGCOCTkS1tzw4eaZxya2flkuwh5F2f
UPkU/FwbcF4deUtnLtb0PGpqq17XPkb2RCb+YKrFqZ8T/tipivqxvgvg0L87RMsjXr+ZXtJc40UW
pUUsdXgDsxz+uGzPhYyMLOO6xnrlJKUfQLMJKK2d8QxML0mHCQz34OquKR43yXVLIr8xCt2ddSjg
hG9ZH+lj9ucyeP8cXxqFwIkEMUIcKji+dwYFCEO4G9ERHty4UYMC9yK60EexgHNUqtjAIa2jHM44
G675NxJaHdUQo6F3JJqrivvJiCaQyvbxRpI9/PzEJi/FDlO16fmzTa81gXDmcQySqVOlQ9p2gO9v
OB9igrGZN/P+hlIypNXfOR5cVMbFC4x2RENutLLXKerzhe3OxPdvR1evbdAWuLv8zqxSgE3B55UE
KxAKO3pJwpBBouhonW9eMzpoRRkJZBtAo5MSMeO7Ec/sNWHZKSeowE5uVyWr6qqpbbIFF3NCHKL0
I7PrE3vRRlariD52OtN+XcyaCbSDvxMaqrG6+KKzYLuAQ7SoSUx7Ll2WF6b4Yqsl5lA1RPBj65jU
WHtTMabcnpmaZoBzNKr5VAA2OBom7RjCdj7dfCVOJwr2EW6gQZOiIRlhgV/7J70U2RNU2IIRrmSV
+GxIAJpMwyBvO1I+e+jILWfLh8qeM6lYG/itKPU1ctkRmaGvmOmSXqWODZDoURsl9uZ+xEKDsqVM
L8LqzK/+yBtpw1fnTYwBm3uWFvLFIO+YiXmUviMX65s8E7fJeF2s9h1X3hIoXfCsPrSQl/4a7Edw
Hb93gd1TNYOt14bizO2lwa6hS9RChsEbfn/njgnbZI7mSm6bJ+Qtkqnvd7m/c6iYBmSNpWUrK8e8
X21uxBFTQ6+HwXtY57drm1q+Qq/MIZ6aw03YPfyctMLO11Xt+g0EwU8ldXzfcBaGhVDuJZ3vQWS8
l5BieGMJc00nEG2nWxyZwSGTB/8qNL6wsBOQQVpXAYiGyzUBvja+4CNwwtzZdVkNeEH36qTwBHtz
OLUfS6llE1oWjFmd0cCdKuhOTLYGarwMoGgbnxW0U0vFO3mkv7WvGyu/W2+IolV1KtlFFftadrqy
2viVKRcSot/izucaTeTiw1bNC3dmltGh9amGzL3qE2A3nvDkyLFc0afFulwU6u0f8W5nFNsVjgGM
ZvMlX39t3Sjg0trvn6dTWZ0w02rZT8OzsjLAmrYXARQDSNrbMMr1r0vAiLaOgoUKcqrXgcThmY8F
4xdUmAZJnBxaKXuZCtyS70nHsiX6huVpLoYVfnZQp6Bkaut+P2Wzm3TMgRp3M9rWjDsNvXGgXpFH
U8Ad/654vLbQPKquZbWwCTU3m5xUWHBsRYf0wEj1M9nYpD2DuiyoWueYvF1eeTpW0eG/YoqyY+Tv
d7JTNgnocR1hO2B2qObc1H86ae+5wODPgo/MoctBwmOGqkUdvmLy3XGYnrpnik0L8e1BH8dDmJUH
LASDDP5WpK3cJx8GDju/SlEbprNFVjud4WjN/3Lk/JrU+R1oFNCzqlaCyPZW1VleYnuwvepxGmxA
X5joctdjSfO9TP9vX1fZ3KBcuQ+WWw514uU3W13Vdmj7k7ACiw81K+//GdBKsqLzQO9y313OYbyv
O5PYFoyryKUiLf7CRl5eQqwsMS7Qa7S2G5AM447b8xLYKaLPSujcsGtj3UeRHyUdptC2ez6eMzfH
a/oeE6wOc2c7w7y+kc2QSz2cGQKICqwdj6RrAtR4csdFhrLH1O5YNZ+liJW8OtZEikO+nVXn2OkO
yPn81/Ybd7FFLZAAnaKVCWLe0CtVjZfk3zSkBeQQybwiBQSfWbG7dFRe2f13hoeFjzflszgVEKss
z4ms3ssx3c4RIcP9Sk7iKaciypGiLr8fGQeiMfXt8qyHWvxXLoLSkJ5FhguXxzqOg94+srOOxeDg
q0seoX25/l2FfvtthmhxImp4uPUCFmebaxnTgVBSNkUxOex4mIeKbuV1DPRI7/R4PNmn4vkO6NG/
WgueTKt5/S5NuIAHop9zqK7NbZD7SdUQ4foGxDQfvJpJUeCI3Aa2Te7lofha6orWO6S1CupI1ftQ
q2ibM7PIS69dQshbc9crWZXAbreQzvtuSTDQHvMoM6AxtYANAiG9VehAMmiecZgQE9b5kQF6Zm8W
36bnSoKeEVYtx7s25SmvXJQ8B1vRlHmNaipfTnIHxMUTFpmihPG0Jzo1ge9CKESmHurYV/nzhobs
3wJqMomH/iaHOK5o4YjgPFQnvIcbP0d1Dg9eh0NTjRDRzqdoZ6FAnsl/5ao3+TAG7uzGdc8avx4O
PQUdH3SBDjH/XNTc6VlJeDkcHObpys9350y0yALRE44A7ruo6O3pWYNAlzO3x9rniRl6d0UVq9xo
glgJVynmobYQiqjZdFrNujZEYwv007+YOeoOlrkn666qHyYaQjPH5Rh7IGzxBx7UcQEMqYDLKj0R
FqcYZ6c9jFQJL5MYOruY907A+IyY0wiVBNNT0IityrtNd5YvCeiFxU2PmVksmX/fz8/727jU0hgm
m6zuDdHolEG2uFWZVebs2lQ203sSDZIyI4YyNAVl4U2ReK+kAcqwxKPspqmqvHj7N8JXRhSIZVA7
W072AVzjY0aFBfo5PPxbJMJHpyJBi6Pr5autzCGug6nHgeGCe6Suj4/gBUipRyTMN9iAiFYvRkEb
xVREt0/wTUPKo1DG7R/tU6WH9FlKyMJoAKvnKWOq1aib2j+l9VzYDSqgphZRKuwdK/Eqvj2P4ydg
SNiP5kAz607UGkr0HDvBRC1A6rk5uEF4xZa+75F7mzjmyEcNuHmgAf1KiD/YpCOpjKzJOCKx+hhI
J196yEV1z4xpL+Cy8JvZ8A6KRuK5WNKxW0jrjW1hPS2Djm5aIDGeumXWzrR+9lq9g3uLtCf96X1O
k0fBqH1LBL/ynQ8Mk4BcmaD27wVP331ofUv53MdpCg7IpMY+twW1P11Hh+5COGmWa1NYGylh9rHB
2OTb17fGyTXxqRuaI4poeKyXAexO3vi50VDpsX5JKIyRxCehIkMQSYnNd536gRhO1gFNmLDEX9Q7
qvkLGRmf7DF0ucwfm1c4cf6tKWIX9zPOv/1gPCFa0RIfB74r9BgpcQ5ks9ch4yueSHDOzSi0/FLd
Qna6ct4CRhKTzmiA9vPcU+adGC6AULCYO7LiJ/0KasI7MULUoa3Y7G50oA0Ic+9U4uTd78TMLR3g
DLQTIb19t+S+hnyEhWXTJON1v4dPWklAY7GuBoj5U+zH/T8wvsFGjqZ2DvK4DPG/vmWa4VPwl/oh
Eg90JvcqMC/DiQFhMHtyinxMZqKRC3goFyI6zFIijUzfhBOlDNqdyoqYjbya9fEf1H9Fy3Wvd39L
1+si8M5n8PdVDdEGUZ/FJhET8wNqER3KGvIEhQjtKCw8Tp7Ia10eN68ueiIkxUHAGQ9MU6GLcvW+
BXzLgvtJ/XQ5ZyRHhn256ywEj1bYjDMU54Rw6L2HevmWDyT+OwtHxfMGoPkFDy9PThmqeMuaoDw1
A08llG8cd1/nsMZlLUMTDpVI1DpvJG2KZ3rmfWeQjGo8zVCke7rpEUzEFcX7GKvNa65ocs3hlACC
gHuk351asatyLG7fFnTRRQEq7Gu56dP9VyOVM2tRj+IdmYF3SGqXOBoIRDe2s1hy1ySl0rXnWMR/
TQkOPc8SVfI9aoS1PNrHBjEn1YB1/dmBj764t5S3OIlEE6d7vCFQNYrbJ5jH/cmzgiPHrMfoGarK
L0+daHOuT5I6KPpQaLRJzwlaqoED2EbruKpcSRWqF+HslQ1hU/qyZDz7OPshVTFQyh/RG7OshEFp
hPlBMXpjMxunU8nYD0XZddD+RuNHrnqiIuo6nFHiYO0aQgafabQ6v+m01LA8JpRJCWXg2oiilgmX
sgme2lgZGgjuG2vVJPZ8TH7FEqNi3BZW7qt/bCNkwGSiDYhPQVXwOde6QP1nOnX0rbsGLhjids6I
OtTcWl5uPUp8CeQ3dNcdTm9VNloi3Nrv7/kGwL6uU9h1Uy0I6RP5QIwRr3qYU6p4TKLDkuwzpIAX
RC9Wm6nCV6D645fs80Bz+qMVUpfZihI4+ovzSOsC1ZQt1iHInn5Fcan/ahmebo82wjpLbuqwZNw0
+/CRBhCCDzEtSAUYVIHBCOOqF/hFEum+M+RQOVbX3Izdh7sOgiYVb9Nela4Fe2IgUXawToc9pC9D
aanf9TD29lDIRDHHODOAWWlpebbY/aG1zkvB50BZYPEs03UssWsGy1YrlgcHaXMWLb8+pvSozCub
hoTcvC7BD6HMiNWWgrwZegwGZ+KX09+ROZw+Z8/sA07NRISSRafas6kjDK+BwY9ipKaroT2QIaxn
bWdbz0pG2S7zjuGK0eV9TOzlgWyQjV3hSlNVsQbJjf7+hs8SKZ8evT+w/0dOiP+ZUZo1o9RmSPB4
u/VdmXXhTLLzxXva+zkHPYizs0jseTydgyY1hw6EvtuhqCDu+YO6x47Uskb7aTsWUhHe5BUD28XY
Uy790+CVRhNZuJTvhjeX0eM0ii2MHVG86xrFXkl2UhZJc7Z5Q//mJ1FCNVn+4UbTiBspqPu4UPZv
sq1n5w8e9AiImskQP6HZzyCHgvNgdxSvkm1ENaeCMEFs5VPIQCWZzz0+O1hXLdUwRhhprwz/lQwc
7eanfZPPldrPzxZMlFHUk18hmz2tZGZDXzl5lvL30C1F3bfK8iQtaVkyhdgucjv0thGu7ezTxJg7
izDPliGpqXtObP/sM7rSPbbU1NeVDN/sEJD4DM4iN6oAtEHpp2A4bfN9tu6WzpO0PuB6Nopi0aHC
3eUZvu13HDehzNgUjTZ5dmh37fcB/JOFZ0dyxN4Ie6gTubG7wNUyuQ4H0mGfK/JKZV0AV/tGK0KQ
3hj/CEWRWgS03Vhy82+Z4Zj3ZlmdZ/hpDpyZc2VBF3fGwgJB68F7b+BcBhlnRjI2IjExLRawtvma
sYUSSkiw374Ww3mVTYleTA1nCEfbE7SU58u1vqgJxdlTTIvRM98GyLVGMZ7+qaN0CSJn/T1lxTqN
3V46DdZeiSqs+9TdLltvzgeXXQv6QzCaUF5MzGlSnF2oZzXsCe5ROBwRV5niWWHHntwvz8LRwSAc
9cD7PG77zV+suFK6oT16+8PGVwq5c8tWmnTcOt+pXv6VZnB995ZZoMEpQItwXMx/rBjYPZv6+9HJ
isRPy78iNhSznQXCVRDrr8lT4bEVHAkTzOhkT1IGZoX6sR8l1fSwq065nadaGU3YqF6OO0bOSfNT
OEPSJZ4cyKZVeKuFgLW1LcYuMeZ1rfPEhVIS5vVpwyk0YBa4/7dnIBvbXX783MEakfDoBhMFGXrY
4SpkEB6qGI5tmnT3aNMfAcJzGZ77jw7iSgb9m/AgYdtg/uVAG89M7oYNwbcB299LDuyR+Go5n6UN
4lpX6qirvgtaw4KA5RrCX5nfhXg2DZjDtp50P2f4UwBBznhH61YuSbU98GymafVxamksxX5sNOy6
VR3X6y/smP5f9SDY91+bvrbnRECqYscXZudZgiGyk8QYzvLY3zt0G3z4mtWHYuqfl1eT3oOTjatb
70cM95nsPi+r6E0XhMgu3YYiTWji5K1NE+G8uFNu7Z4C1NnBWXM9mgFpwIAxyEUv7O3H49uiiq2j
ukB5Yq2YRnw7PvJ+IwzB6vAwYzFm/lzUl90nZDL5F5bMejOLGVQmGxg/rhrM4aAGpFb+L6vULRGb
qQG8KHuurSwWPloAahwE8Q85OEmixptWJXG1+zmaGtGsm4sQsT/eU8O0bKjewYWicpcGfzt/YVUs
Y9Vnj2YErO08o3/xgZ3TVAbKTo2zSsEncgV/Vd93TXUApMuglqlNWImXX7NmCoXknOkzRuDAacbJ
L/p55hNI5tlhRQch1asiWNxfAALt3EbTkf4186yrUpmOW2h/o1fEtDKLfrn5IT+Cf+oEsBKOgEjL
ZiZUbbWoEr1Pe5NdOvC8wDTVL/SS2+y8B63oAnxihnjDmsSRqhllcGwkzsR61peFAbyhMJOUbUM3
7P0m4Vu+zeQlWIMKkhVB2l2kvv9AhXOKNSt+KwIhYe/R22lSeIVfdBnRDPaS33lLk2LM2Vu3CyCG
9TWDVQH4NK9nR8V3KPUlHqwWGMFpfuq+34onqs35UQ/sWD6owotFNYLqT03GvRaSSnD83vluDCe/
yAQbER7gotcEbEKLZ2D6Kyo/wSCJBLcgsSoaKvCbAV4cdSfzs8jAWOXBExUKz4jeNLH1p7vOqgXV
t0YH0hnpdxuLAL8tAOFLwZSVgzKWbmGZHTYvO9NgoR+q+9wj0uHOy7X0P31uJfkbgensnsVMQEo1
edcCF8KyAIlOviOTI4OI/VNjL6T9yc189KYTWj0pWJlP6K6tjDxLUUZTYSveE44W+Dw4LDFDGJiE
CcoU1jDspDbvK1s+LpvaZJgEHMjJgg8jfengoEhwsqqdXN9GzGi5jvNseUIMOU3BsfYBHf8AkWZl
Vovm2go8nW5GAG+HJXhMFyZsR6Xr4oiU8afxQYTK0YEVmSIOynxrdw9d40d483t64t8u0BKq18xF
oIGdu5ln24f52nhlnnyApvBP8Bptj2o5qtO/mDrXcwhTLq6zrNBp+LKG9zeEqYJ6NEDA8GJfVoDi
s/iNfNiAvpGALi8HSLYbs9bPij82a5SRoP6ekxZl5J5IfbasKccXO2/uFJnWXoQ/D4izblQxCBD7
916yavFlgx10dn/SQ4OWMqc6hvukZsIUL1N4V+DPiTPZ0f2jCRjF0jxZKuoooqfbtBq/eKiFwZwd
6QHoukMd/4DN9HG2IHMKp2kiWfhOu6guqWMRypka6xJgrOdYRxPvR6M+IFIu0ONdbDkQ5rXYhbGK
wVXx1r9dh2MaO81ID/ffNJb5L275cm1iICsc7kJi1/YPsBkvv+2/65enz5w5hI14B7MPJRYFSDul
NSW5cc4BZ0CqiSGKpM5Z7QaVBqrR8dnuD7DrmeP96gMPyXt4N5ylg6+KOvHgcGxESDuxtawImLJJ
D64XY35GNAvT45v4ZvXIxSdHIs0TtnHrv+j1nRsOyvI+SSLYebIhsheg2/W6EyfNbFOf1JcKWD80
rWCFnB2a3rhKugWi49HcFUwsIK2EPAl+8T1wVmZPQqGeF6iWjfS6lvBX/gV/ApXxogKD5ya4fdKh
8bqyLV4e2xtckectnIUtPjKqXv/GeQcpbjLxxYSwMd8os4gR39bYvvh/IE6aoe10wlzHLGeCqMnm
cM0V1NBI+f+p0EriTONMIpf2LO6MynudeYFfWpIL88LQVY/WTfi0Q+bScZVGauhpLfukWmzA0MPg
8qK8RIHRSFTN61QFSXzfi8C53nhHVaOW3p+GdsbO0g7U558h7rqGJWO2xKMD9LbfGSMom1hd3iC/
qCAEL4Km0FqaxU5NwlH/6njFaIYjjRxF3yLZTQAxxPvtv2VcFQ7kOkHUiWdDmYlElm59iWTd/2tn
OHb7kaccYNT848XqGznRjH7iW3VzuDd7TOHjoGgWvraCWIG4fG77peQu/41mp9BxmZlSEZwpbigL
IkttXkO2t0bCFgklARe6Y93XdvXCRzmoY+nKFMWq+SeAtvqxvoYWoNV3W9X34ppcqUQKNzycD8dI
ZhHKx481GKQv/PzCxFdDEonEd5z8h9/L3jcHVUNsmJARyR8H9ql2nLwTUL5RCRAiMYHLFg8CbqYI
1IREDsrr1evFZKZi6M2xgmxMzc6wtc17pDQE2QAhjQFpPszWCO3Q6HBd/WtlIspv7LZklr5Vtc0w
S2F37SgDCiElhqnvuFFQacq1nYjXwTbrf22qeN+15QIOAz/mqN3Iv/R1C4kUR1OHpoCKALVFrH7l
w+qv3SaGT4Pn5ajRBD+Nhtktr4g8S78PU2dkxIMC0dnSV5l6e27nGHeK/t6R9vKOMMAjw0uGGhlg
XX9ULTLgIu0dg07M/80o77iD+8fcCIHMlTtV4o29KJe/Ip+UC9kW1oHu2Oe8SSDxtOw9uhICzdc0
B9BERCdnbTornVdZ/UjtQtEDMr5wyVycPcjFmsPUE3u84OH7LcOIpYC9eZnGFKZNHAschwtIfWiS
CzQbX9lzE7x/I35uXh63F9vjWMZr7aDUl3AR8Gi3rT3Nm2r9wP2rS6SXT3Z3PPcTTJaotvhPapmb
3Tn3CGqj2eGYmX+ZoySS0hzQuMfXE2ybaoHhfYT2xF6ZvKCcZQ9McWf3eSojOEaFEFabz3g0jAxH
PX6TrJNWAq6+LvFmcID30DMLm1YJck36jlAU/v9VEaGWMmRETLTtcJuCopoeb8kQcjPuAY1glyIv
jYx5Ry/6D8WogXyZQrREkVDlLMj95u2+wnf0beRWy1mKJ7ReDHAmbf/rh7wGVS/T3dVxRTWut8sq
DirNQVn+KtGn7227r2ijuci8CUYTGTV9nHS8lc74CPX6ddflDaFHZPiEcdbR9npPvPjm+Z2a5y/U
Xu/qx1Z6wQUG8XHYMNtpS8GEpSjGyOEW212y2lLmddR6lgT9yi8g6SWNvLF5RS0+y6s7688bAEDe
w4mgwgHDYIBK47daOTVh4NrgoqOLB0thoafH7B1MjbB+7bvMTdo6l2VcDCEz5FaXpFl1CVbEcdPk
loRwnChIUExQzme9uVX/0qkvX+AX36pDYrOSE6Glw5R+FRqYxDmd9opPpWh6jVsy5lC6spM1COHp
VlPZJa0mJLz09lqgo1YBiStmSjDohowbPSROkjFy+FdFeF5FmzzozZSdb38QHn1OkAGOSITDfMvv
rWNEoXNdj9622ahTXbjFpa8m43IpXEDdBFyxzcNfnKqWVFq793GCTQRA9TveJr8q/MrFv4bSN7u0
YIb7/89btYatI+3gxqF6erYuy0uLTp0gpG09q4ksn7WnpCGZKZUQWPvnGtJ9t5a4o6S4YmE+hINx
x6vFExJF56Pt+b8y0TD9ezUOuD/xNaL2pkRc8Sj6aXsUvm9vSK3j9bGf9j/WbYpNrnhvVmoqZGsb
O1MByNnU79ng1YgwXrMNQGPuw4Mqt29ysKDSiBKX4pleLLLqi1KUqen+gqhzEj71Pgi8yoIuDBm0
RIIWMPRNby4EadO/ZMjeEIYQBxLZ8AR24Cv0phmdldA7hG/A7iM9B6gYXVKgsfTit0VwHTG3UIAy
69hHsy4diqY95u2gOTAjiygpVRCJKZ/tXizIRo6W5mTJMBrRRykY0hRzAajHjNIc3Wis6KWT3q2t
kHV9UplDJYa3CSsy31mgAglZUJ930MK6RynyO8gYXSsxHRllfkC1HSBfk/hdptPAwlnOlLmtRREL
GhqXCrJ8JJJVB074SjjoiaTpeVDtHNvnivqCsqmjUuBVQoMh4/aT0WVB3rbofCXb5OcKwm1xoDhT
BsKgAe0iTgNwYg3bbmO3tAU9PsJqAgUqHPY1oQG6cjU6r0dYRQaTFdwe8ysFTQMU4ar7eaD3KWuT
+BrnszBOe3mS8ZmjfM3vVyYvR0+6tuH+XHXg2wiX8OFP4qiPFHElhF3Q6p7YD9i1+OH3Ck09XjQ7
Nr11DH0sKJtvnQwwHGKkYvo/VABqa3tZkzwJwi7m9oYE43+PIXxYMp59QF4CV6nPTF2HYuCVV/7R
Gl6qosiOBHLdgfoUC5a15CH1Clwcoqtv8ljFILF2KTi5xb8z+B6r6nYbk/xJ3NK/j3PAEdILe5V/
ca/I8JdYFwoLASxiE21QWdtCvgAFCr/UHIFiYe2XpPnn1f4iSF1RFHamjyylpHhOuVIGlL+reuNt
jloAraGjJnN+LOKHzJm4x4wunhl8ikshf7Z5uORjo6yWYLFPzoXEcgX33WMM3wYvlGijpyhOEiIS
HvozuQ07qLrq9GKhu4nMRnvsok3pfHOr5cfkAQme3cDptwdfhgpWWbLsxsvIGIQ2ohrY5B/+q/CG
YMx68ZRRGqy/vGU3+06XhtcE23O/8cyGflbf366jF2byDYAyHnupPneVw6slQvY+wB2VhvS00mKQ
dmV5d3jwoahOHKHWzY/Y/672GnCNzh3+n0zj9XG8PExEgOVYYpzfGX5DgdDjPZvtzvfAO2hoeBjh
EwUwRjBv4syXW+8Wkz+l+K4EL1FANzHpxDqtfEjOMJV5CRtTwwMosLnlHq9nODHvZfD77Mjs6bcj
lNHcmTBqybGSandSCBgpKfj2xXlp6Nrij471XElkC1F1cOguxms1eTG0w7tWHarPZHEgC+vvHHbi
8/qd7fCBVSuTxL5ywM2uIn8aLuSBifaeTBsIYV8NTgED3Yjrcp3uZ414FKe8BXjVDGNBsovHePvJ
A2UlzmRSjdgEl8LQj3o295CA8qt36IXnUVkDRn+eId0BC6WCyhKxcLWT/q54+g0MxpcVa7Jc+bgu
P9AIaJMlijCgHz6KY2FC+J7ISubefXtgv9K10SXRCcll3L6zZZTurrXZ4No9q3dcBtgR22U7hCRL
lLLFP9Vw06iZKhuWr7khP5Cs6K5ryXEV3UUkXrJvPSHcKAReO5htPwmkUAdV0vvM0kyMvHRsQRGl
QEi+rurJb3qaRz97L+B3PPj4PPwYz4bU86V0kUbWCbHUxW1H6PpOGdNxRjIrQOD5ZW28ETQRjpq5
LJd7a0m3xhlrERjzRJkK/dCWo8/mcMtGN4b28Dh9o7rN8VOGhADZvhY7hQftjXYLyDmba343ZxdO
uKbGAqz94LdZU1zqcxiyxiLpWJLqfCHRdaTcqZEV2ORJrNDr1yMl1LonD/f0+oOUy14h2uyha5F2
a86I+UtZ+2qAKawx+R3xkq7MahyjR8INrPt2Av1EIy0DyPkB6yV/nPWPZ8OjWW6ApXvblrbg0onT
B1sKXRAldNzh5cOoa3hGEys+lHZaoaNyg9Zql3aHIMS6stmRrbawkxeZsjM0f58ErP5ZJF5gtVYf
Ke4ci9Nc/l0KsB4MqMkSo38T4nx3fZJglccqA7utleNmXYXJmxJqIrnpSHMF6ky8MfCJb7iRGnJR
zfP/HxLKSG79WbfSPQPTmjE7xh5wvgiXjnojPsSK75k9msbEfalPFDroh73x+sGcuO7ZLzlD1xz+
3XfNGfjTS2vb1X/xSuXalwRy8WG52SDno+PWsJR/X9t8lE7UXZ30FOJ+BSTvnlDTBYXMjsS0yb9h
vXBK2THGu4IqWTtRvbt86+/Hx7b9qGsNYUar8XhOVfHlfr7tyVuUzFeTq6g+ChpIVe2rS37Su7LZ
8OrE8zNcbgxCNts++VVLZSYSlBp49aHloqYjvpCKkF4uk9QXYZk8Lxw6jczFUK0Wb2xLoISrRMNz
G9Sueh/l2aDTX6cWm6RPe2GuOpsljXtHQSCh+zHKbdZ4KpRoLYD8OHYLVTv9rS9wZi/fcGzfIkKU
q44P4dpKHyUaww9vHPH7cfaf4AlBnyNeju2+WsUW+GlB+Kf1lWF57g+vPT1AfV7i3cq6pCyR2qyk
86V0VkCnZITszv/qKKbuWSrghBiJSvtAV3j9T2ipe3945XLxUnPqhcjyjeseKI11vQxJ6jn5CR7D
wn0Fgr7P/Vn4LhQZzsjPrIOGAZ0nRxT+KbODWpk78Op4N8UgUyPAHfNrw1KJcs5/ZWeNV5PSpYW9
IvxbmA0zD+4d1GUF3NlCk/x/0S2E3WVodKu/jL/UxOtjubsPRHiPLbKZxqfo3OByCca8frwQYwBE
h/yIi3tSK32ujJxpOv9YXsVS1rW/XvtOk+MDn3LLYb1EKh1xm6WS/yb9Oa/kSsLJTM36z4NqRbqH
UPa8P4YJ2ATPqK/bp4HZipzv4SJa0zX7U58d2sVOUCTDkeAXzxMvnb55V2u57h+pp1cSGRlIbPsF
uFE/ZKaEU0cqRY/3GGCGcINEC3SFN01MsiNHxNxNzEI3jZwUgFri/+R3/HhuEoi0NANuWqfcdC+M
Ind+uFOz+80wfyU3kDcVy4/S+TDt25JIxQqTDLdRYe0fw/XWvxK1e3uNl9Jkfyuj3yFpXX0HTI9r
rFTDq+v0sRRKlWTXo2rDZFOoA0hAua/C3ina7kI7OqwsPxuvie84u0TPF2w86emE3Py0CwRicJHV
8gAB+eO3Iy68sl62GmcCcmqW+QP6jxRNv95gsT0NV1KJ39TcDn1hkVNvMKRratkaDmrHa6RnzIPD
IA5wzd3/TcFlwEmvGufAS72Hf+CoFFEGnp8uytrjE5eNyK3pka6TlKCRbix4q1UfsJ7Ry7phSMrb
G+JDDiCE9SPK9xLrRYCbwuiMFZTu2dyP76syeF3xyKGIWcU0yO8n8kCMcXR1b3Zsra+EtSyI/9cx
h4878ssaD7fvNfCmmqFWX1FFMkoI9bQNlhdw+6QcxL+uQZlkqXpgYPy3kDCj6XfHz/Vi+SafpNxv
CE8WjqJUR+EeTOFSRSjjjuH3C6chpFjarCNDaz7IftBvjq2cuv+tIkuAb/15J6hnXDCDo1LXWe9L
7j2MPEMu4Lm6JmmOSjz4SzR8m6i+ohV7xVDVbAcgBbTJisPJ0BWjn3hWjhtfhZQTDcDw4jVKDdtc
m42bcjCj/8TN/VG2K4hMWJ0PWK5yxcRdQQVgPqybDyMszKAy3yfMG/H0DWSwBrSRBk7LhzykLoNR
vX9LkMwEuPdszystpAUwfErw23VPa7a4LMZq2xsKOqeFle+34fyNWK9dNQeDAd3BTVzBzRuMYnf8
mhEaSXYcfyb3NYSPEJTvv9xQdcs8OkzGm/NB5+KQdc2SDBHqf/SfzMUJE/Ho6/g0rD1PEmy5eVp2
obg6QrIauqDrin15ZJL5vaGlQpSC2yfJaaoeFOUOT0Z9qUPksVcVguffcnEU2HH0q4KB5c6qq1r4
XVuSQxi2g3JwS40LerZp2LwtkED24fxGim2xvLJkVeMjCSq6tLyXVbY609XUwLEOFV4HQSQe7zRx
djECXwIzm2OHNW5MY+Lrrfer/bHxZ7/eWZIC0C2l5kCqQc/L59RzIR1/8F6KthWFgPHXJhp8eCnu
5/GbqPsrJegXR+4dxPAm+QpKrqaaQuhTxalC6Kna6s7RTVOuU8IkRXRPutIGqif2ggWkGgCiOHZ+
0tzz+RAxuJniKS7nQaAJcKd6qoJbL1nioQGZKs9yhZ4W+YLK+PEeVq1ZS1hCj0jEAtU18TTMxGAz
Th5PNOqt5T1pp1k+k1q5+f2eeAtJ/T09+IDBYnFXNp9YckbrO98AWXbrQeSZIaVDPeuYEv2nqad3
9MyfLd2Fd8ZKSuYJSoSkLLsvYGoE05/h8IlTnv+DhhJVLAGYboX78/XulwjE0Qf9TTHGkK9rjsnw
J/B4My273r46eH7ZEdH5dG09gIcJ0iVvEKJdz+Xj5BMaQsXs2ZFcfBf7K96O305vJEfu9w8vwWPa
6dO+Ms/kDHWUCaf0mBItV5C9XHrYh6W+32PL00f9onZjOcV9Q1cDoIi6fneZlZJuEtTajMTfV8Qp
yyPKTaZI65LUSR7j8106XaBmgihq9P81hRA6uN3pJr6O6SHSngq109hdFVnCurR7ONCIsD3L2y0n
bXnBqbmCwKrcT0Hw/b3lX5c6/1kI87Y5yClEJQNtBLENO4vCPq08Et+1lDY+QnPOyfNc39DpPCny
K4DRXaoYVcdMSG01g2Ep52jGGSvmKLWlZwbRm+rw9VJPYyLVPFco/73KOnxd85PfZKQMoGnj3osR
yGeLNxJnMNTo0QUXifNRwqE8cTM7MCfwsXlV376KfWRjb7FDiDlUsqgBg2zu98X9LPxOrjjDzO9q
COBmXmiF3HmPOOlsb3IMjNPmuzWL2i5BBNMhEjZyRzJ5CZb/uPeGaimr7cxUIJT99ERe8h5E+XJO
V4wlqTHBboMWMsXSKDhUWKwxY5FI0Ib92a0OIZs3ccGt3AxZkVB4pK1uLlxujrAuol5H2KCZbw5b
rNvqErRtTC1L305YMuPPMyxkXIjtb7nmIdcx9wxo8GlwALUCLvI4SKhrDQaprTyeo4sViDD4wVJ2
6Nl8UXtEMEDKHqzNn9Dz62SfodfVF8UF9iddLkzpSZL96wlGJ8X6i5PozWjEfmi+dvaQ7AMhJfyZ
tFST8Rcg5hqSCILGzZ+HBmOWC9HkHH0WFAtBonGH67mD23rsosKoJGusBwJyJ/+1O6C0bIF15PLx
nd4lzcr98ZLI34PN4HMzzqYmVDIJOs4owHtotcUFE5ei2S6Rc5+4hMsEKkCvNsy0xKAWx8qX6wtZ
nr6XQEW4LnuQ9NAO8M+Pz/8MWJ3tbvRHzxzO9pXZ2xZRqEMd/qE88ZD/BfFq0v8EOXuYtVTOBgUv
EiBAYPZGbdDUgRFJuNZrtc0/Q1HDSq1Fg2AQjViclHqijIzn3VR1SP58mnL4072f/79TIsdOCQsd
FsD6PqnJU+fGX8xIIBWYI9QsuqTC+S/1PDwrI4z3rpAsHHJiTZlXE4muII1lDTcEuBK5yOf+UzEO
sFww5W3hw7rZGH5rTGaUkzDHLagJhPB4/SIpYaKlaASpA6J+fNTlsA29Zh1A/RcA04+LqKdbHbar
LVWAnMQZIRG4nk5xL0jF5iJrTfKYlaT3s0gg9wq7Fro6vxtz53Funn6J6C3gWhDOdOHLiLMkV/0S
SRPjiR53CKUtU9zIBn2krE7zwtReAaexbpZyHJ3ysfCe23Vk9shWNfJHJYmt7Dy8LyGiNwHoPJPX
LK/SPjnXhCNPe7W0VNcKXSEhuz+6nrD0h7/AGfMHHCVnaj6JE80rexC9ElLXuLQbqWwCzoB9FvWF
Tp65qnraDJc5YNxdtUa3yW1irNp6tDb2aETAhfGKjf4fALOUzTOS3XTkfhHpDpr1gZSovmt54Enl
q1QHx82pyKR+3yBTatZgdCkHRmaWTOPkyZlUaBIQFA19fI+0oJIxC6AoL+d9Gcfaq1zey870K5k4
rzXRiI66E2HRg8zE8Wcu5fBSj3qzKd0k1KCnQ9789bik6+AF110IJZYjcfEX5VBYIymFwDcb71f0
L1UFKyuc8Vui7gjpGl8a/r96uq/VrZJWb5jgaeXfy24qX6mmFGB7bQlmMVBl1MzO74dIf9c2AneI
+R7HKm1CMQURe5D23gSZRfTaiqbBSRfL+ezvUorvubLnXZCRxcOzxsclEEfffZW+xq15ooqOrDV7
yS4/pIQcj+03pIjDPxdkG+7HHXuctdNGKk8E7GEpeZYnCMJDmFcSgRdogtCpweAvwDQxiZgBygwt
zh0o5P2yDjoqZ3P2AsoqnJ8U0+5Hugp8q/I0RBKJx8iT5aHZTUBBBJkbPVC3fw+C66k5QI9hV7Nx
JCw5ueuOYWodgAcKBLUcACoV2i58MOz0IHnEIJqZAcL7TTMlzCMIiDijGLHa05BdTHOVdGY0n/xv
Prp4xnVHuIHgxvksD8bzOchHkLF67mlb9sJhGlsX2I+OdQFW8aboCwLebI+5E9Jgxdj3R9ycueGz
bWMW7X1W9mBASn5rkfu3gJw2vd6SonTOEBg90Y/rIkmrwbwPHvbmIfPgjDDIA111fdC1bBMLP3jj
2oFBspXtfwSHs6SofBZ5+ParY163HG96SJjdqD8/n1vmBeXYphFSFpMyMLp3wa5rJG+vQlugWOyR
iZan1+CdZ/Q005HMCMcekWnsr7sNer/7V7+fKCAS/QpDzvzx8hXUp/KRQ/NO6CwX/58rOn2Q/9/N
eIw5DmaMskqIyfHXFjyJyaeD8W4hB2Wbd9cLbNUKBEpXjfDaROCKX8KlBTiIxY7Y9uO3glV5rOBG
4y13rkLP31zm6hscypsnFWlwvRksUzBvbqbEeb7CMujIDF7PvlgKQd2S0pwJikdFWAdJFMiyG4rv
wZmzUR5U5N5mY08ewaxxf8AiFUbMeXjj/aZ/XtiIIlYsFZJlO7b9jMvDle/GJb8aggM9VD8WwdJ2
8sj4VSq9mJh2TDmqoik8M81L6P/Jb5mYHa1g7sKbCD1flZWlnOy0vCppPnzScvhQdaqsYoJGbdXq
IKWAlO7k5FxIDf2AU1TlCbDOTglPJYKiCtACnOYCkrjq7FjfJSKbQCD+Jfma3E9rO3YUDCQ0BXFG
heAphcIAl5IYLKqN57gqn7BROYUXHVhnyh/7+Gia7zw8xOztcJOpCLJCjE6qFNGKIAvv3Z+srIOi
oH8IHrrqKYqBaFm2mI4r0HhtDw+KAp914Jr8B0LgCPeYA2M5edC5wm9+fpJ6tDXZd7q37FX82L7a
zDVR35ZCvNbP/0mjWK4Ba//+YyNplRTmDnqZ97N+gOElJ1/EAPMwqVdxwLoMK66YQ8zc64u0AW/K
JXJ5xLMCDMLnGxErQQUf8Fe8PJKNmrcUkXOV3AtsXKnqv36d0VAdQEhNMZ6TRTcjkAG3Dmlog7F3
j0G4JMwPILip7Cl27+pTCj8NQTaMCmtkQb7jGSIpQH+xoZVn3odl9+sXLb2EafGQl2A3FMnNVwgd
Su5z+Pqofxim10EE+O/WQxWIMIzLD0l4uSI39Fv6RG3zReFCjvQga3BOG/1sVJUA21mlk2Ow8+4x
62vqorv4UNH0cmQNfHqAXWL9AS00i8xquMXsPp8a3zGT+56HPwLbq+qvlXIDYCBzFhSP2AQdJEJ+
nnjvOqKQbWjkbVvN9Saj6+qhwiPWvyG2p/Tqu0lni5GGJg04ByaCOMKHLa05CUQGP1LuEDkNl0AT
YD7Tdyn6CzNd/qdPJ/MYCc5G1bnhX+z2p/gpEFrXXZC4Wap6aXalCwpTy4LJLpDBNvPWn4g/PYjB
kQGp9dBMXJSXdLT0+FaBjwGkZvnR3W1ybLC35+0VdCzGyJ/UXhgU8G3++Cmv73icQKuTF1/slgql
0vgpnuZJD5K1+rSMaJjNMaeOZ7Dun6jBOudXV/lG3NLXF8iQnrHEAwmRelJTJqzbx3S9bhdP0suv
s4WbhrxgA5rAqMB+WXv9YPBpRowmhQOxXmPPWqVjC8bjI7PNw3LyjuJqPubBv2W/3AaBYsHkWLGk
ubDr6s3M0jJ6qBNhg6Yoo4j1sWSZuqjCVS1pvys6aap8jCEzsuFHBcN6J+sIF31b4e2GgPer1xgV
y4xawrmRAD0G++pUgPDhlblVfn3KxJ7dL1ZHrJBrYmOZRgRRI7aMRYl30jGQ32DK+pm1kFWsfiRr
5BUHERxJclk876wKeV7bdxPTmp8RuTf/mxuceIIadC3m8nNS0eWda477krc1sb6+YbVT46WBxjCM
AePGlcz0wa3v+4oGGRbp0TOyMPvJjfAj1iWjaTOVuGIsOZcxJESBeowyEeTJb2Cy6HnHNgIt2isy
Y9DZ4nZJ9OiaYkxDlWovV/KPwPPrOPqa/hBUZoAPtTNqE4BeokaYShufx2B6UEVB5vp/a41urj9l
2Ow9Yb3r5mksSIS3OdEszvldVjnqnr/ZJeWtnl4jOwHCPimCghP67TGks/86tyIYIB4WcqxUy6dn
4tPM+O79UGBEV6UKc1jhrLgO6PJG4aI93v0rBPgZfdhD7xKpURpnetrCtE7fDCl19Z/ngIuxDp0C
ubWsHwETuff21hpn78qMngQ/YQmcqVJKIJRIhNaRRpzqrW5dj+n5Xf//dR6qJr/VSqy8NHMOqvsn
fEiwy2N2yfCRVqmXy68rtqETMJIWHt+dVN/1K6rp0DMUKRlubyzWPPoBIhQYlOqheXnC5uZmtP34
oJUAoXH3lRYgguhJcfuJ0IqdPMzIFSqcgkuALgme+0JmswPeC+3klFAcLAYq+DfSo7vyYZQbYa6o
uZCrhyKfISvQdvVHwGKtKwNZq5odmGPvE4Tt5fnfDCPHr8DOStwhV+0l0uvoaX0yP2/zy1WSqcDn
wSEzKc9btUkTQOZsmTvHOWGd0ZMfb86wngJ94f2UbOsMz0817uAiEcACLDKtGVeHZ3+jF0b8VK6E
kYKNdJMcP56feEhi7ZJhwMzrk9+aNC6CQLRyu7fAQk5l0pEjgOBh1YVle4gYfjA/vK1xfnHgQzTe
rjzSAeHEjguXKaCJks0o+kAk9At4hGITMm/fonAp9OEU8W0CBRnNLKd7Lbhqwz+MS8OmcFbHO0IF
cpH0+KLxpr5fx7z5zzVeQNOVBigEIMhhzIlYgbddXyOlOn+l+MP3gNi1+UVSkZ3xSp+O1BLeJGwl
fttqWsi3YlSMJZGmqLQQh71f5yW0dtBrXJxlHG40Okg8axofXXW3jCPvMTVuYtPxZ9UYlOL1+eZc
fQMsnCpoMgD9O5inURhh+Z9eRCIcNhKg1PDqnZpUSWqqL1s2GAk9AqPxmHhfFtzzhPweS6PUZFSe
xN+ctOOAgQdrsNgqSulpCF+HYJR/BpljsWxypo4+I9umW/q+dT2xUyPdpWFkgUWHyo1PGYb7KHTW
OE3lAUNmqhg7T1Zn9EuOfUvBmvzRqJnzI72fgeEtFO5t1do26emeb/jWRvZulPkp4Je+sl9sUBkA
TbuDxd7Q0Vh7z1Q8izfLpKkU1jrYsjf3/8DSvGWtMGFVaFemU4nkmHww7ReELdlaVKhtv2bVVY/4
f+oWTS1Jp3j1kZbl5LYJyFCnLqwMTfdbu95t72GVcP2UGDbCYxYXbHnGcMfSSsBqZIqEZPKgWFhe
OKJmxsixhaAE1aQ2Px6cyr+Kebm/QHnWAGUprZRVK79YMlj9bQ+tZCjRhm8A58dxvdAAo35ktHfy
WzfjW5dpep+UGMNqOXwIwa1WBck6ox264BRmzKhGPjTF3UobccBUt5epea9DWi8A+UhIvPJ4etMN
4udXN5Eljprc7p3sS6dkyEKkyT2TZzN6hY9CpK/H7TNeS9WEeEO6YHh5G19a5mUqvVQV2r94or7I
QhFsPtuvo6uM4eSCvKXk/0m2CacIdzzTcUXUVFTNrMhfh2IS96VRAkG0iS1/Ss7m3apFn+0sVGK8
qaZAMhAuXYvRlgdSaE7roq7H3vXVijlKCrY3qEtmgOZ1ewEyBbjQtZz+726zUF8KkhVpjeqMr5YG
5Mv4yDH2Ti87AE9NM9IERug2091e1uiDJTOLngg2CyHzHzNJhMJdSCOiq6BfMkweRnxQx+Tc+2iw
f405xfYjJzerhvxfojBIQ/1Z0zOzEZX1K3SLF6qiIQcM61eW6GZd4rsz2aZimInP/ylmd5Tg/uk0
L8B7960KD6eiPzMct6SikVN05WxyslsNJOFOyoEfY6EEiC+O/dDnkC6XWlxvp6tMQ8axE+DhKr+P
Ui/rmy8qlrjsAmqfB8l4ufLNqSw1Ud+9lMkv9YUWsnuLFFq9Ij4oshVRKklBxlqHx0XD4FovF66q
imErWP2JW+Cqmv4SNqBKLqUPz/nF27+Ewaup0SWg0y2RedymPaBqKaHCGgHnuaQ2cviuIDz9Uyq2
HKcqWokWsDCrdFTP86RavgADAbgL1EWb+tlfi8VDnyKOOi8hs2HCfkdaENErdcTOgZA4RV8wzwFo
7qlBu+kifoBu+xUQgdwAI+GkLkVRyshnxCL2mP2tNbXshsEJeZMFhAuqLr5R1+Joych7RccAn2PY
NnVyKvxrVTDxdbTiZ8yl5M+646bcDpod1PL+NuHd6CAHGj82y7DMczGdAR+0EKJOiUrbTId7rsve
HeJrregjKoAxrwlmpegYR8JML25y+Uep792eRn98X7ShKjG1iyUO8Wk5SgUddX/xbfN351iYTcDD
UfMCLVhGLNosuWHmp2b4AaplYRpHVQkVMbgLQUJe+gUZlR1NwOQOKKw9PgMEOT40+mAY6timWLFz
X2UF/OLu0/LXUv3vlefzfK/PFL0760STjD/rWuWHCsqK3yAhP3ynmELQJ87q4rQ0y+XvCSmyZLy7
fHh4SllxzAPHqcJtkA1AhVtgRDmC7SKxraGJgH+iqE0o4MuCtY2dimdH0jPjTAjuJGNnSF/i/zH7
6V5/yglqbPo1TUDy8uzTVW2a/pK9fb57yqDenyTjR14kisJrSgqT32GsCyOd2ZBnwHUUOexX34oc
CR++5XVSF+98L8L25lHnsgPMJcmrZOv3FNmCpeKS9iuIl5+Arq9fK1QcTeLf5LWP/mfhtXVLyWy4
jYAY0YgiGYAaiXcDVMMDXFQL4+DrWYtgR0sFHvdYPRjM/b9Ph4n2ThsI0sDwtVywMOIfHDYCNXqa
+NDZQASFy/atDYv7j7vhiCQtl7W+eek3H/Fz/Qzz1cy5lNWSUB866HiMZdY0zdfRMno55bNGpTQ7
18t4nAWC+PlB3EzMoWdm7vt+HJZD+4N6P6//JdGanyRD+M9mJDpsjTIDYWnR73nbjUS7bimYP1K3
anf6nspx1YLVM37hq277l7Lzb/c5wzxD1lR98gCZTl/pPQ8pn5GiuS/M+u6+HPPgdXroTZAyLT5N
AGhVpT6TvxgOC20bWhIrj+7nejZBLTKbahfCudUmjeDpiQwtzoS3Ha915OhHYgBarU/e5KRcvlA9
HSBN3IetraHNmr/o1U4z51aWBfhY05qbWX0th2CdzbvDBJ4Bi3FkLfkMH/76iEE1Nm6AB7Y3KC9h
eOt/8zrSYBKKeBnVSmlCVQo8sB2PwJU2t/3lOOQS7Ogz/naWfRZfZtevcdxOKEFbUFinjfg4FxaV
vK5JUKQSbk66qL4sdjjIU8DaW9FYysvZbx0xzEE38F+Qwdty7ZRq8Yy+QnvdTDmS+VnLJ7NmSbr4
n0HyoJkGbmX082W1smVH+fTV/Fxt8lHlEzGvhkq9+RRZcOV/isVuYqXBr9aaG4fCVioZ1VAUC+Ww
5gMhaGEIdpaHyAsFuuxgpa0YAi/VxyMJnawXUUnO2NChdSgWJXuKXDKeHZTU8aOziSjDdBhebSe7
RK+QfSi5swSU/euh6ui8rpsjHM5kbzVG6zRvVHBPCaXf6Z2MW16yxtK3Lo1OkEDYEljShIko2Wrd
uHhkDqFBujGHTizxAR1EiDMywAddvomqoGWf9MA6F+KO8rR7t+CWe9Ts4+FcplAkUUYDgOSe1fwz
q2qEcYM4VD5HCyMs2DYVFZ15v3rrue3tVPtrmyLsvDDYLHKkERfkFQfDFgd2yJSkst26e932Gn6f
180zLzoZ9OnlE3Ax88/Z3/+2P1QFPAJFZ0gok1+R9B9X9zE94I/j4f0Pny+TbiJJ4VilW3b0Jp9n
O4JSTsui8QJOaz/EyrUkbSbhyh6GWgLDxNE62omrMd8N5jHVNZPO1xSAvwX1En618fppmGe9urkj
1+YJSzWqRT0vMGY8D+JT3Rc4L+30/XgwU02Ba0HpjxYNTs9A+EGZOb2vqJKoPBe1FUVEXx7MZdwy
fcC2XH48z7juq9wreEiojfAamOpxelgboHbInEtZJoJzj7ptPxTmIPCVBl4yj0t3vwVbqUSZnWSg
M0rCNge45pRRb4Z+6D0Tz2MmZDP/iaBov5380cCXMEZYHi2ibkZF6qUO4yHd4h3sskj/YH95Qn2R
GnxpWusS3IRAzcBgPN3yXZY54WJMqIJBPW8bunTk2S0zhhyiZvoBNr9rl1+tAR4Iz7vyny2pTTCn
VclY7BzGAbh7tHoLV4bM2rXi912WbdiJLDBzfiVePerHs2yu//Z9jpNEaxD16J+kg+QGF+484TE2
WsSV8P4wo9masZLu3NjN/hTcAKUBg88uDFvz39oyd5jdkoSxJRpfdK99YBhtn4srces6Ri146nJv
KvPa7hlDNiEb8IfGBAzTECXFp/vtOAEfbaucXL0oj3E2UbmXvS/SN/cJBDZAi2AbtP56Z46pIud+
N2mYI4Bz525v4/BI/LfPnSdyKLb+Y0LsSn0ypgmD7FAQEVl9/yXsLR5bH4dLuyY+PxdiEPFI3CO6
Oon9xhUMWNattX3rk7SP+EgWB6yzh3h8ebQXNl6nU2EfIs+P7r3GEG4Bykl0qlljZJyMkDDELtSc
KScSBj2DvjA4FZiIK/MhWOu9HrPoam5uPZyFTawwIcYiukUCu2t5ENNVvpI0c8phovW1ycjgF2nA
GxLlMAEYzLpDJdgb5gbArMJc1Wz8JiPTKGnnRD3sFxZf6wclYOcwJWa36+rVyOKfbrmXwFFCNimP
c9l/Q/BuL0B6lHIur/I9Q7FNXHn1tUkCS3GmKn9bfX0Ga3MIlIOkDwOWK2fMYakwuCGdkBy4OQGw
IAHw87N3ZGFxs9rJWqA+lofR7tD6ftTGCO6+DrazoRx+ghXah9uHwIWn7G62LqFHdtTYU+rfbg4+
YRvlzEEZB21T8wHhkJnq0N8OYv79Ws339kuPaziNXWK9VUviXY2BfMofrl6zoBalJfHCy/9fLr4q
9A4xlx9bPYMlncjYQ7cMbyMOCNEabGeGqpJI7XfdbB+dyctwxAA9p1Lwp8UDOByzthRg/pXH2l/y
7JxVGZ7FbM2nlj9UqEo7e39/xYJF3UfdDp76xO5MkkIJbwVw9MMvGSvXQ3WU+QE5MHxkZVxVB4c1
KghlSj6cq/o+7r0voLJP/tc3KxcXv4U3PlblEFDhGkDOuksnwgXZmPrpAy66E1al5hPQ6spRdi80
fQAtGYxWrtYaYbxPEQsvaujLN+KQtc1G6Gr3of/Vfu56D+lw3K+Aue8vthsDlW1AFrYif0GE7VYl
YCMceAkiocMh3h0P7TNOoVUNASos/Miv4QOlnzWphKQ95W/CXtKDn2phvcghx2LCGG/5XhOOMxP8
yoeD52ugG6+53ribyDj7NPGJMGlI+73sEovVeGIQrXRa/VsiBDhl/Qp5B03nbXqq6ckUJL+DXuLS
zK3BHO2AnHLIPj/QjC3md3ZqQ9tcK6FwZWsDOaxmE9oyqiKLm96Ch7NgyY1nJSIisUSeXYKHsNtI
O4MyUGO+cQ1ZOzCUFSzGP7jQ10aygSvtb+MVzXi5qRhSk+00yxRXxlSWQDxONZIN/3MkWprBwtfq
97o6gLvoq0K2RUkDI17RHYAeKaBmZCJnEIVgPbKgIfL+2hnhZO92hSa2YkeB6zvVPnW4qcCQVEgG
HfV/mE6jrN+4HpvUVqDzERBWNGh2M2hsRnC75qSQhggpDc2nMSUnzGC+xREd9Mpr7ngfITMC+BX7
zUWqYhPmF5IWvGUeJFj4Kc/8YJHagpPk6JXKvL9JO+ZeHNSBrip3FYVByFNWXmEOSkTiDNc2/mtg
OAUZ/hZavBcK/VuZAQNHAguOi4lvSrYD6Q2zgZu2xIiM/k/WHtznK+3UTi9fnRxGJOpPc1ozc1U/
5eT3uUGO5+y/5T17Zle2SW5hOFbeFAYpcdnAlVglfttTa8j53OYJh5ww0l+VgbwNjBjEphqrsEbl
qFemkmTBWoJsybBM+yI2fkKuFr6ZPKzt+uPdpqS3qiR/vYN5vrl9boT45vUjtryx4P+ThJlzMWue
9A1o8sODbGgkzjitri+c2IXGgmmulnzXFvrdWqj6R6hpJrrCfcv16//mL63O9FHuwZfHKXrGhqGZ
vMrSpqyid2Qv5j92YMrcSH7Zb048X5DYxg7fan4KWLUHQNGjtPZIi7h+Un+ufuwUyVQzO9eDyc8P
ILtrKOk6MQedJLji0TRwGZCcL8b9kJYR+VE1upEZthu0bQcF8payb4dawv0RbybKtZhce5HuvkGu
nfrq7KvNdMTdkwwKb2b+AlEvRAISg5AZG75ErdBn67TpIfa7Tsj0gGKbAOFyoSDOYsEYH2d8arpa
0In/qu0x9qSMmZu34a7wscwtDIPfteLfQ02HRds7KEYFfflzjkjcq6/lXZgtRULQsb4rcg4D8+I7
yIb4Odu4RurhrUAcdOi0yRU4dvsK7RQhk2AI4PCGIEmSd1cewVHYNybnIvnfadQHuKDrZSHwwd+V
JHivrhn7ra88FnapDd2XXLUdieU6ciTxa9mCfpNM3SX81BNdgzoA8bjdqT8MM1xaORq8flPioHSD
z/4Avyh0qkVLCocjVKUaP5Oy9rXdR9Ng/deBOyl4zDN/lHeEM3xpO3v5V31wJ+4DAXFcOif/esvY
AnhzlVJAAxP82vS1baKwh0NGk5mSGzDn3JO+Qb9iWkJVuS0NNsRR6Ksr0gKLt3DF7u4ffGv9sbQx
OYusXVVCEExTkdKXuUMomrniODRBL4Ih1URYhY41s5BiLh+JGc2KJaCvYzJTdZLJbYl88nqnkkI9
psliD/hM6bgBrgX8KtcZfEp8wH0CqXqcqwUmFZUPcSNiYvtLpqkz/u4B5YmLMFg0LK+oA58vdN5n
OrzvIiOMG2seZjXvPfBnqzJvt3/DAM2vISvMf642zSmxKaoL/cHN2oKgcPEZAMiyNGU03BCoxyOK
K5zBaZ46Yy4hObYF1966q3fiK+O2EzaRjuKiNdyuf+TBgtVL+MbeOzZH6JkNOQTry4CYk968ib++
h4zey+2LyzIjEHqewNSysZo5PeQn++d3KkYCtPtNqjlD9rXTzyz/HtSO8I58lSSV4FKhJA4s62Ms
fvM9HBd8l0p6ZSwVx2QXd9PMrXNSBp0cNv8zctOry1K+3euzYdfm55Uz0U8Ig3cVc6fMLUGB84UP
oLuzCUejpPzS/lawatDEmT0p/HrbzHRdNjw+8IzHWcHlyLoALDMu9VfPYm2DR2IUBn+pH0L47aZK
McgBat0PnhQWFSqh3iTpJt0nXD0zsZX9AgD0Uf1t9I3VpzdenZKdod8HPCzjVCFEW1mCCJrNeRXr
9YMIqZOgoxtk/Y6ajPSc1jryE9lwiPXKOCHx6W5Gg4U8kZj4X+6NMPgpa9VMM2Q5X5CqA133pjD1
MVDACS74GGmTrphRXm/DvQSZSBripppgyRiehpO9+dklhZZ1hctAks+S1wvwEMBwL+f/5iJ/NS0C
Ttk37bTNMgDQ3G0uSvtp9gR+HQRaHCG19Qh/QXi5Uc/Jt84q4xoQYYNMt+Mx/Ye0Tb07uvU2wZk1
/dJSOw/j+xRPAE9SKRw7TQr+7LSLJOqGd1Nkx2jOdcrrKgQw27vF54VyEaopV95cM9LkICbdMcIc
GqhZBcK4aK/pHSrL2uAV0AoLHBPhiPKOAonf9H4yH4VpIMfRKxVFcD931LGxERQBHgigQLYS1LxS
71IrJ9n7jAOzWRHctwOTw2TP1qUaAn63qIWGwK/v4rCny+g0YdttF7qdaXy6DAbTuwqY4RhccXNY
/Uum6TAIPnh2PWfqzbhmec7YLz5RcdzBdNDTi3lruFDGIYEowpGnqgXYaqZS8uXJbIEdMBq5k/kL
hSkOq0eQCuJUOAzI2ATF0wonSiCRUa+wR50sJ8IZf42jdQEPER+4zjvkXk9DfMmdFnSuEfpgCEB0
GWL/e7QWXLpxRaWahN8ZEmTuW9KE798rBUv9z90iwiNPMN3YnDUehWdg9wwgRa3fGto+spHL9eUf
5Hf3PH1FRFCjgQmqj1NWXEetfOADsZyKRMie469DD4ocvd/SMxGq5CIRQw6QsCkGaQ85GWXPDVNB
lBy6DbmPTLzx6MpvEFDh6Ct+SludFaelwNoup2dUcVlp7qPUS97K/cnc18PdAs7L0tDVKW73jSEd
TheCUSk4p3SIXM3O6yYFxYW7OIUql8FbxKFBdWWaRcWh7AEuE5Zvf/4O0PQZEHjaFCn2pDmsabZL
xM7KnbaSwmgYyR7d4icKVw60Wucr46jHjW9pAz7pQF+n9jtfSJaXamWXddMMSDJRob4kcVWEc6G+
1gR8yYKX8bT+JWg7Vvs4CbsR1HQh4te5pZcK+lmaQ/pHxPaO8BIWd8NS8nmK4zJbs4jkCsuJEkxe
vFJ4UDmSnZIqkYlyB/BabeI6GDoTX7SSiAXv10QJY8Zov0PRnfg8nAPm3BGhMqMSDtQPg2IwAJ3s
t/vJ0tVVsQLfGG/fIm3eSlPefB21i2gA3zf/22U5k5fkOLppNnkNHUQTa/Dy0B2Hg0x1CZoy4HwN
JrXS5hynHTXpAj38fOuAr9cvup1wc8byWCizw4HiiDX/INPKook0lFMbu15QW2noqGewBcQ6a6CE
+aaYFVqDjHtl4RYI/5Zt12AhlRWsvXbewgcZqThPQbPwSK21suNEwT7UjCwhP749TFHD7wIri5Vy
y2rLDh2/lAqmW6Q8J8OvONXHHGmpIIFqH3LwCLdPIRE9ppyDdc8b67Tn/vvxyXnG9exrOuwqBpG6
WRN21I6PrMxmpWvdIYZAfptBxKB9afGtwYLst9DhqSuVDlFMB8D/9T6Xpjtau9LxVJ0H8EmlI+qC
YHsosZzxqvGJIoWvtTLq6yk9UXcxjtXB2cvVuiXMV7Ldn8qwWyd3gi8dluWvbnSZgkCfBHqVkZ+j
PhNCEbggR1JJ1570ZST8p6hohYG3XvzlGIRe0tJLiFhPXD/UFBcab0Ft1RChbMLFEG9wFzfQjD4j
Kpeb89cAwjvDO+hVOSEVL8aXXfOQffY5Xrc4IUTBHxwE2Bqzgn8qllvwS1H/8+E3EJxjp+P+VyWu
ocus0YQU7YTM4m2CiubO60WzEwROTOuew5h0ymKHng27Qg4GCYgimVt1BtWfbk0kemZPREZir3tw
1kQbtQ99+/hwRnwEpS3qxiZOBYk6onbtBnQmjuwpRCxB0b2PsqDyKyN4FwH7AB5cGLkEpaTmmqB8
t+n5yfXf9X95BounPOyy09WD/TNjVMXDK76avNVBsPJSLUfCM3Vb+dw42qilR8TvMtkKjZXHITEl
M2KV1zgYMdnI7WoH+RXCXWPeoyBL+tAXvrSHoJs2FrE3u8aY7rMIyUVdHml0er0GKRAoQVwBmE4n
XyrEEBYBeh2/k7OlfLbSxY9oDIdTfincbFitMj7KSkp/MSRpYwJBy1E5OcV5Z2cYqvvANw++P9Ap
fRvW0jc2vTI68v7smbTxvRyW23g0W9PPqPHsOtQRnPxci+fLypsPiYMSDUfVy3jpO/kQeMxWgda6
qTeued3Xqzygl7uNAfqDJQpi9N9fCo47WHFZ5CC4ZsTfkndf46tH6X6fGZxInNjRIjU/rutS3rFn
3OuSEoTLZM6I6Hw9PiZdPa0nCDU0FXDOpZYDf/3NLUQB5ulpGWC375K8dW5kw82UxLkH1Gn+bA6t
rtk+bOIP9rA/H3v51e6CteBg7WOOUTXmA3vUj6AgLgfdTT3dAxd02jFWT7kpZ2WPRZcluBxo2nV6
CMwzMicWwRcje4ByG3ChOVuzhm31XYn+wiBNd93J66qdLGG2cJlmdY+v2QA+vcVlRnwTkLvcd//t
/wuyHIpfSLNid+fx1S3LPl0Yx6+BzdUNErHnHhKucSSAIqeSOipAbxoFUmx87qh+elRAn6r9b2Kr
Al35Z+dRqRuxKnRuVzoI6gHMu1UOuScEY3M5dnX0ojuTsTtUo9wABCRltOQCmRbRABGuCvSGyFY3
SVhMji9L03XMJZZ8ENP8MjOGlo3JtXUOzrUoWSJD8jzO8/GiOaTUxLj/EkBcVwOhct2E/cuUFIIs
cDLTbngsKUmVTQFGtPQqVJoFN7a2bBT6XAPT9PQYfkaNe0CgttR2ONjAvwOf/EJQsoVItPwQRlMi
CaQ+jNDkaOOcHziOal99gA/orVKNi0OV9ULaa9uBAg/yNCINzpes59/bU4Suw76vom/33sRU4n0U
GS2iTi3E88B9QspdGEHpCt555amLNQsAo+Rg3KMumdAeGIN5Srn030O69eJ2yN60c5ZiY5l3EtEa
vtIaljsQCwyB0oKf6qRaLqFiQsdmQEIvkQM0I5yibnYPKfkbnxVao3UJaYqg87dJ25+86rcy546j
M7m3KNB09ttkYfbe21VxhjkPXftGMeWjMIWRACK2YbaWU5ir6IcCoIpHDJrFgdfyJw/GrVkBNVqp
evNwqi5kiGrv3n4uUKVf4Aqh4b5/dQrXOGRC08lRp2eTGj7i6NItovujrXK7xjYJx2B2wK4m0Xir
GE6cCUT6ZFy4dEbyIeycQuXt+cttYW0PdV/oNw7S7gOFOFGawO3PLXwXG7rn9ivQeXlxRLz1R48y
CrvnvSlz0eb41ejhBQfxOoBBoH5hmh7/IOAf3yMSyv/YhVyIGmzCgOtdq6bNsL404PvLTnec45a2
+80rZx56bQRjSzjEk0OWajYqs6NyLxFLhm8bbLKUPcAnS+ASfcbrbHARWJjdUpw859a+/hyjpDAC
sL3DIPo+bbNlPu/fv0dOsVohPaqlv23bD3TfLGCsfYzAILVi6A7yWC2HNJIEHxgGfe9nC6s8P6fQ
qDFUuMtVbxDPBlbJitQMspcDsZGfF3bdRUnd+hXlzPL3KqbqiveeJxVHqO61rL/+0uiz5AZ7aMjX
IpaJXUN/JfBH1mxtO/UfXVAv3vL3BNBQoe28enTuKGjVApsJLBrt7KCDZlWNC/9vDCFxZkd+EDRp
LF0Cld3F4gq1+boHr+rfp89oax/ovdyZWybym7xsF7KS03/EP+F2jnvcX28b58hks0VodgJtU1TG
xkeROWkBSMk8P9q2tQb9H5hXo7EVHW7kjNG/7m2wptT6Yb8+bFv6+VeYOEO7OlyCdLJY3nngd5F0
FtOHOnX1fauZCLrVyKLghI52Hbyt9Tkx/ku0/w5fx6lrY5T4LkuUtop4OOcX4zWwcnV67tljUnYH
laqlvFU1/ywAuy5/m0XtZACKi+CDllIWeEoxZYGIE2+kfi+EzcDJAqVU8AvpMdajy6olfUVC3IYs
0jXFuD4yOJHspFhPpVnJ0K9L3kJQFsAzr4L/6lzSYtqucly1E9FYVlLpyeoDNMSUPAdHJmRHp7Iq
rgZD4Smp8o8r/mPJxlgc1jGOSYSHO649/SWVZft9qj5aqin6yBtnzncVseE1IjffGgMhPpyu+wKj
sxg0KFNwiO/ULay/bdMjzDBvzInC49g2kyyUTx144Q6kWyCBCOr82w4XypTN+g7TWWgdgdhF+3F9
7+NB3kb1r43HU02cK8/uRUcLPA8S22NbV1z/PLuqxHy4fd1UzRoDa8K1l59Ww+EE2LHzptH47L7m
27b78mTNb/gMp5MZZDAm/JbtfWFpmNDoBBf+zRKoa+VuSDWiOrNysT6JJGOXpusW/TuASazHHQsR
RQdXsx5UOMdr8Uzfxaw79l2Cp7eaVkfgCTt12nLNALa4DdhR7MVllo1TeaT2Z39IS+NZb9benL0b
BIFV58EkzXd66eCaYZsgKgrJglwELMMxAF7ntYMgb5Z0HbKbu47ZfTH2J4c5HpEgKBzJSkkwaZGa
PtxcT9z9cHt9E2e1yMRvAgxFig2FHkP24y6s54+TxwjFbzCEhPkzzPtDmgGo3c0eOsodmgcb94eH
6PAd4gX7sfALNKJhPK5rsnZ1hLqFbDhHQmbI22Yo5VwmzyQdakud2ALJN+Ah5NTRwPD5U1t8WrBE
m45/sHbWqeiEYg4zKs3HTMNg9bWZ2XAkkk/Ry68bAiZvIV2TYDYH9ti9dTnFSXZr4kwBejudk8wV
gFphHrWd9yOrZo6GltkU23yIPjid0kBchgZhQCq2gFOQAxLgdRT9hE3rJFmqttpr6a+nm4/BmcLl
+I/sArlOsmXEso2PZPcBe6/RPLWgHAMs1apAqcinXRIikU5hIM4+U105vNDuSC1ui3lX/eZ2tsdH
KmQaRnEd3GWpBKRU8qUeKNx++tXHIVjfkw4VFJwes1wG04J1z1aBx/ZYmg91RpcsQXAcNJWrkZzk
ogOXVur6CnEeneAqMo9eMnE0aAb4SsGo50hRwd8IOG/e0h9llc40smigJYMpl3k6+cfhsL5eCPPK
XbR5dP91b/+gOHu2rUROrUYpe3Lt4UYpbzqEVyNVNtYhWaaRsbFsNZAXvXOXS6dtPUCpjgnic6M+
jJQ0smuTkkBpfuovVRm7GZO8EOlf5JeFN47rnXx3z7yC0jx1j34noBHilbRHt+TE1okCKue/VeFV
ZmjZDGYwoP341HgvLvOrp7YlPpRcciRksALzG2uH5Ju3f8g/Su/yeod84n39ej5C6fGHTXTEqOgW
RYvO+UxhPCvf+DfZ1ur9wWPla134YX3jfx7ejLyOrZrAND7ZiHNvyB6Ao5c6AhXTDxBTvgqaO4O+
zR7ZtGSrT0TNq3NXo9vFLy/J5XqCMozdla0Bep+x25UeLxJeBzd8OCeXNsJW50g3am0ooPGWRbX/
XDrCYHh9UH3v81cwo6f3xxgnvVjU7Xi+r2njSnovYc/YH6xI8xjdnFzEPjtA736LaCGFYnw3krrQ
j9wtuQmdpwkw4qB6UpmZ6OvtOj62OnB+uNhRdkzm6j755PUJjVbO8hJncs1lQONrq51DWYEFaDLU
YznYflswA3PsZiMzDju21jaGybberP3EMmSnteL+p1iXCiIgfRBS9K9z9AGHQNaBDAe4BKqKawt2
QSwjzXctjZ9CXzhu6jRlIUQx9ht8Yg3M0pHwtNVmAr++BJKn/o6U5lis/w4kn1uLhUGOwRYduZq6
XqE8Or2XEw1tyNEKd0WTf+QLzf7IRWHf+NQkpaJO4QQUDA6l9zu0l0WbYF4QcW5tZaQ1LECpmDbT
IywnWdM8XRvOVrjdPQRs8fjRs31/VrMofba1fFT/3ziXjogJyES7Jv2PTldHPAmnoP4r2V4yoCnT
suPsbPtfznS5tXzILDkm/qklEWh/aK4gOel9LgUQwJyxdgeJVzUExuOu5gP1Bv3mNaxQRZK2ZPf1
PJACEHLahRvc/Us92S1Q0J1e68hn1NYJNINp1KBBpelS9DD6jToaT7NH17a7/Yg5voramZb6OHUr
leSVPfNG8Nc3Ymtdn6ZCGqbjiZEmNZxzfAyBnKtijYQPnRdcXutppXK7tjHjq+caelIJ8Mao6sNk
brr02nPIxoRf+8nAcbhcFHKLXwfJtFpCHOCHyYBAvW1+CuSjwqmRSOlvfLEKe23ih+vfNLmtZLo5
nlP8GEW9lFxN3Rs8dFtWz7PcP9ZnWw9olw8JuD8x8GgF0Xr/h9NW2zJQSSvrh93gDIIVBXB4Yw0E
We9a9sTSkQmsGjKHpvWIaBBawjuj93NGfNb01nscHzF/zQ/av1+59yQKM+O598HMswrF/zuYgDVR
Xh35T79TIAmo9Yi/D7G1UYoIrO5ZnV31ecGk0wfXMtf7y57i3nW4BsYIbd478hHWOOCG3Ut4k8GC
LzRbKqyepLf+teJfBmK53zxCk9Xzg5pHJsRQbCm4Kdt/o5FUSyXh6UqFokT0EcaNyAtvs5wUCz6+
O6NCdwPPyZjnhTLMfcxKeGk8POq2omvKkHfTy6Qv0N+wGOyn617fz+5wA4aPd15V3/yb1za0o0et
GY5KgSpBGRFPw5xttRXXivWLQhMXoyGc6Qshas84xbsZGef+le6Iao/O6r2kzVPi72Y9BSdb/L2I
Nv9uVuJHWu+ahrvXQ/8imQN/10qyQCVkHro1a5Pb/1/j0f5mSZoNFXVz2iile9Ltr87YG+7ylh4p
5CZjF33ejDRyAl/TbLVVUqyP7tueh45bnmQ8+4laUPDXwhehb0yHkyVzihUGIxjTblOf5XQzBWoV
jO9Xjr9qTRSyP2GJsV8/HIpDdYqAupJjTs/8iIv2OdrwPeoIY6RRzMT6mdz9WRgtrBSwtB9n9RX2
u/nAs6g15Ju5zTUnKob6izbCsQzrZCDGTsJlvCfO2o0hcWKi4kV0wuH31La1wkpSRmyn1cUes1Xe
PbYZjUmIPa9+3C0o7a1eSwXEMqrxxnguDCWgzbDL3QUThjM9McyM1xB77N7I+d6jcfJFTuzVww2G
aJoJtqjkKvddSjIuHMDIHggIMSOTVLkjXAwFAwjRsPqrwp+GhcH69P2UFD6G/CpmD+toxOSohMNS
v/sLmaXhhXUKZEsppWSmICMrs2UQWcjItY3ySLTiq6S3jDqaVquaXjpxy+np+Xjk4aoTiffRVbvE
m7T/6dmlPKxYnyXEyhiOyjB5VOsDAU5u4Wrovn2+cVl9N6iV+CLRGH+5WO+n+In9CDFpcHAmLzXL
KNkj4khW8mShLzBRuDRfeTQpca805BQs0upU629tqdLITEGtSEINlitURGiYE7XOIEeSdIVKFi++
5huhHH8nu+Q4UoJKnIuDQeE0V33o6QLJ5rbvtHkv6k0wVlWOqJRqxoqUbE54AH3QT3T6CpaPqmzJ
ulep+Nb8708jSldEFSMO2/sSbY9WDi7S3YuCi97pbXiKlJnv7ackn0Sa2l0mh+IT81lKb59Y/gCS
bZO2h23XXxqqt7ZAyw5u6onQFRxVkwqZZl/a4sgOlzrq3S7hg7DbuWku1BBpzz4kmip2/HpxZ8Jk
hD+jClMBeG7xG+nYCTknX2OdVtrysR/mOnjdTJip33hom6LpzSft8a1ZDAv3mYMmtmpIJd9uJLmB
a/DX7FPpDjCf2ebzS2rKl0RvMe4fgVQQeDcgft9QZTyn2Yfi773cUZpYbayZWybO0LlfRig0UWqd
mPZ9bkZ3eIy4L+You5I720dyTouhjgrAdN9oPTic/YfwX6ObLLoa2ZD6RCbbgRc72G82QafY6UAw
ApKaxdLu9UwHe9SxMKM48CP32y08Sm6y3xZCRE/p7wl3nQN03HjpuxjsrCyWWNTaYh1VtLlGzBcH
ldhP3mtVbhNDcs1xdzgIbPhhEEdJkyJtHbGoIM07C7ScfaIW0bl0JIXoy5761xnVSZchv8VEilnk
42tW520p1q/rv6pPXiPDolMk0PZfyb8hgZFv/x821NYh9ozzkiSuSc0sw0bZcozo9LzFBusbHWr5
+b445dfkqJnHIJ5ZVZcrbxnmn6fO4wfthQH+s05s8LzK+Iw2cZ02uSyy076mBcY8aKZIV5Njm/6X
4pb8njtAwT3WNf87111lSpNh4/eHZwiy/OM3CnpOFN8XZiHzkxlI8QbUrDxzbVb9mDVJjk1Xjnul
FH+Yc8wT/Zrx6kMfb4fg2b5LMSFdY6F8FBZyknlbNXiYA1rwHyGAOaQJ0z3sFi4xWoE5icFWfMZE
uYEOpANgCas1EmvpVySvowA1KIT99Rf8SjeppakszFcB+uQBaxKPzBRofMiFiWNYGnrQ2jkkbhJ1
ELH0wiNGHYQAinqMC502rF5lVp+zVh9M28MHE8voELIz9uzgl/X9eUAZWh95Y8MjqIwGJYIPCEny
1nOE4BNcpYOxa/Lyi57gNYKhoAmsPc2/C+kDFJVRg40B4zjqrSwI8wTILAY0BhEV5+yltJC0qAKV
epokUuuxmaxBscaZikY6/kjdunTUkn5GoTAqdrkoQxrf/kR5j04rFUaTW7Pj2NK2vGYvNeTv5Q6N
J8Vzd3UTu4QlGTANwivA4mSdC8nDEI9P1yWL9lOiNwxipz/r4q3jkGepL8SkuW+NbYRRBCbmGWV1
vr6ZafWzA+KKr/t9M2QTV4ixF+r6G13dRhuGrw9Ew2wa12hgIwCy2975wkY8DeBgYa9MZD1ccMid
p31FtZrDIPnhyE9G5FQSxR8BVnrvS/rC74s2+7ug1XebsnPq5aOfJiDLNv7w/QqIVLhDrHr1JHc3
onV4/1a9bzFqpNsHfLPyCisBOuyNgov3VA/gSBfnESs0Gj/r9cdmhzoIZR8abq8l9YqR7vCibyLB
ZXjiWj7ucdzq4rlBQecxwvK3uG9MF/hc4oiAFTaZ+1GUTgSoFxu0tB0+tmTRzxHY1FnlAdOJzyUq
FsojCYHLEvByM4vhOKTblGXPDjxY2fLposzlutgBmP+5GsmyFSKj3gN8PgRgEcpQGCWQpFFBhopw
5pbaYJkJQc5u331ZdJkK71hjGQrT9mwikYDN/zZ/1hKkA0DzoYaRu2mdQ2Oqt2vnfp4sAJhW3cka
eCNRZg3HkPpLIo2IQyKszfqUWgShf6gjUvVJNimAqs1stnbDVkKa4qxvo9qTSwHDzXFqRPIdOp7G
B2HZ7jgwS1+ZXTxAdmNkgbSep6fx9xTEP4wMrWgQv96k3DWFjeCEzafWoFE1vgvsJ/a4fOgKZgxE
4v63ec+cUdbKbd+HG6yi143kKCmubHHyTCmTHBE5y0i4vyHOha4YBu/GhcfvOLbQ1QoVBGSn08mP
fgSUwgBxiEvTPw77tka5ZnLxVbr2sdy8OM8ZdW+xGCzo1GRgRrx+SzRfvVGcbyLQdXWjzp1NxCl+
zQHaEkiO1nJZwgpv1hKDqCaJDE4wUMkvNIfDuK02Ka0OhJWjLTRnb2WFNU1eUUXqGet5VHS1XYhA
7nJvtdIw0S5wsMQ41R3AnuJm0hw0cbT4JhvKVuHVswqLVaGs4p9sEsCpTeatNI8Dqp6QiYBSLnkY
+7W0poyNExtNffMCilxrwD1WeSOTv0u4VZAfFoiLYYhlgxdVeYgfMqW7DsS3lnGcklDirv+Db+gc
6esytMR2kaH3RZ551r1mdDzwV7SNNb328yFWCLYIQMxuvBM5zp4R/Xq1vesg72jw4mgiOwmENErH
eTOkRcsoI4Aiwy7MkJyJ3eupC55SuU+WICwXOgEycR8Bjfhm5uElglTTZEiZq9u0EJ4lD0/beyRe
1ds+0iES5zXAk5fCdjW1P0rBOqexp1NQw1VTRxOlXLGXbtjhUkI8MWkqXGuL6UwxpUqMZgFRgvua
iUqumRTTIov/C5g1gdcYPbpweMXNfOfPsSb/LBjwJomL/rM/UgBGFzPd8IcBP1F1V9S4pn1O5zpi
guxOiJPi+yqjPYYun9w3GYzz/L40dHJdVEnJNIA9LbFl9xNYA5/wh40meOUQ9z0J+kpbhPYcJ99B
9FcpQX7Y5qruThsd+d05kMZEPlV7KsmeEG1x0XcD4UCzvou27du3Ml6MgiOUVIoqiMwNyBJZpst9
tfronRb6fmwRJtNo7nLp58Y835VrLPqmY8KS+8Di/qhNAiC1tc8Jf7teLtrMvgaopbmkNbr/JnV3
gwmkERWrim+Ftsw+67afjlX/QdA4jZwjHW7gy1wHWFtv2BffR2a/FoXPwzG8lAxhARZZkQZMEHVs
qsqfYHVD2sXHv+oEiwZzuXbNIctzFCTpfnqWtOdjaB7UKSNkB3sAnkN+EfXQQB9C7cP27Wg0T+dX
TGOTqYNoSQnSTO6XKgEt+uCDIU2w2EM2afoBt++MHZdoUTH3qRcmT/E7RL0qj9GanUVCorID3fV/
DevVRD6KN6r8iOyBEf9jCxMxNr31EGSWrFCxAMKB2PWQHn/yUH/Bxy1y9GqQBQrZVexq0BC9+XKD
iCVCzdaK/6yJjba1MpalHv7HJVmqXJAwW8TzgdgoZmAWx34PkVhQa2+7YSzVoyqcw2Q0ev1qjacE
Waxm5IIGcwonNncmyMwJxM/1DNDro5KGfX4X8HhRWNxgblw3Ypd4CVWWiSMOTRGFdLt0wruwn9ul
IZBua+0pleFuDUPKSEntFSN5KyeYKPM30XDzeuJPjnMAnj+JZl6QIwSKYZcQnGRzPpxD2wZ39KW2
kRdgZu37ojmd6nhOg6xKBwktgpjW2+mz2zL7e08GOTI7oBh2/sCkrzEUzSo0KZu6JAjv+LmbIRLr
3rJ6WEdh2n82sP8v3RAtdT7NZi8HnPGB3VQ0Bz/fzophJ2oW//gxSycEgs8vZ6VqO1PTbQOHBdcR
E6hTJPoRzzdIyxQh+5aChWYa/zoNpPTJM9+TLfn4tZmB/riInZrrJWSk+JIfQEmiFI8dI/3//zu/
0oF2ZBdskkA5yJSROjkXGKO2RKI728Zn+5SLs1dvtRJhBjoU/mdz7GfVPY+44XMwRuJuydnOehBu
xSIBkBUlHhGWkTewnfFcTJ/7V/Z6piW3rdG1EqZhiXj7sQO9M71mgrDbnVUwhBFbuRlVZdv0l/DB
HblbsF0HRHIpnclbrveuGnhAyaJlhjF62cWijK/o/dt0n8Z0w/OBE+ZM3fhNDXyVvJgJxHaAOtmN
ac7HC1RTj7Fmpn4hE/E+bYlB9Xt9iaKXmEtZr+Xf8BI75T7nVZg8AgIqDKLdZXQHKJDHkJR2ZcRq
/nqOW71877aIbqb85bcE7E3rFi0RmhPvPmBmMk/D7QZDi9z2EXo2Z5OV3zFmf0gkga4IwzyAhlrr
VhI9drbBAJw5uCy/TJdPYjHymFDs7ZSAw237uJ8+KXTf9KGdsRscF0CX7+rvSzC9gLy/KJ5v8jQB
oQBgAWSgLvQKv/8+c1r8Co5k5jKtqeI0cXO3QXma/OaWwBZhCrtswrrwA6Pa/6Pue2AsEL2l6LLH
FxJRtCJk+/+wewLpB8dP4UZY6VWk8Z7p1l2nuES/IUW5M/K0TQOhcyfpraOrqff8lLZBAZjA1uHL
6O7vf8QxyqhcYteE2esI8FKXJG124olyekF3oWth5iAgZyCgplCiQSIQWzbzKtfBZ6difs2IQ0ZQ
FtPoiRpFx3hjVG4KIANtr+JbLVCwVDHPmGSAqxWANS3NkOyWKq0xbvPEU/+I/Cx45mBoncsht4vP
ojTvubCBhg9XKaxYc3UxLgEaTU4uFCwDNZGzSzr4Eo1hwQbtaQthUiA+SIgym/F/2PYvQneHF8Jf
xDWB/lv6hiJzF9Ej85OHfqVieFr3SRm/6JgHgB7HwCvz5bFO6RX2CMcBJSVx/fBnTnLPi6lqrh/4
xMC6ygcDGmTRI2BwKHI0RHkJNnuXW0UKc7d/ZZH4+sb8X4Q7/tH+YCnQO7dAal7xguPrx+sM3djy
jTr9FQrgrwHq6WzrAd791tMqOP//YTEykWTW5cMQrr44qigPKXfgF2QXey2Ta8mQKrFPcQViDQ1+
Pi8U/oy9OlTJ36ebdMDLE1CLp114kh9z9K2IxeV4+XwCNSmfdgS0ipO3klpSHXh0RxrRrzOMvY+F
tcJrX70KcS3wmJe1kF8tE6TPjYch5r5sKQ9y3Z20i4VyoecXoE4e9MluVeBg/WUpgYyu3HediKru
6mZ/Px15FXK1zdHv3eHq16tq897IpLLdGmwghPpDxb790u7VALHNNBtArn1ZIzWjFrzVYR8pZagP
rXrBHiAAps4E88brSUYJFjDSdhiPIigDPddjLx/WMiIvvzRAdwS8QC23UD7R3C3FkFD/lIuYQ4Cb
p427HZ5/KlPNdnYC0wKMv0gUf/XGe9kW5YMtPpxGXfBPQHEjklhwNcX0PcIHWu+cs+M+MELffp5y
/FxeyQoef/yRtKMe7cnL6fBdrK9w489Vd+vF4jq8fvwtMO3QZc7xmJDZ3i2e6SlSynQQ6o9tQbyi
bj+Ay9RI+fI0LN0NpSO6Xjoabj5fB3M+XgOLZVqWFJ0fqJEsOe2sVb13YwxjSrQRgo/YG9lrFVj5
NQ049D2Wakuwto0UgvwM9EF38sFSt6aFIE0VonjrRPuj2/FnFHw/dfGljfVGcFxZ8T5g/JxSzfsb
k8urxlLrTD0oxbjSoFBcGv4/5aJGzo4qJS/q0IzXE7VksoObbDPyBAErEXpz0duIz0Uthzeqd6qU
zO20RS1qLpt3BMlger4LrWVMNA2xnLTk+pIBW0G9ldoD2JC0gOB86PjcRDoNeOiuQYEvDLFsR7yN
NOqUf6idMwmQpOqd/atCPlEX+foLbeIk1wtjLpTwPRUsU7/gHFgwtVLpNHo0FKV3x3bH8ARmNKu9
0H5Xmr1W+6iaam1PYq2SisOV4JJCM9KeRdAmmnQOxDi/MjO9Y8pBy91NmBH451ut+hf7wNcTSzFN
JAMbdSsQVygrz1OPE0hWnnMhCirdgthuQ9SThxkH0qYbpCNVFen7eHVlKA+QoJ/CmL7C41iSBhvL
OF0VLg5A7zBQOqoutM2kXqDvM30A7M3eZO5EN15c22OdvfDSBTCV6Vn3FKS/zvWL57jmLS62DAQD
zHQXN0IPPXEstxJxB2EYT6qwympSzbZN4B9WOEKSzJ9k4V6i6EKC0ea07sQltPNUVBMSfnh5g74J
F0AmZxv/CjPDXymoob5VzDuAXq5p9C6IH5i9kBa9cW4FL7c+rzytjLVweCEPm5cZF63DkSmhAskr
g/d4rfCCVLG9AG0o2LZ3G3tYWLwbpUws4b3DS/wVXJzw+xTZXHSFGQP2ftsu36wkPNIoaXP2X21L
SPpsR5JoQ32CCrq03aObP26AUsydjLFCSXycGrH4ekCrR6jq6kITwgPm30/gV5cZUnPyNDXZQBt6
AzaRnjBxVl98uj7IVsER4ee8iwgsJ1HG4OkVbHaHMjRTDr3CM1hZMZmnTvm635J9oMVgrb1vitzu
11llZs8CtZUBvxOw3nWBI7E81QpFgTPyv+ZhV1fPP343FCvp3vVIt7v9V8L/iFireXza3h3iO2Uv
MUJ0M1SYSr992fDK7mSldbkmrI8AomyXSzE97CQmUAd8KZD8WtjQ+xOKjERm9YKx0GVHp0Vi675S
J4uqjZvgztykc5L1NQnTiuuY5RlhIDYjzNmb2TlNjnRL8sYsiBZ9a3tdev2zatqMBdAu4bu3CUpC
hKVwiOO6F6x5JHZ4BiY/wWBnC5YZZ9HnAT3VvUMoqwYfskXrLQBPUkKr0U1ZAaZIbK6LUM2FeFyL
5SxV+Ib035QJuYr9v8UNCbXSTiT7RJnllJJ4Lqy5adVdAkltLOoPTnuwL/xgb+XEKSZ+lR1Eo2BB
KGzsvZ+00J9i5iRP2lHr+u4T1TOD9PrN9UdkGv1Ktx2PYt+WvShPfoSX2F1FfS/XRamk5EIbmUlt
/h0GWH9L9bEzqdvFjQdiMTAWkd8TQpZlNEKtff70zeKuK2yavfaLaGE58XBZ5U/5zZVuHj4YjyMS
1WuteUQ4qQIjsn3hGPH/qYS+kObfom+WSOcwyIPzOiFRFRAgwc52sNbCIasgleqNxo1EPEuDDlL1
/IGVMPblcxCYg+yAGlAK0AlwhDO3m3nSaFx1ICvWIQuVq1c/5J1m2MvpX5pdFoaq7wHnjBlvbQuN
L9N4Lm+oiWqdBPmeJh25fIFEwn05DNUTcv/UQeaa8+AjAa7uR17iq5q3+8OuPEx1tu0Cbse1K5NG
Ev77T8Ew0cfOrGk9n639fwLF9UYrO6rtoS8STNDIwvF0QEIBj6R+NL9njecdYOv84YavSeik7FiT
MCW+4UNiMwLwjSoyGp3f/GHCQcOs4KddJRh17W9hiPA2SizTawfBuFk2KAldcAQvVhHVYGJJr815
uSjxgM8tZGjrvN2ZAStSQS3oNNKuPxLj7MS9NRrf9bJ51Z4GXmGUKuuaGWz4Inx6gVlvEHggE8Rm
Vk1BnTAbjcw6rVnL3uPuOQW27UNjpGm1LDVavMF/AesxC5jQ59xHx8rAOfNNh4BsuEA6MXmz2eK2
nPNqiFpHH1JwxN9LQA5ULxUSfWaQQQsglwpKQ0huRlSwgw2yWvselXOPrVq2ql/9/L+3YIKVxh73
RosJ/E+lNUD8f4zGNb0/GieE37S1PJc7F6tDOxtyF1ILgNxL1WVKOu2xDZYqGHGHSKAwIqRKhYuD
839Ezew7N1SmKEaRRc6ZKugpvj3d04UhAOWHNB/ysSA8AtXfKhUKAVusHYEvPuj/n1WA0x3EICYJ
zqKr+wGIcrFp/fyNpD02V4E8jrGeCwtY0CM21nAsxbu4GyBNrzG+34JMvbIzBFka/QktV72wVpXO
7CodHlgFjP9CO6n1477+DB30peP7Rxl+3myWzCH0wR+fzxA6xe1Hj5RH+rDuvLYIDeWoIX0asdae
9LfHtZXIxFlx/IBLJNRsB66nP5drlmHIBIlWvlMSjc49VHvIjuWihcbBsJ6GSceVZ5fjALEeXXJ/
mQqg2KekkKgGlUB+ccp6+CbAlFB24BRQPQ/8Y/Bemld3xPTe6w1jgh2EXVadBDSZPjUFUZ9H40j+
A3/PRI1I22nAMjvsvdKCneEMYEcSBtyM/Iz3I0RNXrBDdmk8LxNlv/BKaH2qxWjAp5/fyfNivzNn
VlVUILfV/zm3Qg8IT08IYDSGxVHJGRlPa6UMIdViyl50d3Ep6cWDW9lVewqp754z/g1TA8j34ZN/
Qz96sHnGhcjULZaX5utO0VpOfG6mNsXSM8EdXQVxLO8cAOVofKQ7rOvEitq2tGGpm4A9ihawRYcn
7r7JFfWz8UJBmDWYC2jtkUrVj1eanaq+8LTIuGbk8lgzO8BNb+LvxoGrt6ZUmUGxRkpV03qgvcpB
nyJhevziYab2N+1hC3ZgnBkNdy/ugsZ4D5vub07dMR6+ibZjR3SgcMcXR0C7C2c1ZL1nBKQRsJ0w
V6Mb1Yt3A5B1aBAZPctagdNlQ0+pxfypH+BgDenoXK4bJdx0UPmBSHU8MirYyNSQTfRhQ4rVD4pX
t+GdIqrmDPCC5FivllCWiK8VdD6t4STWsiNZzisxqzVkSlY10xImkTqWXrWn6e97jq2ckf2iwx7s
lgHjfAeJnYajHUUA0g1//f4jLGvHxZ7LAhgis88b5btaQW2voKHlqdd9XnjvC1R8urUsvyD1+6L1
E1Kwuawydh9hMT65EbwSgOy7wQhp4OqO4KpywngGCXM+S7HX4TRnJWs4jvelMHbqVA6144m+Q59x
iZWsKjNVUCoSAh5Nj9Sq6ABHNp5FxqyV+8hvPLjSjiqbwaeUON8vS8xKrP+LEXUGjk25m7b7Hkhz
vK1nBa60H/trim72mJuJF3Jh4BTObyM9CoFeUKUZosrNtESTDwv03iMNBePe8jfoYeOHD5jZno5S
0K5+4jhEmX7EqQxj2hMJ+OM31Azje8ZqGvuLJqoKO0xoNgrQOTy5RfEwIXpLTwP/Tauip/28XgVw
KckloKt0QSEjR4pgLcXfMG7IAbvF3oal2c3/aAvn69oBqqwDO0EF0iP2RHVI2BeTAV7SksdnXUtx
Y7xiTxz8lIMKO15ofUcnNJBHEiXaJRzj8446mD1/ICVcuCsdqP1xSTxviG+arCQe/woZR7CXTQro
Uwz1ane3mhSuc03uF6E10l3CDU7IE9k6cVBLj7ecD2LDioQh+BNLZMKjCKA/svaGGhRLALMBXui8
oGiLRHG+4d9dL8n3dl0DGNiUhIq8Deg62lFA7upQ5K/sLuzbXDBrdqlqY+2m8OsMX+0m3Hyt6bk2
eHYNo12dqd/K+FeIjnAPCksBjjXSeM6fcewgbxdmFJPe/xVCwNggBEM/WACpXMcv6sEid8GBIF6I
MA/tJ6rdpEUkWiCrXp2vqBcxKaphWRAzJ3l5gxicQHPEXiiPNppatr5VrPbkc89+wfucN/MXrST9
59/65ecE0AK+0SmE/APQLBO1zCzvNzvHrgbObr7CsHF0plBsw4alUZ52aqWp2qdzNW2MsSKdc0p5
GzS+nlFvnKVwXBUJTOqoGbDyYChwd2XJyfYZs4UDupvy8nvB30GoeyQd14AI1NLiikhl1PKDQypX
WxLuoIzUky6DvicxN9X7lxKgrOPRclX/SaGDgS/0U0qt6VlvnALmz0eA42jiDpSRqssXmKCQjvpt
0gaqaB/PPUtXWJusdglGbUc5YyFB8gUWqZDI3Y3gqDafeiifJ01h2siTkJlCei+Owm6E5ayAwpTD
OcN9SToHmwWrHmOW5h8cXI4nEuXsU98Ts6JjIP4jFpmRCNJpDaGfiPdmdmMvqVS1BBqeraOaC+as
s4ROo8FbBcrnhuk9rQoY6uKBNwq2kQP8YQKVO089JfmlHEyiBql/0fwXnsb58fc7xJzP49BsbJYK
lY61Oy2eGeINKXYvJQUtnTZ81IJjGSI4SOVqZdzqVj9LjDuJXEPQBh4XDPLsFUr0/28wZYC6Wp/m
O4haWsp38EIava6Qw64gpIR3u01EVlaNQ3L9blml6QYcBEPL3kqJfeD3ScK81Y48tcVQsmBqEx8B
zBinZnk3LNIZaRBoLuW4tpno+Z3+ehbd9xQgtwgMx9Cd3ctuKWIEWd3uqFuRPKkXuLhCTH78VcW6
zPqNOyJQSdYXrXuW2s7lo7AjcAbba4VcWYx/eJRkDsp1zM0pEc89hdeIlyWAeiv/va1esaBiFLt2
itPoTsHtwMgrcLilzuW4YjV8wxNgDrEA5s//ptbmUsqddBpFX5WASuoXIwjDSD9n6FOAzJ/7+UeY
8/iMkHFJHhOlml17/NdpYcwentB0bOM7ywcEZ3OXP7Oqzg+Xoltzb3N8jZqq2jMBM747RpKVel8K
5BsvVtavCsD1LCljcBaHaklMNNPK1orbkuDGbNbPMJI1hKGgspbD/mrTdQYiMPIzVsofoIGdb2JL
Y0+DFEZ/MB5GrIRR0/6YteWRJ2yt70+HT66wvAEkb0uhbYuPUGf+nz77SC2LFt5YeTtQ/aImL/6e
QLilWvnj3r5vvhfq+hMesAcR3bW9pKNPr6C6ZhhRjnK2ZvV+TpiFlWKbQBxYTF4Y7FAZMAWBd+GT
FuXcqPYXJHrnocukTnQLYFr4MrQTamz2lSBZbDebhoafmhnG3KChnrpjeUGZ+qjCqJJWkogWEPqn
CUDMVrpojvoftBOWC/EWjbGDERms/UKQw3QeC5a9mlJgEmAJJ7YH+yntLy5PB6xkYYROiI21BmZk
zVHa5IXVm2A9J4bLXe8GhJA3hjlQZ078n+1LQDFA7OQMe4uttxA6eRRldIbOD80j0JrhSHOc2+gL
TPIZkRPcEyLqX5jThNhl5eZkx7r9bvKXG67MOeOkbpTBOuXFrshOH00jJ/V3BmnZrsR+OoHefzxf
6NH2ad1oiapLDK8Jv2JJXp04CqXdR/eICWbdwAINMHHpdXYBtFoD/jFqSFdvZkaI+/SuA2eNRmBU
OxZy1fZI8q0QYsDB23u2n6Up7dVUZjWLq+RmaeNDE3NpB1YJI/dqdcpLTGxVanie+cJeVPKG9+cG
M4nkPJl0PkPXCE+eYKiD1YBzI+OmlRKtN80ofVtLp43i6VJvZbw7oNbokD6vVAcDx6RiDvZoa0AG
4+Y8JfFB7Vr9HQbHM4uGPqda8APvVycceU0XtgWdSKe/4lScAZh8mQv1tTIMPcrBsciDlqdZCqzA
tyU0zpr6pBpAw/7teGbWJ052e+AtIvKnzltUo4hqfkLzJUf3xJxSUaLiUFbdNwXoLaYjgmfrTipc
7hRhHpONBNFlJeWzaD7S8KAtcGOBjMnyaRtRafGJ/lavluGFcSM5PD/KBJyOYsTcpgSakkf6+N/X
K3sNqgLIcYOqMGc2JS4kk1HkAVBw9219qWaafO65x9DLSA90c4rAWEJJgSObLTXv0/t2+ODrro7b
5Tp5eLXgrk/8/bO87+hQUVLJO5YRHPqHQCLbba0JMaqUxIgW3VMUTvXciwDRLtjbkSR+xh3ip/V4
oPGhJHSsrL7iNiAgPDylc1HvyTjfeY+DIKqYZLvGnPOCy+ugGfdvWz/H2Jqzu35vxBJ2NK0fbYxL
JKTiAxTkp8M5b2mbUvvpZAFN9SI5oEdzGlBm4RHIlKApihcaz+mQYnlVzuwSr6hMk6NakzVj+JZ0
hbExWxjg0WuB16ttp8z6gR6qKdSlnYKIowQT2TYVgP4reRGdO79tVHq7S2S3yOIEgSaWOZtWY92j
hySkjVwEkZ8gfnrae8S8wJNGGd/wXOj4APxctgiPUoaXdPPYELFfCpGTsNok0W0rMD33gp5hVC5I
ijYgMgThyYCIasckfS2Yzt1ddALnFxvSGI1T9a8pPrCS20qgPjN6ukndJNKVu5OiELDpNVsZfJeb
rS/ZgwGDtE1X0gdoLC8taXclGNuJMLHv4jJaV3x2BzK4gaK3NveX9+xykTLWEEHPbtWOfo0C455l
TliyyinpfGNEXBOrSMIOjbszsmkJjTs3V27QO55iZFSZ4/mpj7hzF4nRhmjOsGENuh4365ywVddG
zVJP7m1+cPtNsg/lRmr5wocXQatg7BluPkZ5e49xUTB6mXb+9gaO5vgtAFrffUaIHYTiDg9Pk237
huKUDKknzwc8Gci3TT1xW/pX9jcdoOO9UUYStMgPNcYdPXR++gx/WhKWxs3jmN7WFCAfPHERuMiL
uZ1indZATD0f4a7GmeVwFvHHYzJEJuPB2R90dMCcj4Xg8W4mBtEyy6FzGzXT83t8H7RWvP1wYi2e
zEM+Qc4cYmQ2CdxDxTTgUtXw3XVJhJjuxIz2oNVIwnILoto0qyIU6mm8b6e5RiS/1ADheoZ9xCZX
8fBXiSxYrwtQpBIu9f3XXG4oFhq70c+sNri0Qms9Z910P2mcVXAyJZB8eT9Y9ihqZSKXcNaTK1n0
idfZTjq6l16cPHn7WqpiXS2VSjkTSYUWXgyYnDAOAKYBLAXNcolYfArFawDSsFvEI6RilpSToyXL
oxi75NZfTmDhaJvj0SoCBND6bejlpKVA7uBmgKAMUwIt62I7UGrMul2BwR8SmaA14kJmY+4NEwBg
hPDvxxGhwPnXH8Vh4o7a28+RTFl+3ME1TystncC1AcvOXS+OzwM9wy1WNvg88f6GGDnGT4/zJyYV
QedCmSzXToXDJ/7v8S/+XjAO6eyJJONJHKMKp0VbpRauE2hXyWFTy88GFB3ML8xNcD+PwXvYifn5
T4eaYbnEaxt/+48SQFetG00yKozIiYswMEwdf7C07A/FtK62Nm4fQdTXW47YFuZ5T/zCWSN8e/mZ
yEFjjPwSBB0L2Uz2v1EuBHneX4Obub4Q0JiLh6UQ5HaANQ7sVad36OHYrOF2DKirNGlcQ+2mz+TJ
JkNJwA/OmPEPUqWp3Ci73v2WR+xE/cuBRHIQH9tHm4Yxr1rdXmScdU6OYln1K+mJZiGrihr9XcN5
uiLWp2R/+00asAoHt77F2SKHkU7hokTZ5Yiq2I1YavvZO22drZ5usAlvbWjz9qj4H9qGFS7sRw/c
gaqezY1mK4WRfnu1D2j1jh3nXgNrh/0IKdcp+DngsKQNFdcliIkejroXVN/qf6JbdboFQPfpPZQJ
u5XeX5ePDsu1jUevW9TLCeZC2+98uIDuqdfvMkVIiyTrMNdl81hQ2ndKlPoKOsJooOlOQ061Duz+
cswyGV0Mz50LAveACHCtRnCCdRaueckiWkWVZ/oK9zxOE+7fbhsmbt82RfPfTs2a7E1SEFNAnZTp
kETEH3XKdnlhXeABoTDt3GgapBzSkf/RsGqBEkAIhfprKh8cdT9E36dT9boBRZAQunlC0S1czHYK
/ZnRCQtKrbMS0V6RteCLI5LqPP3AWIWkZ2QZ6c0ZyHY7pMvAQQh2M21XiZoB51406/1bPDC///P1
pBXMV4EhZsebL69ig5jXwWQ5jHfrScIp9+W/6O7EbgFSWIp0pPvx4iaGfkD1PSDlgODIWxoob4Pe
/8VTja1xLAXS8BJAAFtmE6/kIm/r6qRdOTJN7XmCPQ3MHnNqvjGlupEqcrFvpmjkDOHNQrdGKZPw
iq+wuOc6fGtdUM9+MKeaTZNAQQSn8o9Fu/mLIGF94rzr5JMitVrftLlBdMAsmAPeXEZGOtqYS0nW
sIf3cOHjE1GvLikZBZq6Sxiw6iAn7OD8B3aQ3oy4MWVTg+E4SJegRJ29k92KDoC0Azo8E7sD5cfZ
KilopVhh+gChEuEp8nxda7kVpO1xSIHxXwsR266BroWnFHV+Oqr+2ZVONtxt0Xkz/DK8qrtVTh2D
YgjCD4L4EpWAm+TJ6tXsOm6ejqN2GvFjN23rzt4s45YEHPde4vEFNTlPNn06FbPjynJw8JXue9l3
viwCgXYl2TMujeyXrAHGvrwEkns8F9KSmN8QtlY6Hn4DqPcGws7V1Rjqgx/AyA1DW8PIJyFpGWVn
w0hHoZCKvPH4ejmS9ePYXc8Epl0JdyBfh5Ze9B+K3+bRKjkjf19Fo8qU8WOT6kwCiRK31w+Ei0hL
oGMCt0AE2FI28e6S1WxQOZckdtHv+gPux7dNmczfn7DbP8IYhA8Vz3z1rH3DaHUAQ42iUR/Lkw+q
iram4paLKq+pg2zd5aaHz/soYduu+YnYUIaISDC5SzaLI02QvdTPkMWLprtZOQlaitHXU9JU+BZA
sZJfTFLl+dUvgxK1ojrVAWiXVbwuDaezo8C4vBdBomsux88d84EzDjAnNtEegddq7sVtA9Znvy5h
db0k5RFBxMbZBqRsBih9hLn86afK/CwbzsD/TqGuxNInfCxSMAnwUPRs5J/mzkV9i378cBsK8LOz
uqu/j9NW8jKCeZomMR05ifDBANIxOq/8lSRvb4kPpgSi6U8JXW2C5PCXAKvqNRkR/HFoodOud1O7
V/AzxtGQu4PAVo2WwLEW7fKkYNvf5jywHD6y990EF+MY3Imdc26K0zOnnFyiEtPU+NlzP3sOXbwZ
0dfKsqn5RmNnIPqL3yGmkojaC82Vz5mvCua2Qxp4fBl47VoVF3Z9EyJyGHAY3krl0NsL6dmMRKyy
bNGDrLL3kwgSAPpsXjf5H1bXz0epOCfrFH1lkqunJkbfaTzm0YBoOcuTAOQ+kFwz1wGfrXYWMZCb
cDkxUQWFoNtQBmq/mA9UozFtRYS31CHy3fiWZwmQtsCZxXc8Cet5S6mxOKzT4F6F43q/XIdLZUvv
MvcdEzGNDqKp9/AGBD1aeZu95xrRFFDcMk1ZgyLs8/t5EFFUCHmfXxAjHgzoBQUMxMGXPHV3FFa2
Ph4/FmDHcDYkuzdMjhsZKGhdenSW4/xJwRw0fnM+wITufF6yBwi0HiDGdiPdHH/DhagpkXt6fyJH
90IrsCM40aqX7qfceoplFt1XQ5669RKDdBEICTelRjve6TZeDKywyl7RE1OIlqeBorgXpDRi1baH
LWKdIrdDCBTsZq6yTszhCoaF3bkYuICUlcWh3beiiptX7KxW9ndP3MpQ7cVArP0rm6tJ3o5L5cgu
uCfuOaVG/8RcP07pIonFvi5N3cpqTTdHeaxSaKLnYy5tssav4+JjN2us3Qn+uH8Tcy+OwLtVn0Vi
GLc/HeXXNI/Ygf9LbkUO5gtmUtQfXRFqDbRHqHYJszLhcdAWyWIUqLvozAHIsY0fO0+s8SMZPz1Z
lul6boCW/96+gRc+HJ0dm2CxgikjOISg2wsc2o3H6kbADRO0QaZNi2SXtj6gnNUssxFyOM/N441w
D/KdbeeF7xmBe3aQlQYIagkTtZUAXG1z/UAnmUrn4C5sLxRhIZbaHiCckMq65p2pvlmdCzfSn66A
adfwZCTz/th5akk3agiuHo3P1O3uxG3GmRNUIfJIYCeoncrO3H4LXP13qbIU8Kc05qVC7XRRxCcV
CP7t9mus/xK1BDBTVwlEV9Tw+fEo7CRtuD5nlli1UKR26Youqinx8RYu7SEzjAeAZoKU9+KM3oKY
KS2sx6in2xNV6q35ecYYGff72HjmG7S6IcNX2D1THgbEP1ls4yYOMfyLMIG6DBTA0ws6BbmMwcb7
NvE8TWUPZdE/piNZXmNvDoRpJAuADE39jtPg/zj8B4vmGT/nz7nwf5+9pq/8n1CaNtxr1VRjYOHw
pcrvW77rpb7R6bSXnCrE1dcwyY/lzFZlZa3OQ2KtSa4dBAJN+l8Qre/dVXwLrekebT1UDqb7H0Z8
1u/R3OZO5LdIqTVEZ2qhfkzSTb2lPZ8ny7n6CTmUfAK1yEhs9fKpDUmsIN6VKd3TddIwuXQYBtiv
q2uepUZWPNi/t3PbFyb0LGSo30iyrvb7Bx5KkaBGyBv0f5DWMXz2zCYUtBRhO1RLF3S3wNuZK1QJ
f0KUeCkgmAEIjvOt+xrqdEeD/KGPTUSniRM7O2mtmOPWFt38qlq2dfEvN96FpmLh/DDO2UxhQKMy
JavRH9n1zM0EwPC/W8ttbiI2S+GZkCpyLmuc3aFLFmmxclv5mVqq/GFxl31Qe40AbqJSTg/Rv5HS
Tv89iHntj51CCepwRuOSH3jz9d0gdg1jRmsyYXTnDEjElFbdgPRAVMBeyRhL6WzyBrvkMuDbL3J/
8RwPkrNhSDQJ6/+nhpdZc6LqfYI1+siUmYS1zIM3ZKLkUOIQs0VOnzatkndOJG5Ifg8ZybMxDLG5
abIacIWgY2vR+kVNG+h6jpDmMM5AsizIQsJLH8v9wn6ss+XejFz+4rgjRDmITlOoxbH5uotK3/9n
AYpFY+HR+mlGmFQ3DKnDrp0f8SISm0QlbGD6LzWAms1rm7i6xDZnrZlRDDjOWAiwzgpvEoIpuTUR
LBbGXIriJWJBceoyaRcETJFfIQx6VkzokPSnfwaWjEZYobcqYK39X0xM2SQbwRt/VCf66YDmZ5eJ
ETLwKAurVlH3zbMCJGHgLKnQm6ZjZqgIN6Zu5oK/OQCu8yDq3yXzNIljtJwcQ63VNY4+yWM8T50F
03mWEq3DOqWQq0yFhA5v4CYdU1W6IeIcVfb4WMzs2pNHHZ+kXLEMkCvQcjkdAJaMpA/BAs/QTKbl
x1oRdWdmnQmDk39PnEE0l/gijx0wJtuQHaA+b9o456mIruirxZbziz7/wq+GycmplvvLZgjSyRmc
NstKUmWSkuFVlZKuV+on8gxZam6Q+ie1sR8ErFsZ0PFAvnabdMYh+ywqWj76mjpXstksObbvfCGv
QgUXs4eYejSj2tASNX8ZlCsRQBx1s8jSXGB4ylj6GBm1/ITtyxhZr75s5cVMgfdGvCZNO3O0FW0O
uCdDiRfWlRpAzi+ntE+QCjmNg/WBVP6D4kDEO17GYQKp++BBq68d1rWCXdJBvXyLfuTEYRI2Cr9R
bSLG7mtgOLtnaVatKiIbVaV36CgPitl8t/uDVQEEVBXSRjDIpi/oTAHO3Ze7893LVoitz4tu1RLs
/LZk0tz+X9bL/HyZsQvSQjpXZ6xExKDFXZvFxi+3IxoKytGUnEdcOLlg35JLpN+NYZ63G9yK258i
H8eU0LXm9RQ0QoO6R9XQaY5hRHW4CUUwV9nm2C2lo1b3vGVTkKGbTvP4XczyJY5LGopR8kE+F1ar
NoUwpP27tVS/P5sGp2HCnsi7A+1SbuWOeV2iRRqFlcCwGgnhW7fUQgRKwJILN1d9+WBSwiOEmvEu
BuJ4BPrcA0AUBg0k7wusuwP6xVoa248/5VKFqcYa06eA2PzJXZFm2OLTe1LZ5jMWnFJKGYZCsX2H
EAb2qbbS4aPhwoqogAv/mMMXns+F9ClGEswkhN2qPleANs02dtXBiZVXUutP0N2K6bEyV1HCkQXk
tPGlCvYgou4rLiTFbl2YnsYnH1nCzRw1Aw60sF6+9etHNroQQKcXkTkyXsgsA1OWGvQI7s3Zwb7K
BKfALveTKXTXHCuKnk6IwaWX2+CatU/gBv7JPHVnvSugBAiYx8oc8qx7i34WoqEip9AYGXjFBoST
pPTOuwigZXKM1fXduWIU0pzPK+Nw0LbHDWyvkbLqt2u/f52PHxj5AW0Ponzol2wHTrhk2Bj5tosw
CdWD95NXEyNmSMNXl0EaWeG4iqKsG0FsRBGjseUdM7sOjBQIWaX33r5SdjmhNLYc6sax6d8MTGPj
30HjYiV0Yxu5Q+UwdLKY0go2pPajJNr9+YYBjhbKto3T88MuiiG6TIvYcUKO+qofkZVVzeFwhvI4
S4D/rrwFwafugO4pqf0h0AY2kSY/J2MJcBh580LXaEmZ0c9B45jhTwK4CtO9yr9DDwchDaYb/M3Y
W6V8OpZVhZQ5u8EUmPHExsB+R2dhZhBWZ3e6ZXY4ctxNtR/9M7gEr3cz+GZlG2i/tnm3HwwZO1oo
ExlIhv1ZvVPqP3L5N7SVZL0kxo90WOE7DvyLilQAfkRJYnNWJQGB8KLYSh314pcFR7yBrKJpfFEY
gjjjOK0CYXaU1ECn0Etl20dnu/OvX42aGtDPsNptIQzgw2+J5IUBYrMMF6dnOa7x1GIUoSo1eFiS
axnmF9UPNYBhBR9IgxIL3N7G87Fu4hWQJU05wAcDMhvt/Jh3iqjMm8IyMT0ZccGT56zCAnNU8/5r
q5SXTJNw0cf1yNsxmcGFDBoWqmcqclXG6uVoQaZSpOWJTB/VdUy+ZS5vmaTIKR9hjAlHe+l5m8s1
jRGQQaZaAkNOHbErePqGGfEBtnP/mo64rJx85w5pkt0RjeDLeQqEIBNBRsQokw7sPwDQ2F/Ej+if
LdfLHCgsVgj/hBUCLGHUL0+CIovkUDDQ54pGQGAoGLVmBLBLH07OzOHdj+ysh+z9dDhc36Cwn5q4
bATEzybdcNfQoPdgfDI4D15P0Dh8w/3GjA7/ABc7u7wm0cbvAVgcvn2ayF4m3Vnw6vA0a8UZbdqc
dWZA/V9D+3L2w3lqDfxIiPKJOYJUS+GrwOBs5HUtuCAjiX3Lm/8sIdbLg1EJ6dZFxJiT3PncgBK/
9P+/X9okVhf8hnzSrI3Wppi7mlrQKKL6rKsvnUfp4CibEw2JnFRZanK3YfxEXpySqlGEAQ5i7RP+
ZRe9lKDxY3XmSERt4rLfymbMMl9HA+FDmueKEYg8v6lYN94ktsrEufcx0GXdDRb6c4MPTgJLI8nW
3XM3CSjRpuHIsvlnXt4WPvS1FMAqimNpP6a9qXlvknpmXiIZiPH9QvkkcmWBQJmsYn8WGwScekmT
7hbkVZUuwdoBaMvrS2i1VLazy1wkA+LP33iHdAIFQ59oZmwt3bYVfybKqa5W8bq2WtyQhpcZSyXN
/7pf9iUyZG9WeAQOMV0AqmQJ9FyAnzS1zbIKVkeDipKHkXxRyfGuVMEUY2zgg0Rm942TJPtFlJj4
l0Ul2ZGbwSJwqq1OBQtcCyva/PVm2csox0cYDy/AHKxgRKH6wwTenbLq6uFZUR70RQGSVCLpogTv
/kYazIqjck5GzOWJg/7nZSbZ2cIRC4Yj7+rHNLLhRTiqNMj41OY/TjZIC8xaIuemMqsbOflPDsC9
SkaNEfhNXtJwRYUESKvVDTGc2FEVbkgYYH8LYAU1T9fn32aQbwK6SeLOBKTOmDRqfUcdv1QvCUvo
knFMl3ZGDC30mTKYSpTshePB3zmijH9BacK7tgVYzrp5yOrhy+vXleNcjaRGGbimmrEQ08UsZKc6
Vu+iS6K5EAAO7oK9b0CGdxua1LWteYsEp2pG5oeskCqawj6lasAh5nZCuZ1iVMqwmN86Ut6Lq0g7
WCXhILFDzx7lahr0pKoMXmzBe2Fl8Au5QrOtB9QzPYdeE/T5kG+nPJQvpqZ8KjXxOQeB/lLuRcLa
l0IrgYACslexUFJ14C9kAC/YdoV9DRHSETFQNz790LYk/PRYJ7TgnWU426bHoWL17VbLKvl380ML
aAFDuwSi8SMoNvs3+OgBf/BXFfHDf5ZC+n5Bv2wiYpxn/6TfPv51fOSVY5RaEsIk52RruqKnGA/S
y3yWDeD9rfMfj6uob2eo0V+XWah7TWq1TnWKVkOzrcykrkP4oCsSugTWxFd38mx7Rjw0H34w5V37
dMpvMK2WYHpoKLNGZe7I9GiMj2tlUCiw8Z4z7wtCshsb5Aqb2k3z94OqAyK83KTkbGMkZG2eWud/
ljn4WCIxnciod26AAf1NAWLQDkiAgrajagcehrAgKCMNT7N31I/gYn1J9iKWLkPGK5TS4FuomSZS
aJujivOE4v/1yANd/XI5CPoP/XBDiQuJrDD9Z+elOpsOy6zOORlrNI3RaIOBbByZizgh7njJ7+Zr
lm6Ydqg+5j8A+oyfmH7zoHROsBxrm3tOSCL3fuWgjdmN8hxW+2yB6Xe7xNXS1nedu8Mmbp9E4Dx9
uM6Ell/QeJmlNIFOWIhpTo2oH1HsFZOb9k7kW3g0ND1sDLoALRoKo8/a20WhjYtpX8xW8jeLHKwd
j6D49vchJYAZzpBCn801psLLACA4vbLPDqUyr2Z/XJKkRGHW1vaGsJq6QMtAvShp13LUTtRAQuGL
gIO9I+hR5jwJAG+fEeHW/Yia8aKzSjJN1jIOm2I2J1OXUNRQPZsVeHId/i0SzA8THdN5KwruuSrB
BN1NoN/M2yVEATF31y5mh0LX8Nb/kVOPnva7r+LaC1CWRKIoQT+ZgxjFJoR7VCRgyIHOWqhqovxj
pIZuY2Q6HRtmy5tU+yDYvJk6hC0kobLqpLzBkucCl20t8ZhB0tZ8xdAZ5WPCTsmWrN8gsX1B7Eb1
ll9t/qPBqxzUsYm9UdtBebRBxZhnbOp1yPdG83tl/Y3qHuTE+yJF1Cz7V9nkbagXqzobI2nha6Lh
uWrZoHvSiSkzJC6b7SYWB6CJq1pbeeAVRpisSO8peHLWntTFypz9uoxfJKsANQfpErMoxkHrQe0r
8yokwbTg6LtM1D6Fpag+XrMQbQgd1KjqhZcQRthmNcGmAizHSDfXLtwftqmvFoJienYEjMxtXxpV
c9O78wT79coeD6le4qOhFlmfcMozm48/tu0rDdU9kWrRgyvDcxc+llMxFNZBtRXzo1gmRwG8WI6u
VCSAQSwG+jvtFWko8PjdEG8Cuyy8E/78/TqYW7IGSNReCRHVlpwt0bRWH2k+djZEfWzDOVIMYeia
sTnKZbdpEmnqeUOXXlChSAwW4NkPPT0dDaEV4frRqYHvpPDub/AvhKsjjFMVwo1ZPZSR5gg4LTeO
DWFflTQ+HEnyr4X8nJyNMcfvtQCAH6ej/QIvUrCFjCp3ApoITfcl4Dh7MoQqTNRAuUv6cYmrGD4G
wvMon6LewKsbyfPIQieI5IWY/z//HMg2UWpqxswvEAX9LEVhtceDTHOP5174rE9rkvX4Mu3IMCvY
SZCGL89YWq8KT5WEb/F+VeJt0q+DrR4jASZiWv2nT4GSGVGUTLyrWvfMPql+ZClBrYDOSMrAKsPB
xTU/mfXQgO6ITGCQWmgn0RJhQ7A5tr8pw3u0qev3WIqB9wrJSDm3oqoOycpOKJ0hlZ12VFoaShD7
Qy+UVGW3x9p9IaL49+ZqFiwt/K/mWlJKIixKRaKuScTiFN//1vCbri6QhCzy4RIgQT4dUicYXa64
E0atZjba6qhIDbCGP5Yfx1FsZb7FmxwXt6I8N2XnNqFeAAH47M3pi2QcbRqwNKKOl1bxtur2S2PG
Q2+A3c+OZE/CqYbmV5Zm0XunvO23+lgJlqsh6Jhs+s42Hm5Dm4qrZL9+KhW2zFfr9HqH28CmSFnB
ysSU3GIglAxOBRePVaMDaPRh6Q3AaQF6O+gsSej7YwVUO2+1jwFeRwvW0eDmZ0TmBtv7H1UvzX6J
f0PVGWRKzHhZG3s7bcZuJmptL9BHvLu1jrcJbUP65athF5rdiD4CpZZQnTnjvdC9jK+d2TzzPiTf
DBidxGG/eROmvYffwCq6A4Ak8eldxXx0ulPnEFb86eefjeY9Os1tT+vq7rYo1NaPsQBwRADZanKJ
goNu45XJfnqU8fr9FXx+bEHBsuhrzXNvyibcQF0wFX6Hl//LYSMqTRIwtSiY92VPcvhxF2C1u2Hq
Uoau7Hb4tvyKTFKNZttRo3mf1I39UnrQmavBh0ELOXvjEPipZmlt9waDHHBlfJjuXPzX4kxfZiOY
jnfrcXLGCdw4grQeNkAZxGGngWFStinYrs7olcLM2X3o8bGbrNAgndgoXbc+HFmlHnUnFINDzlWJ
U6kQBF/yVpFt7MbWVv9BMG+hmpU3+ZbRAvo9fe0brz6x1ooPE3zJ0y9z6+2X1gwJ5l8l1bPolI7n
ydfBkS8zW+MSJRxeR3LVmENM+q+2Zyvlh1if7xKuGR/yasfEpLWEsL3s+0dcOERHvbP8PSNwuz65
PnG6dVQrBPhNJRlMjIyfZ6o1T2dj1WzHNoPbXo12z4ikgVvXn+2Zl496p/5nXuByWKLxMaY78nz+
yB7EUGA8tZdsyLa25Vrrpl6Co1Va3Gut7XgDS2nFdEshVI2se2V2ddMJEMJK9uN1PL/mv6PCZhZm
vNJ3Z6BfuMdHZaOxNlUJLVTpiSDV9Bh6VqAj+8950McEnz9b3Ny0hWxQKuUDz78iNfSu3DXQu5rm
cY0sEmuN0kWDd9+kENqsWF0/AxYx7VvfPcpDcewZHNTkku0GyMwHDYjmTev2MdtbfEALGgXivS2Z
hGVtIKF/5Lq2rXBJ8mZbMc9CN0Ir87JmNlA8iQ25jsHYWAMUt0qhWjN7jDYKhidZ4c15wvOyv7cJ
YSmKdnj9vCfmt9OLC1zDPAHce6IY+f4CErTbP3aB/hz3ycogFyLCEsjiYH7PTYNJymoPuhBiAMhK
ts81MLdhchV+pYEhoXtovO0jL+3JAGf9sVak0o5XcIOAWE9d6Tt3KMORJcIGaYO6GiUxmL3Lb+Ne
8kXdBlAqKRwA5JkjtcvyehXr+3fEYH/EKR9zRrR6Y03u187s0CuVQBTk8fsQjeLVu78BGSiAJz6U
bm/CMyKSrbeiws8Z6CCtoBcKT2iwNSVEL21Jss3RMwH7otTzEgl/Q9mtw2xYx3Opgd3bIFYkjiRi
Yi+z8217/VZpdP2ol+NdrBSv/UoIHJWUea0hGOLDXnf8UHCCgOEIJ5/kxUwMomxUwUoslDUvGMB/
c69rc5+XzuVrc6T9ukCCC4YNS6lNlGtvba8E1vw2RADxlVWybOGG2ntp3Qt6wfOpEts4ob6Y8FQQ
gpmybo7M7jxYtGGYCUJqyLpirPykehfB8HNqeUwt5O0uYeqVuMeXig4+1EQjuWOgVqResSGya405
cPY194/kyuox3ddfx1d1selU7r5YNtT/dO+ptqMUPu+pmgmyICAFwzPKkvuCpzrY2TlKWC8REWCc
eane7/gl8XBItuKb8PWpsr/AiXuHMV++YGSMRzD5IYwfmGRH1uPSHtmgKCkTEz1MmFgpQVTBLn10
eJ9Svj7onRV3uSkAIZxz8p17H5oUu4tY6+9RbxoJ+LRY/Vk7+irReFuxectbQMFFTgtzutYj9oH/
KgRzQ9p4Ow2Fat9XojFgZZBmzXf3VobJLSt4mTH1fGwkUYV1fy1o0cXRMaj+/1anY4uZ/5rLzTs1
/nOHfAurcO3NEpwXFBWBsPj1wPG2MpoEYRLJc598hjt14/VVIz9JuM1xPEq2CAbK3boWppOLrlWD
mCIVN4XVAgoGHxBca9Yyn77mNmSp73zP8giD0KtX4e/AxABiJEv9TWV+rXnx0Lm9wc1XGaurg+Rz
534JdHwbTl6x/gwn4+UjT4QBeEtPlNy3E0GaswLmq7Y14PAe+RA04utUIFZLrhMB2mkQsiYj5kTA
g+Gtu9roFYt1ieNGQYOSJ3QA2DcxdUk1mYoSCtKEdnEDPjfdXIRaMR/nJ3TSXH00ZEUu5CcK3FaG
T6/M3uVfdBWSI5O7LvMNSU0zLPvSgpJmat/ebb4NeI4YAQMUqPnLE7Fcwq+s095vASQHWO1wr/md
kDw3K7BJ1o/2JTFF6fc1O4szEHHVgF/8HkTWoqhp6JsYWiNluZkrO4NJNxcIuej5VCG51TuA4BpG
B/Sq4kN2BASfJSuZiJa5oDTb/PR0Sj390L3MDWQGbYvfTPo5/f39NFMPIwUqYbLBCTTB9kdba5JN
dGYqkYL0PHUIw9dyYWxrJN9Zp3fPU7bWQS/h1uVHBJc6vpvhx9TWyGEpJnITXdFYVJTp16nd9lVp
zqb376R9wwRklM2jL0H+ueV5BsEipZASKciW3ZA3VXZsCQASweQ22yYwUHs66SqJmec+IZykEpco
FcDLfxNy+W1GTmFqm8QX8+P5JyS9QnTW+ZNGcj97z8z1TvsvukvATRgPkqTKdfwy6knSqJJhcvFE
lfVbNIhDqM0jzeTfMlMQW5R/+dEg69uKLWe3E9toQNU5WIsAOAHz80bJkf93xr/Eo3tUZzuSHf4s
bhLF3mPyOUos4ZST5wTrMB1VF5fGFZrZroZW0sCnhWPOEERlx2Tk6IBk5YzPgkDZiHMWJReqETYL
eCMcGn8iqOYfrl+7I0dqMv4mXtQyf+AlAmJpY+hufadIgUK1+T0NdrPKDTgseprIREBhvea5F1/t
4J9X6rY3xCDWBaDuTnbCfGHTqVazIHbrNAM+ZBTuvteI5vFcDSCLg6W2N2svTG6pYQRj11AY3Xzl
9mIvYwGzoITUFAGDit1wqpxhNzzqG8tLv09ur7RvxmfEoG6OsoeQT2Gs65TNLY43zV5O0oZKCkdS
dQ9+iy4/c+MWhmFMX7yh9wYnA65xOHHiUWOCW3ht0X8xjsBWMSYhtWth7rNLyRclj3tjIwvKv9MG
RNrddr3zSUyM/EnxetIaQbEaw4LuRcYoLoV7J8yZpy0S5IHP6nBjkG1mCRjGl2TN3D32/d+BzGpC
EE8rcySaLHE9zr6ng5vABSqIFTLrQs1/Wlh8KLEtSJ0R5G+mOYXbaoGm7pseQNhGtAJdNsM8A8kf
l7r1rMS4AoRh1GSb86ONhVSyhcrixBPowdXWD6JQm6g6XUQL7KY3g0l1YYb0L2DUrbSVsDpgcicZ
6cwP+oFYzhYNAkvCmD+DY8UbK93bX0PG+9EG8XnUbrWqi3j5Q2lsew24WVDS1/oc/FFEGGXgAkKs
x4GdZTReTYF6cdMehAQgOyAZzV2gU1njHU3jHKY5XmZ+1yrGrfdbBhNE3mEFwl65RKljh/0LYkrV
ghzIo1i3BBWgeIJ0AjRb/BMGxJCpMY7ITCKP3Qu1Tp+dwedRsg19VNDr09eU9cjkn1QqGaOwK+e4
QOVqLheORk0Qg3Tl25ztHLQnvYnGgQ+JEBPDidrK09U8sb8akZzZCDe6j6YHPe0dJEuxokLswACB
WrOjGFnKpBrLA8AHCjXGodb/iW+xQkpiqgm4F+Cwpg8A3UvzJ4fCY6X17tOJXGLTQuZdJjUEeWqM
ZSDDf0CW7LnvroUUmeoVRBYraj+HqK8qtvG8/s7+5pZtz/p4vkCsKCGY/hij8yd9AutOeQE16xAG
XScaEzuIqsNyijiUNedGOTUiQ4rmTrZ4pFoZlqdV+ngM1ulFQVALxubCyi4oondWohKzWiEeEMIB
d5/gGQuSW9oInDmtoOxc96sPOq90i4NJvc6afe7KCUq51ooHucka2kcplB6wbBIr17VETUWoq7aL
7dowba89kOBjUn4jt9lQQusZGG4xZQsSKM/5bKo/lDBzYc+mPifA56lpEkluPnv/msjLLq3E99Cm
Ll1wpPm/OyFR9lmvJev46REvfD+NsOj/mgLKfz6g1ltJAOWlssrTiR1RmX8HXeazkCHkKbVG4Oed
ZMwRG/9WnmBWgXkVrZcOQmej8PaxpX1JmoUU+cu4c9UrgSSMtUeX/C4OXNNJUcqQVmXDyCq7Xjoz
QlgdgbZipMWCMUfCHRMvBZ4mYgrntKpige5p6kgaFwbOcETcru3kE8bjKG+wgdIKWyd04bpJbFJF
uMxmbziiKwtHgynK4w+3i1NUIxlYJXDAK31GYFOVGPV+LoZOQRvlORCYKscVd9viDHngVhTT1xNT
k8CSQwVluluj4kKqgZfZJRHmzF2RFMuodOV6oEF2Spx3vqC6I6LtBN+EO67P7GzIZwjdBHBMHxSQ
jJ4iN+xRUwKB7oJn8U1k+ReqPZW/vLY06HYrOuFcSmDk7QmO9+e4hu7y4AL4h4xhFtc+dOZwPJOv
HKCDtnQr+F0FtNBSGrbvnkFVKdUlmyoZPUICuUBChWJc8y53l36yqnMGUWlSKRqjIZKb4f0In8Vo
PeBNCxTFuv4DcjiEs+Lj0aj9EvVNLzMHLSlvBQZmNrIm15r8TAJoSaTjemsPf8tXEb6R4gA3OXeT
qp3rcO5mlihdRqjXKNGsmhfC02WUdmu3Ls5yoyEWLN9J/Dxl7kBgWbfnVlN7QcYGPvXcQTYx57GC
6jw+HqvGWG1rwQ1NJr+yi28zDsZUcJJItuSdYc0VZlOJCNA3wfooUpwmeHfWrdXIXKrpOBf7lROp
5AEO34ho+D/gDuoPSRPC9tYShwdoLDdbIVWIMo+8i76oa0oGYiaP3Qir+ai+7RQ98WQj10QVeGyU
s5QPDt4fax0UpBCBuOfDc3mhPrlhGhBAjfr7T531T4fpXiKusK65iJmmBmBRXit8WYFKEsa3qUZY
hri1ynjYjvtKMWzCRDAISOf/C1PVBZkKms5Vj5hDqVG9rWjsUkOXefCPCHlPtl9evCDp3/cxlpeY
mukWACkVyDoiIaQDWXFIrbig1Byaus5RHdXp6O0k0c/lmzmOvM7Cj8HlABeEHdorqkFcu218juRW
otJBqa5lmSEeknjEDademE20X5eb6e8GawO2Sa472yW5z3jX3BsHBL2x/3mXvSPI7r5D4B+HAHu4
dQstGfgaORnV7msvhuLE8biBmkFmKdvbCtWPmLRURBNXHXsvB6pV5XAs0gGdDzBWHeMU3R1/wBm+
W/+39apjj8YpJr3Jd1w9MyArUelopusubhlBB3u4LIdNaHZGgR4D3Dm1uhHWnmzDKvSNpgc413Do
UibD4WE8syvgcCsSrCYK04HcQq0khoKuzbpeKSlP8OQ1y08ysIBlqApMlijqFZpITDBvFzqAnMuA
9SMtLS1pyzEkMfM9uMIGThRadQvr6rGRZbJjTv1ASWA/3Kr7wqpplh1hkSVqzcq5iOlW7Sn4YkUU
kW65hBY7ipAYGjbNCCewRGXHt64WCrk3msLYrNlUG+Z5PFErl1J4dOSlze4JesLeVTWg7ZdWhID6
lR9XkS1Rk9hyJObWBWpJ4h3HaZ9tCcJPFsWRtK+WrR67D9RvI/vNKlGWLnmdAMnyJWubCyZhQosy
SKw93iK67P7ZKSlZGX22BvCugGLoJRH5PDcyQ6LoYytdLKEOUSJSMo4thA5Q5Pevzr3wwFwRHX8J
WDdSPKXUK5pTx5QfjFI2sPp1EZiRsyiBgkgp7QvGD6zqzF5juHXbuTSBlFVCm8W7ml7jiStDMsjJ
iW4Ulzmk8vFC9riSu+29DKRRg4/TQH0+NBVlDmUAaPCoSx3ya0ei+aMe/pgo/ChNDggdptTCekVn
DzxKkuESABIVo0pJwAsLKxUuU3Moge3HmpTIVmHb35GmFMyhZzgwFR+yWHUKjcu0wWU9MKNHH+eW
zBYIge1Aiph6pWOLmZbG0IrXD6Cz0OH5COcgakg7bdU5LliXF5c/j4oXAYm06EJN+zOlSnEEB12O
suLu4rUaDH6T7ehUbv2o4aLsBvkB6AyZq+wLMVtMHWgB6G3BbAsBax9bs1M3wrnUh+GKh8GrW+Up
rebBEeLLtkOpPYtJZI6Qivt/u3/RdvDgRukDzBHoecv6jk2Ahdl8HIMJ9VGe11ZhdSACSz9+yw7z
iiN/SsqDo/0cijjWvU77SWM9d9MewWNtjx2I8keh
`pragma protect end_protected
