// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Xtm1d3s5ylUZZq0L3sFgy75fX5qkL+pLxG3jN0jg7gfbu6UoKVEUVGixlhSfbQIPxJnE4WVZXzyi
ZZ8ygAmt/qAaV2R7FgE/IlVVLmTWrj+sF9Jx7NTNfOTX9PE5CKOgXGjQ56YyVuoY8qA7PRKaHV9i
5bjrQMGvdv2G1wo49XSNBisEyOlu0ARugKoH7Z+lLpjSoPSnOb0ljn/WvPI5AavbK7YlAErmpXmf
Me39z4PLsdfk4vi2PuKgpjJvTXNIsYJ7sipCScx+pB52sUIFw2qH5aV9f+3JbsQ1T973FLTG3he8
foWb8j7oVLgD8CJhygLRBqVjclaIyL6ENZySFw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24304)
Tx1JEhNfxENYQeIfF6GqF6A/mgVvuEujm3RZRUctP5LcJ9GxX6ikkXRyMrN6R2y3FUCx+qSRIb6N
+h30KP4UDcqMvMNAEZIXYPA1Yzwn3av9q85Zj/yJB3ZO7LBURRvP/POjOoLdLqX8uiksnXFnMG/d
Pg7K2yz1od7vo++dH3gbzg7TVrE28rxKkAyvP4XW2JPevK/S6/t01c7/5QJP8rrDwSLjNrOvHqbp
E4pokcRjhomGGIfEDvpUFhD8cMbeIGecSVsyVptc7ooYUmW1QFV475wW+7YCIJV7f5qMXaUGqxuY
3xyQSILHHKeO3hK2kY+5X8iAUezYoT9xAhKrESj4vDXu2GHCSAVFNqPFI1+E5lHbVGaG8Q6T7Aip
esy5FFzjKsZQzmNNAaeu+4z/LWGOEKtPWy+QZpgMv9ayOLh7MLRSLphqmnaV1y65PPIeQzENae4y
gF3oDeL69tz3iJmvn/h4HMPfOY5HUfqlbaDYE7YBOYkaXzcYrxyl50Afb0/7TWPWm3rOiNGJrnux
1Lu6YzlRoCmwS2P89CmcnKLEM+Xuxuunfe+s3fXhxLZktA27vURrH9p+zIJkohH+UYgmqhVROpbR
pzT3xkaewnq0q0rLtxctvpw9DInkmTNkl5jShreQ8A6QFjpemK00bQgR/fyeuxAHybZPQABj89ck
6DtlDi2BM7chyb104/w44AB08/9OJPv//3K2I/x3YxhtJxrtvzzMTKGNaEPh/e0DdUCaFtXganj3
0b2qlMoZuV/YaBjnVoFwuK9EJl4YSlSuY1JfM8xIFpQxgxycYhnSbGeDiDhrPpMso1GoUlheV6b6
40VPtgZG7Ed1syTm2z6i+yRbQnTOp7yWOGhewTbgT6AZGPASUJfiYEl5NebrMlUI6kN7tDdJPIq0
pejOvmCVrxiTh0uqlBDKATonAj5uzLtDzwRBHmqD7UfYYy1FNa3YvbOyS2GXM2CimnEJyniNywhz
SVjyEQjukGGsTfb3M3rRrG7oNyy+gdASPssn2bHMsIO5L40Wj8aPdseUdmPWkWWruK8AChZrHTOY
TO5/7od6R7GHF2uEhhg90I1ZHb10++Rh5fe1+pvyqGpWEdMIOk+6GFDs1i4JsvZfLQCO4aDD6MAp
dHLMpxSMvK9+ndDGdKoqHdEs5OILYhJ7JreYyWoMND56aZMVleXjPL2gPfIg7PMn/LSDnvSLxo1U
XGfgDVhN6y3OjiJaGdjgmqlN0tLD/Qq79AnCGeRsh30qC4ADp/rTeC4zg5q1VvKlM5952nWQ4Zfd
UOJg/nUZZcBn0rJfxFfFYiVzWkPUAEQJ0zk+sVw5Fqji6fz/4OTcnmpuLUMmdF0cLHF5MPLC4JbQ
IRWbLFuzovWFH1QZLqZhAAmjaVMJJaa+Pw+XFuFgJFwMAHt/xgtnpUz4AcQFamufxqV7aBhKYVKC
WV21d9qnWTubMNcd0/i50AabyBCKuTduZQeJaWHuII9PMtmVE2u/i2cZ3KXU07Dxx6xvEHTZK3J/
NUf670Hfi1k6p5LFPp2LwxeHpkrfh+gqW3hPl0tqOZA0+/SgKTbRS/L/mrymIlYvQVRwvvzwlAAo
TZWweaVCguG+H+LcAdxvRlP2mgli2WjwdMg+hUyJ+YqYD9yU+vZtZSCOM/F6nWi4Do974yfaBRXz
sOJoe4rJOC+4CAmu+sTwgVSYxxY8I0Nrn0mOQ/QijWXiFSVsorTxzCPsFWKo4Gqn9Xgc8V3p7Soi
XdMfdDrtYXn8WrzbQ4R2HvVBlAItI1KSYS0fie3Fovo05/b0xZlfwsQMHDBM0jEtGbd6BaYiknv9
e3F44rDDZCsqmFNkCXmn/W88irCo12IVKlyYpCS5huEPySY9iJwD+cnJb0wVzPt9c4mIchJkfo8W
0+7c2rQ2I+9j8ddxprkn+/ubo85FGTPzZkScWsCt4sTNsSCBy8sHUIU9ePCrc33oiIrj5lyMBCGR
ynr8NdONtqxWzHfVPsCqFOOXvVL06KzVXKpJR8vnuihBA/5baIwN/XCwLcxqE5BtN3E5NqoIAQoR
Pom0SUXZqK1sGCnonbPlLjoVs4HV4hF96mJUIjYSW0/C8jQ6baOb5qbiZ6A95cIUE7HufJYKCRQ/
pGKjPzfpBLYQq5VDQkPA5Ay/HbifmS8/2o/cht3XYm2Qee9kQEnilxnWnRidRT7IAkB7+VH9qNzn
EjEsDAsLdlI+1veYV3K2bbN9R2NRpk2hE5DLG9auYtLmmO9/TQNOq+nnefj0N0Ney8IjTbzGGG3s
cvJGhIrhL6y2SEpCsn29rw49GsRZztvff09Oued6Ygo3qcBLgeHFtRZtFvd4PJ/26mvtrXGn5lje
yyXeS8WqbZqeIoU4vEPT3Bk9eF7BBMT9N59DZ6/mkRMWcg9hsTNqyW6NKAnXT4h2w29z/4fxXH5y
szO0Edt1VzN2EiaMxEuBj2+RzWVtISJjSz/MMGgmxcZkxCtwJukV0QSmpbS/focBqd6cDj64cl8S
SZ2BAlPlWk46AzTwP7c8P2eJz8jJ73FQ/JD2dKsVFkVTqvz161lTsWkySihfSly9+tDccVlmrYBy
RhxZVJSAJ/AVpPFNLWHCysmR5WTj3B/VN0yIvVx6eYo8jW48XZ7j30s0hnUeIaR9LfBQuEKcT+ep
l1d4uPRF18yMGQzNnEHQtVJ6UjtNRXQq8uUtHXg+6dlRI+DZF3JhpP7z9zurNSBDZ3tOA/06l9qQ
gdV/9zJkH0NSGh1bGVf8RH1DJbKBzMJwNlsWuASpVTTsIr7SlsfwCKPHxfqjzQZLFb2ya3imNKdU
x8VyvlMpCpxE6BPGdXosaistopOLk/UFCrKbhJDV8hw1lFUH9aYzapgH2KjMFOYq+lrea0yZNXG+
UIARvYKHbCp9/DUidrep20kHhY14ZMcx6F63mKlf3weF8A5FdPfUVn7XJIQ0ta0mOvqPNfJISWIa
qMf2zeTSej/xv+Drz1R1p2E6uND0y6ZiHmmE/VP8eE3n3jNgtDuWKRagqchr2Pz0ujo7zuBi0feX
XBU3iyGlta/csxYuwH/zGkAxkjgGQCuvme6PsOt5bgwuJqMCzFPYDdZ/pgy17hwrFPhPY+Sumj0q
89wyOJgguTisQ1dUJRdLNXk7DVnJXBTZYLPqBqIGjE3vfxvv1XpFk9nOIBM+JhiRPMTzdaMjMyJL
NH8AnnfdTKy66w3TDSb3UzwbeN6qLnz+9rhzGwrJ4oAVn5zWlJuKXXIIZSw4w6oyfQSavXEkaaHQ
Oq+KwynUzfoUXRtoezZWIE4CHtGb8sjPEZ2SsZPeEgChWXL3mB08x0YwUKY72EKEX3K2JHlSvKvG
99kVdh8p4WyhKRffnJMpRQUJSPk7odTA05hpoRFfUvGpbZtft2Tkgo/nZmdhbCbeb+oAgd3R64fb
p6RhDsVmt+vOTxypsLGNPeTFX0QN0Rmp4CatLu10U3pa5pXmXYNFdhspEkQspqqSCg6pdLuicNTh
kc58rfJG00fhRi0OPBiHSe4CLat8UJOMSmsEaLe+gZV++cgJB/KlYZUczz4k0mDbcWC1N4q+BNO6
kuY07Xtoo0PnVCPztkIGRVZQMM7aGk+4MlxPFkHBfaCulEotoMrUvbhI9KEsBg5dwu2G+UGSSnu6
0IPQvtSVSX44CnsFq/CVSJTN8MCLB9VqCIDg2OpJbMHiAyjpynsWHF8mS5Ze9cQaCToejdjYoyqk
MBdPF6PizJayomcnJ1qiSu713oIDtnnKMpN4F+VPmhtsDoESHxfPBmlLX6jBjVw7E7t6vIuTUeh3
4B7qPRLdaF2/t4etAacArrhdafUXkaZkIcf/CNv7jWp1B1fPbyPk6L9mFfrD0Yo/SKtM6EYI2Ekr
j2Mc67A+kQhN09mkArqWHv9cz0bfF2VLARpkS6oc6ofwVq/lEBzNJMTuT00mR/BvsHDLchwn8tPY
uCIO1x99Iq93XUoV8rIrmFaAKZ8Lf5TqcEGKnGFBk4NbHQhIR2A67UfRpGg8wc1P7pXn7CxqyU9e
tTnk15Z85N0UbOsZBxIDceQd4o8l/YCynJ85n19VrwPshighphyFhHjRYKxN4awnhUz+HOH31aVb
ZjLFGFjAq1aihINUSqjTSOd/zlqhcMnWRVQRfTF6jFTGX0uqIC1UPYwsNe0PDz32OacbEaWko8cz
3u9N7SU4L9IXgDQUgjB+DIVOXn5FJ5JdJ9OLnVJVSwrb0QACNUg2GR2UNjYOca1iVHSX+5/4OCeb
gVM5YCm4OiPkE07CTBrwA/lOq0Hpi+66PJWkvAFVHbBF2E36mcUaWYlSEDeKN7vEbneb4t89yHSv
dM5B7WeOi77b1ojVq8po91gPUohEY7ttRenmcfoOzx1SpIDfXo9XNGxjzXn7PizlSr8PGl0034LC
aUbtHyFogDM+RdBUjQ3mPr07rUNd/IxHS5yn+t9//HHWza/mCTjaaspjHn1Y9Ksc39UzzokqLsar
07Dh7SKOWLO5A/rjsesE+K3RWqa7Mgf4Tqa/yGGSBki8sHm0HmYVXa3MGwBXzqgtz/HSXl/ynM+5
dSwfoepIY08JwtqxPItqc7M+r2s1FfJotVPIE3FXkSFX5XtNEEwC8awFFF7dB2faJ7uV5a24W15N
yJiIl+niuGx/4rNqqiijj70n9yonN5FiOc6TWZM/NWwZHlnT5iovVASidcxcHu4hGzLE8jyvKkOQ
aryfIiM/AIVyD+nKx2ttcnOBT4BFO0jT9DNlvauoh79kLYdq/JUWOVfPnIkp4huTy/uIlZToIEtg
sFJPOcjwghmTMCw/b7UxV0iXmUoceXFf1QLppHPbIvvQ7ekhNjHAkIh1r8frCp9jm436ty2JW9J4
Yt0qsnmrPYaubWsUWj6dxmqchaKFws+vr7kYbpONSQdoY0k8XN6/+1PQCdFH2dx1QBL5PoESI000
/Ls3I0pkujJR3QtMoxjb1F2G2o7dVEk6pA9+W8/WRW6IuYWEywQiPo+GL2p7IxQ18QZZZzi+/8OB
2TbBs9/slhS3rZsT3T2/sBYvG+NJQiW48miuisp4Qd7e3vWi0du34fpTPX/y4A9vfQrlRhdT0kid
s8xwMYhWpRrKO6M9B2oKHqlj8z4Y3Yrx0nUOlaVvI8wSIJBRKF1w/qHFfxamFy5hpWMeF05aysIk
vqqgCnIITQ30mc/7dzGEwljrG2PLo+NmaT8PX49VjGnWMdNn31wbuPSb3WEEAOnQbjC402hHTPj7
Zcrd//tRQr7OQux8dzTqwKGrc6GXBxE5LMrPA4PQeoJugFkGPy2cVjnaAMrR3CMLer3u/DRzK71K
u3I940n5u/2DXOnUZRl8McJGKowJmZAmrk9WwktyGhlLlcJbTmJtsISc18AwM6BG1kgP0bbAfs7C
z1fprp482w7wGKbA+cPRj5/MQOgfoDTQqNaiPB2U7r+tiQuImwZA9b7EmgrJ2eO+GQum8kjwFjUC
0XJ8HgaWzu5yS8Cjf8WxBLSQWLK8ARZW1l1xf24MwDvCREG2mFhJXaNaUbaQCmh0H72X9aL/zte+
1vA6wm+IhUypx3Zrf7lumWMUDRo6ze/fqx1wWTAi6uoM4/mkvtDDMJGMQlcFHBSrwMwc/nd9QSVj
GL8lqsTbszRUYhYITEioVGZ7ls68Us5yGGM+ss4T601MgnUhHIuUBLvqkxwpEwTeg5d44d/HJj+b
i/kvawa57bjNNd5q63sEocedKX5ZJGWmp6N8VEhTHZgkR4sOR+a0a7WugBCY0/YpfdjZNPxu8Skl
f0ychh4X9knDopwSi6B9zXQVHDBVSkS/imZgnMcB8PBOsVeargwJO+XIHZ75sXhlF4HUiI0JEi5p
ppXt21L9lBmYd2HhJAXWqGxHZ3EP4XzqsUjeExt8dW6KpHV0L5x64coaI1irr5VeVBlcW+bVr/Yq
Ywr3ZbaA13GnnksKHKXd9C/SE63Y1K38vU54puR14Cr8bRaFqB6kt96ZRvjBeIEkFF8Pe5XfwLYV
Dd1zGyYlsCrAn1sukBrSge11fB7Ev+VuyCGuvv9tAjOMJ5LvatytO0CpRhmiGp0JItYj6vBrd+KT
pQLEFNf4O2BX2EKbj19rmLLFCwPBC3HWGmCp6eps+31tXJEBGxGkKGVfiiAiG2aQOm9DehJ8IT2V
vOIOZczzjEuMKhRk2oisbqSZpkS791BY8Z5/Cs7pgAgsUV3cfHK5Vt4lau/SvhkCiHZLfxFZvbRx
J+WZe2X8128PtLYEjow51rbBS3aPDF4iDF+4bMb1LrpRcv/sOI9svEWCSxlj8Ux0iKP/+97vWkPp
TSSmGUvTlzGx6lQ1kVHGHyFNb2lyLNSwyNKJoEk2hRnVHrMqhe/BRiXABJk9gkJu5vTg8gmh4FJG
6+7/rwalx5W6Df0/P2VPMH5nB11LKl/W6geoinTdo07pU85cpS5e7ySPrtiUHyr7S2augvSugMaM
dDkewUwgda2D5SO6Y5GNT0qi4x65PWPHJDUsvUyWIiEo1MqOD1aLEEOfzUV4EJ68yrpHSN52YbF9
xMRzYH/+LXWacNzBXIYpE8d7WcSwdCdpS/th63WA3ffS/pQ5bbQXp+QdR7ppy8/7Qe2+fJ6Hwq/D
W6MNKvomV9NuYhTXuMwYC6lFpOCJyGYC5cFeKKaVAZu00lVhLwtk1E1Ya0cgeX61oRz+gqg7Pw0T
L8zOsNq4WkzIGop42AxkpQd67tCYzALSSBtYIeKt8VKBcj5sYY8iQFtCb6/2h8ywnnYFJ0jIPm7F
06A1Cc9dk5eOiyt/65SZZ4sC04SpKFGco2y/AcBjR0kv5Dd/Ss8QlgL7Nh2+RqtNANxgC8q0BaL5
lPdMFKyRAaD4KRxBLKHfLVGep0D8MwqzCKLAQYqPvSy77It0intC1VN5N2obRIN91h9xamxkSmbZ
8bKwqhL2YOdUOI7Ll8C50/nBEfIXkopfzClbkBOpxgGyObZF/RXMFwsWektrkBxyKUvi8Rh+3i+d
pnVgeQ11mMxN7zZmPbx4iN1Llnt2BCq5Q/Ty0di37RajW9JSz04gdkCEhZzpb8sz0xGl5jJOi+An
q/lq7ou44/g9XqSvQ/3Cce/coJpgRq13xFbaso4eS0Gaa8b3/5o8cYKAvAEvZ2KfUKBmrYdSJvEb
IuSSwGu2Zjj+26qPGKBLC9R1cBnJ/vkGbbVPHof+rGAYn6mUfAofMQ+Fl1mT8N9sK+n3Ahr562A5
jR8omuQh/MZprum7/CGu6PDI7Fbv3I+sdZbrY8o7jQkjxCPCyXfCkYG+AvV0w0+XXPfMMN3BKcAQ
GE2CVAu4aX9Or93GrYSEIZ9V6Pix/RKosR9HfcQ9CDV8buYNuNGQItgwEtH6/47qJJNOOtWj3VCR
AjO0vRhnOQUia8UVuwOEfWjCd/Mpx5j5uflPu7rr6wRfVIGevYWE0aN4nj80ZXgpEGyURMcKRJP9
jf9ajEJXYyBjKJeP1pwBn0DtQ6j96BZPx4oDf14qobrBgtRT9EdkwqHGQ68DF0AnW9Jdp4dFiZuB
2GMi4bhQV10Ujx/26QpoxIYutOSTIiwMvUd2oCFOLZAnt/rkCD9ZwrHcLF5l5NXRcKpiJJTyb9KJ
+gPDiXmNBoz5kuKvpTU3fDBluBrxPn0vUKtGw0Ae9QB+s0op4+/K20uR2f1/Ia7+WUTHKXY8jEcg
/kXFrCYFfXgz1MQ04j+MdYBKD92BGFJv84Ip3SEnATreolo1VUgoHvxKlnPDp7NZ9OeDxUsjgyVD
T/XvqqJacyEswIbUDC+CsQnENr5HbNSxmJVeVR45IJrayXzs9aEk57o/HQbSGVa/iPgqnuMVkWFH
N68NVeWlOT1fzZzta6hfG0fLrTlyiZtxV5sH8x/kB+ANOIlX5dd3HWOVs1BOZodj295PvPg/8ThJ
7gguwrP1pGBLsOD/VbXjwMa8MHWdDteco+5KjNrGh5QX9yjoGJxWBFzE/GW1NuuAiY2kfrl6bO50
4ocUN1qh9OZg0/9KSmBbZGbJ/n9atbFSoRnWV65g7sqlyQnJef/Lc5HLVniwKf7g8XErEJBTk4uo
HjZfSBs81YjBrcqQMaor1Ym0CnjDe9OXsqEyEvdiOLwUufeOFh18aK72Yh22LGYbmF7WxYzT8RrL
cmnz/XHMchS7212CEwQ7c6nfxKI7lDV2mn1JbuVs4SIfztxRmNL979T5ynZi6RQ6neJxexh7YUe1
QYuSdIaIIPd35IQvkpu/4V6vYxR7lOVLYXh9sGLjHt41j7U+zEwkpe3gm9jGcWpP4QfgGuJsbVKM
R4t4tqbDHOC4z+JDE1G/j/PwTtnc+LVJ9iXk6/tRxJ31kvRl6aWCoopInZaJZpNF4Ri1g0t9Dr5Q
eNMI6OjJ8TSRIgYrLBBYkweACBMuyZa0glhPC+kE/w855FZirNh9x91LJdYMOVpmNNEceaxsYLAl
kiDFj7Zc+/31TbicRt9sHymvoxJ9CgXpf2Aa3pgPJZsLoS8LQeQfKRxJh/KRDVEZvqDF/JOJB/4P
lCwJJcNuOaEgXsuDJ31dU0Tge6kAaevnuCMo1qlu1AqHi06iFkZKbLIyA9Vai7go5gVFDPDOZWtO
KRX5xs3Zq6FKbFD4mcc7YG8yYEIXhQRdT+Y+QHj5wDD8FZMBo+jEIUBLNJXmXtIE7ldV9Omyk/tb
9d6Kxpjurb5DhVr65aYpPM5OkYWg/n4UsX9k6pTE4YxMVSYHowukM3ITIH4E1KsT47jnrleQR0Nj
G+J9ZGlWjmGuZcVk1xXnq9EspRq2qvJzabRKGovO32Zt7pSQrRy0iImcsQwCmGWxxW5y3xl1CIaO
Huv5uOkA5vQWZT9pevs1TgF7i+sZsMadNiLSmE7vW0JqKU35mK9q9fH9/g5OtzN24oU4kCFo5jDJ
XXwTDIs6LTtURikwbphcPABUdq92EoBoT0PPgMysDl5n7EKncNRS/fiFUZbYfamS76JVwHl+lB8M
A1Rl0+/6JrwG6mtC4P1mpDqhso5fgqh35mdCKl3jWrwrLb44WpVLAxJgz7/vzrnXEycI1JFR64Ng
pVmObgqFARf6UV6cFx6M2+zovqyeehgjX7HptdtQO8oqocvXNDOJFCbVWxbKFm+/zlgg4AJ7Ge+6
jjaXFlup5EJAhhtyzoQSDK4KhIMk7HeaQViGdEMJpeto0a4wMZeIZtYoyL6Ci6FBvbuMcowTyUkc
tGByfP/7frkufM+g5jUjgNP8Xn5IYd999aFliKmWhjgzTHYNSHPKY1k+PCmJ0dqf4wUfcLn6dMvv
2RgkLPABcjfa4T9Seap9DRWSIQXJdyBLRjE1MT7+JBSC7PilIpRqesG+BeS5hCNPKt7Vp51M1HG3
yPhLuE5PeEMFKBEe8qqyavcQOhw09HFV9qBeW2xd0yDaC+57kxEqXELIOBmyvZwb+E/J7vkFyeDY
LGpoaxXmNW2YDYryCrzUMsKcL0tqCvTx4qZbwTNTd/ULoutsQRiYUaxVsCkZLvJuZuL8W/YgiENI
fZIS+jXbRDe83kjMfRBdfZYxw9yf1ZrwNTZ+6zyN76BOH4NWIvKwg8zi3EJ+tdt50G9mONtUs1xr
rMf7AJoxoFJn0TvuJGyu3bWhqwIQrXVox/M1bOlwUZqMCxAosUnu9z2oS9s3DPnXqSrAScPMiP51
7F99X5uueilvGtPcovgaMcOkfpMs8eXRo4g70/3CeoKglHNDDoD36Zu1HtZUtrI11QBq4jxCchne
YsSgxB2VjteHomBzgx4mkvHU3tVeM7GLTN/WtPNt/Jt9+qlj0PT5AETvhJlHQk/VXw8Z2WeHp8wo
4hDciwuXJYAmBSgsCBn3ddhyqP4kOWinIIvK6OBJAgpogj1Pu3J1Q3LPuIXkNV/4HayLLMDDBOIX
qEztovKfOPjIQenCEiu/tOPecG6HAvYw+95U3/tl5zIYW60+oFK7IKqsh6U40E/n7o/GaiGJ5Hpz
CiFBvtvSfveaJqNwDwJ3/jFdiynqW3FMAPLr3GY6UdSCgEw3ZL8YstrrQM0h4X57N8MBHk2/zXmu
c6P5y+qG/RvXCL1MfbKEB/qbnX6DwNMLcjc3FPkt7MdOOGiu/MEHKibryk7QdD+X4qK/HMcx33Oo
qJAgTiBpuuViMBrlnpDWNiu2UIVSHCaynGAQPVUciL5RWYi647o9LBI/iRi3EEP3I6bUVQ5Kg1Cs
0qZjE23HQkRfuT8nG5UyPYPoLS8fi0EWYwtY8VLceQPybfgvh13IHyAQjhc2Y1O2ALILCHc3jGR3
rWDubKGvqMFhEgOuPM5ypx5mClfwO44177x9AKLw0ChvyCFy1X8o4PP/HEINfxR/vED1mssNdbCe
sGqqdPApslaee9haDmSbLhpOkxJ7RlU/YUoqeK61VQR/9IIca0ToUdkdAIzGGxjZmcgeYJw0jOwj
Hum5ez0R+Qd8iUgbGGSd0mSv7csNfKRjJVOgB3T+l+bhIVfbz1a5sJaJLOz3AeiP9nj3CqgDHnEK
jUorHg2CeMgpOu62ZHKpNU4q5iNtjNKMHSmpuQqbLIeTmZjnau5UVWtT2Y+WU0F+jL993R4eerO2
okLdmCHfa5uHSnf0KV3pYqVloZrdUSGO+P/cHz1BI2cy2P2L6TxnnENpsz/n4fsdKl2O/qgib9bb
T/LjPfiq2H3oXzUFQeUUTcwFhi8NelTu9uzqWHxwaSjY+B/uZsXOr1WnxFLveIxAc/PTbP9ZQefd
JhUNbHPMc/Io0JeNPH40qvDeKvAnrfng9Qce/hueV0nZM5fx434cInI4AT9Wq3p5kFYTAV7sUUHu
KViHfZelR2nqOxa0octhGnoQ5CR2y0kfnL19dMW8vKHaX2Fpj6KjNjJfUCmL6cUsnCmFPQ2Pt+XB
kycpz3f9L6lkXfSKp4+gPUL1cg573cKtpESxdn+e0+L+yYRHTErYAZIy76fwJ3Spjg7tQpLhgZZO
rdpe/bbqFBk8tNK8fSL9Y3mFtQgPCvusRpWnavhW+w8bIEtAcvuw1OSM/e3JQun9cULkS8qoSU38
L7th1RyOVLZE2k5tJOvYBg4rThl2GZ0k6++OAA5A7Z9F5zQFYBVy/pDUaXutA9hv+wFk3TbNvcIQ
Z5JD3FIiSqnpVn7wqyYGUvAIIYmilVEYNUPTfpT16xZSrvgDMHsAIOPDpjj6cVLPtrb95qb1ipMz
jOd9rARl64+Hn2FArvfN/ZbZIMJwVrNDJvray2+zXvCU3h0EIZkK3Sx7LKT1JRocAt6GHbIw1fWR
nrcawl30Db0zKnE2LhN/aNQ8i12XqIHpA4T8Kw3A8NAV3rEqcK3zUSeX8mU/hS8yNX7sKl3xBAOR
q8OoDP4minFja4F/Zj7ParPSu+QFuuKXNkcHen+J7lwxOKshJFjY3YgNNeFZI0sFZ4oKfbLx5z2I
G+hOQrS0AokKJQ9Sh7OmoxoR5bIs4OPOXHL7rUg0oZaeaPkxki5F8rWi4T1I2lYVqfaaAs+lTZGj
x6VxgcUUHVw3+LFBhD/8NXb6KRnFNlWu/JFUJWUzFDQp4HinF4NFgy4d9udwo7CihdcuUa2F/Ith
DjMcl/nd/K02zzTloSQpQsPmwWeGYWsfqj3pm/i8YoYRMRBgi4CGYJ3ygmHGpnnZwqZCS5MvzJ/w
qmLHFP2ehCcFWXWRREcZxdXPy79l9vJTno8+hFpfiMM8wmEpunYS6I6/nEUoKXBIYsW5pdjXTgo2
egK1V2XMzypomLb1QBIXIZOhQErdwCznwpUx++tCMzMOB75tw1Ejs9ao3Rvv6t70Y9VJGgl9I1NZ
j+e7sne0a6Oh3HaAtveB0U/ZN9Qi8yjzFoFh5qG3J9VFA4A3DHiAPn8AnpDoy9Fel34ZU9XPf0xY
1DNm8ZscAy06CNlDP1oBTd8IYug1FnrcBfpCYkRVbTe2sD/a0HjOKpRFwaN7DSsujRTv6WWnhM5C
m87471cijWk4EqclbMlGv0ez7aqz+mecNBMknPjGN5iKAWTww7/LEdfYc8d5toqRGCfJSNlJ1ZC8
yY7m7MYhc6QFoK5aJ+yOhAX/eXBTo90/P1nudY/YLkJrBpBa2J00QrfA/FY0P5aOhtjXIi2xTNzb
sSGv4xMIU4Op/QQldpVeZ1fbIJ6/XUrjQyMXHajeAvelA2id7AKLPVivcdVu/rjRsKrIgWCKJbfP
1sQQSd2JsYTwKT2D2UoTLxrD0sPAy994fuJhqF+fiHZoW90Yz2XX2krVqmCzy0cj1JcgAHZ9yq0E
xw25hqjYUA3lXHOB+CAiKLQGFgFYwyd2gUy2sWRGYYEHQioPv97y5LYFppXaqNJcmxnJmUw+x+Z7
iPcsx25FGY7j1q8z6yXb9n3XLD85vMU9+vvGw0R37bOjz5DscEZ6Cp9z84XO8oPB5notc0gQDyVm
vNUZwQnP65YXPE8p0nYpWjkaoBzX5LONBkUp5l1KXNLCz1q4wv8F1F1CDnAru+pls1S4E/7m2Wuk
x86G1ZIGNMD57Xc75hpJVH3hsYognIJKmnJTDE9XOceQnWsZAyzIlj2eFSRzgm3D6W+7iZw7c0ch
IJRcFzbncPTNU2l94HAmT8RYAezgMuga8Y2PwSKbQEbHkp3AFjDwe4PYWW3DYgGcqOlc7N//Po0Z
jDukGEZr7szXrDmwJ2uFmZQKkbHhTudMiZBIDQ4d8vzq7zmKPPDnKGbJlJHeZkmT4xytEcMTNvHy
8AgQbSgkRiKtwxzSpZpZ1tyDs+myHMc36HUV86KTOvQxqnmcB4b+1lqWUU8P1aKMorw6sKxaK6XO
9AivQ0GVa45cp1uWdG8hiY9I3Tw8wOZiMotgj+a6H6t9WiFO48Yw+tu01LboGWBKLiavEcOFoiRw
F/JYwddImao/EQD4OTmLGZufyT7xznYVssZktAql7xHwojQynMXaeDEZE2zlVzgKkTFZNpN1PD2w
gsj0wB6kdEzesn+1s/SRWLVc1Ey0ueKlZwiSbpml6d+D1q5j4cOgRzk3u9evZCtWoFrw4ez0n+1m
Qg00cVJkQkENSkxfqWSBO6qUXNPW6GJ3dqL5rQFfbnefaEq3z6lZeUbbTiescdZErcoBuiBIbRUw
LGrVkNWFSeqYcIPvuczgzcRGO/izCDOhY/llRnrlA82aIWdbmDHOMXKd/PdhAjnMIkit7zSJJ0vT
hq4PYpvr5sEKOylJ9qFrX6pdPDHZfUeQjN6TZx3DjXMQjX7hlPJPPfZORiar4UFF3N851DmSBMip
t7lY+aH4MABxjWJZLQ2JBW05GhS1MV5KpHJHHjdpiNCGyL4LvqsINxk03JTgEQYyDsJv6IumBSKy
wtS2uM3qTtEZ1ZOn4kmVLb0pl+0YdWc0daoBP5h+Jo+PO8V4UvjxL97f0DGWH1Ox102KFRjUymBA
eevaLwkJ41qAJb2oALQm4Dq/XeHWNVEj9zwKZXK3r8vPCcYe8XXkgnS0qVjgtKDvVQ73eOaAd7FP
plbQ2QlQGswrPaazu7JCnI1rtX584P5p83P81DO3aLFLP9AxoVi554mjp2HbNxteODVGoWapv/i+
fZRVHWlb0J2THnJy+Jc2VqmSdVHD4yAb8rbiIbR4HQh8Zlce8BdosZA5XgQc2TNkdxYVMwj+tDGK
RgffHHBVvl0otFFuwUdKxzUsPSCs4S/i/gzKpPO/sbMSMPTNAPbJj3AoE9ooEtCNMvpu4jitOHJp
NxvstbeRTsP/0H4BDK8JzCWe6yABUmxxmhOVKl30nKOejPnyz9kKVXJ+EG0X1f0OAOEha4vkWfec
Sg3RzRoOOIJjLTPi583jWf6bdWGY+WIPlCCQ1QFAUQKWOtKuaGFiZWfDsd1vKnPSTCrsPzZCWDR+
UPFkTOdIgoqBIe0L/dsMP2TtVNQzVPqSWPw7jL1UJPc5hZx7WG2USIw+n9PBR6N1P0BwBB+xBI8f
TLcANbgcbMbRWp86Ig85J0gJFZeXKbPkpn+4j/wGqNjveTtX+liic305hZJUKVrYrvAeFMBaO+Kt
dBpJB8pCejbvyOibJvtH8ZChqjZ/VnC6Q8F9bd9/9vFHx7jJKHWsKbNDyCoNQ9AMRttC8dooyn/u
mT2kuD8UAgY7uBO5D+xul8TgPGXYaABgPAEUV1jfkRVwQ+k4ID94YoIbX4BJILrZq2A781lNAjf1
y6vxdz1qGOmI+Zgwtg6dL3Kb3Evr6AsrbpU03MzC3rG+BY2n9v9IvVteYmwHA0nxQuSZwJtehOQY
/lLkscsrM5Yo5P/3Q8FhHRCU3eMXTTtNGC2CKJ9VNlC8dd/2ZC6y45d8PHrTb3U4L++Dt7505M9O
+l4mtlBANHqtgFEe7/ieg1xhJO24/SeL9asrK2pAV+LQA1IDx2bPuJVts/+qWKIMqK00Oyo96764
4E7gvR9btvTzR1lgcH44nV+jANfExhwRCNui3eJsksflhfX6pyc+ztmu31AuFcIFhkr8YvaqcdI3
lU5OWCQDlfbQL+Pu7785243SEUT4ODGMTLuqwVm+L16xSGT9wGes7nHzBCnpV61YipO1KvcJD0+H
5kCmtCp/OoH/UtPfi4/g0xWEp/64qt5p1VVYP1BEJKRH0t3dV3gybgDdnJuG82UbwNWHZrbqFs30
uJUq9NfSAGFZmn/KjH/Q9r72JShNAFJXQGsnHkXUYA95A2+41CRHQwvTSeNDtp29Aippv2flssFp
T/chCxzqX9RinwClKrcPNjvfARgWuYmgasFRFnDrI7SB6mEPf1ba8+leE2hUD9b5jdrATAgEkAnM
M6/onGV7Rhzmc4Opo2j4Zl0LhOWO5aQG4UQTnImOEbFEU8C/KLvrxrSCViNx49mi511IiNJz8H0O
ObvR4C2S1rqlFOghg/Fq8yBbABekEF3/ptTOtNxzAiZo+rVSIXgy6avOpreq8yG0o4LtUXX2B69+
QFcoiW/SEZCcbEMfSg6hcrLla3r/tpliIxMYwYSBUqLT7LztoYXPy27F6sn435fNtvnm7zH0nn6s
Z3/paW9b98WgoYsFiGoCfatdVygnJVb1gNCKYlnjE/q9pHCsOey5WTS+MqKJjdnDZO8n+8JTnHg0
ffPQNsC9kaA4TQVEcOHV+9/GHTQfQRCkCtvd4eW/5XgCjCoomWFkdH/xHwoKIdkj7GcogbMJL9qH
80AXR5vqsBWFJfONV1ZwiFs3QHW+7JCPI50TQ3hw+7Crzs1v/QtKNcwvHnczul55OrqiHxK4sMX1
aF/q8ob1xbx42g/ngyLdAJDtaYVVHtaoaFmEcdVffGZW/r3AssHcfS3eQvt0k7A6bmdONA5hCpgU
DV+LjRIkunSYNNZMNobVJP9CYzY5mHQEM1gjmt5JLHLXkBmHIpIOdk7cuQAu4mGbDufF4QkgMfXv
tUyJtqDdgIoN7eE79xY0ecTMZ0sn/NPa0xgn0qcX9WvjQLk7heHQUrQ6G4Hf9gTYkxubkTQv9UbX
/ML6Slcu2MwK57HmKB8ycT7wDTSWf3slqIAa7E5A2Eu13CuCwtRpvYMxMaYpXR2+0ltVweceDN/b
MTkzKBMiCoW6TRXQOg36HBVgC/3ExZG7j44pJzvYgxBPt9UD0RZ8Muyau5QrPcUqjsHMOIl2rf7w
PK/P/tvvlVqmScAfuSSHy1LDg9DKurhUYjAwJZJhI8SfZlxUD8pkeI7RPe0qDRaOSxEXuQQEX8SR
pxySbP+lI+UF+8YXBfMqFmtmxPOzZhhodg+t5gF7GfTJrLJ2kEyLHmRBC4JoW98MItPlLg9sS/31
OfLwLA1zzLjIIJzo5hiDFBnAKoCey6gMJBc3ba81KEY/EhHHY8Ek7mswVfRvYywjKK+JUz/u0c6p
Bk+guBLRvZgGkqntgfkExXboNbEbY+0rq1rgTsb9Ybas2Yn8wroBkGRIXd9RzL3rC4YKCUbAQlvP
RF8ZMwqhWF6BGcXCJOhbrgP8BEDMBVMyDzX3aRyIk0YzKHDHDnatamU2AJgayueCnmnfyWIc/xMI
+p08e5ewt02FIoFEojxKIdrcUVvfwCu8zrGLoQ+Lt+KB3Fnv7SBn+QLT/3fm/kjFdUQrYH1+3Il8
GRyk+wZ11Jx2cWnv9B6Yt7t3ynXgaro5DIsOCkthulXqujYVy020lMQyGTrmOZpyH5bkgr0vOTm3
NVrqBpdWp58XXi2e5JLVJYgj0jTA/cYpDP/dKp4MXMVAv9MImNSINnp4sSAW8QVyJ0/npvRaWMnd
jQfrb/jDK9Y2WcNC3H8YGu3IopW2y1raQ2gcHQd3cX/NCFRJomDsmB0gNmvOvWBdRjbW82x6lBNE
+qKIyPhjUBGxG36Kj46oEgm3e4gC2EU63ekpzRAiFVVlSBChzPzNM3rw5iwOddtUTdBazZS6CtO2
+EvIWakQixmG/EzTCBTkiUWVodI4fHQIrTKpb3qJzKX/yUmug4w74Fl5yKiymmvz34ROmRMEkh0e
hnv1w19+cIwTobOk6t19D/tJVmU5ZYxzCgd11Z0SK1i9i4uGnXGGr026x+QLO06Nr6Vy+VYwmXPL
5NX2cesbLFdOlbsK6hRNptX/I5Hn6OujMRUk2QGEylkn/TELrIGhHh9K/8U60MGMs8VlTqy4DO9t
1MrP3c0WO0zy5ZZ9CAVmVsmb4FpvOGMR33rowG+5ppUESWbVRAfiHv2aHsFuIqcEFlebP7aObq4x
qG8HUQjk926zHaejZN6SDSs7EiMaJnJxUZcYbE7qess+rj/sWOJXiz90qnQdUvsMf0ybXtrhwYcp
IkDeX6GJLnUolRfITehuktB297OpzHFhw4LFvPe9HhA7eqykDvs0AotSiqRd0AVv/3cvPADcywCR
WIt7pVfiOVByAC2HAf46Omdwv+6rhnfYqQi5reajisznMsc64c1kXoOk7jclT3KxxfDlMrFu0s8Y
mj+8kjLVvjVcwf4O4ArV+xX7c/x/5l549I3sfoY6lHA3gXkv/Km2sHOwU5LCfsQSZicfaru2r60n
VTX2kbFx78FL2VIQnSF9uQmG1Xum8cVQoHZ0dlRWwKXWGIkVppaJZa0zgOK8Mao9XbX2yL25+GL9
5pB7/kSB3p6a3CWRNnpOXaaS508GJR2nxgarF1uL0KlhgIqQADMpUz8CJEWJuu4zXQigQdA8M5bA
9amZL5+Uz6NIjghJeawETojja9quTUi/CHa8Fu4HjT9U1n+MvafUUpTHbhAMINb74XCug8vBBcEc
3N4SR0Bkrh0YT49LN5bjRiNMrbuNcme6tOkXavyDr8JPpUaf0k2CdgBA1SU3OZQRqQCZN4ZMuLxt
IiQk1tB3StcEYPj08S5AksW/sRH5QjE3Fr0qhSW5BacmUTofbKWIfM6pi/hA+KwjpRoPWYRhZert
3yYWRQ1/lhFIKrbcHU1zXQV8VyI00Zv+HukiJYU71SELgmSdlhs7OjoBuJ+TFOAWQJhSbOtb4aKL
amnQjudRCK8Ef02XyX94NuM/MOh8/trNaGXn32Ov6dJQOKh31WgLp8Wkf3ET0OOLmUUlJz5V+fN/
VqNY4fJuKAuVC5x1PaLMd2th3z9O6is6WdNpz4qOYNNuYjKJkIE8g1p0dr6Vyay2XuGECBzdgjXG
1P2KcUsLLVEUTBdETUDQNpW+attdZW89wFZtZl+bRpSJOITd6hRKI//lIuE58xGcWlFusBptFfq+
z4/gVSHU9V3CqQvL1KIq8vRbdw1RLSvDqDo/NMkK0vToUjt/gMq9VglJYs+FAWgyaaQZBwCV1Vjd
K1qasvrdSbsWhyqI13ANN1YOazNdCpLEs0X5y34F9peBYqiD0L/DD5FAjBBAIwNeg1mdDRhcs1jk
6ahF1u86efjIKKOWUtbLOHkET0KBaS1RWdDq9sRj8VMjQ/33WaT2Q9wCvaeyBYjZu4gtKK9iBZgI
WP5NRCOX8p2sgj4dEpQbobGAqfdbFAhwZTzBbL6Fh1IOVbvDC3h64wA7oW0mrQrAEkAFXJoOJHnA
9zoWU1LX20yVy5zZ7mmMN34WCPBhAY7IC1S5wbCZLXje4CxoFgB7BECEpPIp0lQQcJAUa2X3XmXU
bpTR/XEo/J8FD32VlpKdHljiSKdwVAefTDRSylQe5SAqossAqgp3F6Sg4yxwN+DC/w79SNQfinhZ
H05yW7gsgEFRVEg34Qa+CgkOgJ/p7pL0WgFYXoUwlR1TMrX7t551A0YqYgBx0zZVmif/UHDf/zGg
GrstQnQSoTKtQWSTz1ak6h/T9eej6a9auXTvIzVWcHkgNz6TboQlxB0RiUipE7KZHGYbuCuGM/+M
RYceDO+omfsd2fuk/rrpWi69k7oo8f+FZBJpwekGChV9bKVHDx6bgnieWSJy625++ZRCrp16Q/hy
D8vob8mXN6mT0t475s3JZDXNt4Hn/Nigggyq521LnIZ6IKFmG/3z4S31d/Is5x++QxdpJ19FrHAU
WKiILmhlMFDkw9NxF2c8hvcbcGpnr3wpJJsLWqVmSkjILnj8zAvwWM8Jau2we57Iwdwels7Osh3b
ZHZzz7QE3q42cJcXqspo0PoGdfZc8R3hkQJolJUDjilsldnNAC96l4JzDLf0NEU8yQE0X8on18yP
KHdIjgQVDRVIAFGyBpHkSvdvheGbDOIoq/vbSW2gzK3tiTdW0T40KFBcc7sUn8I/MNxN4m3SbYRK
CCSb3DY+nI90X21ASmbPX2ccmy9dTDrImTDycq+qf9VrO/6vnDIxYAC6M0gUR8Cuf/1LGV9U5YrO
tP2sCKgn3aIea1ksujQ6LdrY0ba8yIiYOGhElitytgLsj9O+rFt9FomeHdffeMKcCJidV16Nf0BE
wC1yMkzbO+yVobDPcB2a0AOHlmTIOg6jq0rL8Uo3mYNga3l64jzdG6ig3iyecoCnTEpvRX5Z2NmZ
ZPeJ8Yb8swvWn8f60nRko/VQkwqBthvbaCDfxaqK3Qy/JLRjlGwJwYbrBUDAEpZ4xZfAx+JNjEvz
MDpRNMyybLTZxIbhpJFQQpAB4936qx08EjLrf+wIlIxB0jzs/M/QsqqhB1cfs1EzzAxKXWZ2avQT
j4Wx+Sf144Z30qwm+Cuh47p6jAvjNNYK0yIq26YK6Y/XYhZc7zo/M2uOaS1y76YAHKRjanaC3Npm
jbGONqqyUBoA8GQd/x2syGZFbdNHurUrbOmUKEXJX7JCsrf2k7peYVps8H01NinsrYKGHmqBqAqv
Xr1C7guVLmYsGR8rhOWxYw2mK51R1cB8q0dBpdOvfR6iFIEKl73oMBYEEz7hJPyh0dlJ7IIq+q34
G7jQ9fVluycnpw9fscL8YcIW1w4jGktbSQJZBSSBigQa4AD9MeDd2Fcxrdf69qfWXLdD8IIqIVh7
EvKRKaZLWu3RwMRVtuwmQnl0J+DCfXYaXYGCnWuVf+vou7i3JB8h5RZk79BKtXy8nKiiiyX46BZ8
gC+9b7oF0hASdd/KEXah8N0LqK9yDGSQsRtsvLXvK8lp2ELWoMvSNqDIO05xPr/Emy3QqBRjDhfX
n7gZvQzR/m6IuBN9nZ2DMAqDLuDXcsmzmpX4X8SYwm5DaFf6hzr2FM1ZKgzw7t+vvq1IDz9j8rj9
MSkDncRc8DG8oABY7TDZYOIPbKxK2bkfP/oHypV6vsWw4G7tiCc7UZa9HzTPb9FxLfhRV1jOuOcX
XqzQw5D2BcX8tUwPbLWPj7LbEKFk7Wjgq2hij8VuqVnsA+s/PY/wWXkKvx2hiSX8B6ldX8XMA3xu
+prc4PvkRCbpBp7fxQsTUNLSGqtkPmXQ4GxMcavfz6ziTG3Fve4iR/pCRtNnEZr5avL9QPm3dagQ
qm38ZXMBYNUSeiSUkVAfRy6NvjCIi/Mpc5fBqRBL/kbi2Wzn2anXCBAZAqKZx7H69bB6ZMqGbX7V
1Jxb2OlNiixAf6X7zL7QpGRZgbqxbIWfxvd4aIAA9c90a8UgH7udTYVQ/OKLH0/Cw1+vANdDDhGc
9TtgThqs8fnqxVt65VZKcJ7xh4VFvRHEu5VjqDEEisfzbHi1sGjoeSUoo/FdOtoM7A9bh0MS8B/x
MgYhkygvh1KRTePkut1n73TOFNtjDkSWENpGSd0QDkdcHMv1dcZ8Iig7voKLocddRXZB+T94grE5
r0MbYnkF8MNHUGxGZJp1qt32wxtyMXm8mmDxIRRIrPKo/LnhzqRavb4Pb6T4jM3NdjThu6k8nXop
yaKNbo8nSRVBenE9Y/j4s1PbtIegbD2cPwtEVpG+SgKhwtD+esljne0aCfXFhlxbcxiDvaTIsERs
8pUjUE7Sg0qSQXtZU34zWkYt6xLeQTnxNu4DhSu6ehY60BwIlOu+oYlQl23n7ECExkIcWMHRSbEA
P/ZTWNgKVx5aa+YPKns4n6ifLM2CH7oLVIvnYzWap9cb9aS85xWYyQhhHglaGqQ4yxo565KN+NL9
IzH8x/cyOaIaWMK7H2YGbuYYiJjC5hD/jaU5ArSHAPCV0Mqw06UjSYq9YSrPJ++t19W555oW5aaX
2EiZqIvLicKqrRHou71Xt1WgPpJlT1/q2gezYFeHPtr3AvZ27RKggY0FIzILg52pHx/9TTK8Rxxa
OlV77acAVuZ/rPwUfYilcMNvYg72RP5feX2B2AkhaR3nIHpvunyvlIJAscas+jyvhRRn1/DSYIW8
WW6zjGqKrRlqXDsXoK5EAlASYz8Bqy1UGlCQgcJDt681UDjt9I6vGSdRZAn3qRYNV06bROQVHXWp
UZZvz34048l/XNxksucVYdeDPFSlJu5IpvE4mvFuorpChqMW2ulz8UG5sfaLjOLN5FxfC+eCh3pD
ITJXusS7bAthr+ie+NxVo6bHIjynW4vF9ID1ey1V8ujSxopXHkPIcDWHPzIvVs+9neq27+RZRmwJ
D5jV5xdtVOy+cP5ucu++cXfBXf6sFmQ1gDhp95LItxVzA6XyT0B+BcmnYrDobJXXPR+2esFzvODS
7bXbcfHJPGMQXR5lXGt54RuFZZLiP65ws35kwrvVkDzhgUfXGw5EKlodBL0GDeWGB+znBEpWORPP
K/xfRyHxXV3UHXdhJ0JF4jZgmzsvhGvQ32tICQ1m/RAWOedI8+eoGMJabSBjU9ucsjwtv5/mc5Cn
FfX/BMo0R3GPLFYj2sHxMpVq/bFXmEZgdjT/mDlm/vPQrDQRyjGjk9G/IxNg0jVBaMlJ3QfHvRqi
382K8yS5GFz+/6tMIziikBaAhg8ok6VMBpmXu7zNg6YXjYFzYbJkTC2hQFM9jjZmDs04WzSfim/C
btuF0RRU8GTsEHIXFNntu7tE6PP5gM/s3mfQotRmEB3M4hPsoTm5PSIJU0a8PXJENdefP80kcXKG
dZVW2L/EOIhp9K7ImKdUYNTDIJBSBXeydv19uyXFgx7Uoh/rEINjsKOCFLLhFCfSi8dW42o8Qqmb
OUbZBYCCwsho2rezVIAAdp93sSyrxb4K7tHZGjKvaKutTf+otXIK0A2Yzu2WaR8Jk7YUKBFVK9Rf
CJRViKCet68BKXjPvQfK/gcmlj9/BmQrES5y0wFi1vbr+APDTNBP/4NYVZ/8QZ7b7BALLX+48fbv
/8Jku9xTWOiYoyvHkM+VjwzVn+JRob/7cfrwXmxuAnOstodNT0+UqfLERvDQshVsxGi18vCUkD97
mLIS18+vS9feJWuVmxhpAZULNW6scpQBOi0TrAmMVDxH2VU874c72cn/oT5lTCmMY79C6t+UnIqE
5SKwTCIif0HYhXZSerSZWwP5r5KSw0YdcGQ34ckppJ/OLCEVsE0CN+28K8/44ZI8N9SawU+64MjF
RWnrO5wM0KtTmVStrmTZINIZrA2hnI00heinV52dRkkS7cJwvU0vEr5Y2xgFnibO2E75BUY7CmET
8do7G0HM5BvFuzUoOqkFronOYv4Vz1jQQYDTPAx5qZ3qoJMbUU6GqgQWmj6CyDhP+OqWo7w1+AO/
Ne0pcg9Ex1oekueS+4si78CxzG1wUFgEjHd+EBsBySgCd/BvpiSOjLbj25T17QGu6RTDOVevEnmj
wgbT5Z9klifWTBHq2H8aUOkqwySF1X56Eu+KSWBpPPpRyw+lzVUic3OepgjKuNZsT+GWkToz6GfI
JDHFKBRpXqBIeraY/s7INq32HwPey/VhFuynwIa569Eyu8v9vmc6axTtGtJNe0bK4/qe4WM5/s1L
J2ciGXwWpGUTz9P9OkXIS+7R8q8DshkAXYZd9DGpNkxzKPj6u9RPixn3cGZqun7xA5w6Jjf8hH6W
aZBZDHqRFLVeXubINFcble+gWSun5N4g7h3zcEFG5awIwkORDEEZLPg0cHcK4ku4RWkyBfAnGx/b
0vfZcP9/l74tWKIxajKQZw0IkBUXakoGvNRgx26ISm2XP8AkLbgLxdqfTRXguXXdTw4I69zPcSmx
H5NQYl+GmgjvhldtoNwgMvTwDn457DsPLKjgQDwFl6yf4hfkaOlWzkzwN6BIJ8WQE0/PhY+B65gV
MjrvwHeLY39JvNEtK4pA15mqJ/n4xf3cWtv5caOu0FUTYDjZe2iBZa5uz5SdF5X5LpCvfNBz9BL8
JEl5vrCWxslv4VKDduK7es6bjJ97ZoXyltpezsCIUc/EavwscoR5wiDCfg3CSmMy8Ydl5ONkyL1I
P54vJcIvrXLVMDgSxFqO2bGZdFCgxQvY9Nzk2K9Wd8epjQXED3OvVMOGWZs87hA041ozyGFQKPSN
/V2EnsPo47MzkuOID2znTW3O665PyNV2VV8Tk98VbZ1kHjI/D2AcBQsNcVcg9YBb1HnmQAcksxd/
qS0OIrfWqwSMgtmUmbJQqiy7zB9RKVk3ojzpRbt+nPzPTs8Q1yD68Oqktug/83NDvWXvrFw3YU17
7RStn0CIYp9g/KL98VdoQN2CvrHXcz01Y49kTd5Cb3g6LvrRPjb9KySiquS5Uj6uThJXJby8RLrG
vRVfxPWThhLU4on2ql2uYoGnIELR37pyt7CZLYlQlCxma/2kurnmYyuxAPIYqzwwonSBPcDAICF9
JotcrzzoMUHp9p9ufVPd6SAAlNamtllL7pDKESHuq7tN8P2mViQTrONMzlT45pQBGdH1rn+fSZ0e
r2GI1OxOps9qy9byIXlgSm68mJh6edC/m5nL6ypE2koLH1GA9bvwXOck1byi23oIskbzz6orZjHs
uzuFkubHUPoLUGTcT0UA13eQ+3OSTtio9bkgFnmVVqjKd77ltIeS+EZ2C4rxvk8WPKrvHl7vDUNZ
QprcawpN5pXWtlNHnh9s1L8Pc0eRLzsra42Zkgn6ryiXZc9Ta5gWMSFVljrdIlMlHAju/WRmvLOm
J/Vd1ag71CVyw/NfYeQXcsESfPQ3T5XnXOb/Kk74oab6bliOBO/HWDmmoVJTNWrF4MI3kmniSU1q
g87NeTK5HZhwqdX4IGfRqr6G/sqF+tOw2Ad7RdIfsxkfKmVYoIAwlkEUDUXU/gODAD/zRRwJerEz
UgIJ8FNGe8kV7y/3R3LzPFv1y+rEvsUi/JIEq1YmgVx8PkdsG25ye0dYZd5z9IJ4tiFPOBhcITqb
1O2LeDe0KPVVctFvqDaR2KKrPQQpfGqB/OJXRMdcnqe2wTNgodINn+Y3XVueouqMxcMVRPKzzSn7
SeYyjqkSxrOhewY2G5Ts1ISHLvY1jze4ALu2DNN8xFail1ch5xFxCTMpr6gt5KCDc/6/2del1xOi
fOhWo22toevwHuy3YtA4XlJUx+BRtYxpn1+vfju3UwhG4HhM9SCYLTeLk8vOnWxuFPcCVDL8T1z8
EY3C6HMGMROuiQP7tOPkinExYZkQmP96+Cm5vGzEcED5vQMOQriZLhqaUH4z8u8uf1Nbg1FBHeH7
XSIJwRsTV58BZO1Z9Kpu5hO440IEvaSdY0FHnLfY7G8rX/7onza+nDskCajblE2lmb+6x6m3IYnE
JCk0t7jhQWVLCESq4Eft2G5hAMGjRhDvfBLQpVBnfZaPeI++GlpQviVIkL5KpU+eBV7LQdCcSQm6
lgWfCVfWad/wDOluecwFBcuOI+4NLHIYL/alrgve1TJ0d59rXYEyAYQCUnofiZ9a+IGISXt4iw5V
99ymteiCSZ626k3fbV3eeQcvq7Vwe7aiF1df8Nz0e1qqceU+66dOemll4xbKmVuOkC+qs/dtDdoi
ehaIa9wlN3mIJdizdUhVdrHd5CoT5Q4c9uvUnuHyqaqiUTw+b3RH7/CQPgK1/8qhIgVpfncdBGUV
cUvDa0dmFZ08MUeIUQawpHc8S+pNnOE9LZ8B/XwMGms+YuZM3R61Wu//JQkCG+ZgPRuYFYI71oBd
S3L1e08+nmq2q/Wx1FkDE6aNH4l30rgcFUmOpGqF+usM/sSzVTiaHiSw0AjZegEDh1J6B8dHu8TS
GLDpL+EOZ03K6pu7BOMZTo5HxIcKHI7D324XW3QWJLE5vTwD+o+j8TjsrSi4zSYhJ3N0jm3JMYLC
DG03vVEkOSxQv/zlWInpHO5c/L4TN6gUNOknkTWSvI8tKeYwywnG/+/0+y7v7xiJrN+TB0+yJgat
7n53abF1carD48dBYK4oqvKpEvd8z8WBJcAvNFUIKsBblr+meUY5XkCY9I0wecLx0YXN9clfaQD7
gbxVr4LxvIahzLvRSDBRRU3i3uUqln6Ii+XFKTmBuR15YuptiD0eJIEx0cJnrVuZUA1N17rWAeQv
+H6rV+tHf5jRLHJl0RP6zo7Ul/J1G/NH53pHZp/9+3Ykr3CZ6onjN0NfJDBVImCl4+2KuvYprUaT
/TzyFuAVyQ/gHdgM3GMuCfxwl3pTY0nLfM5Q2kcoXzootYVnub10GQIYnddZYKW6+uDTh2urJxQQ
PMKgSrsgzRwmylWqLxCarOzZzz9uIytM4f/LQODpfdgn18ybC2EP0iwnnMqm4VA6/Hd7Ug3LKgNN
cdbCr+2FJ5PygG57x/t8MynUInP/if+Qz7rJTnNLomIzgAeQNXH47SffqPg42gHg5ljkbLZJGR8O
nEOzCRwGOOWjSLOPiX7pcFFUIMjSR+e7xtLE1g4oha9wBhx6iW1Ohuidvm3ILjjcrptbMK2dxne5
l5P94x/+htTqbrOKSf7ySLnZDczjGT1N7ACumWJjfhf/ZDUoXbc3N9uWR1T7mt3gEG8rxJYQf8Tw
kKNwqMj7RBDea7iSl5V//g8wkr3TU1PGMwifdqYWr7n/EtSl5uBwpR77M7T0dgOQU88pCFRJjgwZ
n9NLdf+xYeKIIKP/rLG0uE35DK2+KEhnBCx3bzKHimD2Mn7xvWd/ZWa5ow4Iec6oQtfslYL9ysTW
sYlFBzSHnPWcoh9JjF4o0QaTK3mZL0mWNYLePiyjdnFZ/MbVifUYFazSxeqsHqkco/WoJlMlNuK5
7bwrcL7PDvMG/wolNUT84v5UCyEtnE7fw6s9dHeY8wn1H/Hy2VNvy2qd3q28VYS2ytKYEKHSTR6T
n1Efz2mQCS6D07T4wyNPikuOi3mz9kx6ozO8T9Ctc7N5Wt3A3/vJN7VG8IHeuJQZrFDLk8lKrafz
zKaW5QjesHCgHTfzCfggIKiQEUwH19OQveaqbUHwN0VQIFcHUxFkRQMVFvOFUwJA/RWGZafy4Wn+
0D4Og2s7nZGb43uQwrGwNgiDGCpBxVratrA0VwtLaKk7/UTKU5O97lItv2tPjBRV428eIqKx3jvH
DTwTSWBfsSXNsKQcNq1CHzvtiB4KZVi2e3d3WbgcjPmgWtED1k8GtG0TDn0MqyRbKIccb5EJkW6r
PGROCqaNhVzJcTOfFKe+W9pp7LYch3An0fEZq2yAQvXQdpTVvlELKUhnrsM9Xv5nWYEDNDSaSp9V
oIrKEaiKpCFOjYLlCcrdyP0iCSgs1SaEtJtimH0moT5BmPVeGYHpuppfne3YDrpDTJlUxyfy0HOX
JH5RdwMthnvMyAM1lB5EWLDCmZ5BRcvQPmebtjM4JxzwD7n2M44N8aCF1QoIQgHV5TidHr6OIswm
SasxoXdQ9tujFWCcxU9ocmLyt7J+9h89FeN8sPAnjGms4Upxs8jUNX7PMsoupmiAm6A6qBT3MPHb
Jb1EtMPHBtzaQecCHBMAQOB7ZtW6TP1R+flw3jydYhodpQcmZOzF22YCCS0Ou9fyeC2oSCDZuT7H
A3XCKWgnaz07xHqIqxHk/CtDTrG1cgn3m/xjxBz8M7JaBc/788Q58dTDMoFBGnr3TUcM2CbR6KKU
AJa1FluYW/KmW/Oq52d6trxwrCp8KmfNbFzGy3Qj7FWYpCjIFCo/KGfSugGJrwQS0OGZGReuebkv
5EqrTqbWuczGPwEAShNWfzGA/mi31weyDwAz609AxrRKvpCmtxZ0p4O6rXU2+39RL5ZceWJVrmMn
kOKtPcTBC237lY3CV2Yt2i/OH/w5ADEMd/wOx8dSJYvkaJw7aHECTUbCr2NALyyo3dFzB6ffC8OJ
zrkWbse4gWTcgkZIfDzDoA4A191CVscXPExuyXkCqrHieSAjt0W8Z1FJD2PgVN/QIRlHUbKW9WlA
iy2M/xgHTlAd4F872Fa3AiWWu5r6XGVdR3LuaLIRsa4CAGBDYaKgz8/XPz/WFAp9/7fJMIGERGvP
ujJ5bWc7BxtJFKlI6p9oTlnTSKl/NOl8xVaLmoIpez15AimgjU5cPgoEGA+zLvL9E4PidizowsnA
wWf3r4g2012Py2mHiYYY+0aTNkK2Wt8EO7jasCUWD0ZmJDGh/XkbG7VLSGgSe9W/pMaLw+3xRx4T
epd8jddnJND/BCMmp9db9QOt4xMFgyxncT2Ou2NzEuWNuKSyrRROBFtZWLBVG1Kmj3QY/RiiP4TZ
Kb0+XvEGCKG0rDhzSGFb3skxnX70RJyZHw8qUe+2OdS2lq8WSL7BO0caf/2oYp4uDzUSPbIEBOfV
mRj3tSIgPF371844Hxn05k0T4ddaKiI0zvzQ8mVXZI1+kEQ2ZcEf2C8cNvqBPZvmZnHOVhLdXVzC
ZMxy99fB9GzTHn2gGKesYxI60/cd1KtvIUBRpu4VLkzVu9EAjjKRY1tn8NA49fFhmk/l+Ap4185/
F0A73jPNZNgZ0fLOlS0vw8n8AMlFTQFy7gwmZbeFFK/oVwpCzsKN2/PFsJDbCuA4n+PBCno5GxnO
E1BSScJ2vp07ly4HKgPOo/S9+XRDlfgrtY0+BqtY4z9uLLfzkA/11E14Zotxxwq56Fp14E//QEn2
UrRAZ1XF9rFltKN/nKGjqGrmJBjOd76lKb1UHV7sxm/EKjS3bu3jtEjfmjgoNar6u6NnsUEQCU2l
8fjnsI4xZKzIQ7edl1+QkzYzhhGV1zt5lqhaxayB4HCW7H5QMPdS3IDOGtTFf/zim8+orpjS6MUf
0SlinosT6TkOGmwoXLmuLLY3DUQjqDyKI2w156RbTQYEcG4lavpibkOZVqkfSf1dycFzyMbDDpAo
ozaMpvLek3xe54LZkBLUaw32k0nPbUufBI6NzE+HstsPbCweKrSitFk4MORzQJRkMS7fx8VxVZDM
RrYNPxsPgR9j3K/UDz0nwSvbhWJ1hMYL1ZM62tXzvRApeiDqji2uN2G3DoXFV2n+vK9OnhB4fCRJ
daz20pQ1Uu/55MxSm9+8miRYcQJrS0yjsvqJTHvbJt5eHJBjMBgUIsS+VJKa2WBQDqXWu2QcQJmj
YPhotDufWjZRD7ub1QUajHvyVXm2X7ilkIeWUH17ajDLje7yA3KBA6bTc3GQ3YfI3+OPFApvb1g4
sHXrR8+JUcnfFyba1vAHDFk0LDnXhBQ06OBUHp7qy0vtRQtYPR5I/97kZq7BcXvVbnLcbYaJ/C4c
LULzh6zK2ANHTigHk76JvyylWtfPa0rrFbf25p5bZ8EkolfyqQJcsrBOySIx4NwkHxFHRFjuDukO
wqRAfFNYvhdUOCYIUE4xMkLZg0BeJ5mqeWAjz3WWGOvGJDgzFhHq4r0ybQEL0OPqYmndlsjzV0J0
S06bcFGFHQ8EOdz6hv2vJMzJLmLqP60PS2GOqt8mWF/VJSwE4k7Cj26rH8MjiO95Xwk5wulJLXR4
Yo1byQySZl7KUwn4h7Sl8ALuSyQW3NmltSct6M4lK8UiXRQSeFmv+tDPL1iF25f1u/EwPBRtVUhb
LswkXh2B2x69LKvmlkgtqEIlmhwQ6cdgJauGVqxWIEKPvacp4SY4eI7Xgg/YNX0txzkuwQ8I5GcZ
NyD1BcPSmEDNlSoKYAfQ4PIEYgSWuLuwSQHZoJ4EXHH5+KnhLkm88AjyzKoNCrlhfQCJpbHE/ty2
F5h5Mj8k4xLnpS4//mVk52XFyWt5T3gwQmHShJMzy1QX1AoqcHtl5cdDn6KZCvMdSZKYsiHjoekx
pPxxz76GtFfDSMZPbCJVCoB7+DlI+EAWp2SIcgPCGSmZiCT1oSTLNnMrTV9jTmAmsQMhE5MURk7o
sBF5TXEuYQFDVJgTmdHvOT5u7Cn4VWDoke3ozxbWD0wAFiIK85c8TGAmtVpqHsuHacK9xWeLOXYm
U+oVmorPzvu0t6WaObZzEtwtC4pwU/MZZ0/ScbSduasNvwOo6uYFylCZVLJLP0Wfgul+U7714ruT
bROMMJq29uqtFF88NorGLWPnNGZAQDB+TMF/rvIJnkFj3BWS0lOCJ1eDBkcR6qfMEu8QGaiGRlxI
c/n7bJYHovFxpuGxYmcp313bPXRpRLrWYHGpsScxxWhSTIhMznav6QzBPATwZpLP4QR8qT6ff2E8
NX/7riadFnI3PRNwIMhrLrBl7MuT/ULbM1YzUKyh6ce4gOPU8JSiglhm2qR2noZrnYMpQ6d+3mlu
qpIdyX7jyxUIfhotA6xtHJRbN3TZmdRvp9UtsQNluk+f9Xen6lv4NM+KTtlp0lUZ0bp4M+ilB44t
GpDYapWy1USTBWh7cqQnwvXAWw6j4nl6z22jSEcrAmT4ciiNGTnDKSGvkr4nOzDnDHi6pr9MY1dO
pS8JWJwudbV6XRmrBM4kT8Q2jJdKm9ovqXkxTIP4TAwfWXjL6xX4I6msY4MCYurT/JU4RgkaDUB1
wU3No2kabI7qreeT7qrTwdLvd9scNh6t4eHGYaMS8hjkJSZnDdHjx3bupNkQtvDCCxf7dkSLYh/t
f181QfjS8K0SOP8vonJVPsGMvmKIwqF09tn3Voseio2G3/Jj4ru+oWmVQjSgNY0ZkO4YOcWPBVTm
oFhM3xTT74/tCKZZE+Vatq3d67/oTHAAz0WFGDakU2deaUMgVatoTOO0FQM3awQXiwURan/+5BAq
lILh1g5MQ7AhtnKvDTyzqYhIjfY6zImRqu7znlfUQFsByiuBKX5m2xSnetkjR9nTnxvwJ3fodzfa
NpE8V7/qF3agcJGxQMsUrnefZBYLm+nF2rKWZBZNHQn9tmt60W2eJEaYadv6i7L0VvH8DbY+uWDl
yiCG0zhBTD5nQPMi4UlQsSqhFklhqscbVmTtHBKcSAH6IC6MRMbgh7RSJZcEBwDr7z34enmNqUqe
4v5HeyAdIBrOcCOO97lWK0n7bvHKCK4bbfgHZ+UaZ1CcNtNG5v/ahq6fElbXuS3Qyj/lxXC8QoAR
6URXNW7qiOJJalG9FjU+7OzK7VwrltUb50pnidtFJc8KZAFHZ/R6hZ3j5e9h6EPEYCnJEb95kn7l
vxTfrlE70gtMZ4uS0ePTJ1dJxASkERthku2CMXgVQT65opDOsx734SuHr9xqb2jAhOSMHw/fnRTs
UMljNpGXfVQTvGdrKkoHf9E0QSTw3NTfzDrCmsMQ+ePWmcNxohi0OraZTiKOPjNCK774caIU/ZIy
vUt0vTTrlx+s7f1ARYhJ8A9vjEAYxLdFPucG5GhnTmx9/g6JpOU2JeCUFo3O7GJLgm4rCo+8Ikv9
cjLQnURQAd7PL3kTcxfNLpOKv4wb9rmhbEKWV0Jb/g5TZehkTa50fcM3VP0K9SONbSlr+1ogc33o
6V3lKuTmb0jmxgowX2p7c9IlbzdNB4WrBVaqUDvp1rD6yM2Gjr4p9OxGNer065PYZ2+BPUHadKEs
4QdGZg+dcFJPgbYYcDi0O4L9eyi1qVoU4h7shZOQR2i89U/wIIX1ezGUaErZuorHSxovJXmwDt7F
NVXj1qbdphpjkfHI2EK96BMoDbHG2hnUHnl6IGJisjJRJyPRoAA2hf/AI/x2u627ZXH8qSmJdKmf
bZeMfcS0n07bEJ4WU7qlPzm8je7sOYv0ZjoFJzYTvQixJ3RrxRVY5o119+zNEmG5LmVz3rIksPLz
rXoovkv98yJulppFUX7C3bbjHNllY8959u3rE8+r2ZuLSdWKAPSipzgxWMo7ZLif1nadetCvYcpD
tBz0J5QjtzGweJd56izCLyQclhaiey6/nwlTAdPUCGMWnd/crsVcLd74BSMAzj7BwkRIOy8hEQHE
AvzVV0LDKLhZDGz1pqrr8gC6/i/I9u7+c7RwZsC45EFDglezOkbmMkGtwB7pF0enIjhnKmYS5aDX
D3tXtrw1QSWRd+RgyaCySLumfGRx2pUi/Ryi2HUfh4zlQV3ZFYEZv5Z1eBCbNctzUssXnIim69Nq
6gQ4Mvmnnj8Il7DIWNz59SvlJ3sS8u/EXfSBH2ETWWfkmvQsrY3mc+9Nbp9CRK+XSxbouUaLg5P3
SyBHLlzFjRDpzZKciibvtGD/COsQ3t8uNtWEhLhVl+Wm9SamlogBMebiLpFELFxtEQX5xPW+iAYn
SFIaUN/qT3gQud/U7eNJdueUtES1H+u/g2ChT0eXBX3zd2oLtrwppvzEYh5flmlHdeVPvrjUB7VO
l8XjDNsDRCndmylS0zpIwK8J+5RIwQ0FkFBM3mB0BSg8kSWoQ+lHYVZhAnHEheGEfWNiABXf4xvc
HYE1eDl78Nh2ODroKspQoRSxexEwSNNG92JzhuqvOhrSQez8syjxdaIi4u1zP9waMiTvldYXi1EY
ou1eerBiV6CplcfByPquMe9xJ+V7ncb/2f3kg5Rajg4kogj/DdcxC2PGuA+43eMpLl5TrhMyUIyD
4fcKI68L7ABOY1Jl6iONdy46HwiVxrrg8E4ObGA2QtYLjQmAuVDDrFbCu820B2bvsMNmKtIcA2W1
EcEeQN0XUzNk75byhgJmUR21MuvJVu3rGfhAYOLMTNHYzoZAcLu52XarLA/qNqNGptg2pmsb/oGU
BcpfLqfQx9Xbwkp9SMHnijMzHnXdKQWi33mGWsWNnHzFvA92tnkMRbkqM6NLureqBb23pZoh32tL
hqkMVqvNyZFs5Ah6z/sPP1RU65QLeUQqp0HlORUHBnbs67Dcf6UWrU5qNhR1MK9wjqA9hln/R+VS
EKCr++ZZr4xkrAE4tVzwwpfI/MYXoamvD1cfqUhENINz3vqX1asWxwZZEicRtU58XkP4RjGYBeTX
F4Mo6XKO1e9ltj5981016L3crXv+Zy5m61C91QtDJZx7tJfh++eV+F1XkMvj/ojrlT7d2VCCSa/Z
jsA+enWlW0hOQvj7y3Xq8jMeXsfoERbEGpEhKCpsajFvpbGfLrGOheIdhhqNGa7SgX/yaoG3LZJ8
FVaJXvVf/PRgp6U6FWcJh1uRFDdKOJY9HwfnJs75f4MBzX7OfDX57LYkpybFBbqlozAO2OlcUvCh
SQ0un8mGNuXXeF+pVZFZAMqH//vLsN0Vo4UTdXiCcWEHReKVL+gjiXKTnLKJoSp38+OdU9HjqO2x
AHL4Dn6XwdKfKo6EZKKJz5Yed3yI1jE4v/m1SsEv6Bzq+5IEJE5HuOGqGast0M5Ypam/lvbMHLOA
xCV0Ey5vz/qmdP8ixgDm+I1J5DyeaRXJ/ifHWXarF3/wOaFCS60kcmJZIOl/XGYVVo7lOzOH38t/
YG2eFGMc81dT/FR3QTVdtQVXE3jCHXKA2It43UNE9HaC7W6BhHKg5pnoDEKFqgzNxJu0SEdJtbWA
bsDr7K6zgVT/s2Nh87ViaMATANC7AVwRnhs391R8k5q0A0fpIFHK1QkamBlnFrP1HwhrDeYptphg
d/S+5k7fQUSwYk2Ih0vgUe6A8LZVNN4qTohJ/CiwWvpnQUeqHvG1XFUh+nN+CRlLy4yvesBUMfaf
0KY4srz9PK1WGCpMS+w5s2v9LvdTyGH347hdiPFV5OxlLLaPG+hiU/S8uRT52Y3kE1UYz39Yb3eF
T2dKoPP1p/quCEAnFh1oNVnQCKql6z7MHJiPMtHiPjwBGIRJFKDRNTnQuZRz+wRl4laeu5A57chy
4LuHK2dvjlhulNVWrSNOFiINry2dT+GGJT+vpgoaHyrrRWEYj4N5SuOwo+UHeBxFw+xrM7jBYWrI
Li5yv1bRKDuAijk7zpxwWAXPiLfs4PsX1nN0dzLvtN2IzVlvbwaVDs5W6t/cax8TZzg4m748cL+o
VZbYSdiJUEe1no8HeXN3e57CSfyJdoI+48MSwH1ZkFHhwb3fTSmy5HOcA+GgjZjUFtEfZeWS7t3g
33gyR1uiB/syQplxgZfkGRNpwbdq0A==
`pragma protect end_protected
