`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DUDrAHJOO+HRicDCfge+MvjGkHy45+FjO4LTtFqKnHdLxooPMg5vgZDBxpGtCnTA
NwiqNT/5v0c7hiMxD5/9yynHH244MX3pyavJKuUge75AnLL6u9LDPUw0wzmsbopn
6/kNLLjR7I1dS+iLTC7I588DEqYwoBD8iuh7BkAA5iQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2128)
cVOLjDQ/IsU1GVaVjiTuYWBn+X4DNmc/9WMSDGghOJbdFGdDPXq6vwJJakN8oiha
VQucpiC5G53UJDvIrhLw4A53M0lgZYvpEAeQd0Y6m/t7EVa2HgRe6DtVtx7Of57d
vzgu8XFXr2+jI3YlnojvYiNkcZ2T9OxePb6S+6ee3lNnV6GfgNqOAEiZf8Sz/E4e
x/MYEVU4cbeIwahS/2XsNZy5qLo0gbtFkedHvcVi492b/mxIkM7OXRCRvR/E7Esd
kEiGz52vB6SeqxetfGNgAh7ckystFgejPaUH6QxWOCt73xf5ID0Kx/pqf7l9Mmov
tpXEM9GKmBbTSTr9+WNqx0HBhqDImpbd2KEqT9n7HDo45JoJv9wtYQBDTw0JApZX
0pxtSeJGMST1Q/QCcnTdDxZwOy2Wn9x8tJ+yOgCkMyCnkjDQsS8jrLMf8NtLTxGX
xYq+t4UKdGA9dErH+QtOe9/MUAeOicTb4Nonv758D5BRbhS9GIr0pM95DeFCCfP/
dsfZMTSDmS1NBQASLgaY9ivszOXOOe8Pe8+mnZWTGGwK6xZrm3p+x+qMA1P39u3T
De4A1ZVAXU0zPKzN9Vf6CB8cZ8FGCNmw22D1A3J5w20aamm0xhAFLWfd0IEQ5zbO
pRoUzp8QT5UIDCmvTs9drIMb8jC4aSZuWnFhKE6aCtD/jhddhIo3zCbFot3JGGzX
ErcFIM4GpTo6d4CqR3D8WGaaAYQ7fvnXZI3Tl+Qy2AANESjR16kkQ73wbJsqf/9H
sTOWz/o1GmR2nOnrs3uPouAB6IacJDEI6QZ9JBsDwhTk5DWSP8WBB2O/Ido5qL+4
O/fAF9znGes/CsS9rS8/mAl7gm2AU+VXqJTs0VIRy6sghSGn7MHfHu/9NpJLuv4C
rvCcCAJ70ExQzcNZSiQ1shZf1qqa273yhTSuZgNClg7PeH++KNRtTvKg2w2RQQXU
BqZCamE6PPEfIbweeNHuQ6HFpQI5IqBhsfWPK6O0DJQfEhuh4+M1lGyq5H+9rj6h
XVg6uTmoOoJjVgWfvADNbNNQkWS/9KLYE+DgdNEZIRpcfSvHmQrHNYTUNTMJ16fx
R/3qLLph40Q75VvQytdBLMJBW4sdRCLMsayiDUDeUth1KnlEmlcWz3KUwYnX/rY6
VZOpNuvT6LO4GkprhRpj4EJuZgyuDPMgcqAOGWazkEbiO9E+JFEce33mqP9jQaUV
0DFQLDCa7PXANFHMSOd9poc93iThFxXLbssWzOF4B7iB4xQJ+ozbddGZ2XeUT1P5
KBRCatNpbFRjHpIh0KEDpEbAG0w1QvjcGTTPSEk1PypSyRL9064mK6rEemjgeSbS
AFNERZXiLIwi7MggBtzy5dZ07MP6YqxiFwd+jz3YNvJ6A7rkLoesKUWmOjkpMe3I
WcIujlgBaAd9qRj0VzXFFzyIFG5n5s5WlIjdAczbLUpnThPX2x6yiKHkxF8OAlv1
6zDXYB/4STzNmnVIFQMiiehssCFiLlQl8StHsy+zc9twlTrGritbEAgsGPyXEks+
f0OOKcdCkbM8iB2LaDCbYt0HRz0sf+xauYGBHYR5urPuTPB99fHUvx2f3fjH2T+s
0JKtkl4ED8cB2RiZ2vQ4HIreygPrUK0FWzyuqTE8OEqYka8DndBhxCR99T450rzH
fDf4bKBheVf7afOA7i9AK7IUjeLCKsZ49arCJ5/wguveKZzMDWeJK3291NrGOgk4
OlKe5UNXMqPsCxOuMmBjwi0VDwsq6IKRdrlDZSSb+mNFIJCtHaCzza0b/7PPt9hr
PIaX+x8SO8T5ghxwr2dumx+192E2WPWEAv3JSXUa8Xlai6i9IUDVU0QJKVHVQbAx
dYjwYqeFguxFxnbdudj9UB/GROv1kL3Ay/aGL1VtQZpwaai/fwDW4tPPQ2VBnrwL
BjP/KR18A0ArvWcwsGVSkcvsCuZggmgUgkVcS6Nyfc9E5+imps23C0AavZouerxq
xJ+2xr8I5eQdcTJFg4b2Eniy7InmAhIsW8bvQC6dHZ+XIP2+zYnblZ2k66EZzwTV
c1J8LbMbxycjnB9iqqxOnUdIj4SYItI7oZLJ3EqsyEK68Uv4IWb9nNbVM8eR6kSv
Jtp4HWYENBl6GZd8Oq9aW47IxM9bA2Aa6jQcTjKTN+Ta/IwQVvyvzUBm5OCMBjiv
XMd5DfS6XvtLl9HQSSKGfGHMswHJNRXB/YQPvKGuAI08xDinxcgM0ttMr99lYv9k
izQugTSN8tHAINLzXDJ98zk67HiFZLuNdrykk5m7VlcP6KunTlxQN1V6MVxj7F1+
WnmGvWrmPoPfi3+1QmBuCNS6aBqimpeeDXMn/JKq5h9NF98cHrNsQQubn9LvkeRQ
Mk0OXXNLr0ZR5UXDQfnhHquuH6r7H+2PdL7IpRXdmab0QlfJAVYXW/BpqHXS+38a
YJ6ly+mdtPUmqk+RDPHd/ealkTg6KfEiGB+hdBCpPUhZeRfwtxsgn4MJQ/KR6bxG
WU4bEJMdmRwnluTdJEyntVj9gXaxp6fUH6b4nHvuVYMv/YnWcxfngmBtEzDgwnha
ahFn/IBbGahHQQbXHr8GMPrecxiEu/qTXdKlL10xzM9W2nm1qsPACJXu82YioYrc
fVMUsS00m6i44hxEQic6bCpFHm6cod6cixpLUDq2QQOXxa/VMnAaUTV7hBLRICFB
HOAdz5ug0xFkm3C0hCbX2ONTARlG3UrElyB5odvoBYLF1Yb3LR+P/5Og2YZOsBow
Rxw+CIEgZODhPTouRviU2j2gOKJwLgPFGEUM1ZDWbfHogWkMmFTctqo1drdvcjqV
ZHsI8yk09bKJY8Ow8avpAw==
`pragma protect end_protected
