`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j/KrAGXYYqO042qwgogqF8og4SeprEt6MusPRPYuZjjdk/TdL39EY2DiTVQWIQ2f
JjDUq2Dnic0RkaMgkYjryhG8TNjUXtVTHcCRoDp0woXyL6mqgThvQGFRfephaHnm
7gQ+s0d34mcxyn7R1QcC43lQHdkUlBfbuiUQRfkSLyY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35504)
Gwy1xi+vp5EsmM/ZY6lBm4n69IFFU4Ryt7qk6akzztpbK+uTZjwxaRiT9JztaJ8T
kl3AJnsj2/bssOXsNH1Irvy6Jb+zsFlcg8kMCDHxjpxmv95DnFRlH8LwoHUeowrU
tlRWBPdIxLUskvYAWCjLQPJzPXBGWBxyk9PouvjHAHaWbhXzAfqDmiCxdPsyhnaM
DshGhFp2UWtT4ZXdRYLkcxe4lMB7Ug/19DTgp+FHJdsy3TjnySQhsASl7P638i4M
noYjKQR/tzMumEpzld6NJ/sxaqjzG232vw9ScwGtVcGBlpomZxTMjRAooxfqJZfl
7/6Lk/naWwbmXvwbqUi8vfiHf2hc2/SqeMoXQ4ULHtiJXipdFrSjRDBrerNEygi0
kYQ9J5zOAawfiVWZRc541VUn4gvZwU1Jc56KKi4UPRmCAVcFRuQ/5QgTfkRLLCUw
szak8ruPb69zdbCPz79Po6b5ODakGeS2gW0y83PyCfhkg++ObatBsWY+IIC5Tl5n
xkYjjxk/dpoS3KuNcSdldaN+PsYytfg/ZGGg3KgBnQ6qWIBAVGNkDKCPqqqFOFli
ZO19+yXaM7q6p74dTJf8W2me3eXJUFcoWJiLoioPHQcgDLRAapTvo53M25rOoA78
U/iHna58+yDpwECUPlmE5yDGezx5DPwqEfSmghPyRBT1/Ex5FuhjeAUsTWsgPkPT
lJ+Yj5/RtQf2bM58reEqoe/BhhkojuYrGThaIhto7gcc8pWV2mSHNzfzimFbr3ct
zhuE1NDLi4LKaM7p/KvADRUGsxxUGjyvmTBo/qmT7NM9BU2j1PymTWTjB3IRvYcV
ZK0aS0HHH/IOQ0igZ3aknjOtBF88F75fPFVDEt+jewsfgaW2yU9/GOZb9GHUC9ZQ
b5rSvBTYjh4M6r2qYjqeSntDa2d3SyPoPX9kunWhwMFVfyKuSo94emYboKZ/Gb1I
2lyh+0AyZXuRbqyrEgLbF9MFX1XIvRcICFdGuRxr7VWqB7B9jm2++mb5a964Ew3p
gaeHEZqlI4zlF4aALtSrMVwcx6Ay8LfsrM+cky/+y5n28jz3Z9o/oB6F0p884ZSU
aRcT8twFHbWuLOzXceyssVzVQkEOtsTVXvCgPABRQoV0TmlbylzCrPSGPalYbwx+
fOWaMf9X2gsmERZVjCjf5F2aKhDTR9mrHK46JMaof8OIHQYtvbBp/YE9lYXhW4EE
KaTAIfxBnqrEWBIYHU/t7pOHOkYvQXKF9kooLA3p4XoEcsGkcbTiO82ZUTKTgVBw
fTfEnbqrRmkqR7LhLAZwdc9IK+UNY5wUuSZkrqQm2IlIB/7B8vnyKThyHoqmMQ4Y
vcZpI5phV+o4pQQFdxqAQd+MvLjD/Nbfbz7GXAhFN1Ma4eNVY1hCi7+KMoR2KUBI
pGoFKrptexyivYM81qvR6C4Oi5D7m3cTW3zeCoMbLuaEEQy+Gb9b+PHJFafAwD4T
l19GWMFMReIxjS9nU0JvZqfcfLBQdYgpIs2nbC4txlATWcsiG6u9FapGfeBi7rZ7
FFYxPI0Z2Pf7QNrJdtRicA+0KYuULCq3gDD3qPb5O5q+ADTzFVOeHB4wNaJ4mDXN
ihSQ86uBCBmEHvMguiyuEZPnSSQBEiHUCJSpYSo+wQqwSOLSJRVbs/0FRgJSvtTT
jnr1MqhYu39i3P6pYqlmeyJbQIjIDyRqDNbSZSKb45XVZJH1cVNbVLM5t5st+IVJ
lkswL0OqvUy77ED0GLC3MQRIgod/sBTgevBOFqzZvw+NjdOyRTtb9Gvb2u4Al9QR
cVF+hkAS9quhpqqxyvcwRVAiSy3gkkpAk7uTZGllk2Vtf8wvynD8tIgPoFoldCXY
TP8GuqEKM3MY+e7fR9vKAR0t0kN4Nre3lBIKzfWlM7ceVKVlgpoH8SjWk/SITgTM
/sy2c8b4/XKWxmjQmhVz9RS3f7p7fKen8V0NZMeuRB5/vmHRcJAUiboDGiXwAmMg
+/LnNyfO+ksPzmCc8WcSgfAsCMeKWJa0Xh7S7+kWW2dUf9SS3KMytJvjczVVt3pc
ussnQprbDkKPsDL206LdRfna2MN1/qRsAOGKbEu/OkIONFyeSvW44h17gdDIylwo
mafClqKZtOnl37j0CQiSxsbqFC42sQPjHcF8beXD1NKeGuzCdPavdd9QQVkHX7/q
onZYPFi+9qc1TIF72QtM6xw6AKRMkOkp75NP6NEOyMgOclgiUilvjfKa2UOAApYE
nI3pg/cDTNkNUkz7Bb26nkMpKYSrtcwC+rn87D/Scur53M5eB+mLUsVNgPpER/pY
NlBJ07W/RYYYTXo7R1Nw2xFGIIr9hiqHdE+vncBBbf1DzqBkOdPW22BIXy9GAGv6
fcsPUvsbqFJZopH+UqnEk8W0Q7xakBvCXabSu2dsdZReMLzceKe1NFhnWgOGlwRo
3ehMAkt4+mCGSAaIAtkXZ8iKz3QldWN0wpT6fQWMNm/ud1BiopyJIqGygDlpw3iY
i45njQQpJztI0zfPjVSnXNcWZ2qSS4OQ1ISpk4EKgMP1HAHJH3bde3zHTkFqgXu1
ht0uEPQN1Sm9yNNvqLkjqPT9oJMFvpPtPBxDwY3cBv+Aw76Dl4/F5GvYECZidJcp
pGSddDLC9XF15WMnhdu9Fh6/qn1SWnnw5ZFTC+iW7Xrdp2Iwfnt0CWm56TWbKKwH
tTNDhDCjo9s6B85Ya5j1SqY1k2zi5ufPbNVdcz3xKa0ZKrfz3sIp331uoo3aum2O
5622xTMlZlr1S37F2Kr33j1DoYZDA0HqZ8bW2AsVpiYFfAFMqd2rIVmofpGLPdpd
4EJkb+zbfltq2lOZJXL2MvNUaEpC58CIiTKt2G3cmLhbAUEAMWu9mZMWTeww0xMw
Wi4/oW2hYb0636SXSfp2crb7i7p+2NIKFbCMoIuSIWm8lKi6orB7gLjwlSDTVQsP
hIkYYKeH4goMj1HScCJyX1fXEGJoiwMePNjFePPkBcLwTDu2yb1QEyz5ouJcbJ2G
6qY9g66g1vndf3ibq8OO4I/O7XdMb7vSoOYkz01WTrBwZx96KXZkxdULFkUVfwx9
5DshBPRlJcMwrbynVOv6ZrXtW1/ymbKMuFxI+w1OAXvILm6wBMRS+KehJp0DZGLY
aGM1avONrvG3UAlInZTaBb15wIyOiWoWPyjeON+kirz/F0ve60AuXUN+XpS8njjz
SZHVhuhLkLscrPR3jURxkhnHlrWRw8rTg3Kn7kkyi8PI4lhGje9UVW08oPhLnSz0
DBcirl8x+zmd2mRKxKIjC2EYnmf0hiTIZLvpvI1kmWc8FGe7OXu2anF8uqxAM16m
bJLKVL3HN076FVuY8AC9b8GrUyX0jovKrhsZw29y88XtUR1ifN3QCMCgsxzEjTun
r9Nx2+VaGGj4VV2H0zwcCLYSJ0/jVPdnWgW5jC3ApIgtiOKM9Wcf98dw8LLHxGNG
oEVekcEWPVr4uVUMT3Vi4wPp/PjBXmA1RBgGU7D4cxXB5nvOIeXF7/zWS7kdVYh+
PKH11AC4VUbVax3jW2wL/6wbc4ltt9iofqCvDUMBptG/hPBk6VPWVT4QPQsG5G/Q
4dUYXen4NtJhc6++GHVZ9RYCYpFkFT+mlrrI6mGHr1w0Ui8mI2WrD0tYAzAKlOjb
0/iEsKAa2SrsWccIOdPWKCcqnSq8xmnwjyTAy55boVZxk5dKKPytPWz+rnSlqhBB
LfB1hPJXEVhpi+fb06d9M1/fCcltIBa2/cgWnKlcqQdTnymNxomiAck3tqwC87Hn
DPAyLMzpI5hzOpmiumKbl/T38nUS8BqmGxb0A3Z/svJpMgSY0ZoyvXnCVR3D6vH0
tcjenKka5uBBVWMroXhV77unt9mS5iXXKFOhNDpsGpHLJfccTtFK04drKzpxPqoF
3uqJMANIKj6WnDzOTm+3OFWiudtLRdTTS4AY7IldmjEALym3Z7uopQE/UEvXev8q
cVLyDbjpqLAULMwOrv2AkGhtDWr26Rm9Bb93xM4+gUJy88bhCGjF5KY1yg/XhvbF
Eki/AceA42mVUKtMuHj3Rd/Y/Rw26IeP5rsDEqKxjY0nVMLc91ntFfzifofwNsT5
H6WgRJjrdpHIHEJag2J/s9I9Nlbwm7McO7vBqgKYm0dsv8NJ584KNHbv2atYZtnK
5TOSZKc936z2ZXSU7DnIabh1AWAlIG2TEh1qwH0n2fmxjMNjcMJQz6lYlSfzBbEb
SEUFVJcizqtuXk42kacnmx95g7VxUKykI5gYMegqQ9bfcn9tIaPx7SYkrAEAvaw/
xtqbwZIwDl0ZkY9I13F5O/im1NVANV8Qr7rin68FTnokC2/d1WTa5avR+/BDION4
ivI8nuOWZrLCKyCRorI/EqmF2godr1XuWsNdJCr2jdSWQsAwGskpKH4VGlmNkll0
h0+M3rY7Y51j4F3WDi1G1X/D5PpPD2rzyt9NoUX7RmUsnsYLNMKgNo35/Ieg/IrU
QPPsYB+b3Bw7RRj3E/QfJoE9kbpUy70NOJQA4habFNGMtnvKv+pg7/nXWDG31R8P
SxjoIRdichzWCNa65WyfW0IG6D4zeV8WxbTTT4TwT5p8ow3f7SPoLv1aln2/SDnJ
NFifsbc1LjmSbHV6zUWjntiHyELQSXYkwVPfyoMcpYy2ZmopJJXvOOnwnuWHHR5c
97Qqr9X5XNF4eF9HEx2TClRBept/VH1mld9Ar2wKJS1k/xNRJju8l7ZCH//agYJ6
+6zEfSkjQiypl5TeI5ULzbexgUCXcRcBYxz2PSsmSHueTgBhC+cBaspNUCBYYOSz
HmmKtHa51tBaqvUX9UW9jcgd+BMbR9PkxIeE4JaT8E5qjZkA7NGKCfyVBcHb5cod
30Ul58+V6g3Z0r4ZZNzleR7cBBptqMOdBG6YunYHyZ5yzBKGYyfQ2hjHOvadX8TC
u/kDahBXoW2tvpm7Q/UTAO6hhnqoIvxpEd1fY7URcZvrQHG6+xjbyULLtYbSFlw6
8XvpeisViSDXe0f00Cg6wbBbLAXWo2oNJWQy9TOaMFuqcN0zIAn/ggOBfd6XpqR0
ZvVGBKtLHk4R3leWc7qZYN7r9k9n1aTsiyIWMR2dICatq+D6AgW3wTcWB9TyqDJg
YxulMKfGPieoV8GM5dpfigzI4YwMWLftQBbr0Vtghkbk8nzdYYGv5ugU41P2rWE7
6oJbpy/Ox9ybPYzVuMj01PD4agwLKhQh+8oehmhSangyQ4w5Xnye11EVP4A6OS1a
BQ74iaWAeC9xE9RvUUDjak5aJy2gO1RuL/0s+ck5hOvyQdixpQpQKG2EJIrl7ZUA
swtCfWKV4tUMUBezwCIQZzKyQOtQbRRKvSMuV+r3YO+brInyY4DiZQlmOGCeseY3
1DgD/IuqBY5hYM0ovCPNHW1zPkYUrt1+9/DxLoa5y93fDYsox3gq1F+2zcvQYt1a
38mFvJ8r6XwVrTGK3NvSu/9OiAFEIsFSiTUr7WZnphGsNYvEmMHFfA+eY+VJieIZ
MDjw15iK4i/2HTY2ZI+bXpS7MunIoQoqwFcfw3p01Hgykfz3HDiRZtUKvVb6uLs7
tbmRNuzroP6z6VYnqAlpzUdvjqKJV8J3pW21Tl8OOdMlnJx6D+YqfvH5xLyTbdT+
zpIptfi98Z1/WxLAsyYfbMtRNcpZviQyQh5lg5HKuZKiygK7MQCwuDH4yqYCpiIM
AdjCrr4TFpo1Hi4vBDFX+thujN+Evatuvrlm5injigYheZnmq8iOQwJcSEIZa+ex
KR9TnQ3CfMUA1xqdjqfcDhEdkxQBhUWheE+IyScEF+LmbQWl06sJddHLw/oxQAuo
HU2zY4MtcVwn2NsafvDopnRO2ZRZI4NKobinbbC7y8Nf3zH7wFnj9NDKCMc2CCyu
a3wh+W+x8VZMqsTvDT8K7pTM983MERx1fVhqKaYDwwD6l56k5qlBoZxPeF5tmQF5
EKtx4ZO6/lJR1qaedHRJPPOSF14EH8iMu6pzzSDHO0ujok5cPFnQh219LlyspUTA
NXqlOi1+KUYGMQBuHoRFXyiNeyaPKpg1uMRk8c6RK3nTKsF1PcKHbj/T0hoV3NWR
1iIncgquDML4ALLfM+uGW2UDze5D87RMjlbN63dw/i1qCwqa1NccVlGSaynR0TDd
W4NamP4r6zLz9ZyFuVJHL9C7emtehIDbhHbu2/YsAAkYsZu4nPgpreKbYuojdHTE
clNDIbImFsF46gdmMrt+OAGF18InK8/Me4SlNvbp1Z9ZVOuPjHQaHIbmBxC6e4Uy
a245myHgjkWj6AYrBQ7B2oYT70jTAwyo+nr7dnJFRr5rVFWuFKC3AinBtphwRI8h
gtiwQ8j/ZMNd9xWxEyZP2uEhVK3B0OkFV1YhOIX7siTA4n3q7CAVjKtuWK/Ofrul
yB3PWAcZFSO9B9d3YpYhIUvZkhX6oxr/MRbCHDLLOoP/VxFVybdQV8j4b+cnFifU
JCWFdoDL3WV/zGYnw1PC5jihfOSzD+6PwxT5c6TwZ6/x78C5dLUocdITBx2+/bhW
WmGzhDHsZ0Aiu9iJAVIaCgaDCT5corfMXdrdIQvebPpCMluAoUdvqzKmc37VZ3zE
w6+f77POebS4F3x19VquLgqkjr4CBfdFqrB338sHFTJL1ZRp6pqvK8AwbEu2FO1K
tH+q/ljArUOU4wilCt6pP5xf9j+/Rl+SPgIw4+Mt5ojW6X5cK/ZRhS7LQxKWykLl
e3JzZ7Mt8pg5v6JSs0AX5VTEe2cigoh5/2bLI/aryHgYDms+YLrfgRTWRMUJ3BBw
EHYfc7mc2PZj1Lb7zk0IyqQD8mn+Smf8tA4rYORyskOufzOZaGwG7Q/GCHGy4D6q
/OL/FIHJL+3yuhOY8OpXbMwT67Dio79M374vCaiHMixpfrYp3ZM9Ww21rRHQvA2T
QzI9ASTgSgtDO2wjb7whdv1SqM/Vc1weR0x38Qis1nPWGWH4tz2p/dfp2HLuXhA2
sj+10Gkwc4JTr3gX/gp4nUHeNy55w8k+mwmRTDYhduDAc3aFJBQdR485rw0PNmo8
+FfNz2n0lbyfxnUUENPOzQo0U4qwrhhvi2U3egnTZh8s5tNI1yBG/g+S8s4vd6v+
LQebAy2p8j91aaM/Jf8FAgk7vhNT0TouajdipKexXKSznRFCqu7/1K9GuRE5H9MN
7uwbFdleCX9QZ4+t1Upql84eT+M3Qcb+QQRlgllDxTL4NixpDlzR+5Az4e5lSzcI
6PNSYeJ+97+ipKQB/08EF2KPaEoqOiGUJVeF/OjwcyK0hQYDeKEbSC73Z24Slb9Q
hXbduVqWJrj2yuG2vqhvPvDsuWv+MaiJHOmGuVmul5HRWXjCNEaCTO14WRm5ugUU
+ta0wPw7OoB/Fu96kFu55Fk1e+TzJxomhAj7p2gzMobZDr1kL0sBTsPRAFfVFCrC
XD293fJRa71pMpsAGknsRVaxMAkFIhoGSFqsBUV9iOK+7ikegEzAfzhXV8ASSZ/m
YciO49KoQht5Y4frpFJYmeDsbArofxLBQOSXbVZyKjmo2WEvdV2F9GyG1YIkiBpi
KRw0YUknQUpDsoxbuVZh77jF0SYKGf6eG7ZDqBy2P3lw3JG6pW7VU37qbE/qUAP8
7uDw10YvqMTrX9kmRl2KB5HKQreawND5O7yNZAza/OHdGdYVfTDX7/tvM5M4P23i
ugGIlYxjelrE6gmsffQ3QTNb6PhYSwnbyHsK+MRdPra8zXVScwyeePIAkvH2gQb2
e7gDG9W12dUxyeISRTbY08dLGX9qlQ63FHfUaUuO9BHMJC+eykSnYoghAVbnUimy
f5nM2gL7kFDjZumr4TCV+7lb6dWoe3N43v46kf4W1Ik1ZmbxVVq45NsKgOlT8NWZ
DrsLKewdqW6gsLUI5aiOQIOceRfBclPAm9/0r888EKvsO0opB125bEdEfJlNphDJ
48dyEfUvyajmhUMUuc7cckPvWBNfGWaTVRvJiMDm7TgA3EqpEjuS8lSCOZJm42YI
cEfOZ0ctyINwa4fPpPqKXSIuZB7Us/JfEqJH/Msd+O3WmcVYzwrAtHJAYlCXNdKv
jCjmsq0lio4I80ruoSMSkq5/x5iBl7Mlr/msaNNWCTDQTYLJtiejigh20NnReQpX
/Re4tbFx8g78w4nJ6ZDpZVp1RQf17qpBUJA8de0ApMWFbAqGR/vHNerKMtEvJmHY
3h0QUrtvd9kJx+JyYrpEOMwvYzG5cp/KWSdGfBX09KAn4qwz99vJW7MFURNgDa0e
Hjk9ApD9bR29kN5cF94Wn+gQpmEtZl2ahH+ltr7vPw47itaLVCJxlqCHHxp0xx+B
CBvsa3sxcVsN3jBN+AhqyFjGwIaSQkunfoNtkZtyTpprakf35z7DYHSdQJCQHANU
iLpOp5qkx84Er+nFUF9wTis5tVy/yleHPGS3kK1AsaFTZQFjoOZQGNa6eRuB5V56
i74Ph0cEkvBGGua4OrJGaNHqMWJYuuVMUhG2wWeWFGFmI97srQjlITDUOMT26aXd
WYnQxh8R3FKAA33rTYk5QguD/sAI58Jc7jABccMpJOs8eez+OEb2afXcw8KNYsYv
uGzEaYpavw1mWEJlnABVvGAKo9VgGJwaOxLVWdfjzYhOW+kqMsqgWdgeX1nOftc+
ulz9+bGPVGrV/I1RK4YPMteZSviZki1wPCd/oP/RDrpnVzo63ZggXn0G7z6kvkDf
D+bXngWESSjUKtK1YD0VS3u95A3MEiRGhGPiriLwgEXpLsd5aQG4I0FylKFm1u7J
bmihnu/bcruTV5I/iGAJ7kRw0QHcKBaWVmBInSsy4FEzaQyHkGct36UGzGKNbegA
OEiQU2tsfe+c86dgKya5KgHWQBT7I/X89QQK2EzKOo+yGtgkw91YvCeg60uB+kMo
9DkMUpSPsfByJhODn1R7ycC448BB4PnFRlc/XZdrdOfpvIF8uCZfw+PVfwp8dwGM
ln6LEZrjVEcmP2/tDbFwjqJ7X8VGF/S+XEhFLwt2O2TT9ktMg1ls5qScl5A9SVBL
TYQLJaMXAda38srRCGcmuzdlQMQkQ5gnZgioe3q0bhAnRm+nhgPjRI6UkDLQAxAq
3omSGL+QPFcSCehnm3KycnXh8BMShl5XFyisWBnlX7iySieI/Uan1rk8p/3IKOdi
Wf1smnv19l0gJ+OF3oJ1Z86J4f99Jwubo85SinOrPLNQXEAAqMtI5j8zV9Z0ekUu
2/Ei3Mr7nW2pma7/0uXpWWA5gh61fXNWw1LJlLpSPTB0A3XBLJ8jYKLC/55cvm7j
bSTZNuW1tKA+r/HF1Cxt97w4g7Gxpd/5m25A/tb+OpswIGCGSEIQ8P7vW8iz91Of
ZXBP2xhE3weO3uwfAUSwnMBE4y4kQYzcXgciipvYABY8Ft9NX9SGWZIT9JBWDcJR
S9SvAZGpXE9yAyUJF7mMMMDd5fd3+3Z9hVjITkCpR8KrRvwJAFXlgkppSr2shqXl
L/afD+aER2pUJKvWcPGkIA90JC/TXbvPinXnjML3vAtOlYNnxttHOkPRULjG+wEk
ZuY/um23OMzJeA+K6gQEmX8NYsgh5nk4NWQtLzxaa4kHYK3Fofz8rak8bVfh9tO6
EKOXNxYvQfwpRxMNQJx7GN0rvPibk/qovjduWuGc+2gtCGXfJ9E1tA3I3VhksOrL
tbD8gx4WV5WxMxCQpc5O0m5LYiJs3F6XeDDX8utfFa0xhAMhfBj/aQCnMxr5adCj
3umOdln3un7I0E691HSZKMiJKnh61tJlJP5j0xoX2kNY6bGHcj+nna1EAsx/tzAh
ACiy36gXqWwXe9LqJD0TLaY1blDF2NJVhHFDQaF9CSLmg+YdQBsMHwqgF9iULM5p
fmpy97gchyHMVm0UzC0hCtIEXudbY1g7+Cy7e6GW513Aa3ZrYBa0CA82y9r/zf9y
s9GSoKyoRn3DxsHX7ovCKy+b77fCEEHBxLOOihjE+XX5DKtytcDztJx2pGlvURg0
uKz79kwLPQCy04BHeUE8KxSRosEFI4pNDieBc2o6CDOU73wgz4DSk5nS+fNZ5FWX
x6qx6qVrb53TmtHM3IDIm9HmAEYyiif9dHPkmchy6oamIPph1BKWa6Mkqll4L7Pf
MXFmUwqZzUBvGhcO4Gyczrdg7NZODusdtCevx6q5IwXUKZJyevg1WhEkV3yFxEFc
6zDiOZC3nNXewjSMJjpUZdagj+HZ8+9kgmLkF5G7bomivOC0CZS7a3agIg+Gdc2q
MEBXUQvVO16uEw48dL7f/nGSsXhuXMkQjj2Hm22fBSiUXgPzTphV1C3hHZGqJ++O
TjfxTSaffyfeRn7nLaszk7DQFHV9rN8FY7HfSOjv56DuNHFTLFLkAUd1KYHF8WNq
3R/FmZlYTgn1IpxJjZswWCxU3tjfh8qsFDpXrTfduEYTMGCsxlzWxIszdiS/rpv1
ioMU4bIwDfpDEoKHhL8wwU/5/C4BAZTi/ccNhWuB2LcTMwj39dBmV2Zgd9Vx38CQ
AZM8JzYU6qKlDBG78btapVBZEjeDnCC/Tpqgw3uyFLIV91KIrp2lAbOO3c1o+1si
p1ha1fDJqKnVR4BkwgIXvJjd0mmjiM3mYqt/OfCGKj1yt2S7Y0ssjlhbV1ESNTE9
QJcer+Kk+/uoe9LDvkTcGv8oN5HLcxLh2IAdpDhirOizWgqCmgjYd8eJzTyCMz4E
/qfOQaRwDb3Cmdq9FrqEF2u1wETJmruRQ1k76m7dfxCVBrTRV/A7G0FAwXprsH/k
MQpGQe92M6KuPNmVr72qQe0/j9VMAm+TiukRbWB1RBd2kVQqoMPhhl6PoE0HA0YG
u6HDWginljuBSyO22nRa5Z/7Zgvr4/fmNAKqOjit9sR9biqSbAwAZiX2UuN6HynF
C2lsVlZRpF3J6LBuYbBsfbJxsDBgZlGa5djF6L6lolccZHP6l/NFiP1Mu0Zn2Lj5
k1n8tGOUFwNv8DhhbYT5tTeDNe+utNa4QxUuTx1wdzG4SCzVmXfRO4+Z935Sa16h
+AHCy/Jpiioo9LhxQ3/M0dzxIv4FWIXIu2a33/ugOSDUM7IGFqDSDsvxFvbtNXii
s1YeEC+jHf1dwoDM9X772SGldBzMkPmrhejLCcbRAs0aMFovcJuiFuXcrJExzQE4
IKItpcglbn1eO86YNa9xa3xY/z1NtlUP3K+AxhdTYu5YFQx3+DlZNQY9YrHMLYnb
nEwcfK6zXBWZCAi+R9A1g7DjKrqs00A0mIAmdAIFwFDD/siUA6qbxkvHVBKFbdsc
TKewi/WnGvdxNxdxsV2Zj4RcpkFO7iwlYOgHjaZ79hWTfW2X/Iyo3q1w+fW/f6vv
oyPA2atafGtsOfndl4LGUsfiNOgGKtrCjfd6ynArVokaOhFPGFgwCaY/6z3ItqIG
9OjvSxIzrl7BEr9txET/7CC/0Iidc10xgiGT24QOHhZYk/ozTjrHNagHy4GNLQ8W
F/giX40NK2bp8R4SYVXCwL7dWSlz8YvVSJ1WzUXGZljXumVV5bpAG3mQxTmCdFp4
DC+b4XI0qbcPalNfoDbNh1r+oD5I8Pt/4ct44KEc0bSNIi5pt5Il2d+sZb5ASqDI
O+LvnNVQtYptfXy428af0r2KlXL/CjN3ksEsOAoCFyUuv9/KW2AZNaxbWfJj8bmI
xj8vklzasOfr6PA/TsGhNtSojDHKQ8R8hJ+DuZV/C9LsjEm1TZtmJj57TQ3jnTbR
fIK/GqogbPJcLdv29i3sgB/CKGv6jFsG0dTzcpvEoZQH5gl0tRMCepmxKD0kR3aD
7dc8ALakFDWn7novYaT+Gd/ayUj3R3uKuS9zcZF1MsP8tEe1QR3qLfICTu7XHxu/
8ubZjpCeJFBWSQ/uskIetfHtW4xw8geafTFrws1Gsr5QDMchzbU0Hl4p8zzdQyWx
WGzNqZPLEGykU66Qetg5wAQmQ5FvWf/CZ/djDvL/URKKWdreh3mPQYMOu8/4cEb1
Yx+zyHUJcZmAb+BIfcu+jt18Gh3zMWzRSOoCbJENwIJuNtXNiH8kWEN6WrT+zYBu
r/ZtXs1N7buWJKAcjvKptcqT9eEptic36FNjl8pb6PTfBFQNOT2rbtUJneVWl9q7
KF1Olrgp3bH0Av82iDOrLgFpMbSige1llfenHj9x4vPrIMN6cCp2P3TjDxm0Byr7
Hd3LH9tcqAqGx09yVScwoSZxldPAAPhEE0dmZ/uWv77lCLP09HsWR8tO0iQBoxsy
tSeRVUcE7EmLl+xeTjVXmMQm9ctbHpQAw3h4o1fssC41X2aBbHXyiu23hDS4PZhM
t9D1+Iklft4P1eqhfi7BQBSLlwCZbxmLHtWOob0u9DAgWQXTYUwL1vILhTC/n6tg
p+F2KsJelAYgIVbZeSTw16S6aUdML6PwIgSJlLgF3+MUAZf2tTFtUy757PRFysVG
XDbbUvsqq6h2S4irtrHKFH3aypZ8cOcj5VNmixYzCeCcndZAO4WkBrEzzINBjgV/
vZ+B1nkzeLvnNTtNO0XSkMDlMcMAEFFeyFWQEgLgHX4GIuPF/8FFf3/j5FLJx2R4
+VJV2tcDv9d7lP6ANFtFpv7h2znxOIGWf318fcIjRWGswyFyDEUlWRISssS0VHMI
+LTXaa7KqPDkAFTe4woVKDopxz1KNgAfO/CDmc6kFRVXruewo7kE7rNKGOZpGi8j
NTeZu93llvRRDK0DnoM/oq87X4ewdKiwf7ioe6HqrLm+NYVOZTiyciPDDZNbNk/C
82vgTJV8b710z5mo/esOLokguMKVJT/0N6Ew9Kz3KaVomff15TIH++dZhYfDbSZi
tgdjZsQU5Oop4THCjuuUK+vKqLWu4eMuvam268eB/4x3NtpinzTegev5sF2wX+Y/
Q9rKEuqQ7eFTgXEfoAOFhbJWk7uY8AL7vkevDW9/7A5FTnwM0MbKyAljnVjQ0wEy
slMkRRLdvP8k7SyX4cr6hqcWGGOAZXBUYgCKzJA2AIbW7XMb40Vm8DZi+G6x5iQu
QjwgvxqQ6epF6gwXaxhYe5Yg9BxkC+dVPxuqqRWXbwbYIumyiO8QnboyRs2M8ZPq
F932EIj2iVmJaqCsAUh/k0IWg8pyB4A+cR8xdki2qrajv7L/LeV31dRP4bs7wkDr
XcJmZTEETQvAWfGh1oGaLQs5veTCFb521Bo4ZSNeolcn/vAkxZdONmlo5ZzdfJCE
TyNRTvEGrxfNTe/ZLJunJHSICPvswVBMXA1juz10ZbO4T8Zqone7udh+7QCnB1++
LYQliPltAxq72hxTr9c6zO5nwVdD+ZtlRXT7yh5OiF6QrmTqv/9PVyc3DSmOI+Tr
hJT0fwYLQxtoh3jpb3jNVSkEr3cRNQ1ELQA1h3zjPMW2Q0/D1XLo99KZgn/2G3OF
ggiIPORkaNAtfjkI9MXFTY+qEtJr7mFqAOP22ZxiWgAhoqKviaD5uSkmzO2BtHHO
qXNNEz8tGOXKk8tyMD9J4Ql6QeRFUahXk3t0GVJ9jQw/GcPNpsDMql/D+kD1RkP1
ESaUvb3I2nffNcTEo5ymYRTEJNO/F8MXMpC7iVTUuVxYVe3+MoGycmvZ76q0EUfh
iZhmF36fT4bX/vMGA5V1ldawdpEcbUSzrdJ79IsC3IAYj1KRvOgOOYBsdcmneXOd
6uOjW8bFRY2mA/V7Jq+G6muGhaZq7o+q4/T/g1ZIXc8SR+JNZeQdZ0geATMjUuyN
8gXSyBUTw6bImuiLi/V7MsEteFneyPD/9oSLaTVik5l6OL/tlTp/uZsU4igELCaq
W+ltwTEEj5XOW1JW4Cf2wc3OTt4qpIAaLQvo/bMVMN8mh0s4kRkr2Vu0+5wkS1aZ
ZTE5hFxecWwC5AlXOyFphx9T1jrAoGfi61WUPXPSpCMZCWH0R0wJsa9QPBWv7TPg
PWH2W5z19GvVRXF5Tzdc81mSPQXExOh0NLuhmHUCpDpkaPNK4F2YKyzka+dwKSdk
2GdwDnNKQQbbRBToso84A14n7u7qYQ6YqB71Y94F+9DBiMQSNxUoTrMvH0bQooPw
1fVZ7M+NTQf+RbfAmdPs4sjquDzWn4XbGwN/RtbRnv8RFPEI+ve89WD/Twu6OWnv
dZOeQmFhG4ePq+8lIRn95r9ETn1uBJME4y1bUBUb071bcPwbOiiHptGIYUDlF/jf
dp2SQs0Qlw3OSHuSp4EjxEvd3d84tRaM5ipS+shiS0MheLdzettrm8+qhZgR5Xzb
XeTs0Y64NrwF82jdZjHe7mUxLv6SiKEs0QC5QBUihkpr4u3twGrdbHpXnzd807ru
LCdbJaUNECCY7rxuydN7T4TpsW+yZkIrfaLOorkJ+qa5Xn4seu0jarw/PMn1QSAm
6JNHhpoGrWMKQKk1/j/FQP056WBJbKEguOfw8T0co3PrTwub8A2wyCK5hSnKdZDl
TEtXQzG2077qwY9mv4VhQB+jlGsTWfwRx7DQEzI5O2di14XsmCW0UYgMfvFiCak9
0idg8SOTkJq4oM1xoeee0ZUlXYi3oIbucWnbLLaOgebOfM8z3JkEyTDN2UEnGH6I
KtA7LcRYe13cvFbPPx1fJq03PRWiRYWcx+F/2URz3xlIwGjGfArQf819+KN/Vt3e
3sNv7Ep99bZCgsHjjH2TwrQfGVsV1hu1M4y58iQAQYtInLAVZVfWqYcLlzX1BdKw
NoUn7eU1Rvo2UdYIU3I2nhHwSXxbUHggimww/O/hH9D0aWAgFf+A3dgtIH/N0A+v
SzZ/ktZObYcZ3ChMjI757g9mfktIapAMA/XdTvjwUrQttugJ7i8Ow24a5Tzi7Byi
xK0qrQ0fY96kamAjJiuEIUuCegjIvbZ9x13vo5yrKB/KIOSaAZViwvHo+FWY0Vvq
vtIGljR/bJoLZrzsW96x7oLoE3HYMpoN+OEfTvPSmS3Ar9WxdfP6/wdSF8OUHwJc
A5nYUW9ppSXrrCu6j6KHwySEsa1HiIbJO50rD42DAf1hiarXbYAe4Ib+OfOfeM9Y
SGH/XlGXpl0q9uMTSXNer/cQDNaQ1eLec+dI//mwZDA74xGWJlMUJOZnIxhJvHMc
cNgUX6LJI5fgbrVmKtL66iB8cgVacD1EuiM1UqYE8ohb0oiiml97fXGWm5uufHeS
DyrkdKQBRnMgrgfrBsWDNI4Lahq6HAw79z8K91ql/XQWH9wBdLYPosE/f0w6Rn8X
7z9XMrF1KfbBBtfZuLN+1uk3WgPuUdZar4d77J73Oubkd9rcHF1atR3GtQkxEnm+
CJSfx6+VsuSA+WbV0qEeOefcruqRxkW1mNNZ9T7Ij2cJlmcLwkzDTVE4jzMz3VOn
ZIwfLzXI4KvrT8eWykuPE7GZz+c5TLH8PG11LIFSNPy3Qu0rblcZt1dIHXKbDaA6
/MJluhDbUj5sebEFH5ibMYYz+jCYrSCpjlCXYNu4/VLhpS58prkXOTpsdqOLjRuc
8Bry2pTlg9zokUUdIoBazKE5Nv75/uVFndWW3cPRc3+M+KjOqjAYTvBbEA/1yO5k
osnqv5gyr/JGwHLHKDgH43fWp6IbJfZzYGK5IGh28vierQxniINfUQOs/2lyAVK8
Iw+iHdc75gb5dp/EKECNZqDuebvE4de0dLNQq9qbAihiD20ndaEBYGHkfjmfG0F4
PvHLf1KAirAaPqSENw5EjYaYOoeB7BXRyPcw5LaTQpJEWEklXuknhRSgRFEVrsFc
15isJXgbh2LmTAgGbjTnPLGVAkl/IQI7VA2l64yBjXERmQijQZTOwH8SVsQ1yM1B
jeatHe9qFlK3Bn/St1gkr+jdU13BOjscNeKB4CHEtA3anXwoDghBFdOpUbTSaQKQ
+c0A/NyT+fvtidZRCEJ6LBVqg7X6a9xWDMDx1wAVQL+4NtuugVn7VLcEsh0eHZpC
QdxLur9wo+vhS9IlQ6aB3z+uclCEaoFnkwMrnLX7wdiNSSKHELMyZ3nuFeI4SvAZ
cM7hd4AX2DkK/wFiUqF69PaE6f/Mhduyz2MOmVRqJCN2PiA0aIcxqmd5EbCqJK8t
Q53J+cGvH9b49VPcHhAAXPl3nRRFSw76HUypbS8WkST4sSkw35k8SXBHYpZfcKBN
6tiWhMsbREtxL645soCLuKy2fQKt/kt+6fkXQsKU6V1+x1AubsjaM+XSs08n2P7g
QGokCzHMlE51SIlKFl4WH1e1el1tpfL/RQpZBdb3kQQaDidIgI30wQ9yzmK5uucB
gWpLdYBUFcv4YhlD3aSJNqEvtvhJSDo6b3a42q01JAgn20s+AE5e6uyZ8XvHnLFe
SFVkVR8JMSeTm/Ysa37V7ThcwQZARvkEZn7rk1TR1OVTLGOCwaGYgdgj3sAxjCFZ
kijax2s7RM71i95EpcxFwrW0opwjDARoU3TiplSKGssGUVvO7QicOAV+dTMrKn+v
NsrvVL3rtP2uktR8Qnud72xyZurL7WF4we9TK9xApIFfqcZ7aaiSpdRAqWx3lzbI
X62ydK9FYt9jKf3TmzKs+S9p22lXyyxhRdJHgQt3adb18t8kKZXVUAIRq5Uo3Dlw
ER65MfuoDNn2JW5WJRQ1Ph2E/rW8BjNgBPK/sOF2oPR5q10LIjzDv/5o2v5bOvUZ
WjCKiwUsJhhSRaN7UPM9vdZ9wuvfzNb/svLaLKq/Lwx2mPPxPPPEVKndAsMXKlaE
QmQb/gXH8oYbBVRBhJgZj77BouyJgK1kD+7NHzs2nUsyR9Lg7zFg/JcglPBorxeB
wqqlnZ8xTTmQugzWVMgS+ZdR/m27qL4BSnJhgEqVAhEKFAQ8DhjTGsm9NqdlDpsF
WlVp1+Js43Kg5MCdpTcczRER4d6W968zJ3x4Jpznck38YlCHie3hgJxhqH99HfuZ
zRqdPvpcg2xynQFmaTMjAIMF7Oh8w7UN8+HyNijT7zvLKIyYrakdN872rbJGOnGe
HHTysC/hvBW1HWxElcrC1ugikGUvk7hi1G5uliEVK9+lbuXl7n3keIQdOc08Aduy
Y1D6Q0bzSpaB60mJuBuueiHh35oaJyX4hb9rXy1M0uIHccJ8qs4zaeFBYRI/6OTR
R1Jr5tN7yLFt1QFdnxvJ8NgSFomx8T2aJCv1EA3mlrTIhK5MjL8eU3G04n1e+iyj
+EZHjebPXgoAA4QYW9w0u/k7khivQmaMKffRSjdUZw35SMhlNqTWzILJD3T4UaEH
cblwYqwR73ut91Qq+KXFcBIx3r8D5sjKmfQJbMk1p75DMJ/JxmAGFcewurXvXncB
xOSQRbxVoT+eLv3KXnGP5THMsQqw7Mzqt6/qXoZIgy0h1sHGbbRZIxmz3wkSTk2L
4sVxd6DiPT3vVAVvdoQHiPUGvDHzTekDsFq8tlflbqHoZb9nB7CoeSpiv787qD50
i+dxJgDG1W486u94L5a55YTASEv00i0IZc9YA0R1IPf+05JazUdiVDrgkOX044tx
0mjkujl47Xk2Qh2n0Zwr00HeRbWoAjA5RZZ2T+vUllqway5rwttAl8sBooQzaUyY
+Y3CECgASxNwJLp8gce8LGgRX28C6EHRuIBiSxrqtSdBWkZxj0m9qUPSJPb15Yqi
6XASaKBK9+E2K+fpDb6aiRiyLBcfGZbfpLAZqfzVaLHUM9t+UelilAg8Kv6aQ381
4G5/1yNNJAVZMybWtebwuVEAFvn3C+muVByxYiX3Zu9kScl/TRZGzgpCHqqLHxj/
h7kfLx78mq8zqSpxqLCMq/l79+wgepPnThnWab1G8gIWL8X8lwEchhFdDA0O7kAP
yJpwSlwEjQgtHWC3vwQDz09kIGsn82tCn01ETuwbSQG0+JalAXTFBq1F6bt41cTz
rfeG1ELAvt3/Sn7I6uBFd5fR0LtRd7w8e2P/tTqVJppM4HVaiCtzdDXSzq/M/KD/
TWRViNU++L3/OBGz43MeHxMV/xtbKZwvSy+DxXeqHyk0UG6++uybe8mFRZTj2qCm
U0y8OCXnFQYj0S9vQPS1wLtNYNDoMfHCZDCPIB6wXukVZjNX12d9AukiqlXHt9l5
am6HOU8uNcPAC1pH0KXORyZqUvMblofsVN4LdZRsPGaG3EiDBl3PN6Zl1GRmCDk1
DrgpfbKuc4DJq8W038osGGArXVPIA53dPN7zlHrz0la/zrcRHnzqDRMJ/Y3Ig2Rz
Ii66IscuZ1DVt8JFUVVftcB763ZVg4mjTmS0fmm9kb9nbPxPBC0jwkkf5w2vEGYo
9sfrnbVu2HegARyF9QqlZdhtbGMYAMH5uwo6HrpbBDtSgUWS5Hn0vN2H0qhm7FBu
iJ7QanMxUf1vUTB1a6nQh8HiUNX2LSk1QtWCs94ZdthSCdTPswwuuNSMpTyAh13A
jn4h4PapUQYzlnznYO1rc+78XGVJFDMjS2ZHm6Dqduse+oPYhIMwaTfRUi59pjfd
oehEzTjLMQlalXCyi7Z8cxIpuqD4Zi15JEP7QzX9xnwlbydzU+Ro7cDqQ6DiekJ5
0Cmj+BYq6VUr2QsQojs8x5eMdVYTxyWJMnTxudTpiVXQ2M27dAtWghYeBl0jUDAv
pEwgQjgdJhzJMPniKiPoJJv0QCHeJnNVK1bsklxZT/LE50pQgsQs+OQFkJA8/QjJ
9AZ5X7nFKN0/noAwa4L12w45PysubnKP4nuQkUzpPcKTCl+lFt9QVsChKIuvumCe
3oBmHJMi80vq+sKbNaHiCPeoncAeuK1lhfcC9cOUULViFW2AvhR3KyyeQoKmDwHT
qtdGSgKCZXUcj4CI4/eq79tgiy+gYnVe5nVG/lsddOVZtlDk54cdpmJprr/Hr+Pv
ugau+PWsz7VK9OmkrcP4O1OPvRWl/dwcCv/kb3N6h/eS0kYF7QX2ec2NPTcFoqk9
jumwbrxoTB14ZfDCP2gbQrII5THJswtVj5+8A7s9tCvU+5DbfsFccCXcXCA8WsvG
IImJ+xTq9h23CAYvwiZ/t2aoEZH45bgzv42z5MNiZQnmcrj25SUtMra+O2ZMZ9Nq
vTS17H0haqr6akEhAzWP/0sVYr8z+18L6fUiiUndxj589A4RybDPmWoRHNT1LaL/
qa06614AXMOELyaNc3wF5sZFWKnfB0i9Ope6NOqHqq9GDd08ykYM65QkztFcSzEB
lHBAH3S55NCfdM87bpNEZBIl/QCl/QqAbi0s/ISrcePxrTfhlRxbeDkSmZnkgD8N
ocE9udDbko8UQts5Rv/G7PObIUmXCLppa2JDm/GncOaUIMBlu6JSJP4FcGAz4ZtW
fHytxlJysckMc76SKqidlGK6fUedRXi0EsG+2NP9J4cgCvsF3D45/cn2C/OwERVC
8Yq0KdKqW75l955v08I5soWElyXzXdCB/QU3nMchhGBaGEUNfq+oY8lzXVUA26o2
5itNIqxiyp7ay5HMsFCCPsxXBaibyrFKpuAuQLylKbLwDnODB0XYBV//icZ6n5uy
K+NRecItL/Xv0UwAy5BrzwyU7iH8KKY1oIQfxRSZEOe3XfR2DV/gmRCrOFHGhmE2
eI6ob7ZwdsCdp3VoRz246DpLvSzro2GSo0GoCa4QU07GEGMCY83Ee8uPjq1H46K4
N/d5sp/Liy3VMIPqJxXgmh08aGVYxPwp/UFAl2ie8EYC3EfX8WRykzveHmcvzEyG
+GYYeF1To8XLFnvQBpW0UpILh8EqAlU5Us5UuocayuZasCM+a7ATDpqGObweW/G2
wY08F071ZgRPOTC6WtpqDTrZnrBBBN3aLTcntKebHvvUldld5tNIzWFsPkh+Fy2E
7VJ9qXMQar3t/nlIoGZDc3rAc/PDlplY9/+rtUvnPR6WfUXhrnZNGFJUjVwVM77u
WoiMEPvgzxmx21Foiu4mUukHi1FtjYJudTAq8PXnNq/CRHBqIDAU0fpfjd+FJvw4
lZyYQid4UpdP8etEgoKsRMINHh+c7t1xUNdxSf8SCyBwZDoM08z9KBEVJx/3z/5s
J7BCWJ0O1ZDV/6Rl174RlMYa0B+5ZysZ7HLGvuCrK4UrXHCouj2g1tz4cYRg+jcy
z1oGxbUMj0K2dn4bg1kAf4XtbDD803lU+goKG5Cs4pdnw+fmemgQ3naa88E/FJV0
rsDhVBZp2pB7jiruXz5gVYPi5QId+DVfUcjJhkZOPb5UarpeDlEq5IM3QSic69na
J90feoUQMqQdjKFflkAadpDncCJ3NHvkgZPikqFGA7k6Hxy4Y2TMutAxEk8ThLVj
e0a4KeImSLneobWelDipDI1hGsFUzLxmKbon+4tT23QR+oAuowzGxMI0XZDQtXq+
D3FQFwAkmTGjbrwQyCE7Wg046kurWwQ9dpxhlR0ZtprDcYGgORrNEHQQw8K5wEAc
MH58F1Waa+i/6+pPHGmiYcFTsPVx2wHOpuo0RJy0UQPjExJG+3Bhm9z/wyvY4D0T
qlQ1dfqi3K7Z46tpvkeyiFPWypZ6w2i8A9/n7MZdfJCFLJOqyY4c7bZZ4p8Vmm0j
siVB4Z70g+O4bm9Oi38vaMfCZ9XMQBsKGaeUG6AcT20482QZScsKot9ef7N3whWh
hIXnWf526hsGJMfsuw5JU1Rq72oycSrCQ79+gnqCdM5LSyFghf8CFMK6e7fSomg+
TAi/0UxmjhUd/ywWER8tyyu2aIb0WCxRTsoviSrshjrqPWX/FbvhdhdhmjtQ5Sgn
QqsGWsrDrnlZ/TfZe0ONJqyk3mGCzGzL1qAd4DmpnFMIyiAP9waNAZwkP8/gcyiQ
HRQ2c6By9wpIQgw7M/obqnZP/7eM1fDxudUJ476WI1mw0ck7H2gXRgVFjIVuv/U6
Fwgem7ANQ2/QZQRh2Z1grP6m1aAoovi1rAsvbFIhWRj5oL130NMOcHWCG0nELzrp
7nIRefpCvyOklXIgN0PGV+YRX4qhSYX8+6448/iXcTPNoGoI3jbLlqzzgRC0hx54
kWFIvJ+DKaKkAfH1lmvc/ROdoiPX2ziX9pUiDCpgeeAQ4WclEFvyTAf7Np0nBNG+
EBaB6aq+KIXl9gsXe+OnqapZDNkgMZ2Z16tto2UpeWwmQLgzIntkqJ1y943sSezq
K4lj6CRo9aqnbZP45pmd27X8VDCVPhqNsU/0GU4njkLb29L8ZkDsAQesyhTKDADG
ANGzsMQK1v6AKQTkoXf8WKsspatJDaKkdjzshueMqOoqmWvY0Cvd6O6MIAm86bA6
gccbeao70aGj7ShWk+C11PIZuctr4gh9DX5aCzBhz5J4BzDO9OPdEX6zyDDent2Y
m/dG9qLSygjXUFevZn4r6J3Xg3r6+4SnHMy7uGjdiiTD8D3z7Aj+yCUYWDzxHUig
zD7ZsiitXKs0msDYA6KrwZO/vsLhBK2JyeXVVasY9/+sW1uo6KyhraPX8TGF8B4B
8SfKeJGprNmaBFQlsQljY66JWOQtW/LOlHW/y7AENJxbScYkOC4uViYBwqSgGZZg
2q2U5ZTuxuNP2Nb1YZzWZmT7h9rk4f0CgIhz8CE5KSRIeZ1SDKu9uqtFre0z6cDW
Vf7T3h7AjSDl0CuFcE5W6CKJjF58Nse0JNZwcLNjloWUJ2SJgR2aWjF3f2F7dIeD
07ZwCyTnLAl2oWOWIOkRUFW/Awm1+or3qV4iov/v6ymlr8sWUy3CMgxyflHeXeW4
UnPFXO7hWzuYWR26tTcV71UJSqUjtrj5Z5X884NiKBoS+bVsrC8ED6CLSaDunFC1
g4+4QcVL714aii7Hsmke84hba3Fdq3MblXh3dLi6jom0gyZ3z7EW4P3Ipc7VbfAy
7LvRS6P+36/32gbxZpZqElM4R7q7K/dGNMwSPHo2rZyA7hnIG/E2D2DBJmbgnmNw
A+uW0lcTMceBkKtZui10jkll2BqlhPqeon8vPI3k3zywRpstK8oz4Hwc5h22afUn
g8nAu33odt1xKbK6A55LlD0Fkcxm3PClfYUFHI3jCkd1oWeL3hYvZeo9NZDYqTRT
KJvK+AlqnJJ8bOtY91uGzkj2KCYDHd7w4sXU/AUfxcNNDaOT+Q0sR3FhvtbCuz27
Hqd4LGMGnEkOwKWqsGgvTQVacvVAuemmX3//ch6CcOovOYiQAp0CITGpnp/adGrk
QoHpi6JyUfObRtB8HiR0F4ruhVaXu2M+gR7I0EfAna2dukV71R9p/3W1NTONJeXB
zh1VDjg9i5Ww2evhXC9Z9Wj36lGSA79fXih8UXMNrXHYMAEu1qeYsMack5tW9YCp
R72EFWMv9Fg65dHNRmlP7hdyXlMPfWWMMBSUJfyWsCYSjODtLIRFA3OHaKGvFbfF
ylIURQyaatTLL2PPHFPD0H+KR1Lw5NH2F1DJGPDTT6SlxCaPVRBYwisMQWR5Rly2
g3Pl78K9TfgQz38kagqreeh2NAG7r26mCdMQRl/iTbRnAa5cxuzA2PyawluOil/h
yLaPDE7mVlohBC93+vDedoVu0BPOqxfoCjY7ok+l5k0thwI7VhzFPXTumSC8ZxIA
TN/ql5OmQPiDQD3+IyYLNAGYcCbTd42MwniofBq4yc1HPldx1ByTOV6zxLVdi6TC
iZAX1w2iqvQ4pEz1UNcLPoT/5UM3hKvY0lOvZmkKVQ5LfDDLtH+JbBPI84aKDc7P
28RFabwJ4B69rQmMvBMuvjatfwMNG5InFkJZQDEqHbCs021FXWnby56ZKZEBGOoQ
tgMLQKoycLMuflKOKMjAb4FdfAWdBCUW+zEaWFeRwOS0YPfYH1vHdWqgplZcPhnW
DkUs0Zbl8Tje7x8WoL5hAe3eBYBeRfB85soBnMqSR2ROAWK9nU7iB5QG/NH95DTm
YTYxAqTkbf5taiqjl9KTZBydNCH1ObV70rreoVJ3CCXDv4PO0C+8q/+n4ztVn2FI
WZoH4oSXjlXsTj/pyJO7vQfuJM/fapWGcMh0SSjXw15wYy9I4/69ZDfeBHrt5yUU
Nf7vZh1GGEMaFeTWhjRYHJnNtFfQBMJqqNUIfWsEeZYqV+LOJMyEQDZlO8p+iJEp
CQH8K3wzFgn4o1mFeTDRNu/7+lSmkbwVNkoj1mJU9tdNlqx5bFJEq/bwrF/a5GLl
3XfCxJWm2kwKfU3d+u3pJA6tZ0hm4tmgYeQFajQ+Y768HrN3ftTnq6TaH1nEXlAY
QrooPVfPLuwESRlVzYYHQltafWVgBU643b/LCkxcwdlltKlx+778b7TxpNsCFt+9
wIgbsGZqpC3kohmH7+HiDiT84dQ2+WIfYvD8celBhhN21umP7x5qUbPSzA9qfGd/
pRAAOwVY2zRHutcAJ97Cgzcb6scjqb4hFRlKriLWXPSS814n0Dd4nbZ3bWs+x0On
UF+7ToE1UqsNBx2XbyEH+gejNjn8ja0tpjrse0DwoGloNFVsU+zF1VfPEswdkKR0
D9zyqh+Xxh0iYc4AbRGlkiJuYZu+RQp18RpXpIYSR+hcj8w6avIlLKN7ak6+dma4
DAyJTnkWYY+DCLbLCjp+grJ7YOC2yhPlReE+aeG+vTkne5GF0Kve9Otz30ztA9Md
NZm/eezA6c2U2iRdpXc5liHe2H4Bo//0XdKocKf8RQx5LNV5U07a2+ieaJGLFDKz
YbOvbE6zPOytznFdvEhB9iLKqYzaDcxLvcWLds6xYWM4/v0jl2r5uulnKZIrWvil
WAOWUfjlCUrZzqT6Nrz3U1wzfHukGXy/vPM+CQpFUrU9RPtyvtbCExLeILizpMZQ
JEib0GuGkLVTB+M9TBbPtyueDF7R2QV/aGAi+YgKLXEbzkmIuYjkphD20TUjWsI1
GD5HENNkUc9DbM4o3pXpNafSOkb8YJf51uVFb4FP6IJu3si8GXkhLTV9G29Dm6O8
dzNaOamcyLDKNIEVM2NJS8xNOlihkTAQAiWX5gaeYmWPqcQVD/viU6fEO9g6igMd
xik1ksU9WLEYGLQ9i8gcFhdtLTf2Ip6FNyXjQGmu3GHDc986r26Pge6DMHP7jqYN
vrSIt0rPC6Fpdfbc39oj0IM8cV5CXm4IdLB169X2oW0+qRsBjFCY/WdE6s8EyAec
1/P+L3fTrOSHqn17Dy2M1Qm6YGXar+YKIri+Ndsghg1wN3155pWLbgvKYSAu9szC
33h0x5kf9BsxHy6TBs5PZNA5QP4nr47WpsojAIotPoIBmqkao8lAtald0Ia/5Fkp
rWU0dViBIvUoiCL0z0Ygwydt5yG9C9ypKfHr5CmoVLklRQR+9atTiSQ+TLoS6mlj
RQGGUM5rdMyxs20W7zonbDfgr2/dKNAPt1Qtaud0imo5fTlXevq7yU37XAM48eUa
c3aPRVlmSG8eCwjVFMNQLTtwfhDukY6fbPhvOY4DaXe6/vi3gI3vbGrWbHYIJJsu
Fj0kGbu0RQRRmXoVJ6mCVd34vC9ExBl3i9s7/CHD5H37Y+DbuHcUYUzyCXukWInv
u+XAjmnMjBK3SbAQryBkY4ePxlfF7FLlIP9N8nm5wf1foioI3qEygAVjU+7riATa
k6Br55uUEP9+qWxuK6hDQQ2nmfSKz8JAp753jUWfoVYMaY4/pbSM112gE4CorLnS
K7/XqicX90PUW/Z+1Dv16qowsTZPBXiLFXoJee8eC7jDLbNuYXRfqNx9XY7y73pL
rQw6sS9qO/OEj8keDezA196rHLO52HYVhrV57bOk2N1Ibl50BiXG9qbzQMO5DnCZ
xqym2P69t/CqWjNWqxd76Yl/fFKK5yPzXrw3HndY7qze60o1TyXzbUfMSAX5nvfi
E5zPdST+ebyOuYCSfujj/UCWrNywwmqTLofCBUpKOIMATCs0nr6UP1dpXj9fb0me
Yb5D0vl4RstWjzBZl7ojPoeF3yYdRrf8ih64NrKyXopqUSUnj4AH9dolgJSEnJ/y
kc5peR+Ug1/v1bM30nYPc37bBKIZCi+o8KPTHDw352xgXbUWOOx227Vv1/tmKOhE
pgyI9bYVcegHCNJKG7a2LqXpZAdjx/9KAwQhAF9UTLo9IoH4iDE/vZiruXchHonS
n128pq3fYl5F7O4hc4hGv9VG3Jfzy1XT0xQu5IqDmTOBvVYBYt2BwW1j08z11vcE
kSZelyQAr+epzxhVZnWew9jCwXryjVm+l1zZKyf/VAtFffdAk91K/Tugxkpa1h3k
RO3Yu6Tdib0FfBcSmG0OM0bAX4BIfP3VQ3N1ejs1b47aAJBeYEWC8pZBdb5XMPIj
rzdTw2PuhEAE1fGgMejHiyYqE28SJ1M7qXdSsIBJKibZO6AdH3jVCet/Kb/ehfjU
S3waYPXt28s9gAIS4rBzImDkzdJctwPcUnrwCchBiYylLel9VwcU8NHEBoA6ejJM
7Xiyrs2x6mH3Im2MTBsEuijrYZogwFTskUgPcPwcO5o6lA+tLLHZFgs1LvixKyuC
vDyJMzfoF0KFy9SLv7YGmF05AjzA8/TTsGTHEBskVSC/HhHrGeEbSiciCQi6g3hf
6yWe1VAzL60QC0++P+VEjfD91LuI0ZfOHkUwmZZj2kqFb3WUcrX38u9KkE9PbViO
dkQMWPzyzOERg5pM4AdARhWJ8+6GND9Aa3iVuoEIE+qrnxYWZlJ9Jt8IorcQYf0w
cxqqA+jN/mA1viCN1Wij3WHv/MZb9GqZE5UKl8XaP9jJgny/NLElZN1IY1Dwxwgf
Xx5eGIL3OwNdH1PPSDvWuTkbQQQ+kMCKMTu8x8yoTPzyZ4LIBhKRyC2R+NOGBjjd
FuAyWKrp9fLj2eMZC7pv0/llYx8lgMuUWfSVlyzBexm6P3YeKmuY54emns7IiLzz
ZHhPpo9c0M7dQrbW4K1u3gf/7G3qrGSWiLChpPUE/Sevpm/AKpjldK/lHPfZUPh9
Qee3bl3NXqdjd8MW50AJrRn/QE9yM0PI8ly8U42SMEGqYZfdgZzhWOxdB7gDQqth
DAj4VdsVslg8EBi0C1HbtNGi3ReziqP4VcRBnOzWDHG7HqKaFajOSMMKFy4537rM
xgbvYXeNhl0mvE5Fw2Yggb1xYjk3wL84M5DquB2OwAEuaTLH93uFq+LF5oSgJWKs
Ewdx54lISezqULdgGDitFHuJOomlo41UcBy9qAKv/H6e+4YhusG7PWTwUlSur3U8
YD3Cp98gNP7TBMHhXohxukGAmEUSgRpeWnKr3JASAxbTOboMg7fVfEQCGaiDTuND
Jxg1ofUscHi5KHl5YW4PkmSMne+wpdQ44gQxugdRozuFbXUXBrEArL/HZP/pxEP9
0Yg+UEtFoQg/5nrbJiKInvqaZlHp5g7p3wXVdb3//2vn2U3i1D8WgSMMDlmDPOVx
5CsNFf4BwxwgP8dDRYiVKNaRPEwwvmt5scrTAJysPsy+o2taf+5PIkymZHPnuqid
ayYATgsbZbdLJDMpie2rIIcBBzL5rV4/b2AK8rEfL+F3M5qfWC4xqLmYU9JZUrdH
pD9nFBQKp2pMFlwD8+NLqBCwlyctmATYTJXuLaDDPUt8ejh8dCGq3CzsYeSXApgi
mp3nWalfBqAeqjsb+b7/CoLmnYroz1uGO5n87OPMNA8M7KaQXomkIGi6ekGWda5f
sHPQ4zSx5LcZzPN0XNrM39G2MR8f8Oi6qE7VRm6PeLGyP4cybKq3j/mxFkhGpEXG
8qpKHz50yc6nqcImUNrhustoPDASCvdg6sCKb8eY6SyF0/3LVYB68Q33BN07CJiP
oxQAfcMdOh0ivviAhQVs4TCkp1DQ8KMLR4d+bzpa2izB8xTIe1N7LvLZ8G3dEFhF
fqeyb/ON1sYY1yhE0xvaUcBqc502UR91Cdex21vCqg+VG/l2qiR+9zXgaCib7Ptj
o7KdG2MHHMEknwNAwMWug38aRa62Rr05UY1Aowv3sqY1B1eOCSlbKnJYM0T/JHrj
xjk89voBYZNc0JDqvdrkVjeMB5F+P2Jlh2Noto+GsjgUMkMeAp4ibFe5RaJ8HxJJ
/JtIMU/TJhbJv2P5ToSjgCl1URE53Xvb5OK7bqWhlhppfdJJaHXInWS604rq31SQ
taYG+O+OefFlYB4sVQkYRZF6BcVsNLUFDiz3okHNKtrHoqCdz0c6sKTlg4Zmavuf
M0LiCGg6QzK8tQL44i4QkYsDCnDfG7MWbqI2tCucnRyOy1aVxB+ZOEJjweyG6QJ/
EwiaeMuMuxo/HPQuV4h2QfMFOUnph0rveNlWiJSmS/4YZw3USUslVgPRQx4Jyls5
BQpLC56sZz9DDxtStGLNkgOAMz5ukA6YjFaBPGr3jcwUgsbIP4ASUPTz0e0KEDNX
BKews5dagkcXXMIGDuaoZliy+AYg2p/V5JHA3e216po8EKHLXQBr5qHLALTT0lT2
erqi0HS1tB4+PNda+EfbUSNVUaZ/QnGUNpYJhDPf7Hvs71ovc7MzIRZIg0qhkBll
mDl1Y+XcadNkYsBSsNs4uWBhs+n3vLAPmaddvE5R2FNOCPuG/Tkj57svYcfZo0dD
VCxC08xgpSF0LAOXPIAsA+0KNOVyWVIVS1wfm98JLgiP8klKjc7ULHzfigV1HF3l
8ZS0DDm7bFnYEToBqXyyd8bLL0MPJc8KdMrjtY9z6jCJFrjT6zQNLMzXvVZKHedI
aUHpAaydcwvyy0PX7MpE56gbULt+btftgQmmDkBPrbVpntj86DIe+GH0Rzg6KDaw
npZgOBjurtCcPiksT9k/1n99aIH1p9fvTR8FgmhendkBogDZx6RZk7e2HsyLraNA
I5RF7KEH+95G0mcwYTYezwWq2ccChLYe4ZSKF/l/rq6l6fc5PdCl7LOp2+I1hXcn
a53O5DaGSEwrWy69wdO0WXC+4teD6I0ixLitiI5la5Mh1acduUrF/IEmNHN+zGWt
eUi6+g94nIJ2vsVKbHeHwjqGFUsu8t9+lAlEWfhTayMs+wvBs9fOogNd3RnUtouX
vF7mzR9qIdlHvK81z0gUOCxeu5Wc7SlGNzx0Fvpjc1G4gGtdY6mhjVpVTpH7nuJC
+pct7qGQeCbXFlxD4WGxLOjkx5T4vodMTQLY2MVAlKjSWR0WOrsAknsWQxqtuQTM
g/oHtzMADN2uc0RUUxWaoLu+uF3M6K+500zdVGU5+WB5PFWn4TgTldYDdueTPjy/
hda2zrnN0kmciFOa0FaWsT3S7Q2FEGWvlNNGI53vPwXzWBNCyjPzaq07e8aTQsHG
gGzW38bmJZTme7QquI3fnhDauz5b8XreLe2cBO5RCen9MZKK8EaZupuqQZSU2+Uu
x7Uqb/asW9SwViT3+HKQiD1+v5CPuvsK38u/WrYbP6eQXzwaiZasqp1nPMkYVkfs
f9gkfwS0st8WHXoJVt+COCt3CPi6miHALZaJRif0xewr1ZQVlNmyH+z1Uc8e28G/
VKkdsNCY8SmHzfNp8CJ+xCeLn7N1HwZQUIetPvwsarhDllHcKdt+kaHZiqtMit1Z
D/Rjglg9jwIT9D7YYMaaHKQ0IIv2vjXvVhd6ZO+p0qN7sBGl/UUbmLa1ffcuIN7W
od1wqm5jAa2H9K5iMhmuDOIkO2fss6kTex2h9jaubnxQJvuoOLYWmpPp/AKhAcZ3
ab0/myL5zKv2I+gQmXGZ/EUExpoMhhZsHEvhEuGAhkkUyQkTSPG8Q4S5CAzm9Dd/
/TCpQW8iz3ZOEjZhhiN291787cXa2sHQuuCfEVxMgWW95qMANCATwpxPeMDLoqkd
Iov8F5l0W3+IfsfXpwU5Kg+u0CP0zYHDRgZCCECBvOfnWh3XgoFebHGDn8BHQpLl
qSZIHa4VPEu0Rx7PS69l7UbmnTPD1ORlKOiZq0wpWm1ybTznDIHK4LoMWysyrHiJ
3qIYvj3vpw9BG6veE71X+Y30Cd4VPawneKDD2+UGiAUPCPlA8WW+8M8L/OqCoXAs
T5JOKB6RsSSc+3im2Aq+nklFmVAsSdnkHSoyl15pkiOy59nJYVXAdpNs8l/ATvlS
txCRVUlyCD0pAMUriUHP0PVUgWhpH40XYoDz3aQD3g/8B8L3QvP1qu1kb7mC9Dza
BXiBTwcImCjrGZxWrSqH7mbF2c8FigIOPMzFD+/kZCRIf8cAqEsf0Mzm0Vv0vz6r
0FLag6dhvzbutey31pjVkFINjaQCr1QMvqXLIlTuLW21NLLMLUaaawlFQ6+8Sjdd
4iiHaS35qGLOUo+wgqFCanAGhALtcjnV5wOOiYQTVJaU21kWl5sf1mYcAEvu+3sJ
6CIgLFBzpFc8smw2PW3CwYEPSJc4ph8qqyCAMzWMgOpX4w5hMiefqH57EmsbQYZo
enOiXi0FnTcncMO/js5J1JQBhLC4j+v13BSfKhQolv4jb3HryPnuyDiop0LyNhym
tpD72WgKcPQOsjQgcVPhS62eAJrrmPiCtY4FIMQu6QGQi+g9ZekAZ9KJSdQHndaN
Na3FdDblfoMWPClmjFbD2g7nGmmx2+UXQUpRuKznhzJp/OxwNKkcqqE0Hw0jY4FQ
B4gwmt92n4Pw6kDEGUPYFwkMz39SlVjUM34xmfmcBJIJ+jMkBm8YVE9S6IEKeMEc
h7cOsmOUTaEQzCh9481dBncJoypTgqj5w25ZfY0WPA7H9auSHJjysHyD+VPiPLbD
lFVRB2IG6sQVDsGQCV5S/44jVKk6hjHg1VJLo4JrfQYKann/8eyDCWmrc0eqSDGb
XvxqIE1wn1QwiBJBnYmR/VCVXSounG0lqGzB4uYNUwqfwDU6ADK/PclkiZ2VQWoc
zYrf53Wh8fsZeTsSGcZLIFzUabZ91jLaVDOIYRcYubxXYCLTpaExyfb8Kmxk9vm+
gCzEvmnbUX1vBYF/rvPb4ucIe/HyidqQM1hIh8nWQn+/nkqkRdbVl86FraLLhgdD
hb3iN2e7TrAVlN72CO3NYUFX+phlOB7BAckc9zoRE6UwZXvkdJhluRksUYoC0lXq
AhJ3emeZsCSm+v/2uqEyNUsYVjuyPOvz7HwGOUSpVKXUGG/U+oss411qSL4+d+dx
oNc2GfodGIim0Lt43g66/kxilY7nU4eKVWqWruxlubEYMqAoyHeiDKnyk/tHns/c
LtRyyrnoodvcriXuLAUP3yL2PCdkCo3OH0n9v6e2WQm/1I6fjkRoQQjWgG7QwzWs
ofL5J5MT7BG0A9i1jIHPyTsWx4n5tM6tScj+qDu1aaIed8EAJLjYr1/g2evYK5IM
sYY7jfbyhDUMeZZkjwDplBTVkbTR4AH6v/mw4Ex95oZrWaQHfm3Ko8qVOEwUvMh6
vSt5/SEjwlHvibZFyCnIa4PKMclxireU4hetDWXaH1mgecLunUkaPMcXMkYQwkae
ws9qGcrmEule72G8RJFcj3zr+14ObmhDFnzt5QgB5mMUCKHvu9j+BM9Cw8vn5ggG
ED5Lz1mOYjeAL9zyvvXVwzhi/aMkhd7LpRnRO3wZAx9wnwI8OH1gKn/BOivHa31O
wWxwA4/vb5zz4KdlRHyiRtqItoQYjTsZnQehSfmzmHdU5+9L79mWD4sEhnZDt12u
75sxoM2zU4cYmdWQe80bRugEUsEb/09YTxeNPiovZRPP8FUj6uwBePeDL2ikg3AV
bGVP3ra+zTAdM8dJIGzA7CU2q1SP9gucunPbnFNYTjWew0wP69E4g0xdL6gRSWR6
JyvUXJYIm4bG2vmvo2whmE/GE/iPq9UTB0+wZHY26Mg0nVwqEpkN89b2K4Tl+c63
bFkY1hl+AFCa+TcCaFA6bTbDKdvkSOXP7jJMaNatHvB3KgVBS8dhpCBFdD56jVjI
dF3CZ4CZF0PNYiHNVi9BvkwyeQuOklpK171vcG/IGsWau6HlHCgF9LzLz26Z7dwQ
98yIyZFO3K6ynkM8mfCx8A2qGKn2PTIKdMsiyjehf4nGH7sjPLuJ+0axmYxYGBi5
ug4XAWrcRQd7NFQKkFEKGKVGX98eNZ0dgvtsZ5GsFpCXQl6+YXa5GJxdX23DWryF
zrXOXNtU9n9sRQJbPwmqnU9/QjF3tSLvov78iB1dVeJbr9Hn6q6Lu07O57z8sW3V
iMVY/0rBVkaucqM8lBJQEAoNl//h/Z5PVReZQ1Pw1TQ9P9Y1swK2S9U5Pq7yOLg6
+p+BxVyEHgWg1B86nwnaTxLxkIKu/G2sNE2uL7frLQBg1k/BPU/YU0gTLHV2Oe30
99cHqDG7c6exduHwnxdb8aG/FsWV3JHO/tbYtjef339Ulu+4kq+VjyST36FdxZSM
SSthyd/k+AW/he64hTY2Ni26NLQFQlcn8qsCCFDqE37Mw2W1IvYljqxO49THuqbx
bEkUG7Snm3L2olwUrwWfUn+Bs+ac2sbWtyLvHP3On4hk2C9bQ5rqfIoOz1whVQ2r
ijGq8U2J93oGXfu8Q/nv0N7yh4EKwkKpZE5j1Kl+d0mNorjPDiDIuCW++GpBZUON
+JX/UB70Ftg/UNTFooR/4B+YQCrfrvIuGjmJmpyU3ZsvqVulpVKf9i3wObap2ijt
oQYVkSS8OzYR9mYDZjx0CgpCPu5trhi9gFNZiDqHhPff1SuOW+39PH5GJGTzr80E
Nw7eZiJcMrQNXSVjDo5G7AgIS6hP8FAPznmofcR2fQClJDjQ1btkrbroAdsp1xKQ
Ou7Qd6TYpoPmUu4o5tQbYog5Bq9xb0acZMWy2b9tT6rpbenrCT6/fkyeMBBBewFu
3i/xjxUpbIlZLkFqvBBt7AIXZFbSNwQXXsGg6sUc9Uk/OBxQv1HmkbRIgVS5C+1o
w7Mjzpc3ieKjFLdM3XNbnHqL8NcOi5N4woWLlo8Q1RCo+voxFU/+vgguO1Is7yeW
+y0t81IuO5Zxr4SmG8zw+G8ybhP2f+lun1I2w8SPJBr43cqpnKN0wXu5agjao9k2
OSKltG2McjrBapgO8XqH0wf+U2OZ7hHAsy6o0Tua6WND8gLfGq9+ri7RQ/j+wT7b
jRLD/b9uFTpa1mqvOmm++I/tdnNRsVgv/xNm1hrWXcUAWP+6hCwQ8+RHheAszi1V
uoKj6ZFS5oEJPmdespC1Cimk6afTuzT7D1Wg3tkbFcHKU8oW6siMfHcILTpuCJjB
VSbh4ITtyOFkqj5QkuXFka9Y5a4qiAs9HK11zIOKnUTIvouTa275fHV9HQuYc9zX
BL9wLWaDq7++YvnHsK4P1ZgqMaoW9lEYM5JgPeMR54jaWo5VlM6Sytgjd2fOq5Ma
/ZA5cEYgZ3XdGThPr92xROcqOaS54hizti9An+KGjFMLZZ0qyjxqXTIXzloOkMq5
E39m1tCZ1aBQE6/KODtMGwWJGb8QczDGq8rInwyfRqLL9qw2am1XilHY+N0Nfw6C
uoHiVt8nOVWGYaONZT3ca5Xzj4ZiMT/C5fDyey5es/qtyJNl9rY37Xr0bh4+G+7K
/b9eH6gLDxEiDkWm3C9rMx7JFrlO3tluXWJF/iVYGlbKrUHaNeZX/Ck1IU+iQ5C0
jgi3RYlfjNmVNYkck4E96/rekGCU8iqV6TszcSEz2NQkotvPPk6XRjH9nKfdCNS6
xrpZqtkXfFH14eKfWQ+jTzHLtutAW4Jh9zCZxrgyhdJJvpYIAXgAwTW76w8Y3vpU
Z2p+BVyliXhrutDGceFeUQlKT4u0zzaRNjY+jb6V4Ev9PrtwAD6V7q3hSJje1oLa
UfQpFjwA2524brHH94d7SO3Z6y4ZqLHmFJ77XyBHirXXjul24Tcu/QOW1gcrtLWz
puvcLhDk+WbtLf3Pccx5xN3XV72GtrVM2BiwNgMpaTc7/DqRo5Ck8+9CxAQIHYd1
HqC84yn6lvEyIYwT0V3APOUKShkH3zXWGbin17zV4B5XyWnaZIZsfIRYnKtB0nh8
QqhQ0OF5nJE2N639yfOYiXjMACPBseCuZq3W7bL0W//IX63O9n5IKn6sWBIFz75q
vPUV0jElM+1Fvr5/lrXAnfX9FmmK+7+IH614KJhlaOhGPl56kNrjM3LH0AoJ1Pai
VQ7zLFz4PAxN/9gQ4g3UGPERapLv6rA1aIl8QsrRK0n+LCjqzxPBsEtjEXqv5wDp
+MQGbwdPFbNlst5arr//uuJGKYyMQ80NK5aE4q7Ys07PPnF3VyPgI4pXpVO5S5hv
yG2fprnGVzGIwkf0AgVkUp9KXJiYZ7GN7r7gKaTwxKSHdwCLamn4Uy4Lb9XMO0h+
v5f7/myipSrskQbFyy6s9L+Y14iv8wrmPPW/H7cUJ8mXmd2swITSmI0dGHPQECuM
LLu9N/89JM7kUaT+xfugrMN8dT2fiydh/yBj/LQcfO7aeTZNHyNNadHwFd18B4zL
ZLwtfkEgpsgD/furSPGG/Gcy2SprVNUTBkqODe1U752Zaf/kdabt1T7GyhDZXbyc
orMnkixmcUb581+JLjS/6hLVNOTkuVqduvjDe9ecNOUqkcmb4keq+JdkRVyWDd2o
jhewUZ8eWNSy+0pRAHGvXEMGR/WC9hP5uYt1EZvog7A50iedo0c4RwGJM3Tp8TNb
VqMErRKIBWu0yV3nHuSUe5OmaRgMRhduqULUfmam80ETiMx4IYAAghVuoqaG7c3q
zF3ul8g4urfEPt+qxQndNGcqUx296SLcxuQJNMbtzPyrhMcb7A/o2QkwIicZwyl+
4hKjGGEcYkCLcRe3ta6AtAhC+70t8MpaK/QipEkIxAUO+a0yNb8O+nwwVHqlBzXU
KHhrw0Iy7EGgTYXDB9bmANPlFZK9iBCvBOtTvOifi6vGM9IJ4DeF0kGwnPcY1y67
dcgBvvJ4852sj189gaCcZIwUe4fIK63K23HSvYDuQK11avF+k0bpvRahtRjxTN07
zceyQxvkNEHTK1opkEzGjqgU/J/8DNZ9PkU1JCg2tJsiL1NZCglk2n4mIbGY8pKQ
hAkp8iAtpJ0P/cdkGGzr82injWjn0QLg3JXP7Jy2BTFf+9des0kUq9zn6hnA1f02
7AduEeMSrjQMVUxZNAXZQV28RsoJHcJrV2XAl67jfToFgN5npTToO5r7gHNFtWQP
QGs/HHa7lcBn7ca7b7AvKbAKjhuVccjYh8ONMS0EevVdjOWV/uZt9ZDUdMtRrFtM
c035AtMN3lCugmcaIBYyZQZrJPIfwLzSgTf4GOjvZhPCrwv0KBV6oUsvwRES5zUf
OvrvNCURocCOTqHVopr3jtwCaJMxop0KjR5t8vb+RcpqyGjxyP03ahquDvCBivaB
nQBHT0VVC0A4esZ0by0R2zKw1o0ziM8ZwkRNYyYZQt+F7aaT7KIR3fh5isg/5QFB
rupYJf+G7RmE/mex+IiIl5lLOzzDAIGAgBGwtQ7KUbWN71v3WkmG4Rx41ftHaRm/
O6VvJ//RFeJdujSUVlnRe5Yd0PIrhWdPLwf7ljJVNNT7Q695EamREerIBo29N0OL
q7Ok4CQaItnE8Mx36DgYWnqL3YjANJPYdq5L+CJw4UNTYUv9BuqQ1/ean+ft2BOf
LvUaL3NjXaGvf0BdoVZQzPjYRqaOLpDJkW2KoJBWEoTPmFo5U8f6uPMIvrjiRuDR
cANVkcGml0iDVWAoYrfru13lTBT4HBQwVsis/RX7M0IiDhENJyFcTBHbSBjD9t9r
XZCm+TGksWbqREoVaYmr4IgbL/QpMB6TiKPF98KtvCsM6oQMBroIZYm6BQ4WWI+J
memmrypMETQVYbCvHIpLmqmEAQtq9ZC/Su/N5CDc8JS1leWpZtdo4Par2Oo2TQRg
nd1F9Km0jcSUB9/hWKhoa6jxUcLhf60meROvNoG4Opf7EzTrdoZ7aTaQl5sPpt9f
ZHC8PT5w4zj2b4PKUQ/Qec5LjJn7dgLKkfrA2Kzq3E9tY9K81p70xAcKEMj57UzG
uO/VWm1trOD7qU1Gw+Yw0UCoadPta2AJa8Ped05u5+GqRSaM1ItbAgngzCja+wW9
vfaYi//va88hEbRgGRbLRvzga0MINVK9+Tgqw6eWSzHgqo2CMDoNdSB838S1gbkO
OT7dFEkOzvow/77heoPj/4exj6JntLIqhVMvbcE5hhKhQkOridzifUu973nMyxAB
8UI5U8iMjuYKlrxkzAUYlruu4kVrm2ZM7XXyzuAOdHzncxIrQQqUsIIBIqaVUJ8y
2AMsgKaK1VH16YTrSBbiZece+vV8s8aT7YsMsBEsmNU+jELScCfFKisSY/l0A3vh
Rvu15CnC7uLgh3aVZlUkbub9fhEpTVodbm58QlSJ08gtUcw0WGFH0ViOvo2yuH32
dZE72ffnY8sfmq72MDIM66N7rdm3A1plIWpg89/ebLkNZuYElDZ8MWrQkZUmW3ts
OQoihXDo3rbwy5IG8U4NqnobcEZNF6fYaqL8rteyWG6y5ETq8CtjRBgIpc7BD8pG
Dwxkck4PaRfIloYcfHqTRdt+v2asDBmD49A+v7V9TEDpN0HBpQss7TDLnvb6l6F6
DZtLp07qWJ0R2+YQVMqGOUK8zaoCUeZlS9ZJCWyZQYiqQK8aimR5Gl7lCNJ1SqmY
+Qcxg0hVCXYO/OEB5iOOTL8HrBF9D+8EloQcgOtfniTvZH+KxW8YX6CM8IlvT4Ww
bFNkM27lCfcdIH2JjomaJvZqXK9Us/4cnn842TwUWVrsSraXHiAlJXJ8tcvphTpv
fruhaj+tjkOFGdeRzvsf8dwkj07YJpGtwMqIaMymtLsNBb521aa224ib7RLiyfei
E5eiKimVZA/1bmTW/B8WoqQwUDNRjMK8o6T++jZq2kDnu1sFgeqdslOjxsvk7cTJ
AtpCDN96g5MRyh/UVrvoEP0b5z6pMyliLYWwKINCs41ssHasNfjrRq8DTaid1TFr
HJNtPLMML7prhY2jfwPD7IFsoxmYri4t+Gq0qpwrXRSGLDZhrOFhdTWTYx0eNHtl
43W8UbXofwejHM9Wsid3XAVxm4NkJPfuBWCqitEIZYzmZwCer9hGWSSL3+xBUP1s
n1pGYfXlGQ480GOrTNXT6KjtBzZCwAqAdYDPkSS730tC3knqUV8WYEXK0M082fKI
EsDfJwCBG1dE2C4HZqMwYrE324Uk3YSyDHz9XG9Ukg0KITxyGTMwtdbkylGbDb+P
kc0kFpcJyh1KIn5ZR6JnBQzWL1qu59xHHY4b8oYmUE4mxD4n0KZNMJ1qlgBzn2MM
HytLMyLxy+DDjBXv7WaVo5iQQoyeDp+nLLbKI+EorLzkoDo9so5iUK12KE5hwewd
rbOCFpNn0/7dZQ09Qj6xoNCjGs+MRj8rMGe5fkyRxl9+nl4g8pKQR+5T48QpiQuo
VZ05VrcXQAws2StCSiMwWm+w2I1xFkOFyUY9WnGPg+ykafAu5rGryrrrNJJ84QDb
QCNXLUza8Jts2kiFUlP84JSKNJn7STTYi1tboKWInCFLkUg5k8gl+5fBW9NFTgC7
XVdT791NveOXn+eMlnaqIR0h2t1durhRteGcSXA4K5FFFnvTFpyjmYOYwTAyL6gZ
j6+WX0qZKWSdyZcEux5mGQ/BZplk7ef5QtLXboHW9CIJaYAz9KC1T9CId61HqR68
ctKr93CzOSgGALJmmIb2+3R2+hm7y1903Bpzr0yAYCslSeZ4DeWzGyOiBelQT0ww
EPve76ws+EGVH8iK+1IXr3fPvYspg9mqazZHMcUOfV7bT0+auHSPBbvEUF+GpC3t
JZZ1uYfHxBL06/kJf3OYhY3ScOEDZH5uoOV5yIbe0vZV7Xh+d9O/cEEt6muxoulV
VYgPOUyLq28SmohCLm2pkA6faF3tRdxw2X1ZVp1QwoqeA/5Llg2NtTmI1F6tdPq3
8ZQ5FOUWVIe6PLAKN1pl6PZMDIWFYftQITuA9RGg1kGDLEA4KaWmHLEv+wzCYZ8K
rHfh9j24BbapvEfeO9SaB6nxVIpDXk/iGozZuS875TMIJC68yXbjckSp0cuZW1sJ
1EJeDsLXja3KzRNzp0ctapwox8fx0uQQomDwUptOdtlaauQ+n67i0XC/PFHDsOu3
XJlNVfte86+ohmP8IODUG+VyCbqFw5I0+BLTlKsvCD4C5JSJdzWUyi84KhJWhAoo
OQouF4wt42Qbq5nReM+O00XicckPymKRK9gKjktNlEIF7sA2NHmdgPvl4aFTComD
88VYRy5TscsmnFR23FbuAWvEHKQhwybb1nqgGLJQcUfUy+9f7XdFWyPW1tBz8MRh
uOz63MLDrLxHJWPK1MHG28A+dhQJQIvULDOuq0lHa850JfKpyGe+xuQH1/7CNk1B
/GxkuaZGEyaSY2z8hSJpBWZKiFTZHQvmRO4Vayi6y1K2BWyg7T/3k7WXmo8oOnKD
0oVCr7cjxtAhy2oNwWa4TpeL5EKLfK44VpA/IobLp2Mxag5e8H7Dmi5z5tFd5Esk
RqprDmQ5L62YtAFsA8vOPw+cJTQKfdCU7FdFcuQUqUi1EgN2+8/Uefe+/uyjizC1
RBGrVbN9Vk124v/2pok5jrsmXTuFKAUgWBcHKhj/F/J8XZ4lJfTrvoaMJmI920uK
kZhu8tI1IcZ2b/o4Q/tbf0ocQV8dMuX0KkHm4qsHvQ6Ggk0gXAl5f8KC3fos/oWb
ue0HjIWsSDi9Wwl4D6UvpRiv97VpUPSWtrFc5RlBhYBCL5Lk/63OHV+PkQduIEmn
2NQXVa6g4S7rVotWSIXBvefi5xSLpTHWCbleJr0I0HRABIUjAPdyiU7ttRaEreAv
js46ThpYs1s/qZa/m4odMnhakRaJ6CP5PFe3Nc+B+JDdpqweq1BdbCE20V2pJ1qz
ae5YCuYQ22OyV6JCGcm44xKFFfpFAdoFtG2WgQ4GPCjrtaYVf/AkxQbRcwbh6ICP
B7SFNDa6F5Cn/MKaxXRLSua6av+kX3iO5/xIyaLYQ9I76ojeq1WYFxFZMaozp9sD
FKGq26itE4sFPr6FcF3hsfLTBkrs4ZIh7Gvn1kIdm8Vf+6QUNXNjM23IPmpiWiSg
U8tcqXGuEIZF/nQWoQyP8I0UDE+lfSa6VaqBg9A6lvL1I/noyT5KFUCF6adRovDH
zlEoy5qKg5Qs9TLjsvYD2ReBAm5PHQmqZYlHqjAXjsxc2kxf67Yz9TfXdtiGCYNw
Ofs/ILlht5hYNkW4FkGl1Nj9e50322mjNWVkBYfRrVpzzRL3KA0AhBzl5S8IOrlb
N3VSO/kAInHjOcpwR9R5L2y62soriAhUN8gPA9i4cYjrFwHqHcVAp4snOfey9vs0
efG8AzNCme1XFQT3KWw4O9eeoydrQ/8M7JyW+96r7KfZj1psYaCKayhY25Nhio6o
59ZXMSdDFGzEnNNOsEGrYW0HbWbLQ/105UFZCRmMYs+rH48zDeu1vvIOfqIhNBvL
qHQMeTTLy8FQkrcCJh7p7oh6HNz9poNgSmd9zW7NUr+h+rXCPsvankb0Ade/XCmz
lUg3ZAUb9Nh+04LMaAAK4+VzIYUJP55dgbGYPVR9eUbc6wBxHQzWslsLwvMiMmDd
4xMZAJ15UAVe41O8JhE4JaN8Okc7/V+QHUIWW3/iSVF5/SUzUO++CoI7+4dF437s
iaigepr76R1FXvw9e8/FsXC9ro6BFDW48LrcDnavb27i+ashbHQm1mmupUT7BOGh
XvIOU3qR82FbBV1DWPZ1gVck28B7cdH/xDssPG6wOzwU1TY8r6+a4Xxm5QTEUwZj
6b3TtVltM7yK7bhMKbKqQS3EixRWzUXtM6FThu+0Hf9CTztmwgwh3L497geXpkQv
YkfqGFWZbQ08hrzhu410t6TZ5SO5t0d389b5wXmE0IsvBicQ2elfVUt0d6yYWz8i
zsnC6Sdo4dHGZVZPTyOY3U/zJ8H9SENSGn2rL5ZUV855b8ApjLd+cCOm3BwANjw0
Rx3EkmwNw1ySeR1QRRty2RqVwVMooyr/Kt/jXCrk3imAIbZeyjZpP7bNKmKZaUEn
y4eNOemaK5KCbvyDtAfiBzwRaQxtq2Wfzdwy/xv5TSJ04gczHyErRk5dNbM3yn5X
6gsMRJySAoHsfi56HvfOb+VaLQauyCAQVSh+cAd5LcQs/bq/yHBZFHenippBP5Kv
PnILL3dCY7sSznEIQzztyXFSsEJyVgiRSHc5Pdf2al3cX5/UMis3EmlAeCA8X89H
4aOD8LpBGF/qjuSb7E70BPtt0c51w1VdczL0iTXbIbzqbHnGqvAsVg9iVNbKC03v
/IcEZyITn26ugWJnbnCQOs1MUbjVpOl0CCSrMMSctCjo08PfKbjtP6nSoME8ggHV
YM8xrv46vOlYRSxyh6/NJDZhEbtfRyn2hLRbaPzgL9flQ2R1chtdFCfhKaz3yrTR
0L4kLc0sYRWkO/2HiACF4yZhdkoqSrX5lhe/7i2B1+MOjrJ8PrWtugNA5LUcdbS/
ryN0tll3JdBPB87MVSBjfeQmmRoRxk85eRloq2chWQJ65MqN23JWit5PkTNYFfro
C8ql7rCoXbc4t0LYRSK+ZQyTg9/iV3KHAVzxoiuu4lIh8TW2AKOj5256SKeoLZ4e
SB7/PC7Nd2Bd+xLQQAAPW09NQt+DLleDqj8lhrbZ99zY6i8+bwCCkTTgYuDOTi7B
UwX2T09ikt+csn1t/GrPua6W4Mgku43NUEgNJxxvCrOdq3NHig/4dlai+f9CUhJ4
rD91NCOew/2gksN6Nibo0vsMZ8rBiivhfoiYFWvubol5HzUHNM0LxcUKagK3TBmj
ngfjv/KFPurGfv5hJZ+WeTmu0it3odJQIN7OvSWvGQZMDSzrODFEWJ3rjWxI1qFM
yA9Y6N70O0BkzNhdaUeShiIjrZm237QFhBE79ryX2NJZKEsVJ3PiYRdUwJJ3zULX
pbw6noS+HipRmp2L1pGwuotxMXFDVQN/kWcb+MZoeUQzcwwuG8/POE5KyGKOsu9n
cZZEPMGUXEy/uEIt4mVU/pVHGbTVNwwg9pMZzV2v3mc5lH8plFzH8KJVCDAu4w5u
VSRkX+NxRKiouEH9SN8G25VYBQqidYD7LteXScP9Uc47/Bwz77gfzpmkSbDpm0+I
Eyt54qlyDxGwjVt61eGAQQE7DmkOT+5hRXWOTCOgJFdSZKU32Wx6OylsRDw6v1Mq
2mOi0Jfv4P+0LOyABQgUqZcCOy914u3lZA5HbJKUtK3ECVJJGo9pPfMX0SVPeyNd
I7u69xfu/2+I548ix5ZWQvBYOqVM4/bb3KRZlL/Q+egVD4GOmhI4w78sfAs0OpMa
kEUa6AwnT8BaPE2dI59yfysurs0Pu1aH1M3MxnlWjHlZfjF4g30RvUEvEGWL1qwJ
s3i1Zyjqa8R59Ot+rwDp6RzifJmmhVlPQS4Lh0h45mp6QlZoM+jOVNJomgdOqhaq
p7/P153/l2yYq9lbrnQTX1+wzboX+zLMt3IhvsNO3EIQFI68Zuu0rCLivITjsrYh
Ku1MS7hmFTQFsyZMRWXf3YrpKt63ZNmBgj05hhLyasNvhf1gE8Sm6q0H/ckwbNR9
sSRryN7hyzR1MmfNaBiDbuEcN90J56lLVCH9vgW81axzY3Z1GKHE01M4ZwdWsuhI
jyo4MaFw8ARtJNMjnY6Yt9tLyfk7cFu/wUmNGXwZKetI8LyvJs9yA9bGsbzCnm7p
Mm0haV/ZYbY4Ktpm8keHRnrW+zkEXsbDl7NRTSFtSHLYxNyQzayuMiDtrEZ9V/A2
QspeZrY+oXCpYS1xkugFEk00AfSVF1awpki1S5yPcdzfNToVJfXyTO+mk/qwreQE
Vg5dO9e/0bKB5t7E1/Ot+anv+qRUW9e6T0gfmokOoA+stLiCLFmBwqTMmvt+DPH+
QuGve172LGh9LsCE+c+7QT/0jcc0xYVXamJtAgff4DyB1bPO+7J+lYdfmzdQvwAt
Tndsf58QIrTypyvc5RHNgIwJ0PDwEvKLDJuOSjVQNio0w50+QaJGVvuh40sjYLwM
H+ysUAZIvis0x4ClciEKO3ffbQzgPHkqksgGN9uRJvwDxBi1L+6GKhZb2yg16xAb
5vC6e1a5C2YiCS0nRcHcyjcsl0WezU0qXYk8olL8C6mWZ+bnPhCI/OHGv35FCfya
bl8YKCJxOikLkJWf619XYRxJMb3xDTfwiJd6p3GfR3vRg2vQBk5YdRN/RDDicjwn
w0vymzyFzxj0ogdCG4vnKIIqSq+WT8TM+nmv8pLbZum4q2OcJQ/TklcCiWw5dNMp
QhIgmB7RlmwQruGAhTBGUjf70hQUZRGd4qJO7i4aFgPLeBFEUnoMKbPEMck+y7EM
rWHFlJKwzra8bbEUwisiun4Q1nesBw5b6ee9gnzx12v1n5rr9t0kDfyhcECzaCn4
aPhpdlYpJGS2u2Knq0fup5sL091kI2eJK/+w905amgCy3Od4MnHRb2k0oBUtSu5Z
/UOyd4bxynWxfEU39YmS2/dEPOPtkSbfvBy7iJco14Ugcq4UDITSBDFyBmdlxjjq
+QtlKEZGJbcme84bypG04khC2HaoY0g8SRxiVMtMaiXImq2siflOaGGp7NTrA6/2
rGGgq2TI3CCIjUVC1gFJavO/KGEkTXOsISJwo30qXBmPNaCcav+MONHka8maBPBr
EKp0euIFwGNwyI9nkavj2UO/HWGEmf6X8rwHnA4+Fs6BJ0YU0vaJFX/sLSvLy7Bg
7jO6ztswBl5GKnFV/SSInGVDy0TQBtwXm2Pq6uAWd50V3cDdkEcD2SNnNr0PzUzg
JZdIm33KMAs7my4JjV8IjRGXxfkpvcCqgjDBUH7wy549pwKxcjBYa4zgKdP+QaFT
Xeh0e9iSixj0pKI3VfA6UaCcvXhQ3sRmGl8tbybq5vfuGLyAx68nTJlqTuOrWWdA
V6LIlxdxogcFUgLUM998fAmpkCDTe2Tv4ju/tEEk1kqT4Ptd+kJdaR5RXwTSxluH
+IKFem6Tf+bksSm4PfR0tWyRqGneNwgYb4dFQ8m5422uPIWGKnh5kSALXrRP76+j
3spfJah4/e5gro10JbgDybWMhhrTdYm8e+Wx43Ld/mfsfI2jg/LjkmePbNoBl09j
hpDp8bnCI52IfCv0ZEH1OYx6iZVggwwmbr6pQcdzmOmWBSfz2PGHNx2pb3MdZgm8
ZBVS4fnLI8MztsgvPy5jC8BtMdmokLMluSqS+ZuZH4snmlx6GBcRUTDXxyH2tKhI
CW1jZv3/nw6mEdiDM8NLE+WI8rn3OGb2wYePIc8PCKxxvo34e3bIiG7tgZLrYNgs
zsx+qtjcaZtEKvl05a3P18XCLN1Tmp5E/1ZtLEte1lIeAwYkvPPPW3OZWDXJAzSW
3q5wQmz86hT/RwwAo9VClaTWlxalVIGzgWBecvnid3n6Lo7OGwKPNMknF/y7aifR
d8uI+VatTexwdHwvrTDsFPerkGZWzl9Y77xoOp+5af4dKkw3JhRB63UNZ8ljLzlo
o88TsYqppuaVu3itU+zDlmYjDfkOWr25to7l/J/KYv+maoyfrKaSzPEVT+izo9NH
YNUSU8iKuUroDVKQxtawn7Q36JxCjvcIyAed9JfqhD8tcKIL37/oDLbrNErjjntj
FhHcDP1yd69O5fTznvlEbzn1VmBTkMpEn2a895mek7p16U103CqJHzgCgEX69Fym
iTcAoyTjiK3rEg07f/HGqQZYW/hxH0iThCNv2kayGGakIOkmyo8IZTUf7r1bDPPF
t8tIugPIFuTKkgwWfZYl7M6zDmi5VQYBDUOa6poJDOwlkpIPASXlIXwnQpdEJrpz
V+OLoyLWo4/VaobiSnPWUZlNH5eD+raVhPYCIcloKfn82345qpVEyUJOV9YcrK7W
R9jzySSoHm31bL3zFOO5fIj0S08lHx1OmU8Q8QmiIS0OkACzjfOjFrQ0dr1s+rkN
EW75KwqiKbGG30jV4OXVSogUSKDAvQMjixvArCwkGpT2P7EHSSjgjL8OMlaP1sky
yiWtkzxozCeSW6Sa+7UUiyiTbqVJwxTAUzkP8lUd7U5Lsd+qPE8i8/ITzmp9w8J7
OchJVJTSsZyWeDEY694CZz7puxKMbWxta6yQt32v9C0RHvwo4PeWci8qjrQnC0eB
dliDJaXwZjz5wx5UR8TNngxv+oLWSdh8n4w1FfLfuGZ8ysFt3GFT9/I0iIOHo4fY
8qdWUXiTedFLVu+ePdpW1Y105r++UDdNvBx628PG9UdsHrKtVSylWU3zDyyBQI+a
D7Vu4toCNayQFhGe9Wo6jGGS/gmSmZfnN2XvucKaz0SNBK+mVBeoQFCJIVqjSwMF
uvcipl6HdLMLyqVY1p1/aqJvbmo3tXT4kfFHY1bq4+EUdmQXK5IWFwZzpnIqADG6
FgVk9SpR5JjBLx14gjrzO1YrvoVVXJHehw4/CdeXhL4emqbKGMibaj/RFcCe+P0H
yCBSsMC+MQbkffsYLRqDmq8GV/Sy0znlm8WzPsANlWuateXAMBME6CmZOq9Rnmor
fNOvtn3BgF55/5IEB5jW4TUTdAsBPWNRokgZ8sRcFWkBSnJ5E7Bcjx64+Cn39Wz4
Et7R0743LaCueyvDtf0bNzke70kxwZDRgCXUbeI+QwylSkKcgAmbZdf6lBLaktoy
lLgbI6V1y47sT1WqYmWyHhmn4VjypHFoVGg6ypR4jYRVpSGuT4EDWTpt7q8u9IFa
dG8USd6x2sTmtyylPyriu0dP7rATgngOsdIZXFyXIMiOzajcaledT93vCLQhscwh
xqCp6nu5wlNpxLr8ezpKrKjmGbAAc6FBSqy8Ld0ycyEalJp3dg9QHUGt97eoUTeB
Nbh6oiE9RQBd43G82feCRJpSDkypNlnahMwmIrjib+KZFKUmkIl3Pr5O45Dh23BD
1hLXuoq9lBEE7J2jpI4MlURXCP7hNOsFjP1Y0qdjVPxHnoKP8IuXBHVAr1l6BQ++
ZqHAD4EvPI0J4I8rK49H7B/glCs8PylfsZQ64ZxJieHe2EUdM3jZ5y4x2oXt4+TH
YUlty84tlicYzlE05bnQft7tQ70K9rzmu9jX5Ifw9F8SugI9LW9YUJAv3464c4Nh
aHrStOIVndeqNm2PwKFB3WA4daxzJdCHHHJY3kLMcB1owIr/U9+xXTr63ZuomPnJ
2DkMo0O2Dgg6uFyDeEn0RNKxNgVWwov5wwsQjtecY/Ad82YzUctkgKmQkPNqr2w2
OAZsFD4B2okmjsXDNW+1dIxA2N5Owtc59a+molt563o2B/LQA/oB9C+QC0L48wBF
SpMMpIMzb/+nurS5UFUvSGWS9A50nNEQYVi5w07NvDmK+KCmqTuedmNs0CBuZ8n6
em9LocWwMhqCY5fuWOKRI8IpOcixoUX8delG9sTgEucWZh6iBjFE3vZ9reBkPOw1
cYphK5dCPAGWpZUclAvpcDLODr6WMVBcW/QsoCEldnmWSwEEq1xA16H5bz3cQ4gw
o3MaMQD1eK9T9XIIcarONgctnUXd+H6co06xomioziovDbRWEDeTQ9o2xbQxKOQ8
k+TmuXhjHpzo/hK2rKm7kdRwLEYlaYYJbj8ITRAGvNE82iFlV3S/dYEOEqGH0Lri
tnWOhAtSWIKr2JYnfm5kksd191Mz13wOV7UBus+Ai4Kk4AZzPjCOlvm0xgTwTqPR
hj+Vr6FYj2LSQXsJVWYPevy8mz4KuFr3176cscgU5Aufp0A0m+iABOnO+FvwTxdu
10aRhITjEKYxVeukZe1DBp4v75EJpP1UHaJGcREl2uqqvKBfdTRqd1COpOhhRgSu
lSTKCST2cc24NT8gZa7nnJ8UfzamFovJQZF3hpFWld5rDt8ZYiCjFzPRkS7PhpAs
SNkOIS2SjNocJzfJxVhH5DhmGPcTVc2hL6HFVwnsk5/PouMt85yW+C+d1HgrSWcb
HkkJQJsXriCYDxkaGr2w/ZV8nKL8TIMgbwUU8GtVbPg7FiaH1M1Fy9g0ID0iXKE4
FYYdJqGTJbwtGYUXnbGEUN1Cgr1lw38btcTlrethvsS8guJ5h1wiFrvO9t6l/HiM
vaSRFL7IjMgL9+OTmGvTUlx6kWBGdOaYnDLlProPm2FlkRb9E5mgNu6NcxAJR0av
0rKpYHOy2Al5FyfNdZPDyTodV4/YN6wdHeT5iRp40u29GyQjYreewLtgm/GHg2pX
q72U2DdT+TLJpEaxT2eRedRZf9ive9nH44wjWCYy/+Dq4CrtwqmYYPFZDDKrZDxj
fTVJ2LbqEy+7/zzXSVnA7F6R/FNjLlz3UVY5xtwI5QTVuKjwkl+5dp499nIwlMga
mZtLR2WyNDYvhlbn9V0CmaC4iIebeqgQSiruhY3fEgCGLW3N3/352gmGC5z9DMG1
Bq6bT/dLGNZAmfdS0PQVWI+UaAQev8WF0AldPjQY6SdZ9t0FNqhuKiIL0nqLvYk4
+VjQWlKxJir52o4NNt7+rV+A0Yj7hmB9iOb3Uc11fAMajgo+0a11icshrQCFmfAv
KN44nUpg6D/gJDgZnfhDGF1Lwd/6oOb3MOzb7THXjwtxi7BHhgOcPOPERQeJUwD0
QqHMDR2BiH81QXA7uDDSlX9u8VwZl00hqW8P9mzWEtz6DDabyAsyqZa+kDGMzHEe
469/PcQUfbkNmRAQjLsrop8+o/1D9D/misFJQJSUJNlmJQXvyvfTnsijzM8d14Xq
d5UDKaRGB9EJUCOfJSIQmowmUb/WsHJdY0ahk3M1KR+ulvbNcWjvF+A+i1aDmBL3
LXF+49Q78DvAPdd75OpzecrfH1hl2Zm66unuB0ahX4X3hZwYrmRIdOzCmEcZlwyB
mFTrlfh+LCnsUcaoalGSLz96T1e2O9amDnP8PI18vGsZ81n74GiKLew97fw7FEni
FhMGVd2N6WnPax8y+YQ2FoUL+tciGnRwhib4IOpICXfTrBxfnBB7E2Euo+g5YYO7
tBxeZ2crw6G6Mg6xTutYoKCK+Gh/tCQRIEiDLcMB4aB6tcNSLKwEPXNOuMCS16vj
PksggQ0c3S13McGqlmGAiNno/mcToGsPuHgRY3iGbMNdALQLviHVyhXcedWywswt
ooHkxfEpfLjtMTijXB4qBrBp0gtPsrQOcIM3+I8jcgHh16rUPTwBNpxfaO4LLrez
i5XdNzHFRdpLdai07kVfwT6oG1GIc4Ku8Uo+DuSemqdWfy78aXf2VlXBEB6Q3oRi
SO9XR2pG1+nqUClNlx+8PWVarItyr6//7AtAD4GRmPon+ZE0Jlr9lBBGn5NdimAd
Rq+LE9lOkCOZPlrHd3WQHKH1GC+c789iQOTl1VmXn7polX4ciemlBxGV7h/MwyX0
mhcZZapNR39QPdpO0dvY295ZzqpNWTniyZLWUwmTYLQjYb94W96RYlRT3gdTJVkv
OKir3ldvOQM1G9b3dLmmjbN3iT5HS0GitZn0xLz5F9LvT2xcTxOoRih2vDT5Lc/R
aHDC/QR7jFumN/IZgQK2s6vJ03dwgcSrIEG03giOWcewBSeLiJGozHcw7KfVt7Ej
EWEVFHBLrjpIvPdcXzyrI3I28f8zF4g2IYT7lhhOb3aPlBn5Yn1nn1jtIrnPN9LN
vSt13LceuhuxcGQnV7LTwa6VDkkJMOAX9QFTrFKwr1gz0ZxUbf+xtXAZhlj0sJj1
PvgZ+KkAAIdi47HUAtxihbni/QKEXPrvSNGnhfbVYTQNh1Ut946IAfyZoHLpHSaB
XSEZtFRor1qI+cUbk15O/EKFiQzXZj7clfT6YkOdcR4skojTEruAbCDJ0BGJ+gTI
vh5mi5TQXDKNeUJcZa3vDNC5LE8SzQ67mTKTuqeYdL4UbzSEZtNS6e2zT8D8YqWf
KZ2O+ZvJNon0r9m6qWey1qTP58qP3PzB2itEJzr6dSOb97PbUsxIaxiRfUqVaGvA
XSaJIDYvh82TJI08TuVwp5I1FhsJKftqFYhXyuSe2X6XPEFRkXQS+8/oi3xnRGh3
5sQ3Tj57qYqW7Pid8aiumfkYpcFs2uzu8r6QtRgKrOKcvNCDDpKb5XV3G1h8qBkA
TS0NCNg9gJGlpfuof42J0vwZDC3kLLgkfnwvaiMO6DZ3NQAiclWXyKAL1ADUk71Z
r0q33oY9L27+fZIJjdcdT+/SdpXU/OQn9SmXuYoWKne17iZHM7OKkjhE7pr20PdI
7JFJjWQpWF/NVTzzGxaiDhP0MzreZw4EUhU5NPcZODypk6SEqw+4+O2um/9ht1do
GUTyYbI72aVLLDJRcV5k5vqoSICo/G5KgihzEEDy/c3MNapOReZ1kMDXDySgkz1c
z9zHnc+pX4orEWII0OMmkdFoXK7G9UCx+vcURiZskJ6MwQcFLFzCHtBy/PkXxp5U
9Xc2Ps3IMLP8Y+K9qNmyN7rVLnAjT3/1L0U3jD9HixnNkKitBw7EfQjbg9lGw8sH
ZjcpWFS7LetMEekLhGeTgHHPyk9kyrhRTh/7AWqPo2rU2z+dYQrVhafrneOya6DT
AXGlme8G4eCSKQMOm9TOtWgjxXDQGYdNsL2I70mTsy8wcvPq2n35QfeIIgaoJxiG
tjhWcsitknl0WMjo2dlpItHTJoNX75B/qKcLd3ZQ2xcATb8zYyNgApo8qVZyLScH
OQr3rmsvkb+2PwznmvoMcl8ZS7/sB4RSVAu4HXUP2r0weW9y2JoMm7A0L5ZFetbm
7qx5QrV/OzqAhi7zqcx2WMHLmSeHm8WnwmpVn78Os8U=
`pragma protect end_protected
