// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
k+r3rOU9Vu9Rs/jkSJBmxSI8Om/YEUg7A/POqv0Qc58sfNFyokJ6F2C0KUTOhoGl
Z5ucbDOpuLgfNYw8Y6Mbj6MEmnn7Je8TQBAeRE68xx+ERzvpDH/uaRt04ede4wkk
xMlxMXbZQJ2+6Xk1AuH32vZnhkXyJTGO61OENwQuUZ/PYw6lWApfDQ==
//pragma protect end_key_block
//pragma protect digest_block
wVEyHWmzk9ExhGq9XLR330ZYA+0=
//pragma protect end_digest_block
//pragma protect data_block
QAO4WQnj0qctBZQ1EFG0QD9vD47S9a7CoF7eEXVx1u3k/e9fFEU4ACqhsaZ5vsfg
AvNn5xX+eAFf9q0w+gPCZG+fjtsVeiGbrwO8DD4nf8mjQbsLxHz1T+7MEJO+8CVd
16mGz0KUOa3j+Kd3tKCkthJbOuDDfA3/NGMz+wKXFrnxuDki2iXX5f2HKIo8uf2i
wVFoRI7HeLpv/W5kmqyzKMAFcox55bBaFrbtk/VtGTfVWUvcu76Z0eewnK7xhB4q
2J9qDGk405SVEki9jbRlFGggS3BVEhiFSWnsM/F8+vRak1soyxFdRnY/pkp3+xaA
bt6tD8C3wSg8+DbY1MObcEkrHciX1yOTy/2edXOMeOVuB+sNMbBp3Y7WTZjPhjQM
qXulvSykGWs7vtvj6zZHKs2xnGs0ogdjpK7kigasWToAHkpc/GOhXITD61Fir6lS
NV/FeKIRfWY0Dv0j9v9bPwoTXWu4vkwnbVK3E16HTKhD4RiOhcwX1mlGc+r5XuVN
jid3JzDcaO8AN5iHt/E67F7s7ZrD5cn1f5avueOqdfJpA1rlF2fVLCoyLKdeP9t+
D1zxNPLwFTSk1yQdHERrbiECIT3RFKvYbAfBVekID6gV18kFTqZdSlrL/nJkrmyj
0z95vg2HwbbofpxRtIR9X+mVKasCsAZfMyNluBjQu6876DiuYEttEq9KcPUahpjF
UQgqTfOanReP0SJUlMnn8wIzlV3nruDRGZLXdkGdRnkj0iSBmW9nGuyr9J9mk5CM
1jpo7uL/X7lrPYMu3yd2Jw//qp71BdpYaf5BLv8TfObZvPGhAb8hqQCAfdk75OZf
eEMDOF9N+tYLwsusHZJBWikoh1jEeAWR0/O2wjMMmY3j1uyS1iBbr1kuGo0goDxq
Gh5XPMigFDmSKBb4AvipMn+h2y3ZyZLq+UH8j47PocbDSpSqvjM5k6yTJhDpm4jv
AT/OIlfDumKC9FnRZOgsnjGtD78DhTCPvlxcJ8rEnjSZFplZRT8uafvzYm8iGOlm
HgLmZ58UTJSlciPSDUa4fp8+RCjp+MeAtv8k8zDcwHIFDEPYlca1uHtNGPBr4XhW
JElC5uVbUr0IWl9MisjX2JphcC1BmthOIfg3ffAMT7cxe2R0NI9NBudZUDM2sX3E
wdC6s9uFla+tFqrECR4zAyeBD/a5T8z6mw3OKufcrig75w+fZ5twJ44998/Jpxj+
qaZOsuwa6XtBgDiHYeYPl8OZWeb6y2f16YzyDGY/izMsWkwmZha4LVqzyhzA1REC
hE22uA1/BXKQD7g/R9zf+4ddDvOLey1VnJ0vWIiKmeBcNGLunUOv+vrCJ2xtOBmw
JzzrAofhDTpemwHkEPPsUNGFOKA7qyzn2NIS03aefHcXRTLynAfQb31B/35vN10p
H6nvyAqWrbbjB0CdEAivqoWnWCuIQhpuXm6Nlawn112z6go41tT9xDpWQHf70asR
WnUD5nSbTyrFUnJFL4NuYkI7yzS/nCIUQpBz2YlqudzO8br7m8Gox1TSJY/wQ6fN
TTECnoLI0dAwIKmvrTXe13WIMFrc+hZ5cjropP/Mx+VGw2ew9mzmqGqbwuK5g+KZ
/FK37mZA5jpwfkSVy3PqWa2AX5HQA0DxJfYHHvMaLoDPPCKf5RRxBIFsEmT/zZyK
ZnJs1Zwz1iC9vDkmAazVzS3ebyqUrmA3EMgJ0U0c2LxebxyEV5zWO5p2nGiKIdOf
XyJfFNAbYEMTvYqZguh1Q6lcgp+uUG+yeq7xlku1NskznqwlGK5s+i/yWUpHDoEJ
ixpDTxmWhcWoMxm/n4DyBd1aS/RFdLrggyEK6XNckM9lZ2T6ZQ5pPklpTaL4oOUe
jc1nso5PLpCiy4UWbP6peKdtzMTV+MupGPW0hSiHUJlRZ7HBvhQ2acXLw7p3H2n/
KMjoRMnc8r6MhywrIngv/8ZFeJ5K4rGCEh+FNwZtt0g9w4tRS1M209VQ71EKKlcr
cBXhngwALgkvXmpkedkfb/Wqh9oFPmAE+ChLa0WLwDnxKdA3Ef1Se2hxgjqxi2Vw
yJAPlfyAJVhEVz/iZQijPfv44zYGWqqthRs+ZS6kQ1ichtnztW6cfKVUGsHIzOmG
kRK8jS0cpu6Nhsnd3jsBOptSLU5V1KlXQjKvZ3OGORD2y1p5xAI23czwa3AN7FMd
Yg3gi0OngCF3x2k22ed05pWspwo9LZqqJVaP/z9mONfH0o99aq1vQESS8jkAvHaG
xpTwaESAz38NIMg3Zuo28Ti/YivM8xhZHhD7mWzMJfGkrurdHoQByGcOvvrUvFek
tCBfYkt0NHbwRB4NrggMVeaQ+coAjwSzQIg+kSq4l3vQSmkrvdGjbtDYjsUJSh+x
k/X1XDNjQ0aKFkPEREcF6bnjc4Q5LUYY/6InCTEDoOELw6salG0ilDgakRTkCUJ2
DkCpUKd7PHOwdTJa6i4wGBuYv+47YY7ePzAPVohmC+Ea/Vb0bzGhmL0/cxfQv6LS
hlrz55XGvRUIoR3c7ZqQ0ppGsfKq/wZj0ACs0FExQFHGFNmJHv34ZJxIUb787KlG
Vx+ad0N4vcmxoy5VNQa2uZ3pkd53/riOEcKRhDbKMNgXM5knVFymoXWZvLerScHT
H1RlSvg92zmcmczcHgBgpjE0GGtSNuwqdkBG/Ncd67unzg3reRJchZ1SY7Y4Ngc5
6WqmwE+lW5GrW8gvnVgFkdZd180VkY83uyk4ScuN35Tdi1nfTXGCq192VN8Zzu5j
YODCR2bxdUVs7kM3QG9LFezU/QqfJwOjqMIj9/RAhybnHIqJWjpTRDPxh5fX7FC5
jxaXOW3QU7I5t2R/nru1mV6CNSSrgzTa2wVoOds5NK8Q8otMCb3CxtdGgDgURG42
iYWxRo5gHBByDwZ9M8McDpFlELwRd0geo8hN4PB58qNZyuUzaJVcshnHc856vgza
Hz5WNpeoe3VvhICInYZxTBdcneHMkDjaapqhJUZJ9khXVN9K7FTTjbgUodwgjWH7
EfWmEB2wqjQEpZkBi+5Xl+mXynmAdER4glBmyn41QyKiAIm6MRCcI1D3vVQsrK+a
LgEsujDoRm2FbeBlhbSgpb0MzUmtzPaCuGLY0sB/e/RBAaOBLxhbCooH3XG/cs/2
DzA34jPelKMpQJrJGiGTSMuwREDfEnvYkyPO24KKqrp920X0fvtepFzKmB0ig/zI
ZjzjpCYftz/ukKq/xRaME5ssZsdqLzylEbVmpku3a9StQF294BObiSqsMJTnLk3z
oKD3isknJ1twdSBd7g95t3ukt0VxlB5XzweagXrfOM4V0ZMi8v11s7xjPOlm4JcO
I0FxLFvKDTd+a4Uj1hSgVIzFUNQbNXhF2jOaxuTFK0bptE8fHxXsocSmWAB0LfJF
F1p2JyAk3hplPApxvFyai47Vj0bSxyL+PLRR1LK4/zPfjadmuGYOqpYyEJgrKlf2
LO7tulf0E1Ew8YgpMMCYDMEejs/t3MtjyNOLXA3pq1lvcv8yK+XwlcO5eZcvF0AS
LUUa/hhSDEb/TaG+SSzGzVS1yTQPrYJus9QJd0LaDmjV0wfpNVoNWxckSeIOS7Eq
1GwViIIPA8FKrRepdJZr9s+wDJ0IrJ6QdsKZtSjx6nAaCLret/hqbjBbb+7farU2
tZSDMQ7Q0+XloV8xmb//NvLTGkz/9HlIuIluntDh/KPqrLKEwhDX3XBzKY43S7lj
qmULAQSgQf2SWjVmITYOhhrMBuQwOlkEFTr7lT4k+6gFse5HC5pFzG0JVKuFfVN6
LkunPGzrE4TGdRGR/j/mTZ3cYm5wmiYH8Kle7FPQCKhvaprEBHU2rVPRAp1QHUOx
KqG5Xtx337l8ob8B5kd3SfqyavKmwZKPdZPJwkVMfkDh/JS74euyzO9Q6NRqKWK9
G5j1H1Xrpw31kpWhq+ndrtNQmmOnkkaN0TPQ+fchyRRBR4rC4zOpoCKFYrMGHRAe
riATf3xNtpGQKpjhjyo/f7CrTD4rQKX74O4jrl+Y4xM9cQEbTNcOtY2UGPcewEII
YGH16mZ1+85bj5EHMDfIcrAaxTrSb154timGccc+HPoxLKLhG2Oc8DDaU03HUV6L
t21O/HHFw+fQIjTk7u1d+nhwh0a5xlvVQ1ASo/gCzETzLeLrdfA/v9erFfykv7v8
2v+VfVI7TwTeQ+tu/hmSvnsjHMF5fXRd5ThE3HIQZm1WDPQ/oaApJWinJni2kxn/
1znmaF8Wz6dKeiYPg55rg61Bx9N7CgaaDIbeG44v3r0NjYlV2u6imbkEXuckEDZI
egaQmg1nPzTJuf9BHbwz4jgdyWDpD4uTznI90aQ2ZR4xZygaIQiyPlFs7qMis1vK
lvnutCrbudmiR2XvCyq9VUg6LBUjItJMMFF5grBSEM6ye9ZPEuIGwJrLnafPDIRH
+t1erDXanebj/ke/ckJnnLL6mUN9ml/ZcWdbZbiMunJ0M7bnJbjilKrKj0Ng0QNk
qGToRZuXadO8+VlnQf1p2008WtQr85uhD4S1lFYjjECwDveCE02y36z2SuScGOMl
PLvNq5haddz8/kYraKxlaMcN2025hFbTNeF7iLGfoaT1INC9qdhmm9obW/RZKlD7
x5YR8RRtsZ3TmT8XWgdcPkxKOSuSTvRXWVdsDGy16n+DRYK/ZijwxFcgT6n+8flk
VOmYFzya0vw5JAYd+AviCA0OupswqQj1b2R1dCjeXS+U53yOvE9ISoP1o26U38qu
04LlxWco9+EiOXyYRPMsiSDJLDkfPoKsLxHbxOeSoFcHDsNkO/Z1DxGZzaXfZDsf
jXJhWJOrjcu2v0u9X+3oxgvB+iWziJC52T2sMCL/beR2FsJi9nAo/X333ogHwzJB
b/ktTXAdCoVe9ZbnfPX7/PrF9RC2ENlEK4RiwTCyE+yqPGNuYibsRVvR3IF9Q5kY
b+JKq2ya9+j4H69tqRc6Da8RIqMtp1msebhpCTpqc/jBRgRM5RsTYCPmbjy+X3/2
PYdWE5quLrLk/YUUjhaUAkTHWL9JJxpjob2MLOHJNaqdBLTVg1P51h79BtZX7kC6
Qt+wvBg28ZyxGRKS9oCbXuS6HYtNc7NF9UtO4ALpklZRopcMOM7RSUhFeFlyvFy1
62c/A5CqQ5bKlp9nzaxTWdNJ6QPxMdePGlPOEmSwiTg0Xk9x9lAvkajgH2fwfN/u
cwpTdHHprPFGyPw0gikaw85psXO4B4xxqzQ6M1c6eSop61roucE5GMdyz3h/fpAE
xIXWu2aEb6A2pedQF778+JdQ2U4e9ACvtFmx3bbDOZPgC3xy9kY4DubNwVlsRZSO
u9OoERApYzBPIlryZnpGmRtiQciwxvcjLEmxgORR1vOWLaT0jADEqXsUskP7jZvN
rz8do7WbOU5MJ1FhaJLxqVTgzcw7SiAGq+00kxWG0hhCoBblyIKZmvZbnxCqTArx
N9XJUP1Yz+nNLL7+X/5KHjBY2xWDWKSHEEkkWl/YYyFMCAHeXvhOxE5sTyCUvUrP
SMFceam/Ls/vjiSih+MYMquQ+nL+8Y3Kpqc9SP7Jgq/C2SYHtOeff6Aq7lYsD9zf
ocVqaqkDFpG01PCC9aOKBzhxefRqfiJxrqvF0nxkgbT2atjb1IcrdKw/aQzP6OZ9
B0FYjHhQFkywmYgzQ37O0nch/1CPWLlT7IWCFWE6OnT72NBlk4f8kC9KKBcaTrRd
3ugKlH48yQTRD+LjB7pLmDTAU7/mmNMWTfvpCma0OVAbKEAxRenkrsbDyzNjOhJq
8hGJ5U8S0gYLlNv8zsfxuhSb2e6OOeZ8GnwvC8sxnKWYL7moWF0PiGFhq4LMSxxA
79g+4sI7RPSz5U/KlcvftoE6vDuPeYYv53FPv4yaAAHuJ3MZ8Wv6SoFRhuMcU/xx
vbHL3SAduk6U+5Xrhles+8+W2j6oeQHP5wnRi9+yVrx/l+upta3FeAJ/rrMO5ICG
xfK1f5lWXX3fkmoZols842jG5MsQWhjoYnhHi4XJdWlWsIAq2cTmborkg98c9/EZ
SgS56hLAnEN/a0Nnni0NP+IwjAhq1EIVfTQLsa8f+UW8AES0tSfoUTVLGThYTzLs
fTcU3bI6OAgsoDQio+23bW3QZpbPpq5ltFsTbi2T4v58Ml7ou/lgVaTrXsnyEdW/
pRnsIkiWqGO7Y5iAfIGnsxYqeKELw+QSQkVl+Gw9mjHkyWr7iaH6fkV4bITRl7wJ
pNep/zhYSOaIM8CywR7S5m6fPxc1NcS+lWZzmKJcFzTMFBIZ7vQbuRRdmO55qUii
+eJRXgilegPxvcEIVuWwC9ht3y6VAEltym5prhw5jSo2WCZhll/CZzoXWF/4SprD
E05wGiEHcRdKuNaA7mDj3IxdpGo7fGLgHY3OGnEFS4n25Q/ZoBKoEpXmxVwrFA+x
YendP1ruOjOc7bdwkiyRm/yz/zWQtpbu+jOPML1KexZVX72Wo+r6reuBV61Qrvhs
+HMdD0jjgRvbwhgsVmT7LhKA7WcqPwUISWdz4l14MAsew9AV+zdlFLxCHB/pP9ga
cCag6moGGQqOLN7ZtRv5NrqcdD8uv3ETwelPD3TjTpa75Qd2QSSlYp3iM2s5fl1I
L6l781IwyMmxmbBnZrEpYlgXQYLzY5hDvHysBzAojKEifCBGLhWMU/dLTytTyWRS
3L1ePjkM2IQgR7gJ06nDBbwP3BztF1nEPnq14bf4S8IEYPKi9W3neMRnrne7jaBP
yJdFPZ4P52fpe780OZM0RYrkdEBmb82lm9SgAPW2BjddrA9+lq6CFIjbrDcUFN0L
I+Ls5rBvw6ljRKx0CDOTLEf782nqBcCdqyl3K1Dmt4RAqBhWDwJ5oo9sshcdrb5I
+8W9vEjnnMCC4kOMrgKNMGkQgtumREdNOcXLjXd9TRAI2uXgEqZh1jhv/s85vaIO
Sq03E+gwqoJgVeHZyIt5g3WbhMjdHLfevMt4AjV+Q1Hb36orKNlxNWz/MQ75eMmC
qjSEnaMxBXf8h63sBzP7CW+LwPqwUe9GxBrfknbAjNFMs3awQdOsBdh+WkCJAaq8
7UaGfPS5KDdVSkJWUg6upQeOaXlBPIKC0nCVk8ymmIZX+OH2uGqOsppf4c47ycJy
4ezzahldbRcJ6N5d6s/HILfSk8zqcQCeaYIwlhskTRo7N6bH6H4Ji0ad4VNRiGGs
qe5x+MLgOVVZ/CcZ6oG7aGFeHN8LvTsDBsjwVtwbLAhZ2H8VC9TJdiW4xdWy4SCH
vHnJ+1MiU5HZb+Lwk7y36Bifv0Yhxygqi+XmrNkMqqBlphD1cN/gpEbVN19EGgxV
CijhdXW7MMyRFlVwXf7LYmiXOCjWzpks2Vf/UDAj81RLsYnX1olU8C62fGjxU/lB
5Nz5aFQlo2yblC1r4e8js3kqBo8qd7xcooeEuYhK5WrPqsV3MNtdJDi9DTFjABFU
1TKpgtMfx9nuasrIudgGSsFisVbKTQsoyKD3Q5IRL9MWjIUui8x3kSh3yo/uvC7q
BVkZ+aZivj2rv6el3HVWzUQs/vC/yQDPwHkYni+f3btZJJwBUf8P6omPZS9lhcFg
H8xfxEzLCOAU3KneMb3REhV1l36whpxpIw0StTDJYb/dC2CS4IaQFQSVTsXqr8JQ
JYTvCesWpOMyMPqhCToE4+GXrvCRH8kEFjpvOf9VLsKnzeoi4Fj+E1ZuXVwYYBMy
sbnlyhr87E9iON/F3q38+iPKwX5FB4LkuMkMF8xmQtktOyv3COvMQlxwIJeGJXhc
SEu+aJxkDS5fiW2l+gw5OE43/cMTLzgb2q9ihB2IXZgNWfapB3QaV/hPNPR97HS8
WFmwd0cnkjdGY7tQ9h1JMN3oca9mD+aLsjLLwwzIWG4q5nSnkdSJGH05rclb84Xt
1QbOHuyDzjS9ppx8t9KrEllF9jYZVpABXQH/O2gar3YH/LGi7bQiToWdsPSfe6r0
Pbp/h+xI/7M7d5qqJ1hDsuhF9qsgoBb+K3K9Adr+JNwbXrq4sPhs2kHWEtsnLMrt
Zi8NkKEe7DQ2UZhhcF6171xWk3jbfrZ4AuJeXQ8GMBGJbJ+luw2xDPX6GNPaSf30
g+Ik0pV3TyYtn61YvsmQMpB0WalmsazwdpBkpsSO9sII0bPcey2gYAxF4yRIbcIQ
NjnnmwiPghM+fsx5+5R+Z9PUlUkwJSUEFY/JaS5bPihEKhe0O50KzX86ay9kEAkE
Fsuqkc+JeJ8vMO0bV09Cjo/RYgp/F1lDkH+xH9vq+vuJdxRx+VopjSHOIeUkz+wc
mMy1+s6zZk94HYceLrCbE//jcFM8fzIX5o41P8WCr9s3HxQbRrTqcdbedc+vGzJG
Eo2sUHrPbFQtf9cx4QEpb70eCaaU/9t0o7XPhssmZGHDTZ9MNr+BXxkGkeaQ2P0d
vfMzfbrT0KPmhH4i1XZcA0mWYlze0NNqWY3OEhpSZ7sVDwLzyrWmc+OTKZG6QCq/
j9fucY6m8tQ8VY/OysQy5KBCROgEveyCXyFyWgQfdOyRgDFeW+PbkdLy3JEbwO1w
XT5jX2IdTF8HyYVWSta29Fs4E3SAJ6tM0U4p0EUvkVDjQJGgQ+I3uST3Ghk+i0a5
pbKXtfWdJmZ/U5NhsYwIoiCSMITprF9FTWxI0iygfQuKcb3tkiHq92NLTjk6q2vr
Y2Pl7rNs/xyYArw/0E8PXaz2wZssHRF6rHyja9SIBMSfcV4vHBfuJvhAPZAFwLy5
VsQgSO8HkmUrnMYuS58Sv8hLsjro19G8ztOsBCphghoNUauVpI/qAdbJgfHXtZyf
CuTwh/o/Leys6CnHi1ix8TtYtgG5LMtsLcQTCVroAaHlqAIbvwqF8MtQ/wT27CIe
Y6Pn1UbaAISJS4EDNTlnnWwUGF/DlCA8SU/uayEDYGrL3ZAeLnSs0FYVDsm+GhWo
OmINtrEa7z9pvbpOg2gu/XQgwThqOpePk8F8aOw7yweqfHNa8scYeKJY5hJEOBTM
aNpVlK48YwKsdzWp+CbqfTDQv0f2jFTT5JQFyAxqEOL4T5x0zKfP7wkTBfKRFaqU
ysavwENJgrCXmZYlKwg5nRCbI3KFKjAyAW6a5oU9c64KGDKsYleAByWmRMU8B9wK
j06+zUPB17lFyxbfVX9ls/B+QeHYdysjb6IR/i+OLdvFv/gcH7Mj6XI50xusA5MY
wA1SlCcnQNqg6N/01jAATTmfGknJuKrrONN5Qf8RLkMlPU50ysKjUOtcDOoZcgEl
yAFCM4IX0diLEeQp03dDouvZ3fuK3W/IB6f2jtrrlHcE3QJEuOowZMYAeiUvAtQP
FCHru1FV8e55bbIeTJt0hE5G6rDz1snZaheljRgHuxCJ/3zjXgmNuGyhigu1Gb/c
uCgvodc55TduwJJPy8FGWxYmVztQU0Ynv5sJCopxFMmwjtFT2OyZQYGSYjCf6jGS
o1MirMbM2oZ1w8tbguz7Pw5x7jAypuyPbcORKG60LMdL51eobyfwYSQNhtLsjT9j
XTpzU4PToGtsYikN8/sFokXL1RCBXoenidDc/rCOamaHYXv6Oh2e1GksPAEa5LMj
XCYgUOOMesGatS0IxCX9XXFUHoNF8EoELo0+3/X5Y1RKNzl3Z7yOkX38en2kjw3F
kG3LPXCJMJidN8DyovMMu1z5D37B9yjmrp6RvVl+Y1tmgaWtnn3otNlReSnKiqWb
gUWFJAMdFH+R/OzFO8c282Bynj1UMU6QGCG6choyF8WmAjLlshevl23D8fh5m1LN
PQXUMtdzUt9jf9roYRgbNHT4pmJKv5fbfJ+np53xPxXioOncurpAzqBki/3XfwlG
xSCbbQ896+8VS0QfdxAGSa5VVyyjpbCOlHZ96IkJrbn180m+0+KC71m3ZCegepJk
FuGES2X6C/LcidtcTQcKfIpQ1z+CIiTLp79EmmI+NDdO7J2qBmqhgfGQiX2mboqt
VYU8AJy6hu5HOQmgUl/Y0gaBMlP99rnvXviWo63w3g/x3deacl17IBQr48yy+Kjn
ZKKAlc8DIaWeIVZn6RmtFMJoJ5WbvcYE34N+YxLx6oMmcGaeAoCQA+BgIRpWsC7X
gXr0/SE5S7hyV4D+UqTD/qNhsp/uAetk+OBI9CVGBpyol6zKomVBT/8wuptED9/h
rFIBl6107eMDBgues0Jd9mT54LBwTe0YFz9z1hUZBcyUk0LYc05kuLgz3208veS1
MXqFVlT7a13AFxF7mZP79JMVQ16rKvn8X5NaaEm/TUnWRTsugaue/usX5ArBHyRO
5MiUC3EoEvd0XW5fQj7cIB9V4ecB0DuSnPAEwHAS5fdAD+nmZ0RYmZqt58CStHwi
U4jq2b66weH0b9rzV4S5W6deax9mGQ6VmFFBDCRkLcdITWEDReGP0Ge2ef03Iocd
/S/Kfodv0CmHCmglGEhWlkbM0yy1H0arU1TLnMhNdt8j4AKyQB9gZyx4U8Nxj6Q8
8YnqM8c89s4VyFifACOCKITMKtc971pGQfgKXhb0etAunpQ6STDvTcBb/Ps+BLgV
/sprrutS9w3jY456ypsaF/c6kyRqBDDqnwwhTFf/az+sMfZExEZqq6gD3dZ9LTTS
lh8pbfH9OAG5+zjsrUpMvdrTHsFdRLWE0HdpnGL0Rg+r8hTjtMPBr0d1zVOd6j/u
8Sg/ddMsKHH4qaUAe/MiwBDwG0Azuqz/DdmuXfNWb5OY98gfsLZbHrmQKPDEcmOA
PDKTtO3Zsr+PR6MjvDUj7/g76uYdThn/BbldmPry/eWfMuqPh2aAUHy43DuLs2Uh
CNTUWEdbpGWQ8/0FYFKT8FsU8kIsot3OCm4mw0UPS9Nt2SsqfmCV6jv8GTcXLAYl
JIsf7vIbDF3/ARu6AsKT4GdvJRojvmAKvTmvQJv5aPsap52lffqnjzrCWUvQ3O6u
XCtKt8a2tjybrzbeWGmlP+VnftLrCp4s/XqX6KS9GtwpV2zR3HSRzRQuyFmZOYWH
8r4MmIgT7bmii3QK3UP6K6dG0FwlnhlM4MSuYRX4fmwVp7mGtjCtJVDzZE2TdWos
Q2paDTkepmPzbz9OvzIaL9JHET+h83Y52UdEiazUV0NSw43Job+QQSwTwZwkzKR9
ADFP3DbMBN9VFG/hjZQCa5hA6tQwKAPFKJB8kfjtWIx5fznM25JqJKndBpfNxkjR
2GFcX/iowCKNLpNhcjAHHWW4Gro0OqU6Eh+die4rutVgyySz7rOOBhCWhuD5N80p
MAYL873tcJ1kGi2oVBfPSGJC9vugggq8jaw5xbCWJu+/2UJWsBG/ZPOP2pjKF1S+
SvoNLaYNNV75Xb4PJpirgAbEejbqNEPbBwu6U4r7DYKTGOySGSobsyt2ZpDFRIi+
oFrsMiDX1AqqTctG6K4IuVk8myqVMUDqSkB11t6e122DqR93g8DI3038xh/wC7v9
02BCkk1yig41LcvhMceQ58IKKLoFK2nCoyOcXUN3eap1jAwkhu9ee0d4/HvEeq2n
yKWNsvjoKW9ns5uul9Pc4AZ03JXmnpWiQTmKrYTwXFeuEro0keJHayWrufgvWGWz
3Pqh3kuLNVuyMrhkPikeygMwJtpWdRipOvC5le1J7OJ7tzQxSq8Fo+KeYMmE1SHB
PYeHJiX8MWjS6k5eK/itPMBBT4mbVhHh0/3Vw0PkNNGUcYTa7xf+/dumA5zv4/dF
WkTs1ew8c48X5MGgcc0zgXTxETt3JWY4eInn3Bbuw4KcdX9qjv3JCC5SfbpMMfGL
xfismAhFVTsJlhH0PVBm8K3hU3wWj8yyLnKbqmrMZUfuSpMsJKSn1wnBsHez9Ovk
nkkely7YAfpHan57nQA2biEJE804zuQCCRXZrzHcNQWXwE9tPX8jC6onsJEI1QwB
PXceSYSMLJnaKWwCbSB7vjaagxWWlgb+PAJGiDqAZX8LffM1B1oaZsM+0kr8j5qv
M3JJySMKv5YHKiG5Jx2RDZRAcNfmUCl0YBwG+GoHty/mHTAgydjr7Pt86lanvcoi
qUoUsRFn+wgMPGh6ygLCYq4m5kp/JMaw2t6UVy+LS6FmR6ju6EFkrJ7617I4XPiX
GLEIDEikLoukFgq6GHTXifGN0QTyzurM011VuXwlr50O6vpFiElhCLHMV0THZMeX
W95DUaZhr6GNP+XDLqsUUVlOnF0Ir2BMYWJJu+D7hpMnXc6ie8u3o6MHbcmr9Iwp
+SFDmauOfuXRdBQxkyaEhZMBIdg3sIUC7WmSuufL6o31FW2JbLLY6stD21mUtedW
vfz2hQ4S4Z/sOsNXzTFR/XMaOeu2X5jQ2Q/8+Mt3p2NxSpo8NH1xjBo+9UZ88JR9
9ibSU3b1tWYDoofA6oOIx5Ys1E3mibRSKPwMXySZWnvYPZxGQpWk5Y4p6x+f96Mw
Il8tqejRCAOxBJ3lfa3rUjmn5WpEWV8nQsbgHkkj52dBC06pODtpqUS3iE+gdTCq
7nsy+BrgcJcSfXT64FDkBBgLXB2HSlh2HFaWex7D4HMHqWLBsuLcH6icNitWhp9z
Zv+zvrpZj6BO2ad+z+XvyUVncoHptD+JOoW9QScRSF4nzPImo6aR+DJUf9KpzdZP
qeYRUDFoPkuOZpe/n5+fZn2p7k8qUV3R/EVpiA32sa9+Kr8Quz37wrD2NmaZEwJN
fUQUfzm8XIFb7WcQavX+TYjTUjdYR8bTNZcbgV91QvsJtwbIvaBHueq3f5fHc7Ns
jUplaKz/35GdU6j3bUTV4qjE+XRRfTIdtFx/TnwOnZHRNOcb066uRM9LcUIABf92
nyElhBOF1DAG24g4Aqe1WuS9jK3zD8QTlwwVaV+bGkphPNZvUFjrSCXBnZQOFg+G
yfeAwmBDm6G7Ex0aomF+dlq087q74PtOC6pa7IryFp1iwnoQAarGaVnOs6utZ+TH
/vmU2d0PTAth8lGlqE2xTz92HQmR04bNFasig5LW/GyUTODfGE5QIHEVNrpWXsFM
MaaavbdkfC2SByw/uHaBvE/8zLRILGag6N/GjjOM6vHoMiP9o1ixWeAauURtCc05
DCZJ2+EpA4kAJwds/ACzN73KGbij6FNawTGWJ0xTAIcut5tj4+wBbbDVrozy8RGY
qBnbZRiKgy17D9SYjeUhHJc9/knKVw8d2yqq0+Mshe438+SE6yA7C/9Ffm/mdCEc
srOV5msBh+t00ZMCVlILKv4Dqpf475fJimjT6lvJQQtPLBNyKUpbsEbmqQwwfSjt
Y8NT6zR44YvsPiMiWxs9MRSh3cXFmQOGuDCLJvDu9+JgOkAl0tLwvIBXryXnfuXS
AYv/ykJ8JEv5wDR6rBgcXNQL0/4KKjimVGIsmYEGC6LrsuCjY/DhZmgmr4SVsDqh
tzKxlR4ldovs1eS8VFAeMzfoj/5lwr1WagltxS5t0sch5ChAHp3biI3Vz3fSw/KY
+squFHSmRUzDPAwiOLwo5dIGBEgSxPNjaPAW069Tw6x8ig95+HLZfNsbcaW79dNR
Mg+9DxUctzWIJ6EziAmam2kz0uCbdayeukrtMyTiL/E8GYbdwPou5rm45WD2qod4
t7MdDmHtg8pvyrw68vHtR0ZddHXfOgxi3UaDV/8lr94PoaUHwdPgXAzwQOZ6Cld0
hkwUuDsQMI7Yi7dcBeetMuwVD3HEdWiLoYFKQZIzD2mu7GgX/r/648bjavLFu/h3
L3jmnCFD7GGfuDGShYePgDuFV/BjBC3zROSaCxsi7iupoaWdwjXz381l5Mz0P55c
mRW6mnCGXnoX7CMy0JrsIZdepD7uzccAzVHJUAcoTMF/uWKZU6UNdTl0xLgQkqkr
K4snz2SO+Lt97NUl0AP8r8/FnhJgLkV8zpKvPAwA6DJy/TptTD9LG/5ZvNf5D4MA
/4A1PcKc4eCQupILcugPZbxz9ejacSjpMIuMAKR7w90Fnh1kQwPgxA8S8pBz1zUp
xt6SLSDyVrI5UEAUTpCon97JO8zEy0z8w7mm0Y8M7h9qpNzgIj+MdlUmSGW5ke1i
cOeiScmlyKw2t7QtQyzdGVCmOvz8j22K1JPd8uSoOeYmMRZzFquxrb53fLuBN7Ei
ah/2xCp9DCiE3sStyh/MqbaaN94lkrV6g9CAWq1CzWsG61cb1Ie3Y3TjDLNMeXso
Xdbii13YjjFkn0y6eJl6oG2TvKgu1V25RNQar35ge+pzXBo+YiKY18R2Yf4hL5YJ
3uO2lt8lNbNSXCksQi4FeuRQjbOhyJRuzWWyvSTD3lKMb1hmxQActYdkz4/eR0IY
9GBXtESADHy9ppa+goLkXKgO7P/NvBpleAqZdk07r8mDAJagBIlyYJspERYvXdFa
69mwdm2KfhtPUaUvUwywBoOZWpcAckqtoNcuhsdHuUhdX8qDWTOY998YxDg6lHZq
FY6gyXGkZmFsZrkXRAiAdb8TRw1E37bhETj+2BZHEIN5kCcnd/D9WTX2F1Uz00gW
FyQN6ZOwGRUp9Ye49LvyJ2pNYTEw/rVk8YqbVFQwoUrwrWbZkPfhknfXuLj70rU3
RxMS4qHpoThrcKNJYVpgYSPkiFw1SzYsKi0PYLyM800O1SIyDkCvP9NGTu2XHzwH
ToqMVXIGRE8ZtfFZiuBGdOfwLRvhZ73M+85lmreswQkdoDRL5be0sCSwMKoVeNjZ
5fzKWVPcdpjVba+eZ5zDKvR7DpoWenqKhkcFfG5t3lYnc+est65ZNdm3F4LWjUZP
VDE1is3QNR8lwMxy/gvAPZfdopMlW6CRZPOIfyaKETXFp/uNKWLPoS/r4jXf7Ij1
vF0lxx/3nbwc2LrPO6FNajqxcqWzFLne3lvNUToizjweNe2Rttf8kpSIKLt0Vz4+
9psqTC46RfJFyzIlapMRiOF3NokakK86JQaLukbUtID4/TCxhv67OnGiuKMgWvzl
MFs1r2NCWy+orJ/Lj++RpBSGLCGDTZ6K5jWEbv9gnS48sKfJDXv+Y2LdBjdrKjbl
VoMZ0J+4zlEorVO18uuRYrVNFiQG/BSAcbSuF2KwJuhAbuveI1i6AvuZfSMC4ESp
hhNGO3KG26MzR4JLac7liXHDjdO3DIQFS/f+IMFvt9m8mfTBeVKTaJJu5zm7f69J
KlzzoqwtHqLDeape/baVvnRAkymNFhVf2MikmHJzKxT7MYnySG8QY88gZQyvY09D
EdgVJeaSjHnSede9L5zhfmJh9xOicSh/tgGsjD0A6UccsUm5m8W/imAf94yWJXCH
EBE2vAaPvceK3MeTbCcFUhVrq+GeBJmeEMZTMRYXziaTPAjOAilxRD0e9hVxPUZE
wlxGxs6htKCv1GYdMuD7Lge6tUh+RGCARNQAMEfA63uHY91XbcpLOWH7z+9llhs7
wVE6noXpHDI2kb3zsYE7L+aO4Nvf2xOaMxQ2tWC7fxGmO7o0O9BbWBjvm9KxWPx9
hvcOiQl0OC9FacJcy70KvwZySYhb9JI6+6sNb6mUqmZsYUNpVX8YajwaDA6p3DoY
H/h2vbbsTwngiTQ5DiF9S1rN7yf25dM2FiV0+8MyOj8aHrMoLKsoxXfnXQBB5AQG
xf1jzbaFTsF2YIO57CGyyYigpHm8+nyDjGpaHPn53SjGg/YL8xidVtipuS8Nlq5u
mYJrot1YUyb49o6hkumTG0voU41GN8+g0qL7/TC7oWGc34VZBjiOpgDYfKPrF/xq
JqtRL13ht1VilI0OLg1Uc+FPJI1e8aayHPTUt4Rsi+fI52UQuCW80+aD8mFporrt
ZnEMY8f7CrID0p1IEZRZEvofUvUgkzs4cMsibjZSkaD5NqGCxBcvSpbLozoK9cuS
2LXMDzV4jQXZ54yvw0dNO9Gd9XHthCVK7cJV60H8toGBypigr4P+sasZ+uxj+du9
YeBuADGluJET7EOuTw2Uf2c52o78q1hSqZL02UQS/cG21Kl0ak1RxT4qEu8TLpgv
SFkdlZXM9cApnTJRy/FvbeDP7xU/Ns0arDTjeh81rCSWSYhB7h9xWVkqi5md2vyM
xOLEeEQgtfK5QzTeOZyfIYsToMBJDQ0EqLIlJ3YiO1pNd04ifA6AdxqaKvHCFeUG
hwM220jG+LH7pD2UhyTZD0uFIchHFJFyVjcYS1LB9+bWX6annZGtjTBhpkFN3ikr
FsfySaaM1lkfvx5x6lx6jYoiqysRidcr1YQoeuD8MNd0U8AvU94UqZDk8PPal8UL
UjXMsgxz4jDHFPZrTLn3incTPTKxMmN7tDYL3qCCdW+d2mwUw8gHr42GV9efK/vi
1ftANcxueRfd/wk7q90ZBr/rPeWmnrEzn8/f1yq5ypL8Vcvvmdr1Uttlrvoh2XoS
TCi8oobVFiEKcm+hG9icHu7JS2Ns/Jow+4fHthNiBMXsb3D/mbaZbVY2rUmVV/rW
GQ+qd6hJEC9FOUTS+/Fm3jyKz0z06H7xn+C2OsYV9czv+uX2dLiNaii7sUESrMfD
uu+rhi2wC3UCZfBJptO/q5zxL8JSRxwZhEtVWiBQorWmpcFI8WbFG9cD7lA+sHz+
R0LLbC1Tg7KEd3lVFalJCKhD8ryiIHSLzoEVPn+A/NFMpANl40+l/QPoP2+6nb9R
UgOjAf9UeUDLzQ3YaoTerc3OF+0Q5Mn8GNlWxSYNxclrUjKt5zLfhU7aJsTl/+q3
WIBcOX8cJGEaYv+KuxHYtRyx49VesGJCc15fMkA7vl8kvBtDJV+bzg3wmV4Hy00M
xvZFmdCh541n2+OgMp0dEFIqCwlJWWn1m8qtUAye3aPpeim2yRjT1COS2AX4FBzj
9htKYKRW8IeMvs8LhkgWWMleY++A+ENzv+xuNaGltXw6YPKukpxWfBfgH0duaMAo
1gY++CsYddHBlfKiJttyx762sB2GSYgaBOgT8gY+pd78NKl6sjijo6lGWme25BQQ
VJsesxHKoJaEHKe0mXuIFeS32AUYOUt1vvvUBrg8HDC/05qFx2UExmK57FaP+YzJ
nJqaNwzjJA0wlFlqAk2RxOfaKMJC54iG5+TThVg9D45+SviYqMVJ+1Us8Yg/wUVB
RR0FDnGtY4FhTh3ip8CFsXLkxb15UyCWNSStxlO6euCRgtyZeS5UqBDCFwtQdMBE
kj3S00KQg81QJ9qwrudkL3fwqJeVXPeag64XOWZsEc4csGStbLRkx1P/O70WeLEy
krDWEj/rlla9y7ieFE6slN3GUU0Rn4c+TRQQlrrCHb8Ivf+Gke1T0QkFY5SYhkIH
jvavMUiRRX1HcBRoWUhlTQ0LCxiVkQbwywl6K2qG6Ozp8KGG9ssNU2v8MuMx/4fC
5UaeeAKETgUI5JnEUK0L/P29C9zDLZXggASJYrww8y+mbfsWKtZkD+89znpjJbjW
VdOnxifTa36wgSbgw+ihVqVP5lIAC6DADoAag1EJulS09rg0RZ7JhTDKpHGnDxCf
t8PBHrl80FhflqQZmGq4Ih6sJUHRosxkz146SkdPfFIMsjZZHsjGL3p66Lazu420
qA3QZ9JhefcNFKj7dVii7wl3Pm1KqSQKNyOmPhJYDgFWhcWo0l6f+Yv1ApfU5AqJ
+XhCrwvpAz0tGem6N+JWYqwAQwR6wFDU8dSVk63Y7Pd8kxjm1uvYo6FkbIU3rPw6
uPVay4ENIZVPh6cWaBf3rqyS9KS8pK6y3mWl0Ucm+I7ArL+uQkgmCMo7oMc41jL3
5JiVCnb1/JIAPBk9qKx9tIyyx1lDvJJwTs0mpk+sRHf3Kzt3YQ/20zVMV3z5AbsU
3JwWKd7yFHFApII0skcNkegVUnJZW3uA+Uc8j0ujtNtbweHNWwMVSND7F+eyXxcp
+LYvfQlwvc1VBuCxJ096H+X5UOGMsZNVwZDSMjTNg46FD6lzBhFaJLCYjHuYXoTm
a1SISXz+WKONTGUXlVgVp6p4Bu9IMzDelXyfCyygzkf1OBpUJb5M4TGNm3Gtx/6l
KPNiCiuHxf5pPnPek+lf2S/5l7BAK06IltWHOoc3Z37YD/MQGjE9+9fcAZclRDZF
zkQztWWXl1IIeC/EBkGVPGhDY2QzZKD9VZTCNst6C8lTeqqj6aqwlfjbVWjYMpDa
fzCwuzCN86zbRjzAfRSV6n6z7/qJLumgifsDyTDEy9Pe206UrPPAz5b5jF4rrcF5
tmRHOQAQbs62g3ZCaMxF9IowD7/QmcxabeTPjfrdEpFZQLMNgVIVNPUg+3SErkX2
YUEAcTpZzFU6zh+olIN9nl2rNRfqS7rFjSkg6HgHQURmXxJvUBfwb09sHAy67Fb4
QICUF64Bp0vCzX0we3DOru0cla8FMhV+ZzufRIcTRZ2UAbbsdNJSFepebjj2ujWt
YcKSCMBHfMg2H69T48KY3WhKkhKb36sQzOrX7t2825fSTyfVVpYWgpG7Y3XNPQwl
fgSPDbUXGaO6AZo8RN7HCBsj35Xu73OWqc7143Mhm0LQsbc4Y8+kDFr5VI7JRYtj
qrD8/b7NMeQhJJxo4RmBQhmz3yYrkqLiHoQoM2zN3zJQ7V8Mn8pZfZog/NEWK7lY
t5w61bWKIDAjWvOkWo9qwU7iWxWkt7M3TWz+fC98TtyXLml0dzslwWtcygsf/PfV
o1VkibgH19AFR4AObnR30jj0OqJeBaZy/X0w7l0FJVYk1nPuPNJmEZzKmhk2cCzL
icZz5vrNFam4yu26s8j8j9Fk7QGzv8Cr7kbPTglD10KXNt6QDu2Vro8SgPqd9tez
4PjqhsYrG8gUxP4/juNRXO4rCYrHpGyIYP2uYM1nSEw1bPbdRYSvcUz7JJNEOJr9
FVnqoDOtKAxVpHTcF20TubtrKBwIZ6+odv2hmu9TaeB6/EQyCzbEY3Qd1nJJj7Bs
77AeULYGMEIwgdRnH76oJ1XZitkA8Q+7xLC9xnY0DwULA6aOg3vGX+N97e7jFS5R
vtKxp/T6I2x69BeR/450isbyguEASzzf2oOnPQJeWkjFTLkAVghtRfdlq6pJsQm3
DzolxlCPcSCzdbAJ969KakSF2hpuhQWosBI0e9w6i9hbZFRs4Ir3jIRaBDZjNNrP
5Tqs7snjDoFZaEPT98RxFpI0aVp/VB1hVv8LCaoywQmICZa+fzvbx52Tyto364mV
PEJVqmNhLIGhFWxl6iiAFxtHYNEkOHM7DQ46E8sAPnMxJoW9ZE84aU7dr5mq3X/d
EpWamHsxrEBO6TI7WdPOEKq3hQpYxxPCfDhAW/Gzn9nx6jXClmgaqttcloD5zD39
jma0PzT80lceLR5ZCAEI2CuS0Kccy651sp9co8EEAp68wWr/aLdSxEc/igFynnbE
T989wwAPnwK5y9TFO3S8iDaL3fz6Cidfb3KeI+8xeBUMaUcVnmYll0URFY8VChrr
nk4TtgnNss5xTF+MYljXo5AL/NhtJr6uGZd6906OeFAfxvcZQrY8vcUgFqf55DbR
E5jaodMb0bdmG7qZFZFNqvXX18IoxcFNOPdV9ErelPK3gukGWN5K/zvR/vQ8dEdI
+rA1btZ3FuDGpyHErpU4tJiKRWPAbn6xdS1kpi0CGOeZ1h3y8hT6geMuKav0ihgA
W6gbS4ZlnNQ0Vk5O3lhPF4O9tSL1Od7+C7AtbTtevA5q2+neJNviWUms25P717X9
rD9MlCGFjF4lVL4kRr+ym3w/Qsbtu6kBJH5PItABxyxj/vwn1RGlU8uMyBrbfAe0
uaD7lyg4ES+5uLyU8/hywRvPahCySDsy5fEv8r1BEJWc7p0hD+ZbaDvfEY1vaPT/
v914g489ckAeYUYw4mIU9isCGr7tecEu43WHrhPGZYTuWW4fqfItaVd0GEuooWHa
AM+64LkGa37ZLdXiNEp8mBJxcUUoBvj9KRaYGcpxAkylVT5+1Y61w/R9NG0ON8ZX
slZ2WWewtR8V1VOcmHtLhZtgWyeRdC6cB+OBjY6bxxkoedRXPNvuihuWIbWgrjnm
t9FcaJOPHYtcFR6B9zN7uNHU+E6WEHPadEqQ/UgzTzz74KJPKNxPEqb9sVvD7r1o
Tp8F0hz+CP2x77NX/An2D+M7HST1sqddWdKXvvOY0c7+1mDNIn4yCpiJJTFrrtUK
fm06MaZep2KZXPfTU8AAgzeiizJqXrrXbwE0UjxfKPyAYp2T3EpK6Ojk8MSJa6Gs
pU9u67gVvMX8EKw+V3nttH8+FIrXm9yqTmM9Z90sS3fbPIY6WyN2bSbDzHp5CmDd
PlprGb7gJuXW1e5ng5EwRQqfPv3ezQmrTAPameuXxp+NA8PeofylXhpEXeG3nez9
ahusFJ8eVgHlpX6B9gsSJxwJEY8BP/wti5ZntHYliPNEqGUXbfek0JQJfcfzXaF8
t9aDhUNOvEUS0HsOcBFR874d/egIm2TEx0R5AwIySBcB1Yh+hZa/JQtFafEX2b4O
8H1fP+AXLPx3EgED8wzqeLpEufmUMy3IuMRyRnhyIyA5DWRqa6Y7/Vsb8cqhhMee
PgZfWF5zHoB0QmNku0KQrhxL+Gld7w5HIVvwLy2os3CoKAphsDmlKhWEbJWSFC7W
vEfw7Lzk00TeEl8T/THaApEHEphFd/hhI0Hrcf9eUwvM+m4W7ygPVQs5sSq8AcP4
vGRmSoExhzt0egf+eRcwgjuoI55xI5QHTQJMcKUUtXcy6grM8B9NN7r5c/VNIYW8
NlCf+2I/CC98Nvl1VqvVJqhkORenyRQQPfmVnIzBMDtkkb6txIY7nXEIygxvexD5
hHNM1Z4iUoHI/f+qCXtLJV+6hnHzvulNfEY/BwwAt0PguMArJF6qSGoDKuNCXHy+
gPTb4oMqQIxAOMNpapm7ZlBnQenudvFbqvWz52wUZWzo/vXxxsKFlKAVFXBHpmvH
/Z3M7OMobcyv31j9fxBnf8J5Z/sYHAO17wY+y4LXdVD9213iIWZmRF+RuOvcJf6b
AQaY7I9fowjvL13/paWt4h4DCsM2doIC0v0OZhpZZeUH3C53AKZIhMCX4gLz/5Zr
ZVMUTJMWIDIcjecEkkdFonVqaAQAsWyAAsEpWQkh7xGTkyuxmJ+/jyHwuOyeRR2j
r7L5IzsbyMN9C7j3YmONE/qeKWv0ychydrFHLI/RRCYzI0mDOS7bRrSliZ6MLI8+
pVMYFNhEKHBq31BAHnrs/7zRE6tlm3byErpidxyYL8zJm2nmKz4v/VRMifwB/jyY
NQuS6cASonXVDeWGu+3lN4t+bChHTuVQOGvDelKfXLbWejk2mtJyoOhQ5a2caEYk
kyX8BwUYTL7ug6Zgi3VaQEziGl74r4ewgAmKmaLEVqFAeckMglbWkqFlNuXrGBce
8Gt7l7s/fjlRGGafqzR06P2vgoIdsBhcTpxIPVumhwEKMmQtcIg4JE5SXfeQ6zGL
BD/CNHdyIdcI5Xe0WmV2+npkbNgXSGhxVypl7w4KSiAHh0WheSbN/2J8EM/hFHVL
beXxLerYOG9SGgDT0SLoYggiPHx1xrb+2a3xre8VFdnLlcQTOPtRop4+XAulU2Ut
Qe9Vuny0OhgJfl3+/RNAzdz8qeQFqTHtD7PrfTzkg95pPg+QuihOzKfuBkyuTBfF
2zw5meOHoQ8/nlzrqTWAgSB/OyNAbKpgpYdXorCHnN6AS97u0c90THizV3bfUrLc
qn7H8pxbE+qpg6ggU40jEr2nZadpU0n18suIXhXYPnkf7yZ5dzo59twHSYlAvXMR
WokTnVpNAh1lQvFnT1YO9h751pLRmb7qtOTr8N+RSpkk6ujQthWsi1z3CiQSqBCk
jZP+snd97qDpfE/fhcVeaOFCnjaxTdctvM1PxDbCDL/CxRKHFB6+hTrSeDZw7WR9
HJr9NYZUCwnpVWBmWG1DUBNtvaX5i09oAOF4eod8vsAK9IVSxo49Vl8wLJlgmWhP
BUjcPHchHq4K4sC+71e6BEN9Dy1IuY7J3BoXfHxjYOYNSAmwx0tXD/d26vOLxcaE
zKfdSZVvU7OntyOrGGTovRRp5F6TMudY3eZA1MPJ+quqlxW8lkxSZIq8imE8u6gu
pt3ZXKJz2IazSX2LHs5Pv8uab+o9j5uNRR59rMP0eD0vPVrR3gcsPFR2J3CsPI1O
jk2tyoj69R0lLq4WRS7hPFv0+FM4vhlzmfMbYsCFAulGrHAsNfXmuBN0VED9reJt
WuORDCRNzc7En/AwKaYd/jzSDCa/3WaXP+A+Vl5SAqu6+UzNKDXb9JmI2U+VLNXA
MswvceP1WVFb3Y72t5npIUm0xbz8hWTe37uPgjQeFgbWOh3ux36xqDOdiWg4XYju
oaClLMRPXdXjukHll5QIqbXhfkai8flFKylj1WhGu1swnqGb4Jb2yJYqulKp1eSF
4Ka9ZhiEClw4MUfmUJjznNokfBl/Eu3lXDVQRax2x2AdTQ39go+57nr90LZ9GLBH
joWjvH7yVcTrHxZKcLBX0J3e2X4GSON1TJS8T3YHYPorYq+zR5VVIPvrUSckF2FE
Hy0iwWGCNqH0HKYtCeHP5jqbRGJQ1EZEHfFUCYfUWolKbNHneOzNrYLT4bgY05kK
zfL6+48xpLUrCYHfMu/NCQt8nKhgpWi+TR8IgISYXUNiGZ19nzRa0uE7KSybwqz1
+YpCcjc9mBdZuq/qAy7VuyonPF1+GIvjt9Rz0s6pe0bY5sVrCfZQVdUjGhwLk9AK
d7Ag/7MlPZRRWcwurWSWQcEnh00kpd5Efw/79xEFFjoiypj5FLVNwbupesEtHbl3
mdQwR70GSv/rs3BxsZs14gZx1x8+7wmUyamnXx3k8biv9q1JJOYaOyRhQxBy542e
9KwCtiFRXOE5QHM0lb3+q1vW0fevaKRFNIJ/iqN6jeoyCCUNbVRHClPnjo269dKk
tiYJP1vjfKOzyz5moDRdgKZITuj74zhKCx0oibISesPFtGSRhAB/sJl7PwOgDFDm
iQeG40kyvzTcjncOuQsd/Dg8Al1GWQmP1BsocKX21BJ/1+s71QLTV5vgHXq5mn5y
T+WPeoFv4WgtKb+2PUhNNy3U9sKloQ1KHIJYm5UFoSXJqh6Aymg72/TV2kV0QdF1
nyIe23Cps4HoKRst0uqBjbFyaQAeirhUgp14c7LwjYCkNuObJDrtfl3pR8QHvuNx
bxheTwbiFm2aWADmptTN/oGatQNvjizzdB7940Auvcn4NDaOZb7p5f1kjvlpd6yW
VQCoxHakl6jWIauBXqRM1+fU1jNzzoujq3ok2N//YBTy3elkRNNahvHQmitStGoB
mhj0HfydjH8SKwgUOQdTDLGxUds06QfADYMt60OXMTO7cAJeoC1KRiGe58o2mFjx
NF5ballZhvhjInnZpP8se1SAHCGeHD/F0S3FuMEKEzlB//OPoPu0bnHSE9Vpw+FD
CXYiktaTMHmW+u0XmP/D+0ttcmS4BcVPWhyhEwhmPzIxTM6DIf2SZ9LeiB+pQwXX
gZ9w28eeghbag9x8Q7ieqoFG2MLCvKpenGu6pupBA21U+GezCxPkvcOIoLtEWifI
K+2klVgk8vxVpLkv+lKt9sIzvkTxBAXeBM+Xq5oWx+Hz37v0S9Wh5gCXr5/uVMEG
bkeQ4FQsoIitmbKMTOL39UseGAVrDubh7DBH68ok5mSiyMWHtEBZomvWHmbmW2JH
nM8XQfWDkLRjBwwRoqu8f8xoqcs5+tHfOUKKjI9vfSzUjrC7aRFN82sHrQ7mdkMU
eb3r0bQSBJemjSf7pTt1iW9sSgOrNYontOWz2IbQmAkWbx22gHrGdAYh2oE5TqlF
brzK6CKd7ucFMHHh75btZjXuMzwFsYjFaelFzGDzJ+T0UUUZDFLp0Ag+zrVwdJDW
dbNUT0iHvl5GN+KgkDQhcaFR5CT/dVnmkyhHaXwpGXdwhKXSKLxLfR6ZHamt3LDj
49N94LVNwhOejESWahc7Drp/Bmr2u9Gl7IKRI8Xu3KxcMdmrnGY8WKhogc4O30l1
EUrhGR13NTxjIO2oPjidSFuVTAiKd+cLTyVr6a9mQw8ZkBiH5nGr/+AudSkjtjvc
KndUvTCiWZhEnb5+NNA+PZMeoM/1JusAX5ebPYsduXwCbcY/ybkJgmhJ5YlJ/d7q
kt5A+MuqzvldXrybDQDqngELOHhGueiNIJ1wyiTUXxqvSDWbQcMHy8CYhVXRy/l3
CKvnMuPfbmUlTHnfhwl4Vt3Ak2GcLIvXPwYQxR6gZx5AwXJL+fe6NaaUlqRfdj2i
5TtaZpumA8fswSXJM87ZePa763/EhO55i8A0GKrRA15eG2+EzwLNr+32+1Myawzn
g6SN4tpE9kT0q9V4/Zj1AIIWeE6cxfVX++Vfde3ldHJ39PHQdcHCgKlhl5wDxju/
yfmYL8u4k7PKLWkFRxbUv0ljS0Pox60NdBaGU7fmnt6aSgEJ05bXEYWAKy9eRWIJ
NgDFjZm8kBbFquiXPyzIDF1OJvdrN2ct63lH3TscmMdS5usYZDz1XbOmSystWgW0
MOUnzLCEFglRSEWlDlQ7+Dz7Bo+/PquM6vC+xgVTWXiP4uqa1WPWe3MAjVDmQv+S
R8vDJPZ2hU6ZGoWSLt0NOE2zMKJvHJZFpY5xWnCJF+EczIeMtZ1r/OkokxDNY3vg
0d6kQaNX69Xun6fqGmIajgFzmXmF738Zop45TGrIPB4F/HUxz+aFbUXfNsyN+b+o
q5t8KSYNkaRtakidDnd32ULS3V9zmj00xafepfn8q9I09qpGKisi4A/VhC6+7TId
anQjsMBu6J7c5Q5RaLH50QsS95Bv3CoIYzA/eqMWWzj0qNfdJp5WZujzUxikrt4t
g0aip8VrolcLqGcREmXdoJXaumGP0Mt9V9w1a+BPkLwW1q75LL74PxdPHgg22Jo9
sr0TQItw8OmAbKccXGzssCjwkk2DddvyRCxS2XAqn25eK+Qmsa8W7ZzmPl9Veuo1
xPcsaX/zp6oTUHmjmGisA34LvWUFSR9gyBu+GqZc6bmln/zJJ9DMgig2hftC3BR7
z7PcI6fm6hWNEUxSniAGqWRfCGaqQkenT+oI+s98piva4ERno8sOQdpRqa7hehUp
uElZeFHxDtnBKU2Ht2ZqYO/HqL1Y7dRW5RxHIpq3/Hp1hqEZhjfkUbQCcQz3Kz/q
CaY234Ko7GgTvG1ZhaRIEkCBc5VxlSawj4PlnU2BZDzr6YGvtMv0VgmIbG6PaJnE
V2/5FBa26kpnN2WX1bDXxsbBMPbbfe5RaoZtmzw3fwIUXc44vBnDKFczOiCClx+d
c804IV5kOciAknWza4LhdCS67IOSkMMwU7HZjiR5vky/swUWZKeANOVQ+WdI1rel
4hdy1ak+0vianA6UTW41FEmcbMHSyRdq3CF7IpMb+Zrz6P6OcbRs+uiTz6x8XHOP
80itcGrwlwCyDeQbJALtwySgQT8SmXbABUS1cI6LSX0w3yiLCv4GIlQt2+aBzHCz
wOfpK2bWFGBQX+ewQdGT45A7yvjG9YX8UqQY6pjwgxQOEO8mupwprSf7IUizRNp+
mnvNuicOap5j5WqSJY+/tJN3A/UHRE9mBVeWGWP4kHv4JuZxmSYE2M+QTx/nInKg
YKHAYOxir5DfI6xSjXUvsEDS9a+7YM39mupqVLmTeFWMt2ObkovJLmbb0xs8czMW
nHuq3Q0d6Vv5k9sSVEQFKJgI8noaoLBz2Xp356mWiy+ZwE38EJEUGyuA7Eg+gnCZ
Qq40gMZ90B4UV9aQbHnV02TFOlxLjrHecOt0mq24OzvLbSd+aC8LiNFfvqIl7ZeQ
6+zEEnuMCAZ7hPFLuPg/PHXGMFwF02545Yent2rCXrZug0RihZnLnsJezhY6AG/u
wZmDAThgl18lelGRjvpG/3OYZb/mpqLKDFvQqGz7F3SDpVAMVGAPehiWSBZsuN5l
R+FWf0yUVvzmerWl4Et1zCQO166BnGSIbrib/ITbVeqve4vAWgRrV7T2emPDoe5J
QgLuzx1mpb03SiveDXXYro7V4zQJlT9FtIPlNF5mHtukBbCfpkc5J8cmpWXR01kw
5FtVMZSVry0IIiOnyEoPHN1qemBLAiV2RTLHU/DGSV6sGwwKSvbzm2PzBne11cDh
iNzPE+WScXOuf31mB5rz9Q3o1vA7JBHN84AtH2Ihvxu807V3bELyQJeg9EhL+PhY
Hi9dteBzdA/XF7d2+mdxP9yzNTBP1YyCFg2IP1DoRSnVNri5WGe0W+yiDObTWZWA
fOLgw0T06lz5ODkpKJNCWtKDvbZD/o+S4guUzJ0ApQRzsl1pvg8STDMxdOgB2gXd
0Q7rii2co6U18d7nDIHiuTGjuI+hbN+SI+cxBu3jbNzCDaEFM4PACjcb7xWAkibU
CjJsFNb7Ar1fW7u1bJZVRiz8/RwlVieQ5fzuZSoqgjku5WkvHo7M3/W0QEEuyGMU
JdCD4yFn62uDSS8qDHnKJUQ/fWhvCWI0xfuJMjmO3qXKn1QoSnyuj6u6R8r4H7LI
yo7HdSbcpahvAQ+8SaEe9uoEEkr/v5QnlBNVQdk94duvGuRUhSzON+RAD9heqUnr
5VlEdVJ/6xq9YtLlGaY4Vj7WxdpkG5cqKdayySneKtZ5cfBnwldZJQrecCWCe62F
X/8+Z4jEywt5O2FLSW1tEl6qsoLfg4JnOuOGgKzYr45Rv2+xQVBl2j91fQaGQYdA
MM9epJ3g9rDQpgIeQcVvRe4nZp2zXzZdIALiB/Quyyn5XR8fsnFiSdVo9tS+MSau
XV8fUvGckGQB/kyYiKY8YGFNyToJrL9STPTUz9v1z7rXMpohSo6/NGaS4jiL4Msl
CzKSxQoA9rsAA6QgSwr6/r3TYWO7zIhdHRPboRpGzUQet7BdGLQU6fQSZ3BLv0FT
6x46DIZr7MwqTGXaoZmBkx+mSCLP1wJiIHWqjZce3k4cgaThhJ+/Omg2dcBVPFFD
ms18sd4/yqbE8MxdnR5w2mHBsUyPTda/s3i7Xnix1C3lXfxYHMz5mI+o3Yr9Eaxt
l0utBwFHgNrAoNobo7b1kLPzbA03PHKGdE1uZR7ZsKygcZQtsCgPIH6uHtDNM02a
AeeZ/Vvfvwqq47FI9PMv27N/YrAuXooQmxUNkrsvpyYjUvwEgr8+roFKMLGzGZd5
4rtuDKElVLyxewPtlWVjO7RaH4bdoX4b1gWsqD5yB/n5ss4k4AQ4h9LeZxZRTmHy
JgFfSyj8PYGTh8KbaTJlaQTpo5+jfwbtdVpaYt+fLkD0UVOrk/DGiJWtTHurQ4Qw
na+VItbhKBJ3BN13fzjSHVBUn1F/5zVLyQr+ntZZ1IkKbL8l9/lIP8tqvSDGz/Sj
mUS6w+Bpm7r9PV1Cz/LXUtJh14Qoott91RiAqoD4lOEufit/hYP7B7152tu0J4eB
RF/EzVG67+QyvNyPPqF5S6sfw4pVKbWAJaxyikuRBJNooXb2UHBnlS7DlyfN68Rt
EbnHbgfYi7mwSDiDRiTkCUq/HBJqIEpaKj6vWR1xjI9WSsP4uTAAcKINY1e4om0b
n9iQN8+qwqfraivDVeG2dnCpkKiP+mJ3KUNMrUe4cswbadMbxhMWDs9k7MU2GAuF
ePrxPdgth+uBfO9aEO2feraNIWqSYPPb/rvKnEDqvdQ8SGLITcznkLRkv6+5u6Jf
TS8bpVzi1hZvAsbpts8AcaiHCNfyhl0kG2Y0YJnDuwF5U/4sIuFD3xCZGbCV9F//
5Aiq9yZ03sb9/heAB9y/RiGTcs2e0A4xop9GGGbOaGB5NsasWTqhCDW5yAUMAvui
12yncAlomV8crjkzIcyXFSYnRPyYi+d6x1F//kjfDqLqHsYC0j1VVUYy8fJy74pa
RPnOsgJ0SChtdm9X25KzLTCRQ8mZu4XPVhk3dRpodn3ienSGWvEp9RaCEY4SXiCQ
zzB4+Dx8Crl+54Mnnrhbe/s8N6Xn5HbaJzaRCo/mM8YSHzDd9ozTZv998pSd+fbu
JIsENQgrHxK0pgon5Awqc8AI3Nr1Yr2CbOlzKfqUluexfF119z88ByKPXz03TKas
rA50dIVH7kIsmEcvG8kfgPEk5NBHN/PExNNHkFpZPSw3mtVYQIITUneBwC+ZWm4A
sgQCGa24K+fG0j2cqmtka6q5c3mgKdZhWlmTyr05moPzwgfmc4TpBut/MsrJf/F3
/Wc8ETKXsJ4hMT+5yeT3o+URRkmRxVlmjlGqs68ihGvniY4HXgu70eLZ0OL2X+lh
c8NMHTe8vK4FvKao2Yocm9orOJFDcxi6GJwarKDJ768BrNsM846e9G+y21+2SQkT
toKxYFyjwN1FhiQqEFr1rDeAdGYJIbOx2daHX9M3Je9990n5ZWjktW7x23XZ8rFB
vRR4n2IdzsnFhwXiFCIZkbykVBr0C35ltNot+fuhaOBlmDI81Mo8WB0RFPv4qgnQ
/ujTzcV+D9hvYi/cbL3Z8eufWTCoSQAhri2zdNrOcuE/XIkLXimsPUL+ir8mcpGc
79JN8P4ONEBQ797obGWZBnCUYWxOe7iZaVQm7KW6Giph/Pg5Gj8JLg1Va0EFZAcX
1opNjUaEOwjYR+jcgtTYn+1iRii8+rShd0eux0fXbB4NVzjjDQl5A58K93EJjS5t
xZDhdY6p9tes13iuOdzJS2c4+AAzTqnjjrymJTSvCr9MrYCN9QErnDNdwNyUfhRM
CMWFYhxq/RguJ9fxouQLi3wagv/VUMBaj33aeHIS3SIxNIX53dizrE48NlWY60/W
tc/pMA9bNa/RO5EOyUpSqjQUy2s3R35loJpsG2n7u+Xpx6wGCvkEm3JYPo+Vfm+O
/kF94CbN8l8cL0o26AKtbD//1xNsQFYg0eN6cCcrWMQOb1rVIJm6FzWy1y/QTOSs
SpVNHtKCvY3LKMyBB/shBpw8SU5hfUgvxtfS/zQ94CFcu7F3vpoa9izOr1t4eHsN
GdXeb7lDopu019cyuKR6jJqBZaxMKdpsJIsfxDte6XB4XOkPzfg+cPdbQSvYDrbB
fGj19TWmJrzXJ2vUlkNFNaWspmB44YDFbD0CF0CtIQ15TeSlHU95HFmRWnZLbSCW
p1oU1+75/fJdd60mjllvxj2G3lrwtoY1r6uCoy/fWy7UNZ6pjJ1+pnSqVSuTf95o
uDeQ9kGstCes5EZDkVA8fj6EjmhWAQwGJxuDWOqkIJ8DUIrl0oDlc5K1GKolUWM/
xtfqjRV8hebGwGIh3K5VQ15asJNieTbHiFBHvddRZZoakUGSpTadbGiKAB74jCIm
YWTr9Jo5ssE8gEd9e3iYavFR01aqwPEl/v3XcJmIpm+w6r8VRR/TKxBGe1PxgM8G
6U3U3rzxVG8gXVwRLSMaLoxJGxrvpy3P22PlA4BqLmfBv22w+T3V8lc/hCCCrjD7
faDybxnPJ3X+Qa51FlItbtG+n7HfVmTQ18ODPB+tABiq1Hdqvq2ahp6ECWMSEAiv
D9nG8ariDi6u+qhWz3tbNwNgggzJ0Z9LiES0hua39TDIWc45xLEYBfJaBFN9zewt
RAGrQtSB2FrjVs4P4FTUReDQbQ0OCkUhDlYITqEuOVrNUY9Kg7IcjkhsZtpqGpeP
aBjrB79cETFDyoI2PQqlkYqQdDP0v5rR/0Kl8LW4r6kIV/gKHh5MVZ5f4WMpXhse
3m6zOI603a20zkV6FmAoBWNS4yUPL7v7jj1fdGPVn67QGwWIiV06xI1wc0jdg0OU
HcYyVBRfAZNX1/UBPboE8Xm/YqYCOhrsj/wkVcBH+bBof0K2WSXVm2seTnQ1hJoS
cDpWRZplnUmR2ebcVAnrdaQUpNeXiiTI912KKnT8nwbvVYxU6bQn26ZviO9d60kC
auXoJ/d5Sb6Mz+DujwUtuAwAMKdA0TDBC6FdRW3M7Z5ME9a7wP7lvyYDSo94ibpV
SUoHgrRrMGzeRYC3ek6AEfzoui1Z4t9mA1AIafkDBXMb3em3TbeDuxhbCOSc4Rnk
DyVPXMZpiAtkRi0NnFXul6A1fZh+ENjsBnSco9YeTEzZcC3bFAiAOrfPwDAWrW5I
hDoNl5ed2NQjoh1v9Qgqd7Bw7nMvv4c0dRaHb3KYPrD8EGNrDJDh5LgwZqa+X+Cp
ec1L3fku+Z4qV9pePtcEQ1dKBcRL3RuODeC1aHJh682ILtJ3CwMjts7J88sMvs97
Ke/U0DBL7+oRfTsT1nN4uizmINl9C7QtQ7Y2yJb8g62OGa5m29Vzmem+qHGbnVzF
TsLvV8RIsXK+xTEEW+yXot1BUam+qOOWb80PRCKNuKPLuZJRoHer8CgJsaq/UQ62
3JQMdzpIBt5yBQ1Z6P+RfpQIKv5x4sx9TeLgXKhKITUCG9WdBOKLhqd9Vm0QnMIK
tqksp3knjZXj/8reO5Xeoj7EZQHCiXCgc12NpRGENoTKDuBmfPWAp8yeloiUlhG9
nxg5fTVu0Js2AXoJFPzNeuA2jEM6wxz0b1W0009LnYHP/MBA3ecOMoTUEK1rYLts
NavjS9ajA5NQuMNv/VEfkw9OhPljveFWYdEYEb2T37aBscf1vBSszgGFtUnkqWtm
m3Bt0PtKcgbI11xGNdeBUhgq0OZJmj1aRfLXMZNnp2laysd5AXKyEByuOlUXf08L
LKPqGDQFRas9oUSI4r/Xx/EIINH2+YZmWKvPMd+L8XImElfHwzNDl4e/2qhWSCBE
p0k4q93/2FuDUoiBImFB9K/mRqgKUU/JjaBEykLJC6Oa9F28am9bADD/ddyx8I8L
Mt+ByP2UZnzgc1Iv4e+bdFxnyI6ipkBAAuF60w1CUpdUnh36i7GuuCBDCvb4RJmM
q54yZh3Zw0B5jnh4aecfp4QSePzqHcrVRmJaocwEYFLpF8cGRm+rY6z9CpLEUnO/
EmfaRZpJowhgsiPePObqBoO9OIXUHhjfuugxUBuZa/kG4h5TC5w1tnVpRSYbLIBi
3VUk+T9nl5HQ53Y3QtIdJ9QhOfy5uC2Qoa8fwWsQlg93vK0Nwrelt2Ka9lv3243F
2Ef123NUenskBt7zjNJiZ/x2W8TwbasAowiGMCN0jcOSmhvTtJKQ9xwzzmXSWXdt
whursvNVsjYTLQxYi6YXQkOyZSFFlEYYLi6eBrKHdMFOmT1nUaxMEHj/v5PKSFhp
RGhuyVQlHLqpSQ7W6LCuzOjBsIbvzymx9x8sT1oyGMP2FWxZSlLaMfR6WVxBDF8D
ycTLP0zxw4OtFjxNqILbykrIQsccr/2jkRAX5e77JyOXk8gidH8aHrVTO3NSdhFO
nMbhFc4iD3Xo3qJfZ7N6Ndv+XhPY1Dpd3Q/ubqGi6UY7tDAdE/jTxTUWJk5UWyII
DOTcZvaNP2mNObuAAHItbz6A/2FwsTMh/HnQa5gn/eOzaB6SFot399Jfzh20tLrF
JNRIZ5Txd3DFka5yScF0vT53f3q/LThCwDhcone1sRLtqjsic/uVoItLQC4WsY2u
sZCSTD6fAyE28iZdcvMdz+C64MGZ4PD1ls6nIfD0iO6OYxx+p5NegKmvE9H0++BJ
/N299/iAkgQM2TYwllN1mLWyZxvvi5pNXDDARCDyA8TfvK2Kcv8akXR5sJ5jwxCU
yXrrCONuoxTBZ3mawC6bJtzuJTkSwYREoP7obutm2PqrTTWQTlRG8F9KJvMAhDCp
eiSKKiHqJVGewI0T3a3xn4rieTagbsZqD7jyJKyMhsJMOiyTxdyFsORW+u7QRlgr
puWLG0BZotIQSJPHa5hEsNL+qvRlLqBIp6dKjAHFEqnmGFWwGNOaDfaiy9mxZml9
i9brZk7c9AZloQLJQPuzkg/6Es7ee/nJPh4Dl9X95SkqnkV0MpnmJSEVo2Y4uHIS
NQbFStjCpEQ+qtYADv17fykK4n+rmfyWP4VuFVeGWirgiR5w9rlLjdJW30pNaGVq
uvhw1/XmLdbkJrpc66g2ddVzu/dbin+moM4pOOtBHPoc/o21uSAxIVJz3oWps3QY
ICZDZHVAqOx+ODgYTTw5E/Tfd9iXLoh1Px3PGIo+EdWVkWG/0DSjoVnZ1zR+op3x
oIjNB6OXTlK97ZGN/HhLcjgeNygJ+UkPA4+jsW3TtPzZ674wAuc0uTfGaCiCIR+x
duWRA3wJvvU+3tSoUKRuo9BqYbDWGjxmarYQ66qVz0bnVr78/xTIk4K/Yv5Y+m2K
fNBr8qsiT0jtd9h0YRuYbbhDMigrswBn8D+KUqbBOq+/ZqlA/0U60TEDKEqmvTe6
Q/tnh3nnMobuAJT1qtoWjFbzOcZE0sC8FVu+s388CXCswQ8zXr425D1wACHDvlK9
p994E9Ml2sX8oUbDivFtEqLvLDd4BowMNYxSLyOs28H6GMRVKyhJFZqdce7yOJwA
pZJCzFBGdA/wB+2KS09J4t3chJ7X8R0k5Bkh2e6UWikGTV36gvMOsNFO4PQazwv/
W+xEn+v/nI1XhsCIkEciybj6awR3Hl8i6jF2ZmE5AyfuNwcSnkB6TCgAD7WR+kXP
I/6ko7bG08wQygiXcHpGFqGHQK+ddcG74aaASH8xYXeuskDT05UpTAj+DypU1Yjy
JXtMzK/m1s7GP3whmPeGAaZTiUdEOXCSWKKeocVi/S4Vm/slxVOgB2tF9Sn8Pj00
SFEuk5jqrtAZFEhAreCboeXflU305Ic4pR5XlPZB1j7YdYzcF9qSeC/4eJeV8N2H
WFwCw93srzMxwdWKKcIBAER6bzROhbuXJ/NciOD7xRfyYKy7dcT/2KStC58nOIbs
mALYi62A6cPIPKujq7kwkfK1MKANuoYkv8FCcbVdCCGTfUCTsteZLR4Ut6ChwE8N
IdHX5uccTpgNTMFrfYT4AoNtkd6rX/uGeoMVYghK7oa28fCujBPl0k/jkCNFzCd8
A/snoX6BO0JA/L0TZVKVt4NLpPK/pf12CZZ+Wp3eDIuyIfZSkr0i/9Eyd4YjLj2J

//pragma protect end_data_block
//pragma protect digest_block
3m+E7FGIrg2MhhTtDZo2fmTdEgk=
//pragma protect end_digest_block
//pragma protect end_protected
