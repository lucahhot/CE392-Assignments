// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
bzCLD6cIy+ltmFoPIMK5AlOd2PnKSUKg/44E69+cTXqkxU9CoHJbBsiTIqPEciQo
nC+cvoa+pywY9rxLxG57k9zN1lilesd5DKr3CdfE84NrBEEwFrfXAwxU1zSQHEl1
Sy2DoJGXEdsn89aCVKiPg52kSdlFyiqKchDBMTojZp4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 22960 )
`pragma protect data_block
dpJn6HhBuEti3wK/c6dLaeNh4BF/trZUbnHqP4O3tZOpVKK2weCPzqYWQ2nXxEaI
1n5Yf260HnRB5fZz2bA22xKQDNBxkL/CWFf9gUdrz//DYZbj9A5ADc8lkhRE+fc8
1DIAVGTdxjb7U0zA/dvm51apN4/IGIgxNTD3nozmqF8iaIZImF/A5IM/FeSsQek4
ddhYDqK9eCZ057KDutcGytlr8XTGXbbqqaMhGc5yLOYKLwIeNuIGBd8+J7RiRb30
FDuWUCxVfkd0tW3Iyrv0LhynEkj+vpXPzdMzcg56CrEz4Im01JhD9NmGV1fYAnYu
J7feCHoBJDOP0CrMseFQmE6zJbovtKXeB7cBffmmpwaFhNiDPKdDSdzoIJUXEI9E
Cz6DD19Vg04qGQjtdbnPy26SAQaYPJEEW+bB7z5bmE4PYjqgG3IcLwR94Xz8tHd0
VOS1yCjAs97Vix4OI+5Tad3g3m+cRHy1ZmWgj374JQm9e1WIjFb9FRYCxrhAngjl
CSMGF+IvPFXGWqj5rVUONqb7wKOhrkNLa3FlynWOphA++NYR5sqwOnYcSQa/cRGn
97M8xrw+n3nWFiDfj4KzgpGlrnNzbT658YViSFE57GTf/An2VlCLMu+FRvJGf5Wi
57hna8yElCNioBk+BVQPD1fXP4QCiEvfYs+aGDwMJDwxIKMTiA4wwmqYF9kusFrO
bSFglMQEHeyVjoT27cmYVQhm0bFTht+HX0ZY9fAeQMBMyxtdzjewObb5RLCmAlpM
Up6eL4RjUbkIrPBOsM1oAqRxyHKljRIwL2TqrJE92i1B18HX5VzYkuYDpVBOGgjj
FJmYFgWUuxQgipoVIenNFTB6PrXStBvKtvqeZ1o4vuDlGZH6X7AtZHXNJubegnMb
FaPFLOjKAS2c/oEqUWQIj2lxs2JDsLtPdG+6hClALSCsN6pJG/PjaJSi5y88Lhn1
ogOC1zq/sMW0pOIKksdBOQrr4d8kbkn4kWfK5IhdGEdOG2HwoNfr6Cj25uKdyCrS
yu+Rd6ETnm796W5E5BV8jpCoEiDOUbeai8pURXB4EV8JpmUCB1I7auF2ZEXTznle
gmoG5Xt5eYz1ahQVaEAAzelB1t+rrCQ1FIx/mjWSW9nVung4+QXLZJIEeCopeyYa
B4Koe+MRl82OlY8Iz5KH+r7BzN1R33QCTdz3ebbRF09QFubrlHU3Y0ugN3z195ex
OKZP6vnC4+/4wFOtfvhB7TGBI0UNcQpi2uGrBbn17ei7qDlhsfVzq30fWlLtepoI
rUy0k6IfG6yul/dmxVUN0UMN6Sj27aUcV2zYKmr0NtKrZKugXCRIXaDW3T//PzZN
DG39sPgXTpnJJ6/FKdJGrWAMUcEk5vyFXPrdoM5HLF/sXSue+65qHSiYPK8RvZtZ
e2oZXBfdO3TwrstQpD/VhLw0lnIyXuGahQtGp43qV1mjwOhZT9srmKq1BYSW4yNw
ejR3nqQYRw1dOxk7HmHxcR77aoUQgiT39ubfAs/aGLf/Vz2Smnp4pDIcK6uO5i98
VqL2Qh+NhDwkaz62r/+0t55yZXoH4STbj4NptMiyYtfbc/Nj392pa9AAWwh96zvB
h68wlNV3pTzl6Cm7Xxp4PWQUW62sT/DSU7nklwRmbEHQv4UXrFxD1gqzjikiWaJN
80xtbytoreHmN8qvSiU7QGcqDWrZHDn9anJ92miQM2dBhCXoFOATgAWmQs3EUy9E
5wZAA3+Gz742o9l7XSV7PEnm0Wb+7aFGPpRmHD3Kx93mvtCMvVH6Fl/haSH5z4TC
h3E3EyhWSuNPM7P5jrePVwfPO3uYiI8PfY5apUdcpy9ljPERMoG0vB88ZUx9ozH3
m8uj69rTb3d9M4dNFCIjFlDmlBQF8KsP6VKBfoQG1CZBMbRENklzwbnqgmCC8Abi
fy3NaVw9KZ3vnex08+259xl8mXFG7kv6gJfgz6CgbMQPDo3MoPIeLnZpP71iyLs7
DXqQqTNiSR1SGLEJ0CBidub94rP89/bd/2E9GwYa4v7OfPlS4+u2ppqaprxOz6Iw
uYuBRyBH3XK6RsGvX6+Ca/Do/WE+GCuuaDegPK70q49InPoTkV6ZDKGn1rz13YSe
eBebLY6VIr/oCwdiyi3DauO4iI7C5lFm5y3LZXwJub5QtMSvb+UA20889m4ZH7QL
o2aZMpKhDVaZa4QN6e9xLmsP9CVapONhCiGHVw//+XLcK4apGvRzL3I5cm9+n/Oy
wju8y1VnrLQuC1xDNEzKon2pxcxfuTVlkwGE/m/YV8JSa3dFAikiFxrqalwBKxrN
EvGj4bAYYTMq6bdOeKFS17z9f2N5EusN9xG2o0pXuwD8lvvVMM/Lcd8ug0nRTBTf
m9ZXByokz9dsM7SvuXVNAitB3b2OGV8PcuNb0Q0TrweCDd8yjZlAbCuXERp54n6t
Qry4CgNiRrrRNpSGYLklAcbdx6XObn6TUbAfY0n5USqytgK84xWjfXAAkwHtrczM
xxi/7H4PAozndH1k+4KqLkiUXzdpRVnNyLjZNCqUVq8eavBhFe6auXGfhFzm9B3D
K6vzYO4bOfP0A0ByDBN9PcNHexlwy5m5EFRe+PIuyLQldJVEJJWyOVP8gaholQ/B
wfVO6cZw4aF42cee0pFr4PDYFvGU2ry5y0SR7C7mh3Lv17nh1XiE7yN5CnOeaOdq
uEggURgLIXn4vtWo+LysSKoUEhI69xHxxzFZ/hLCPUt8Mmlxlei88xBG1Qhjzudv
OhvaNt4cWJMXN2HT/hHgCIDEb9LGjBTN430uxP1KL59fU0R4pZ4rIzOD3g9H9CRl
YEgQI7hfriHdCXrSeZyjkmTAR14lRWgF+OsrAEKCyU9LbO4UkZwhq6/qmH2hgWDx
kJ4GmHBiwaoZ9/Nm/gKt973xOHuDXOtl5u3sxrypt7PdViWtiX033t1HDoF1AkYn
n93FeiEGsp7K2QiVV51YSNfRHw1pVr48WU4cgwIkaqsnbZ0BFzLnnFLvU02eevO2
gTZxHrNDfrHFikdrhua+snq/SvgPZ/fcO/JjFCvgNOsxBpmQ2raBQRBph01ubV+6
rHIpFa6ptsR7bZ+wHFkKppz4tL1voy9IY1VRYlXDTdjwnekib6cxEq4KUuU8h1ZQ
8J3nmg1ESGxGtIuCauRJNsZU0ue4OXyHRIQLJ2NYLLulnap9funkpmhL4xCNWK/U
efh8sIwp+OUaNBGVFogEg8puH4nqPPQL/70oe9ij/dqkkqjuO9x9qMCwF9pF8O9Y
VLNPbteWaYehjPCr80tUtriw+CmxC7UMuS37VUOFnkDa28tfWV1uqaHlj6Iszhx4
ckTBOHisJfy3Pus5jbaASTePQuvlPvwzQPj4A2pMn0u7gxb4RRo230UwVbLo81Bu
tFViXFtTg1/lNpoTKtH7/3qE/HTQUBje9xXdUUHkVDuYB9mapOS2r9SWuXR9sumV
qN7W02Qeb5gFktuElKehOm+sVeNTAagbaDKZQYoSnnUvkclJzg/PPMi122iHOxll
csZYA+TgbNLI7t2b3K61l/OcqhQNFQPX6jFRO3GpxV0rQUuSxNoWAqyitfSVwhD/
9ZZ+zWSQCbS2bbniqiynpLcYwcR2T9HowydiQdbtebj0QjRiFWhR3S49eTljve3z
50iDMysIXEcb6XQxp0pu2N6bwG2occ78jYIIl5ySU+eqWWzhwRBxG0UcIxcWbJUz
bNxVHjEyV7VcwrKwMBn4cvqN8F09wpsqWgzJYYLE22bupHp854dymjUpy+OjcaDG
FOLyUGtMOsrf0MLCixFNIHGY9DixObgc0AqrLlPH5ViDLrGBYf75b5yP2Vl9bDqy
MC3ErfBqM5/weHywiPrYk/76bVGk2nlc9hGHHQZVcv2hdHus9Y3I9fcppJN+AalM
TkGctQvEUaKXTXNnuXuYpuEgJs/nqvYztHBwKZzpkls3EXEJrY+54fhFvIy9/6AA
2098RbPg5tNVw3mXEnZhh/mSJ3C1uikalcQ7a6LlaSnj3+//6C9NoipPEiqmbXFX
IZ/q7rnySPDByKc7RG/eIGzXCuPD5nrrZLz2sQwa1/7tNzKWbBL9HzNmN5iCXy13
/y8nsaiO9qmuy+vJzgj6RRj43lbYSjrag9NLNxm48aqm1MUyCEsn1bdyfr8BQfHg
za8Z0yQxabjAUxJct6FORJZ04T+t6lrbiOadYT0NsZ5XQIH+msfNGg6i7ITheMLw
KahTjwSjdzrzvQ3cjlPADN26N3p+mke+XxU72MoM5Zkrz5cSnqtKfrHKoj3G407s
g8Z7eAMPg4Bb5bwy3QceaNiC8VUSpNoQeR6eGCd1AfctI6Ov8RLRNh/mSxFOB95u
/m46GLu0e9TaKmV77QmtIAz9ne6E9/+6Pspqx5DjwcWBsSFnjqfgtnAkM+pcEp5F
BjvzsvlzsD/r9VLwX2eTW7D2KHhgm44tFYmWvv6Coap1AbF71Wujwuslt5acu1gn
OR3zzN6hMyqjo02zgXfFqNeaIE9Iwr2hECZ6JvNbUmzvZfI9f2Vi8Rol1KfW+s21
0TEppRKGI9qu4rxW5o9J9irvSPaqz0aLhfxDMJG6/RX3aTMZsVacB+bYqfF/2R6U
zz8+p6iecJMu6g7FaHJBFBD2bSiSkZgf6gde8hPSZoGtpjOWIuGXEAMVhDduejyC
Ta3E2T4o3b/Llw77qvZMinkVpQ2PVOCV1Fwr+yypXvkbvyFI+Z7w7nvht0kpM3VJ
4kb7jd9S0dMhwPD/AkXntUdjoNRiEXQ2cVigfAEjGXViKqlkZ+TVWhdI6CJWAnGO
j8Xx8Mk3MdZqfqi9EBsVqm6A7x74SHOBryzO8SsLJrlCARWt/NE/rCcRERI6V8Q7
EMvaKQXrboQeUx0dRlCdRDIqqruVXuK7d+i0SoYNCqUuvdJxx0KS1ot5nf+JsCi4
z+L+h6gaeZBH6p9fFh6+LqqHkygO4qtEoB1gaLlTS6u/Z2px1K5xCN2Wjc+bAJng
eWDFyfsbcq+v1wHygIMVuQjS9PuUb+ggDtCQfdl7UgvoXJEnjlYW/m28zOmWnCTs
PFUkMpiEIzPggYIyyKxPP8oQXtCDZFltN8RPfkj47xfLdtoufKtFh8KULhn0wNrC
A2lEG5te1lOp/SK2mK3x5+WZWv9gC09Q/1pY9UuSvRK1Fxis+1ONE95hfx/Qu9LX
+ALmH/w+TcXGhX34ZHCx4SGd87p8bS66Oo8wWs0g02T8CMJIuo8gcJs6QtrjyamZ
LdZFTWPBJFIYwxMOn3ZVHk09MRciG9THpB0w588MNbQ3v5YgsLyweGNZ3n8NlsAA
t1fn9TTkShMQ1RJJDkjafA/o19n5vXIMRGrvdlcTa0gHDrMZVmO1GE2dWJvSP+pf
vOu121eseLS8jd9xw2oR9YU7deA+iQjMQ4x6kbrbt6OvNXYSv8SdO7KxXvUAKkjG
nmuHQnZnWNkX5kXVUcSnLey94d9j1Z5s1EWGXBuO6L/B/bvDDW6C+rloCy3IThkA
rioT4aHorfDTqsNtfos2Uq9hIO6qd7Mrhw4PLf1pqdcC4CMCymYtFTSqj9dj/U/W
7hdu7q5sQBK0/9nxqg4IImIPEI+o44zbGqKiABEbeisplsaii0oKO0NVXKRHYDKF
dx3saWmYaB4c52PozDBxwIkIK6H1UKezSLUrPLnPTZbqyriAc6ERHaL3KhwotYM2
+gTv0WRbUpNCtAQzc75aLHrg3n8vvrkqbwgLWtKpU/5TNDGY36HDErjyp7HQqO98
mx7xF91l6onB8uxjQWBNOSidp7r0BWlHyh1OoMWDCjTujdDAD/UzxjtLZLFGHwBA
GMSoCvP4foNd45snMz1yYBFzWjeoOvMPIDpVXuv725F/QiEGE0ligCoOKab9GPkM
9MfiHxpNr/jnu+bNkrYjb51g5pyMa6oLY7Cce/eTRu2MR2fkIZITeCmH31Yc+6Ax
jYSSr8qmYbC3FsaBC32asACcVJ390HlmGp5hCTEZRqL+LonSYU/CEF4duQOQXQhU
ee4TORqZIBk9twnudIZqFx6VNjmfsAlwOHz5iHXCmXrnT0v3fwe2Gl9Mu4uT8A6E
/nGxEb4dhTnuSC98y6Njy0pN5BJX8TyVfg0GOOKUqzN/tHltcjVv1n4Pxr0GD4h4
C1IHZfCWwMR+VbdBtdphIjGLV/rJe0UqELnLtTz4VTEv71fPD+L2LAvPHya5ZAhE
tE8NIxbr2jY1lKY7jqScBjxc3xCYR8Ajy9nVcN7b2sb750Mr18lJRCTqi0QH3/ia
mmB6c16oi/UhegfHgNhVnsvXRzO+YIwwoHA49efW9CXeMw6jgkdrR35SeKbFHrLf
sFq1Xxr7kmbLrVZdaacyOeoEWYM+5CSuu5k5YQrRlcyj0OC2Oe5e4WjDUyGzZ+C/
dLHPhypUN+xG18PjNjDnefTYOJUJpVoHVbB/IInjWMtlaUoi1Lr7S8sPCWZqAuCm
HFT/Sxhl3XocF66qZO2BHCiiSFMldue6VBJGpak8Wph0rmbD9l6VOrFVIVldsRdk
MpZN3FocapuQsro/S0DJkwCQHJEdOViRlfoV183J6vIqLSS+i2dvj01sPsB6jKWq
/GE9JncO+SNfs4ut/7PVG8a2qHbXGOpjHdr76yyiXkL1ArW2BuUrwMYrkNagvbVf
Xx+x8HhpQwpvR4Mbz3f/nhb7CZ0PrqS6zoBDNFvztssBn/hAEi+/w19bj1RQDUUm
yGj46BJU/McRo2s3/xtIVN1JdZOXlBYOzkfjlF7Ya0gdtwnWhxNrW/wEIZNcglrQ
zoDx/rafpuypxVwkC3vd+TgQiq4FhAQYr0+e3Ex3+SswSlV753jthax+4wWH2KPE
0C7MkkO3MPBG6/uT8LnRcuDHzHwelUbB2pcH1Pl2Rc6qfZrEb6NTu9EVfnHoJRat
nn0WGM04uS8J7KuJaiWHQKsyaup9J28gVG/7aoEmJxH/pNrzUPUcXxtxl43nRKvQ
5lcMtzwPCZljewQ1rv4K6d026FZpcgONONPqE6LTyxFfs909m1kRdZ5qkLD+DlOU
K5KAvk/F30RSyoYr41JS0GZJ/sfifORe3+ze4asJ5BvJvBtoNvpS/wooJWSErjGz
oU8TJyFppN85nTqH66FHd3PG1gwsncRq2exck85GTU0QOxQTHGl0sWgVsOe/WUTC
G89ww38xwcjnm2hRHRaSI72lM+MSLCRoCVtNqHr2Hzhm7BwwXRzepkqzoo4WatIy
nppOQ4EyhOzJ5kQkECqtDIYh/SdsFdi8d9crGjyGMfUksPKub2uDs+AwfAmfoUlN
fXFQUKfsmrpkav0Md9tVXxRpBTCjTAcRWPFgQl224VW/REz7+W9ftUBrJekJ6WuK
4xMrXTtoogCC3U9toSEGbGvmy2gOmuNKehUWTcTLp5RSA8FanGv9wt12shPduxXu
e6RfVRm6fZh0Q5m7uNYc3thTUZbWgfoZAZvEHRs/FpPqcaiN9cyFFV7lDfNveVhY
oX7FPKw5W9dnuHOKXPmDyTO8zkuy2cpF5U/lS7+ydK9wcAH8bcbd7QiQkIIGvlDM
AHgIicqVLpd57gU6pnI9UxC4409iHBz4bcbgYed8Ahzl6WQ+J5q7Lg93rKfIOU+3
LRyyT2ohZH5QgtBbUNdkaEujWM7H214+7JRTGFr3yP9ktQSPit0aiMfEPKy6eScu
LYAspqFuMcSP9xgQe6x4usmli3MNqzu8cekZpjDhfLYtKOpCMSwiUyeDAj0B0pBc
TkokcWeFal7Ikt/xgOEKcLbARu5okSBauyhDb9EHB3x46o/a7AWKk3vjXUJeDudW
kNY4kui5abhwLE3K0fDbMjKBrnuWY1JGLppvqL3h1uDGoPzK8cNpBXJN+d3+xPU/
8XWKSP/NR3Knlpu6F784Vbsc6qzyejfoeB+mi0823v8w/wYJnwiPmXMgCENE1MNL
D1u822Xrf26kuIpA+NIWkVjL0XhCshje93tL/MSSI6wWLlj+78HyAQwqr7CbgHZZ
GbCGiZc29MXLJvCEGpRg+JrKZT+ShErB5XKbtJlzFq/xOpeBFpwvg1oDM20g8NqY
4Fqhvo+muhQ/QeZAg2pX+RNbBwk+bImXjAnOqpDFLqVv4LeVDPsYljI2YsKMPjbQ
HyJ/+wWGRfLJiYvVA+TSgAICgTuDySsre7RTkokB5punkq/8ybaFKuE05eHppKOP
/9v/GdL4nyH0/9Q4+Ls6SL3wr3xct41l9mJQbdmwHzsQ5cEIvxHhP35p4gZzTnGu
QabZ4nNbICtEyhwA8kHctqxoJf2/8S6tIR7jglXwCAztutMSOE3KWCU9wdRr6dDq
Bu/zIT2BcvCgBYKOrEimg6bPPgNxbBLWHXwBVcm23oujxY9p7g0rHmZpZFVDyAXa
1EuZs1yTjkFgI+lfTFqTj32emBOMBNS65oRtEhftCNdOl+xn3N+44gKpKAaLxx/r
bF+K4S2CbPqYr5MXyLo0fED/BjFhg9Y1NqEl7QND3CnJOtvS+v/SL4hhDYhFbzbV
j3hi7ul+8MInu3/zZW90YgWO+KykUouY/l/HeqK099Zw90eP04vFQ3/0juZIwoJz
HncNj2eIz553M/Ru/X55FzLRHR9Dx2ossTwcaEavdsidTQa57b195aKLI/UKkfF6
KTqWZe/UuxkG8p+tmYQHMIts+GE1s0vqqJqDSDnGv5PccVFGWx01gCP9dCvalN4p
siRdCALkFmg4v8g7jLA5llnKNqGrrjwBrie+9Wv4JpyEXRtySyQ1QxuhGmREkhLK
lFP6JMazxdAlAl5ahfJDAGb8Z3AFyCHV6egEnrWOmAc6vEtrmr63+wXgI4C8SSRC
hidyXk3FHk2uOkJQhFJD/S9j7/Y9RDvOeQ7bo2qZUS7uufQFvtW4PNnE2C7UZ/dc
I19OCQgSjK1WRPXtH11CC2xDzhoKlPVdqJDfqxSI0BQFpdWriCP2TMJj+ka8BskV
dv9PgNjhDp1bBxZiA3hb/88DL2pxBEUpatsnzLF3GZsajl25XIQ68ZXGm/QWcsi8
8u8btOn3a39wZoKs9ltBHEF7HRDhyPPuwlpMPoNWJ5P7wmNzjb4Vzdk5vC2UiSql
BVnB+i5YW6rjgoAhhzqnUMs/s7EUKrjBRd9f6p92z3vjpA0FdCeExvHoB7lIvSQH
Ih6ov1wM9rzjQJm63Os+9GK3hhuEpR2linevlZ0mTd4CS2vQ91K9To/muUQFLtSw
5IHAzXlGNC+FMuJcpSteG1jm3y75PsTXgDTskjoMcVIluT3AOTPcxqNWMeMulGEK
5mX/4UW/qSjxyDYK0f2LVvuitexwc/PFmoViSLxxAC1eCMTIMIMe5FLsjx3dz++w
lpHEmLlOQOnHItjLBTgS3JCSzMYLFKiRKvumbpdWm1D/pND65sEIN6MYnSS38XEp
fv4LzONC6rCqTDS64po7DFKEcwUY+XBTxqaOATy6dYA4WOseNwAyu3SKpZ/ZVHOI
fWRSz66mNtaz5y84FXwCWWWQNW+8VEcYha70BxEhPYISiOspB6rfeptFtCeLRHhZ
ZZKWTXrG2bGMWF2MOBGjCQ5ET34rBfn8i1ydlKjOV8ny0dVrgPIOYqt0LSrZj6a5
ODTq+PO0FvGxOUTmbaM/G1CkpzaRY1GeO0z30QSJbRG2si/ykMz2/2wu+Ms0iz53
lLH6proZimhkoKuWhweCvLa48PVFyVgIn7Pt03lOVIX2U82SAus7B4Ge09z8iSR0
3jFZZ1rG6DdhkbXdPGB5vYVHCI3xFmoljxkP0jAQ0eEhN5CnOwnY1yatjp1qZS+u
j+lD/MqEjGfCrX2KXqcV6kmb6/No7nn+zZ7J5N8VHjaunK7b42YRPhpMeFKBmIpy
zWJU6eEx1UwFig78j93ouuUFGL0sMH1+zYm7S/hkmFZrEidCvN1wXDwTEBsfOpTS
+6I7UfUaoXfHyoeykG1stTfV9zEpmUPyt1Dc+Bv65L+vpYcB/7vHYzsb43O1QWdJ
QUMoi2tIvxTxG00xwJ+dpUworzHEqtbhzXbQNXTGo4Ufdh8rjZdx8XGXZphgG0wS
xYwVrXviqSfcrzBZwLHs3yy0tfqhnffUsJhInLhx/SuT1ZF2USKLHnG+JZxhNBmP
oBXmvZFCTCcY2Jh6GAZz41P+bt4RCU75tz6m6PojikEsCY5sZ5FyQQBCx9eJfR4l
Ma3nGKtTzORd6ICBeJ5+/p7jYbt/HP/A8BmdxuzUt7Js9gKDykcKAEJsRQ7xqc3p
GxOFlQHvcd2pL1L2E0XbFnTn0eFUV3vJCvxglTYvDJwtFkGSyxsAEAWu3Pxi1q2g
Pbcjddd33r8DHJ9Aeo94/S7elJqTwMYGxdn50RGeEq3MyVTfyeSNy62/VmJPMyGw
TXp+tnkHE8IpdZEPd66k1E/ZbQI94LZTUeaj5/M75ZCzjNYUGVsxu9qdeORHGxEb
ugWyYcDYk2oBNFlMB2nDgoBx9wR/J/ySMccvhSMKrzBIvnoSsUwp3BKsOcoxvJde
0a38FthHE3KPogeDkxfmxeoBbWH6C5maq/S04INZ/it3YI05qzUmy6OQy3UbYCU/
By0wtd4s0Fa3yHvCE8rs2K9ifDV4Jc2oUHSCJO6o3wjd4LB7KCh7olUqoCmYMZPd
aNePgiZhITQ+tikkGpfL/EQlwVfi0ZppM84QSg8JKGVXRofPY9cdTMLqHeyc3E4a
lHc0Kl9udK7ukYZ1LtOBNVhRPNC9OpODj7CDuGiKYRPaNoRaTEFAmltFMyeXGuwF
mLKixt6otSj7m5xdI39MD8gIJqdYuolPYIcmIkOyeO3319Lshb4TZeeCc5BokwJH
6slsB2YqYi01WbqYFWOgXKf9Y/XIgJZSj+HakPNIuuASQZZqnEeKiMaDloDXK9Ml
Fc/sVc9bD49ZeBDh1sZJ9nK2StF6IwFO1AblmkBNFpHiNJJ063imQlJOGnqyJj5n
qMMBtZrVtdlIwcxkyQ/pyJMwTto00fhmjSfzJ4onXjUlxzVsueiotT4Veh7kPEi+
Uiq82o7rCgbuwpYfWl4I0+M5FFZeIKxVAm3ceKYYsRDuDhi9B37F82saZHEEmRfE
oei0bw2rKWafO2O5bXoAHGA2IV3QF7lyb+C5+TNrkW418h/otY6cUJDbGAA3HTnf
OJz+RmCSBMdO42sVNqEYYed+7Jd75RSA68ORlnPEE9gQz+J2ubxwmeHTH7j4LS6+
Pxe0ivwpKsson2OT6No31nVbw4xrz2JBb8ShxmxTDS2dFXTjsQ1RpTXGjCsH6tji
SFTknIlc8QR05qMar6GqSpteNrzOIovoTsRZLtaaE0HgI5zmmU6DR7r3o9Y6em8A
GD1hhMWKKIcCNx97ghh7G3B27ulIE1pahBL7aQBEQnHqSjzUWu9XK96foiMaEOlF
BsAaC4d0h3RYhDMlnGIxY4bW5AIid5tQO/fFn9GrtJBwZU7x22s+51licn+PVFQX
uUz8LiDUXW0aKsrMYSNEnnvIrCMwDtNKlhzrcIUcyV6HxLpFkER1MQvuKAyRascM
XVo1JbmLyi7PurR2jpm1zd9Y0g7CZVmnbmVYl0jHFtPqee+1EGjHyfmUeJCmM0Fn
8bxo866VKQzeD0DSr5eXjOT0m2hvxjLZXc7dT4aPHqD/y/chqPFO2lh5JtH+BOup
cpks/I1+oDci9LraqZ9cmLdLe+a4HgwWLDWiL2oSdv8MDl6vrrQTBoRJHqZTHwyj
fl8h0bbx3T0VGL07KyM/HlspEsy/h3xGaeGJHcinKCiBwjgB9N2YCCGbbrgVmFx5
zQ6qcvj6Lm9lzCoPIL2U+4tO97WxJepcEVeZn1VH4l9caqYjDV8tdwrHvgzjuKjl
Soo1BuQ7MNCrlKLlBl2JyFq/2AMi8YxSiKL5CgeBnXaT/U4P/Q3QdfkOi6Jbabdo
E8DSDO5PNjpuUh9hdqLwUt6tcCHWNhSa2OMFyUlbkL5d7J92ruHXG8bzMcK6rizL
d7xAz762jt0Lep6FnB2pc3GLDGQkXyI/cy+zTXm4QTOMC8X7TfhX9sZmDcxzsr1j
5Xg3Z9MIQa2kpGGm5mT5vfpNayjXU+L8sE22ZYRxIeXwtcxYvbUt27QNUyFu5Ysi
Ph7Y5/g2opgy1kQpamI4jRMTzvR0cWjdSZ0wUc9Lz5tTZm1ezwmGV85unzAuHENQ
qio3GiRTEugz1rDFPeGd5GW/s/ZZ4jBTFiH4kMzRasIFoOAT1puUxrrQxODyw6of
bHoYNaTp3j+oZNKw9DX8Ia4/oTh+G7sC/g/AoUGIu2DWMFo8I39L496AKjU8tppl
yBBMUen45HdUe8zTPx8GngYrIZVXDvrOOp1COpp1rno27aGavLMjBwXP5I1FeYPh
hOn83GJM9IVXlkX5GHmF+dJllop+nfxtT3zcbPCbcWtiDtFM8f9g8CiNVXiuwzjq
gSlDoLeJtt8xIO+Pu9XNOwxLiiFTIKMKy8Cwglp1ez20kGgESst/naZPitFrQqRW
Cr4BQI33iuJVGb/TXQXNPXBmjDgQ5LrfPpsgPWELtgczm6EZlBuYGpqALdWI0kr3
Ql7HXT93VmGbgJ2G4+ZMCE+//ZI7Py7czQjj/k4aizD+0WPkGOB98D4BoaZSMlld
gENfUX0yt5ScjI0fGRX09pDxmZyOM3V/R2FThXVbFX1GbJAOB0hza+zFPtYjygel
9hq+yv2qoIXAeY5HsmbfrVFlzBPHtTonM1hokVwclR88YJs3Dk198hFEwwBB9pja
j3jNCH6i/crb0H4cPJ7t42ltiwMDTWBy4OE/cSCm0q6v8Kidqbxuku2oXIBP1H9m
ff0/AibeBQ+/H/lS0o/SoQ/wd19+HqCtyxUTc0QqKAXd0hLCisyAvJtAgHQ92nqY
cFwbZnq7pZeyC615umikJABeD8jTHkQDrs65b7DRGEzKweb+nzIcqStpB4F46tq8
FrUeuVxgG2Un8Isgodd5r1yyaoZjRwprbXdoR0cTD+O6ywHciuOf2ts0foD9c9Sw
T8VaweuSjHLMv2tmcdLnGfDydjJvw9EfoltyuoWvrHtMSp7iRnpr3wri345CyB8W
jtg/omDwhbi9SAETfU9ON0+hYubBUEZptiu5sFf3fXY1zqLdG+xYVDIB+NuhCVlC
7pOWzn4AGg4BfRDSQ6XBfrursO2BOz5BF9e3RRa57LoIExykGLP8ua4rNwS6myye
WtnBi7GPJVlh8ePwdLUnXr3P3ZrCuja6qM8yWXEG/jjrCiq9293J/vTpnsI6/18P
Lpj3Y9vy1lxzzPSzC1ngMRZWFJKO8fr5dJFBXDZPIaWurh8TDo4RiOjjAZkgS4Pg
5HoTYVS3Vo8aPF7s/L92DEyxb0NJuYESPcTplbgPUfoB/QI7DMoNioPKRqwrWvQN
eiOGqNvtx4nhHiRnWcsKR/QBDNNJhI1PzKgoTuJUezitpUrIqVIw3L3LM5hPnWUg
Wxbfsd+PVyL6OQZ0L6cufB6UCtqvzkhsDuGES0PmDZ7xb1dAwEucRWeRiCnLxvhS
795vAMHjX+c/xUA3npORdIhDusqPb6+Ktq46UWSMcfOCdP6U2l7YWZspZGa8gh/a
tCtR3FptTerlXcb55kHXX4CiyzGfOzXkfnSW2IiV/mzQpwprKFoqG0KCAB1t8/bv
HscoISbnLwLRxOn2fz42e5y+yN7anHXZtW459nkkuTOha1PgH+Lj6G9ny2q0hnYY
pMtxhSbl++8PdwWv4kR4e6X7ZjBvO2nfuQojqae3c+PNq+5088IS2mZbU/vFuvjy
0JeCVdZh+C9JPq9E/hGCNoi31x1nZ9BuGVXN4dCAHcL9rgVVf9xTN+0g4cva5vg3
SyXlK07HVVt6TwPTfrBq99UHdxrGRkhdBZtSexu6nG2zRcjeCnNkC1E6nZKA/ZUZ
+rEsY5lJlckK2atYhW0+gAzpkYEEjqZ6RF+YPSDDh4uXGGT9sJdiA1ZH1IESXAlQ
ZhMCwWl2tQQGEVzfbNwHQIX/FRuMaq1eWOsiypCFWoHsbCWREZ26IS1+dZ69olz4
TJz6FC41l/O0Y10laVfspaS4/XRKtIw/8Qsx0yT7yw3K+c6H95SDNnZT+ctzHxzK
lgdBjDPtHvpyg+fD7336BveQuhgc6v6xQNmxM4t4uJviZvAkF4bNQirjhrD5wmC0
uFOvnzNFZVf7WRtXAwrlt0IcR0Q6azla9dyzf+Fy02jZkSeV8YXNreizqusJCDa2
lgiqftxvBUyRQ1etFWBNEvWsXtOwmsXb1mGq8w0GazcS5O655D0M5oUHycvAEsiD
4CgyTA1N/Uwha0TEOQ8YsEBh8B+20KEMLs+nsjd+FvBuLOPJxshwSdFY5YtaaPxe
DxpTqSJUBXViwEKSmhsYmK+Vdrio+VEkXizikGxFeZR8AbMYAMMu+2BfZfpN4Gtu
i5MmPhzgaCBh7pt8B27Td6jb//wvf+rJDQWcLBF5+XBhhvcFiabuiNHWrRhbQPtH
/IbyhrqM0gVfK+uIsxxbrQpKFGYz48gRyMP1SBtfN5JnEtqHuTJPABbLs+ym09Wm
4Q1Ixc3qOEnGubdsi8kVv6pYjl9ic8qwaH5ARsfVX2k/xO3ei0RdSnXynSS6CoE8
ESmV+M+iBaFtzG6Nr3lj9bdlkeFJ7s6iQ8lI3Ue+KB51seql/RETkB8YzxH1zhGn
xIvaUHQGjaE7XdZDywChTytjJTpT7D61cyyu0aSGe5HcHEb9udQf8h95R6yy+RZ9
rfgNye4VGATaWLycTkJIQ9l2jZL1C9lTR4VLKMPWZWlqob4p5mO8ExgZYp/rMsNN
aRaEtrtPDX6If7iqAAF15eQRr1N2bNzr6aZtsugv31ojuZODSVEx2hufXLKh33R6
weDPoh2ZHPYEQxcczmxFR4PX7hyXNLCFrzOWdTr9+Sq87AvyeHaJRkf80+QjOZbe
xIFbQHABTDhXiyPhrrTVRcPWVw4zLfzDvOGOlJFA7I+nfOCba78Bq19lDNiUUAHP
UeL5wkpEXeNBHLPposbCr+gEvGv1SNeMGR3h9DcObvJRCa7gmDrFsz6+KUxeuqbZ
2zvoxQOBX/sxicEIDTfPuAJJKLElFX3qkQU+OruNDKjJh47J6gGKn94tDKTfCtKo
TEpFGf7o9dYwsowtlviHJUUfPDOc1Jnlb7u9w8Wie9wZTyyFV2XwJCfQNyUTHU65
R7PSkkINQdhqyK2NNXkBA4uXC2wMadTdkNxaIii3f+B11O4cSIV0flf7HYjW0Cv1
9YzeCpgYw5reTJjw71bWt0ClRYsK6K2Xe8t/SAveZhrM4C0rtjnTFxrqYPcfT9xS
PakLdiHTKx7sf6SLmmiyxIXJ7HL7+XRY5RVJtVsPTD2+XP0doPN40R1QmhZ14JYR
oyQ86phNbT8IgSIZXTEG2zRrikjo4baD2xVjwz1Tgapt4GjZL/J2pjyC4qskmlKe
8ZMK7FnkLKz3uxUTKocynbzgQxgEzIJvgbkeV1xns7LVUNAVxMF0BEi8pyrP7yf3
Tlft0iRc9m1+htW/foRfc1DRI3see6/ZnS3OPJwyXQ3svURF5Fa8HhH6oNFXKm0m
Bx+uBF9YiwAthj5oAVuSH6EULN9/EZTk9yxWwZsYMDIPFmJFohvTD12/lNY/MG0b
A85fWQxvxDIpxiALLjS1cOI5p7GpYndKrjmd4ZO9qWDwP4ZVwdk3L+sZF1Swp+tF
PYwfONTlwI1Hzaqp5BK41cvoUgP1dlz9czYQKkN3p1amuirihuogbeZ8xSWT2wat
Z/2Q6C6+5BJF4fQGiEFY/eVcGbZ0xqX32hUzxZYoS0vm1A6nD2b/re1pkpZA1N85
030pJ9Murkg/XVfUfeoXpfyPaK/hazmjfi14XAa6GuCdQksvoZcPYJBLNTkvBhj/
JLRJtkOS9PhQPVXOQvWzgTZpTBexMsrfCWXim2zrth002sPOy3GnUUUuhSlEp13V
XQ8FS8o5+kNMRx1G6JLE7SpXh4HD9rgZX2RMJ/TnxgZd6eSNnNEMTCJsdIVcvomO
dzGoIOIgTvn1phEcRcXspVsSfXQE1iolIFyg9wjLasnTwm57jLhRzvale6qLPSdY
qoiIy3t4IWOKeWrY3HLdtSSPpW3GCAG8gPgfMjIE+N1PWfwqDE+Ou1PBjPbFV6ex
yrMWJxRPDfxb5Vutmg6GUORhzyECtBcdKV54JRPiNKfN4trnNI7MisDzR2zhaPgT
quE9ddo3xlH49D678/L0bXMMvU1kAZBRYlodToU7MjUNWkhmJZibE9OsNWT6LljJ
GJhPcYJ843zWIkbgSyU8Y3Ve/9kh+DHmhvWBYeM4pH3CNT4RltTZprxelk/arubP
qzCw30PoqY7pvhrX+Hzg1ZlS6OUsnoRr9XVCjFIUwqnNLwnVXDoM1Y2AJ6ulg2Mz
Zq9vjbks6KWX4gPQ6vkPIfCH1SaBJbTFv+b7RVJaYtI6UayEq9eB2ImkSyMlXyl5
LczA4TVhfRTJ1kCsYZp0le/GlI0KGroTXcQIF1s9+TNAmMi8YIufboue6dlPEIsG
AAAthPxwdRNGPwZZM+P5N6z4c9iyqB+ZauTedM1bMV3Unk+sEj+Cykq7rFpVpU9a
JEH2E+cpLwS5V/DSuEVBp8bqdzUn5UaHipE5Uf2W033x63nSAOca7SV2oU0gYm1n
eovzmwIXjRdtga+wQxNzb6YDaZkWr1DKBw/kBnFMIq3SJ96sG4/7oO0lXppIC43+
Bclb7+x99nScqC3In7FDhf07tAM1RQngit46fSj1HIjBJMMq7xvpcPPb17Wq5O+d
IG+zcjgIsCf9wTOGvF49pNG2BWQSawPYOh4nTfgw2Gl62oTZ5r85uXaSYDn7t+oE
/KTBWoHl3YMEr7rcalZF/ciTC5heAeS2b1LYWpQOLO2vCCERMaRiAc/iFFeXTsXo
RF4O2JvrpiCUSuXjiN+AE02+I1DP7AysLSPivgKJQM2VD5NbbfUUDuRKrqhrhVJ/
W1RI7rh8+E9lJz0c+JivfLNwZeYGIPk08/dfQwc9arACvBf4X+/qoxjSTCYxAH9q
Y0kMEhqGmFCmRM0MbBb3xWV9SveQ0UEUfhnWv9ixQI0wXZ7BGQr0jStXBtBaHKX7
e/Hwp6FEld6eIDtK9++HNXrmCBXh7ozyqjfk+S3Ac4XEt+9QCCBXrugwsRuqeNkv
fzW2SB1mYtTQCrBwhXX/WSsvfTfSX/BEz2q4XMfBgkxfONQQ5R2TTwt6hgQRg0ak
a5EBgfsU6i9E9gGtGaaaU5szhJcwPTI1og/h3bkH7FGvGoK5iLCF/Bfq6zoblmUP
oOtlrQib6Qjdr9xbs71CTNYyO6M/aXYWbnEJdd0fWfC49V4VPHXSpv4RZ9eZQiAN
2aRA4qy/XzU8b4VpRSe5FMGoMRONpg6u4YluyvTOHluPtqAUOvRVgFUvCyHFv7Nw
dqX79rO+jD1P9zKkQrv4cImQBMPYk/ninEkxKKy+Jj97C371MD3vRwPQkymBCPkY
/dJSZHctKpzh03DQaVAow70MydqWVMGDsOlU/WPWPO4bDqmemqqkoE2Y2tlD7uZ1
twfQU6uog8fWA1scVKeN3Eaza5kGQLF9zvZK6XYFv+cITn0aYCIegQxM3+PeAUzO
xxDr6bu/nL97jkHNQH9IbHfFPowb0U+BfxfGuQp21d5Cilj4gWrnYAiqsVZvzNWl
fBGXKZcxlur0yFDL0QRcY84sktscIeeKReKhXOIrYSn2cy/OygCvpJfstPQVx4T1
wx/bqUqqqqwgv/hGjF3YVVDKxtCX4E/eWxlN7m1/70WYKyujBkEWn4dySykeiyus
zttEb9GRd2XFZi4YANFT5JhQTptDhnqXc8NVskKAJ47Maav+DaAP7JNjhfvrsrHx
Qf19qptSF6mAUomatGLhhsTHlTALqye9A+cpDX+k81AuBKVy6BMla2k8I96k1Bgx
798Ivow178A6Yx/5dP5k2adk7F7bIXnM+Pm/faCpFqjfADcUmdksZPlG5YiysF1u
x+JKmT0xs/4xcUNbs7F9JJer9j8bVYcG/2EHxgwnszlwhXIqVZrD2E3TrF1c2lR2
gzuOtQTvlpLKYAgxgNDBoDB5IQofSKBs8sZVQsiOd2klpN9W/PGK4tOABLvKCYoh
0SMIh43/NJEmj+BbcaQ7YprtwloEuy3BGPFIsLVzU6+OLQkxZNBodC/SjlW0+P8Y
8mIfhyKl0dvFQ9k/3GVfQGvUJkQ2Mj8q5zyitzo5BILghPBVJLDBMSs0F47nqpsl
ftrGhxrky98Ocdff5nw6n+l9rdsht1DUHGEpM8dTlXgPLTqvRFywpOBvK4F4woim
XBHPEg7jiCnhftI6z4LWCX/JKtbMN4GYb1Dii+3Wru2IvOHSB0lenacc1TrI/ulg
EQsSs0gni/pj2myZVJQNIQJ2Hs0lQHS1VuX/rYC6SDoRHYDLToD9Hm7fF/iiKAmS
P6SNdnI6bxWPFSRn3/iVbYd6dY7TZQDO5irbtNovwPghvoIRhuTkxtYvEaW5AybI
M51YQQMMK3OSEZkKbKJZbOx1pRu2QwoQUvKPZuYJJW7jlhTeaSG2Cb4lqI6D/sRE
jKmousacuJ7xII+ZBy9BaPkciDxfT/f5QkTl27e5HOke7uU5Pa7PwTz3br73mX3U
rntev+vzg2cs5MQHAOVVacBO7Gy++TL6m+JN2DGpwKZVqbQluspmdFG1zCupJ1TC
Xlwy7ZOs/t0pdABk7tdxO+9eAhyEhnfsMVrv2Mj0HGyG2srfp5gAIBPT+YtYxVEN
85i+GxaftMHB4Fm8UV3+cm80kSVIKxL1Vo+Io/KK8GkTq5ZWQs3mP5IoRvP3WFI4
FppFto8RLIcPFH7i4Nd5IZY4+jSDxKf3Reut/46dYtiEXqVUF1GpeagFp+zsU4nS
B9x8Zs39CZGRyCDSJ9/PSy6d41DIbW37XMYfqYvmlnDoYJfdGOHNTFQS+llI3g6E
8ZUfMxxK6as9PNP2dutoID1dlTHVxTIX+BmiWhVlEpmFWTDzM/sql0+1CKwU2u/i
mmIGGkkhKs+alV6SOKyuGs9jGKBH7UROSZoCcyHol00OoxHCHsI6yTPmKhmzFv76
7Zo8bIWpXBfMvjPgMcai5fGw/4jTEN4TvLkxQYnMUCdp9DIhLrqb6uR9Tn0RS5fF
OF+wPGAzhmsJkvG8hNPYlF197dJP4+Jyw+4paSemgO4a7mzvDzbapPn+8STTOA1i
JTpUrvjrahQlWW5YBdG90GFvyGhbgWqsEF/7VYsHCKBweBeBMBKHJhT786bDKmth
NdBDa7/sIKoJ62vKyDX0TBXGd4/4rEXgduDmon00jmVlNoLCTGyTISGnFcZRHEDb
Ax/7Va45+IuLE+JSh/NqOejUSzpldWHA7acT9G8nnuyCvEFH2/Pehi4lhvuol92w
DcWY4TMKYn+TONX1HVQWTRoyXllsTxHw/NmOJz1cMFSGBI784pkoe1zrlbCMw1CP
e6CLtd6ksYipwa2rr08BAjjnvWyMR0/Peea5IL/8gDpux4EM94KLB6QkIN9A6jwe
huR0I2i8wtdFL3lEq+ZCuei/PsaSzVBAiUS31fchIwl7s0BwJgDTVSP/azZgPaCO
A+jBCVfGEQ3Q8S2/o3LGXuROYdt0H295FbCYIWpvYSB/8JZWkG3K3oyb4RUgPQlh
EiZQ89nuKKird5Dj50FrZgKRaS7MYSF9bRe2HjlG7gLr3ec88LPykF4J3fxHAJ68
FRhQ7uqvgAjMSlsidnb5zvVW+tWeGMZSHBIzRGjCFo/WV9PQwZ3dKqpUlsLhnKdg
/c3ukcCUPvZg6g3dYGBazQjhu4JwO2XNnaR7DQYeaj7WEqUxjuPTDPUb5bj3pXN7
Nyq6LLho1KiCmcQR2jF51O4XQYeLiEBrgf0Hf86JxGiBm81tb6uoPCy6gGbMTbi0
p4hIp8/mnCBXdP1zXy1AKe+YvL0auCb+zbC9slXsnes12XuKd/W+r8RhM6jM+m4h
rCsGM9sNojj/1H2ng6RaFHCXmeX8DejoVt0ML/3VDMXYXjPgN2v4yBOI66DJ9P1v
uZM+BfFyJBX9s4YTEnPJ3NCBhm+BY+EkNEK9cguoc7ILAJ6JxqNr4T2f28eLxyUX
6t+kXS6C1cSB4m+eYiWHygb8M3YWuGYxW7px7xnJWJAe2B1S0sXq+XWbet2GCN7k
u1kAFW8chZ1Z5fMgBZBX8K7mD4caZB8St/rSp9NkCaS/Lgd22mAR5Un70gii8aJj
PFTrZv1u2MBjW3b9maP27B4bqvfVYjEwkX+pWVZFIFaJXDLfcGq+F/AG+92wRU+4
oqDZScFjdcLT8MngoNppxtAIPk/WgL0dSKPLISLiMEInFbzFZPrf34ebsADqdQB9
TXiSGceW1/4L+gV9zr4/U/WlzBMhQORE0UOAukHan8QaV1pCrKzCSu8ebPYwNhH8
9vuyMcVY/hJN/1lGqy7cwWWAPqvpij9NYt69QrPYJGs9RkzWjFuEoNYI1KiaFGTy
Yd+4mRPo3DZpFqTGbSHQWBbcVOygQpuYjmz7OJxkNU3KTd0rZ/AjtQadWO9iAcvD
XCTu6BQnSiXj7F75iquDhlN0D+8kxLnOE0B1igSpJh8+KPkOjr/GsH1ohsRy0Vlr
raXTKqSdJ/Qhe5pBL2uXYAVd4mnF8dXr57VPVFPQ1kpwSIWkH3GS1lwJgOtbcNOW
ymFwTjhzOoMpiLPg4+HXabF2PFyz8oTUaq8hDT1SceEMVCI3rECLGNn64JIRwDpH
vanDZxe6QlW2pIDrFLoFZ5PKPJ3mQCuJOBpjHWmUJzDBw6DbvVGR+Vek20EQxA4N
vDy6/Ncl1ZtJu0fpFLrRQb1LXpQxnOIGTy/yYiysxqfFt+ieT7JTNhviuG3UQ5W4
VWw2NMgVaN7GDw26r8nr7L5H2y06ctn67SoUN0f0xdHlAB9kzP3R4yapZIUtWXqq
KTg5kAi1AKAQJSzgVjss4o7wPq+exscJIecfJH5CIgHo8DKa9d58mGVQaDIV7+lL
sYdTXUS019IO7LV+Pn/Yq4zZgJQ33JEjhx++/LtDgV8oRPlZMAT9GAuIV+BfFjLH
qBh+qzv1FzN+Ii8hHXfc7/FNpHvbsuMFy3IvgNbJDl53nF2b2fxGIxr95MoPtdg1
GLj9pPObjt2+bb1mP0A1jid09uUsgONQC46ZKvoy34Dr5hsj1+ycBr1CtnSUiEQ7
zhnRRpYSlWbRnSf5HWZiB2raAnovvXoMS00eXEDbNsEWPmnmTPq66NNKPZ/UPGh7
culhUvwsT8+DfPwmc+3c6rMAFBuh7tr0AVeeFFJg6E0ZT771woTPkFMlWrPPo/Uk
NiUAChsXokN2CNo/Jro6vg3wir/uZ98DpIqVhzCO87DH89955XnVFWwXwiAW2kiD
7Hd1MfBgyK7fLICEz5V6L52eRESD+Jb51jW6gqLv8IXfbLp8Vv7ek/WD8yqEmLxu
9uvAYuihgZnMnJ2PFsJzytifDWWoR03XO01GjVv8pfAF1kvw1UTqr+pFf+xVUfeZ
H/b7ov4UgEfOxWO24eijm2d93qnkBYz4Uv/xflO6XovHOiDVs4/Ijy648uLowRmn
f2yaU+JP2eNi7Z0fyPA5YtFerXUOEsgzKnTyd6jB9rqj8MI2U6UuWG2TQefAGa/6
K+Fsz5ycm/ItJ1Srez4QEp3tQR108IeRD1XrwNr6Y46US8FLFFlOXlHrFdjdcOEu
miyc2BlD0RjPJa2Li3LdXmIpSLENcs4s0l0/oAgmoWU7GeJtpgrWCDLDKIQPFzsm
jxZHwZYtqAaou6nzp7dpxqLjquBmIURnAUb8rbSdJHpxmgyc3guirnmMqR7imTta
sQ6eMGIugBZpRSToc10nnDuNN+wChy4/zy71qg6B1V3eZiBQuIbtdM97Nm2kyP3x
bRbACR8EFH+mpCzv1YK9zaJDXyMFJG2Vb1zdSH7Kb/QLxbfIX+y7YzSlAurPvUK0
/shuLM6/KIOVppCDfXM+FiJl9FHc7vKIxj8V7tJt+/nkfWW9IA2zKb/YBF3ZfEbN
6Pe4bv3V/AQwbPHb7sX87ke8ytXdh+WjlB7nOfrrXI7R8HfMF95fRtZUcDcS8NQZ
SAN3AQ6OuLzGjlEZEZGLApcuoCD3ErxTO0dG54vT46oO/Z38ij540YfHcV/uL2+B
R8lWDBdVyvIqT8Gxw+lFyygfs0ySojhuPnO7GbsjIbzIO55jTy0tdgcdO5stTCmr
X2eVR5VQ7VbxLWlRXUTHH/cKvtm1kKjO4YtlJRgW6amqmbCXv/V6JcWvgLrftKn2
VsOOc2HNF+KrMLb2+g8N0G5K8Apx0YGXc2p/gB8+9P1ozijob28tLFmyMxTcS7UL
y1BlndwN24duV/53zH34E02qp9tmtWWkaTmO90Oqw3jxgtySZFLsOpXVmbtnLNRr
21CM2+SaXGPTd2n4nuPkVV4l06ki1ZAN3H27gX6bu5RH86b5tompQrFUofCs4ONJ
lGgfkCjEAxP+Wrid96JpOttU2n19pP6MyO11Oq79CIpDs5ySh1x0qZ1ORzPjG34W
fmx4IIl/zf8uQ7oLAICd01Ib/XCopEEmv0hukmoHcZfoGiqtUQlNhGGKdJYOoqYM
lvDLUfkq8SUU9nmENhE0KpAPwkM8rMU/0g/KCT4CNU8VQkuRhdbUwOivqMaVMjTy
SH9c/Fy+iJZuwx1TOKeaLVZj3jmxyWL0AUxSTNs6do2hgL1r9nz3pAZnRwtg61Bx
i5q/vzBjaEVcLdbX2zN9L93yQBLWzf5ityp9HC0FrYy8xiJUg//DRsP43Z7WQrlL
8bcmr6l/659uar+VoA0inzEppuXwqJPL0tBIgDGidV131GGh0tSK4LOgC8jYV8/Y
vsxwWvW9JiHw+3lyfFBkD5A9gQOGh9o7Tp1ptnbSHH3ORRr1pHJQYe+CiK/2WFgD
1mh5uKP2V0u1+qHPrUCSLcO1yBYTza3kcSkn1uT66zlF6fuJUEaDPhZfWd1kkrOC
5MZhm0eoCPpMxc7szi0a/F88YK6oByG2kO+uX4Tx+yc9hOPuJHBx5uyddmAmMOub
KAUWqulDZlG87lcyYPpFxR2KqEUdJIRcH6jTTe3p7iX8XDZZELm0A3iMT98rxHwt
QB5OhM9GOCJ/Kbl8U9cECBDFxDDbNHCDdv8ZH3cYNky49Q5GDmeLKJTE6WsjitvN
rMiMIwuzNjBtzeoEOnxjtOO1ncAayy2zZYHRKTJYNpG1K1lkIFvv+qR+5Fjp/Fyo
kWd8ckPF7re45/A1VDbusS/T1eCJpK/xRkscB01xMAZV2Ro9HvzlkcXQf6H6Lytf
1GRF+ARFPEjUEym/tbIe6sikuIZnDge8WQv/HFqfZbjHfe3jtiKGMVbRQC9iIjON
SrjO7iJ7PzlEPex+BVe+ggD35fvGOouKXu/uDDrTq4X7iPv1RvmjXd29xaVAmXX8
lCLsOfVoUZ6WF0Fbh8pKdaPRftHwXmISGnknjcjB7lxYwbAasAlfGd9KT8fTm3gd
7sCh/VdHAqIOsn2G9sV2B4wZ9WSBBULLNk6WsLXWdExNb7bjeMaq0944QZeYXG45
pfmAwG+0Xx0M4KKuJMk8DUdw835PfTSqEnvbA56z91jGlMSjEGccNPs/Rhp6bQ+2
tMo1C0FyRD0NQDri1sfKb0SEoP97Rw8g8SrDRCsgKciAPdl+vFzR3o/Nemov+JLY
Rro9MdTaD5+yZtmM9dOXQGEsIQueQM7iQ/OXq+fl9Gwy150dPQE3SnG5nXSJ9aPV
rrHG2EjZfp9+fGVUtbUp43czfeKz95xH0ih7My1rHEjbAASVHohny24CzuzYmX0g
+pjv6xz1Wo7asCb70y4Z758FnkeTpl25A5vurv0+C4I0E3j5KE8ExpTvEXbUC8jN
GVvMAD6TtlG/EEKRzxQ440uPcWjxgiXF9e6PEWkP/hRE2pkHE73CkfIbIjBS4WUO
N3ZVrTlKVi2M3saQDSi7YXcJ4lINUViLuplRYKWHnm6TX5L0GwJuj0JOCyaBYk2i
25d+D5UhnU67rMqVWPcfkoDOGWvphUQ/rPH9xIvKuy184C0nx1/CpTi6kJoHZ94x
bWH7PKjsZcL66trZnZ/84wfot9wOm7eaY8PxwmvOytL9+E5U2hp749FzqaxMNR8H
Pu7Qx8K72GBrLocSRSPGfU5nwhMV90vphxlzgKBubD8uugN707+14bR3YNN48yjd
I3f6E1j4gyeb4jH6i2eFzqZEhcpcZafPsSRmSPwGIy8O8kXXHB3EQp4tGB4qsb8s
XdW5DR1qsfg7H3+4zhHk63EKR9zohsDovFqIAxq+zhZ/E2uHJbg0m1eQTiLdsDCt
pwKVjY8gU38gFEZ/ipI2xkmyzKNpwPBEaO4CzREXfrfMQYrBcHb9YnLCVg3EhLLT
TBi5il6m3YTW8KRJ5ms8B+3+xvkOQw84Rjc2UQh7mHbHU3VTRRFKr4hCJ6KCONrT
pvE1tTqfUSIUz21N+LoNo7h5F0d2hxWnHYm3Soc/zB6oD0GZ4FsdL1wKd8SHSOVc
CdCZiFvb2TSR54ZqXuwGpSbtdbyvKlxf7Gxrf5Ys7sR01R5VBr8i67nySZQEmMMK
kqcs0/KkmfTEvoV4MWE65UupLKzBYhjYfKrgvpf8VA9TAX1ezyqUGcFPixx9OBsv
zQF/GgGE/+0A/k/wQZSgtV8qyRbUTLgZKvvCN6N5c44bJL+7cj7Ow1aZbHcyKmbw
HMRIYAS0Cz6TfBJLN/Rq8EI6F7mmRCzWi8zZNzNAOt1mZiI1/APl8gPJwv4jvcFH
ztn8YpsaPHKkbxbt7NRjUFsDd+yFb/HYPwrVCARYye/2Y0INd8kt4TIU/fwdNmt5
Lbv46bXU8folW043TQJIQogHFArzHE1y4df54QfkMCkaKR6Pfy8duyGK/xN8HSx7
as0BbiTaVCAzLDSQ7s4PMBLM/kSD9jSGOfDJUhvEKNE/CJ8tiFOiyveJubw96bfI
P6QVU1urK8WNdIY9U1MHwO3L7vozm/Wllrr9kHgCveZ8CwuOPSUlRjth6Ip9YGM7
/IAHkgdCKcwbxSBvUCEHB3Dq5LuwxXk1QrsJyGlAfT/V+dw7MejPmczmrA8AuZW8
TGlFQx/VOuQqvGdKe9yNKMwXqCuAtKjYefZd9cRAMN6WZ5+pCTe+PO2O7KcMMu0g
3eKzyFx+kK8ZmprG1zYdXLynZJYYVhXQ3mHSdmayi0Rvu30e6Ct0axmN/wy7KsWs
FKn9Y+BgQQgRpq2dI1GWCLg7tAcyYHqxPzTccKj0vlSrwHGuXdHEJH6jUWqZ9baM
jTCLEJCWuLZHPzJ/iCIyKbUe2YbNrgIoBSYBf2G4+c1nKrJ6TaP2966f7yXzHuta
RHy6lM4iG0zlcXENSnpIWtuC2OK+oC7yJvOIjns6lf9BZvPBRfEdYdGwPhgKK85c
fX0YAifGxXJ+GVfg7atakc3Cdx5AZJXIZXJpfYJyaMx7LoHZBHfvQBm6FKLlIJmM
Ry3kQ+EocxLfgTE8Spn/w99x5CUMnxj8fFHEm2J6H2T1jMPinLrz7fZQyv9Oc3Gt
lZMRJkrvSeoDNLwbqbzAjp0p3A4qRMV4Qn3B08s5Ng8rwlTcoMpJ+oklKnwVcfd5
Vya6D82CxLUAu2+7quCI/MISUtXzRp3Wx+SfUa4Q9zViGq4Lp4LvWcOueKkVE80a
oPz6OAnPzQHvwujtNJUamW6cjLWlMU3CbvfcaXgWH8lnk+y1U2wnKUC0VsbJVcIb
bsbTrJvwTr7r7i1ylWPfESCDIv0Pvm0RcL2m8qRY+BhNVFwkivp3X2Gfqv6d0t2/
LYM8Bi/Wv5CUVR0smQj85lHndjKok17Ch7YMkvTBimtaw1QkqT3DCtRcM9w6XT+F
rNM9ueelwPy0pO9cJ1Z/KbOu5iD9+9aRqBimHs7B8m+GwHdNZPhmwaRIuO6APiE+
M0xN4gx9d6j+BI9Goo/q0x7uVrBFGMYPfchJJqmTV4acaPtSSMAhcETRgP/870by
Tvne+yuHtfnYSip4Lvo6Ozuk+EQxC39D9Dv/TIsFJ7CiPm99dlC118p3czPmVTKp
dkOXiCGnFJh5hjbZ/U7yJWhjcPm8SvOu+QjpPX8U7Xz19OVsGl6as144XLLIHakB
OXjCBsua9z5Iz65nlR6Kgm802sZMDD6ZqZPApialz6ovN5t2jv0i0g7v29QnSG1E
P7wj8yZcvPzbMALgHTpkjfVl+KivS0j/U2vPc8qCO/yp7Tlz+cJ+xODFbRQ8TB6n
yWTrVe8lkk5OStyubtFq5mbzjjsqKXZS4k+W35lpQqvYUcZRvtwXvMK5MXCnh/bX
T+a3GdBkh6893gcBfA38/ybGFK89ktPu92oHAbIw7LIIjW14mEUXqIA7QR6xCHls
pLO69a5QwURVQLyaTHyIQxptCqwIwA4rwr3ekO9TcEcRhgUohCqtx+dJLsQJ+F/I
GfCONIkRD7DK0WX1nbJtxzasqSEqiI3llD44LjrfzndK3H/IiiTr/ZEB0IlJlEKQ
hjfOpGpM9i62wR64Pphi5Kfl3nAlGdh0tlWNijLtjrxNMCHxCb1y105RmXXLiZ0v
amyr+DHPDQrV8Tij28eMv5a/JI53etZEgPI7+abeZZJcdAaMwt/vnUYNehQrEq56
sdfrEtW37du/yz9Fh3zeUUfQfCCB8ZjJyy5LRI3jr4LKi4beNHdWfq/0Kw1xPhzg
kX4G5fksZVmiSA5PAGd4ltJNX7ap3EpruaJNHMcuKfXKeDNmCYcEqjQbEs93EI5k
2jQDp1cBaIguPffIn9PJFq1WjicW8TYyRGs4PltpQW1iWhuc4/NmZRNC3N5CaTjU
QR7vRhikaltWF2fGs2Sv1sKS58BnTGKnEI29fNnhPW+73AB9VSge/lcpomCEAJQq
xSfv+1gYeFghor6VTc9AJZaIE6onQFQenyAnmGonfZq3wTwiuRuoTCl816t3PS3a
C9zdxnkzkkSIJCzEAeaUEw2+Qq2h4mX4ynGw+ysYvPdRtE925X0x1wsY1CNp2EnY
aR0pVANNL98z5/U3uT6y4yLRuDPcriz+2G2wbc2xdqLm0b6Nf7J2HZN1mMiWdBOU
aqCEgMxtUV/JUxjiZEMppV9TJEqEixQ+zCi+yMHds8yWV9Kjjr19AP4TJ0pV1J5k
XFUTlReVFlzdY7rFK0+TfR4cGsY9fC0X2Ze7qz2ZFN35VcSRjzq1DFXX1RD1NrH1
ShjpgfUOyTEGCtC7Xr4JSGJzWOvRarfgsQFXprn+sYVeTF0CLzOXlJUhPpqctZ4p
HWzZUEkQk2HZcPNTJMS2FLJuwXtchglUi7Fbmf+2ztnWDKKi2k2Pt3rh18jwvMQS
vU4DkbMCR5iQk0smyWb8YeRAwL0JJgzpu+yDQwnvJFYemBk7hU/FxlcI5WEcpVwy
BDafKOJz6BzH4H0Td3avn6SpNL1fHBYB1sVe1YsstQV/cnWaB7GHQZxINug1Izwh
rajq9bIjayT5wJsxZf/OG3owy8I8MhztvUAYK7gTVhIDijZi+7HlRvHIJdTcA8Gu
oUaS7P0q70tmykyhkufuVgKUFW7aJY7D2EQZvwfEet1U8jUY103epoatFgqgXhe5
tVnfxo6pjBzlSJ/gQq3LviscsHW8XZJSJ8hYbIlVJEGHM1wdFp8xeJfo1kScWevC
CiHhL1SyJViKaUsvH7Pq4bihgoPohBnwuwa5uiZCUJ+BWe3ub0qTvbZDbFuijR+y
8xTD5RKelz9eGRFC7VWQYV1/vmGH8V9AnAdKHJiDweplpomwyZnf9HZ735LuhrK4
6ElZOfy6XFdoDI7P+3E6RwY1DCxB5U+g0l1VT4TlRuzmF3OaiVZoqhKrLhIF88CD
+Z4ATX0wKMF9R9UkTk7214R1eLxNQ5JLH+m6S6Q0m4EetzbRQ8fGdY7Pn+TsM4D3
s9b0kH0bTTuEsh0XBRumt7nvfLVsfT6ry4nm+bJrauxz5SEqd1eZ/W19m7mBlpBB
tR7e3lybASX8mAx8b7uiZ5Gx6uVKMNcXNm39loo1nGI/k+aM0+hu7tyKs5FTmPuV
dxQwvPOzl5MAM6Fr9Ocy+2CTmTraZb8UpipRwNLeO3ZAub1qEkMmscV4fPtGVBzl
d8RoqR5WvZZfEK140YHYEkuKD+HtkOhoUnLOCPwSEeyFqPz6mTtvCIh+MBUs+gSI
XUvQ+SIiAwSqNRygr0frCPKCfnlMYo899dMuFL97AoyOkFng/cAw8nHWI6C9i1a8
SIcqiLzbduIyA7kt2B/0XQ1P0s+LIvrw2SWGdsknEgyuIvPAXsP0zmc/KI3uy8zW
1dH8GooBafzgmB+dp6/Iy/eihppSuaskO2Wmp74Rnp1Tddxk42Z23YF/XSnWILeI
7/NxYkxjhtgl8PWXcPzTmu7GghU64f0JHNixq7PLKgEbU6BQFDI4/tyTXc12m8oF
goFGc7Y5V8KxqBjhvnUipfvRdZnXNlsuvn0CpLtxj4x56X/bDg18+4FjAUlorDQN
hUbDIIkXneMJzq+ZJ8BU6w9uNB8IwW6hw8qr4AC4hdzpoGwEyvMjgbwKxklpuZ/B
EcfM9jyuWWjOSAhO6yeGVHAszbbrKDn5qn3bkTy5ghKGI35qOoR22j/u7uD2pF+M
i126RxJn99Lg+MfLG3Lw0VE8fvpIwrzz71Z7UlLCeKE0gKYuCiTPdrNQwuhLVdgV
WL3Gf0GwbQtNiPuNi+iaBEBijZSAKH9oIkFhN2dmlsk9h/tryYajrkPNdowC3/di
Yi6dPdm44eDk6DMwiN8CxjCkXtsWRM0jijiQL/T/AU6H5eGUJNJj5Aie1ZuUkkz/
9DszPT6R3o23ajlcN6XCFMVd4xVn+upIUTlweJjy2KBpXQLFvFjW0ekxhV24V2fj
r82tIe1e1zqlvxc1QG2bHpo5fzGq4OAobhN7cGPtWpEAIqAsrmSND0X+8ub7afRX
ZGvaDkzG645CHRzucZ1palMu7Ll7XhgCfE3iVMa6UbF4W9qp9m8nC/C+7fXtLJ0I
BEGCSKkQyi6jk7s+/JFwQgoBJ0+QS0jO3NrQ6LoOUTeKb9f2JAnDolaCKBxiIQ03
tANH2um+ln3e9Yhy+NtTbjtD9g/FBRYWktR6cjp3VQACAXxGZA2ix7AwEaEMecKk
hRW/oHUaLiM189yWFqdSEBe9g9KE369XjIoglv/3z21UDEaRnsJ4NGh8lDwWRDza
xBOUEVKOOTd8rMjgCPuxPCkBaiqu+FTfBhANM7qBKiH5GQFBeSlY9gQI5DLVYwxa
50Te5ybLTFsSa9kWWWGvyE7umrP9AB9cragkJL4zLg1RXpq3VofFbdd9UQVMJOu2
bLNBkuBLrMSRBM0n1JTbWI8kgjxCN7pnWfbavLgW/2C6HBR0NH5Eh+YxFXm9ezTa
yloCPJVUSw12SSD8bxQJxjmw0+hVsnKxoOPn+sCkchce0TsD1gqAt0+riX1Vvxx0
u48YRIIdrkM6jopMbUeIZliGkTRSQKel3Ggvw7U5/i8BCw0V5d32sURQpI/BkVxM
A5iUP1dqy4GaXY7NWSEB1ylmn9ipF5V1HlRzzyjohGbddJgp/H+v2pF9Zo/RreZ9
Uf2NQr4cZM4xlvQvRpgchVaaQ8rokCKGNB9Q/b1KSRIv6MyuBlmrJf6yIa1ToGhT
V3VMBT2+EG/L0B0ZTsEIx7cBY4GbsSaXhfUWMsbsB6nj3hdEvFL55zsl2iRPtf2q
RdozghuV7h+g9Hp9Ln2RrpSZlOoUgeRRo6FcQEgwrXiPgrRDr8Nn1KCD4yxmvyCx
8+6ZeXZ22IbhUeDqaSO1r8/8rl+NAk7sDren0y+WR/QNYDQGxOnKkG1pdWWUdCdo
8ErbJPawMiR0SZRodC+qK8r2am5TjHyNpfV0CPAvlyR4HYbHNl68SveNnhO94bZb
fLpRb3tXdFEXP17Red+3ahG/w3dCV1FZsK8x+ZoMt+lGxzClLwKo8vJYr9HatcWj
tj4ldostuwEeTfU5yKRFbwSQ0YmlRBQLL2qmJxzrAtl5k7pg9o9sS3MBUV7Mr7zv
WqNkjl49hzMMV2L/fWrH0l51DGFgqVKz1zQQyCcbuuwxNUjWrtOa/3oUK11q3HTj
REd3p2QDtyKcBwtovvYUHAlhHCEXxSjq+PfN/BrdSyT75C8iaD3G3G1zmMxPTxwJ
P7TfTNou+KZgZV8zJWXChh9K41J7f2X1sUoYxEWq02yRfMG7AAbsyLyEvpxkLEM7
uMJWH+KV8CLeNRokJW3SR+C9TQP0J/OZiT4U/QP7PZ1KcYj4kXQDU2IlCW+qN7Bo
hyxfsaWuIB0qUxHKQl3QrDJ0YLOjVAHz4t/teMRTO6o8l+HGPmjC4YklEHddEn2c
FxGydQndPYvFWzG9eZwmJNa2Jw2K9RdYQHPqSibfF6lyCvQRj/gvHO2ywVARQihr
nnHQzeX1a5q0Hlw3NlQ3zMINfxHOYwKDdpLROs0zIkaTeY1AYFs9bakSjnRpFK2f
lrBA8lTyAHuKiYJLaBja/c0iKGpnBMZo0nJI7nuq4vWNtdBfPWNKn1uIfV8wI7+J
dVqIoxndxbZw3mAbYNnF1IERDgz1/AY/o/Zfvfvp/IRTDdpfJCBSMsAtE6MueApX
YtOI3iD/f+H8mi9xEf8kAw==

`pragma protect end_protected
