��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�a�ȝ��M�(�A@�=u�R�%���I�ҝ�r/~�*'�{Z��� !�>�]~�c���0�lqg�oKD� _�8���RD(qK��u�oneϷ���V"��*�	�O�i��,"1���RN���O��HX�4�Uc���
�ω�s�Ȧ��?�ɔ�zi/E� `��Sߺ�_�(�&����`���'C��L�d�۱6�t��!c��Lc�7�<"�F]T���9��n�x���ۮq`M�+�㓍���pBR4�i��G���"��׍U���u�t��xu޸Y⾍Ιa���C�%V�(��$9눓�{eo�#~@�����KK�H).� W��/�\,Ǌ�Ҩ%����[�N%�հ�52<��,c��ӄ����fav�}}�^�6Y�>�Z��6��	=��E��i�~	�V�B̒���B�K~�L"礳��Pc�`��A1��f/Ѵv.oB��6���]L�[d���V�W�)�g��e��Ҽ�+^	�h�ԧK��e�?���o�`�b�q���%�!�_:?(֞c��n_�j��f ��91����Yos�{�Z��qEdc?H��#�y7��e!�Jb�d��+��4�f�*�O��/��x�FEz톼.w^p��u}2��>Fu#��w��x����I���*r{#��A�Y�@��2u�;�����+.�r�U!�	�$��M��H���s	M���� (:�L�6���qZ�AJiҲU���EF^�
�aVyP��R���O��
�pqt_֫0.D��@�߶�}�͗��|�v�򳄛[4������b|ܨ���k~��"�ͮo��i_��4�;0[�w`u�����K���=�8�,V1�FB@9���,��%M2��Ҧ�������K�M�F|��Дs275+N>&��;Ϭ�,�M��Q{˗!�Z�"�z��9�a�B�OS!��+c�E�����~�̀H[��U���*���iĳ�T d"A�n
i���e����t�4��2Xs�H(297TY�N��4����Q�kŃK�v���ѡYౣ���.�E�K$|��r\~sS�a2v��+2A�ay�T�x#�C��t�H>E��m*dP<���}���۸֌d��OiHs�um����5"���޻���}�>�!��t��r�C��Sy;/j�d������v�+�G��k�N��~�š�I$���mѺ��?�u��a���?�s:��p��h�KU��x��r��5�s�]��z��t?m,��Ғ����������@�gMC��s�^��dQ�~��d�����(m3D���������S�O<g�e��*S���C�=�^.�{��M��vP�o@�+�a�'w���De"t*o5�_��S�w���o��Dr���<&!HM"�b�����ɑ�3ٸp��PE8L�1	���w��@�·Ꮛ�ܹ�7�R�H�Ʋ�{����R�"��B����,�@#*,10y�S�yt���+h��N[� ��5��ڮ,j~�gv_ ��u=�y&�h/��<D�h{���ݼ�t������+ї�!$w����qS�B���Z�/�J$������`6Eu��%�W�ɘӽC�.P-:`���9ت��SHP�T�)�
#X����,S2s��SB�Îc{�!���:m���:����ݓj	MO_�а��y��oX���ՇE(���gc�>B%������A�8>�Gz`਼]~�>�PR��-�܈�+��ke0?#rOz˨�{.N63��S�y��?'�'���Jb�s���y5�9u��@X��X�X���_u�͠ky<̻d�͈���r�ڍ�Z�**��%̨f�J���_*n@R,],û>D&{D�O�5��\�9(v[��ۯ(*M�qz�V/J��5��F0��ubW�r�uA+��$NX��0��]"��8|���`^�W�eBzTQ��)bnW���H<ݓ���O���r����5���"g��aeV�n�}	�|����k�<2v��]���|t�!�'�|`$�,��1�d��S�и���n�ȇ6�\S�a�i�kB/qF�L (@�X>����#�����۹Л���#z� ӷ�>�܃Ay�¹���V��ǀ�r�F��S�{ɇ-�AU� �&���%�4_�xV�~ ���B�(�IHSC�k{a>b��nGP��lH���^�+Uh�}I\Z6���Do�����Y���D͘�v=�@��d�v���M�	�OY�E>P��:�],X�� U�्1��r��1Q4i����EB%Nn���ч��[�	<ק3�Uz�u���=mP��͏��,��3[q$L�P�rӰ�=2>F!�Y)^�uh�d���N=�;�3��('��?�a��=~��o���j�4aC�X� �F8pÅ�1�ؖ��5�%5�E� �NH�.h�ٚgg1��vke��������L�&�?�h5-U^.�Vj1�:'���ô�'9iv��`/�R����C�	=i���>��ئ�

�r���	bd�Y��[���"�y�4؆�H�z�w��,L\��x�}'뎦��U�n�$0�K�(�&��~���$���y��>�F�^)#����>��W0�H�p�A�#3>�D��҆�")�	ʈhڦ�|K�?q�P@u��^&��x<��F-q�^[�!��z;� 6+�����
b�ZT7�c�|�H��?g8�w`�P<�Q��Np��/&��vᘳ��K�M�w�.9$�2s���qF1M�j����`K�oz	��u��`�fM�/џʶ�x�7��ysb"�����Ru˵�\Z?��&��U�UmuK�z/�.k�sʥfJ�3Ǩ��+�Ov"W��|w?���_��$��K*�^y��[kl\J�7�g�T���TY)�����F�������!q�U��3�� ���#�ŬP��R ��UVxL�c�ɟ.��kg�I�O�ۦ�L�*��*�I�:z�;�0G�5l�&��Is�n����%���m%�L�������h�*C.܉%�?ų%��Z��4	:O�4���B4C��4ؾ�R��wL'ҹ�/��u�乤�2e��+Q%<dS���f���nI�&,�C�?4)������V�l���'�/��Ԓ�J��N��^d_�ȉ�ذ�$��l��`�*�J�lӶ4��v�h�h� ���8D.�<1�q�˥R�k�a������;J��6g:㡧��lyo� V�"zB�߲x��C}��56r#��#���K����Y�V�	��W!U��,�?���m /�\c2� ��cޘ�'��M�b�<�j� ]��3Ӛ��j4�c��~��CWƜI���$��b�U��"D�d~ǀ���
V֟p\a���IA�����T���:`v�r�ͽ_L��s��OF$�)!�� �ݒDx��������s�e�O`M�$�#.�B]����6��\|��~���DR#��u�����x���k�?�N�VRL.��m�5��6�ȅ�

�N:$)p�Xv�����$ؔIN�Z�H P�M>�1At�H�C�5��7� J�+eP�M�0�3��_�lx��q ����!�SG��@��.��#]c
L.G���:H	hڟm�uȵp+-���{0f1L4�ܙT��`Z�(p�{��V��a����
9�Hqj���<�H �b�쮭!o�m����S�ӈ��� kÐ0��}��`k�FޕU-���qb
�'^B�a.�������zp�8貰7��� �=<4m@~�w2�˨��`e�
�SB��jR��'���z�K/ȝ1$S��5�]\���߼T0�?��V|���9��pJ
��8�q�-�s̾����.�(�M[f}悚sr@ a���i�^30[z���&� t|}~��*I��8.������P�6x�gИy��pV�dB��_2D��h���Cb�Z�����_5�WN�X��/��M���&��pz/�Df޴�PL����V��=]�2l/(��߷6��L�����z�]y��z�N�b
!?�EN"�#I���q5�~�tT��l5�W�.X�r�n�����!�;϶����F�8���G�����q�K5�Lز4G{���E��3�Lz�#3���l+v4���Ï� �9 *�A��b
VNpN5����m�!���Oer����N�}���ն��I�#�]W�\&b�L;�B|��T���E����3�vn$�����t�Y����N��.�x����4�>L�U��M�&d�\���[�4
)3��$�\��y�6�>��v|欪G\� �f᭷���;�y&�#y���Y׎4�Md��0t2~���̸)*aц�� ����@�̭v7w�NQt6�k:��1A��?��F�<dMxZ��s��(�;˵B
��w�_;X#7~>����r����̀AfY��x�ڒ�x���T�$ihv8ռB�5&t/�?a�]�bF�1ߣ�-X��q�Wk�EVnꔇ�ӧ����s(�v[�j�k~o��؎7d�<��N�k���+��zp>BS�"=j8�CvX��yq���:�xz�^�~�
���}ԍ�`��m���mDq��^&y����XU\��r��5^�h�H��1{T!���J혝���"��@+�e� �Cz~/'���$�>c�.%[A�r����	:�[�3Kw�Q�9��bS�d,`�o�#�Q�r1�s6h��yL�.<2�����_M��kT���G�P ��G��)T�s�`�wkAE5剡�����X�ӎ���*lN$-X�.o�v��91�e�����@�����%��k���0WU Ȳ�q�RRq�m�1���hFf�2�~^��??������"iC�<�D 
$�/u	]V?�}����\��u�����pO$�^@b�S��X/��_SS�L�#�z�Pll���H�N���9/�M��Gl�fJ�^�զ�]Ƕqf���'�<���6�qo��:�j��5�nݔf!����|H��\#�eۏΝ�SS%z˶��5�e
��Fd�T��ɸ�������z}�P�Y"�;�ޏ�]S�^�4zY����-!ą���'�N�+3�5c���*�2����j��C�z�Y��Y���CU�|I������_��YHЦ����������о~��Z�����g��~��B��d�md�>��L�k�%�7�gI\r�]���?�/�f�쥙��M�Gc�Rz�{r�L<j>�!`�5#u]J��
e���s�n0{�cջ�(���Л�,�����9��a�O��K��N�Y�9Ϝj��oGɗEP��m�}>��^o� �=�{����K=Vo��{���x���� �rӪ�}5�@ pC'����a!�� ᤫq�����xK�'��V��e1��ꮖ��y�Q${��9�9y�^w7�<Y1�	Fd�I� �[/�}��*�6h5��@�X[N��X ��B4�FE*w���N<����*Nn��A ?���� 6UFO�vV�Oo!�,q�����`aǮʓ!e�8�89b�� [�0�$�W��v��P�=9�p
Y�]�ԕ��7��l��(�p*�������K�g�?�ݰ��=A��徴@��:��ב_��z�U���(��2HA�hϤ����C�Y
�Vw�Q��"�d@X�!X��n[��^r��~�w�� ֶ��X5��ǯ�rJ����ܐ6Sc�����*EC������ד���@�����w��������#B鿄�F��-Q���à�����7�F��j&���7�
�K ��3��:>a?������w���XJ{�ZS���|�@�Z�����+rr��c���~j��He�1*�jwl�(�C\o?U�G)��Ԅn��?��Q�]k1i|D6f\���ΰ5 �R������
�>=��UT���%���#,����P���}��4��A�֑�7�%�aT�=8=)�3�C��3��'pK��?Q�H�M� (O��5m��?��i[�������f�46��TN��#=(�sp�(Yf,$cȠ�x�J��sbp���b� �3;�_uxH�~kagh�b\,o�;B����4��k��Pv1��d��95��9q/P���{ ��"@ K,h�]��:��p����ɤ�iz��5[�C�x#�F����q�������y�WI�X����2�#��;.b�MD��n�lo�a������6pJ��G�<.�%d*m����IҡT��,b; ?�J)~�������܀�Qa�g��^Vp�C|q/*�1�m�:;�4������˪��}��E���'�z�D�v俨��-����R�E݋:�۱NI�#�z$�ֽ��G<�hs�y��ύ�t�o�4u����.iAL���%��b�Qf�f�U,��ϩ��t���Y�/������)��1�~U��;��i��ZƎw��63�� :&�Z2ǀb
��"��"dz�9isq+��ȝ����a�A9+�
�sw�R�9Ԑ�{�mn��=���hE��k�2��lĆ}1�����s�"&k8�`�7��j�����g�C�͖=���H ��۔����yM��=�N��~ʪ�ei��D�pk�i�����f�`kY7�+�ζRl�d��uR�4R����-Kǽ�{��{���(ԓ��ᜌ.�N���ge��(�v���(�g���W(���W#փ�"5g��$��ʥӾ��
�����M�A��ݪ�6������OS��a��0��C����U��B*#����݌�-���:X�!�(���Z�F�oD�V�6�����l!T�B"
� ��#�p��yF}L�����Oq��r����^`T��X,t�B?7ŎӅ��k�&���N�&{�D4j]�>�{MʻH�*4`I�Gq3nh��U�r�`�?�Xτ?���ê���ìn_h8����<r�7qlk���D����G��Fx�7�zlx�f����ͯT�(;��4���l���Ke�����3P�j�dP�쌲����XӋ��w��:���✢ч��/r�/�2���Y����*Æ��of�Ԯ �9d�.�IҬP�6Ӌ�(a�p�"d�IF����������C3ł�Ϧ��vU�C��~�`?`��
����?d��Q������[��1 -��Q�� |��ʀN��ͮ��]�Z6��d RԼ�r�C'�|f�[��X8q������"��o�l��-`�pXs�럀��[��b������b$_�ظT�D���� �cQB�7Ij��uT�
��Yf�q����f|�pȂm.u]X'��ϴQj���l�zw=1�l	��F��B7�7\����������`t�aW��B�������&6�)&�	���9@Id\i�5:���}ٞ��7ۤ�}����H�ő<I�R�[��+ܔ�|$�dO;w��$������<1���݌wS����a>�'�\���H��὜`��Ζ��'�^�L�)��]S�������I��4~�<R�������N�V�}�F
����/�}m�Ӟh�|����}g��� �%�Z�߶�WSp]EM�4��i:]F-)Ј￑b�6�^W�w��ݲ��ޭ�#�(����
;���p�����jƁ�0������A��X�9��Bi�>x�e�)�9�Z�O��]����K �̣��y��! �ZLPB)B�e��!]'�[g���+[�z�g�@����l��?��+�$)| ��P羃^����Ku�H�4��h�X�&�7�:x���zv;-bGW��b �W)� �0���4^��t��*0mO�-�o�tN �9�p�w{7~~�F����I�	���I#v�G�f��	�W��ƙD�G++aXQ~3@�ڒ2ǜ�/!��|�T�����#��ӈ>=��[��3�f��nQ����<�h�0ˋ�B-��ֱ�J��%f���?��<|?��S����
�#4��}���d�����a��qd �,ƐfI�p�"��gfTh�����>��B����u�(o,ڪ(cXz-����3�.��,����c�,�	Y)}��VK���a��h9'>�g��l�ȫD�y�.�k��#~0����"��[�PU�UIc�ʘ��ku�<�]ɯm�V�p��a{ۈ�Cҳ��~�˪��e���&#=�w/���*��F�����ċC�*P�PҜc���� {:�92�P䰧ӥ>緺R:�_!�8?���togNA}��U�@4JS�6�C���o~ã�Ji�$���z������)	��%�#G���~����_je��Yo=�!�~|m5����63"���P��C�i�ۇh{#��lZsxS�]����T2�g��a�t�_���EzK�Tҡ�!�Ձ���& p;H"��QjG�Dq��b)c���ft(~���qr��$�H+�-0��|ʙ�k���p����r�f�����tt�|�V
3�'\��[�DŇo�ax[�r=E�V/�(RFJ`�V��o�Ƃ�^+����_x�14���ʿ�_)��_����PǶ!��/)-�t�s����\��XTĕ5�_H��L�6��y�Ɨ�
�h#����ZN:���2#������_���Y�k��]dZ= 9P=��>�>�r	6�����~uXS�K�����j��������v���B7��8���'!�	��I�B�壍,�K����%B�5�����4 ��@C�/����s~��(z0.*�h[�k\'��3u�)#�f�8K>wI�>W#W.�;j�eGsbi�|P���*$��U6Cj���J���(�A�m�[{>�%�qY�Z'ñG�pkn8{�P��S�ӠF��O���#iwZ�8���Q9�l���
�B�: ���ؘ(c���3͕����p��l�(>�R��P��IO��X���o_��{As�[��/ }����������as��e��1Ȃ�Q\s�x�)͓ͯ���_3�NŮo�oM�+�K*B�����"�r����^SH�Ǿ1�"t�Y���ߞKJ����i�����	���١ �������M*|�V�U�Gkh�@��mQ�V�oX��o�R\�����n��y.G95�~n@:��jS��q��T���w�-z<�m(8~Dm3)��gr;���P�%c�r�����y�����oas((�,( p�g���Ǘ��m�UF��-,�j�JP,՘UR���08�TR>X��k.@�*� �Kȱ���}���P�9�ƫ?�Gz�A�+
Xˢ?���ci��-���{�@����]�G��msܔ�F�i���A�)hH[���A��@���u��z�X���o:���.��x$���-�b��%OX�͉<=�SE�4G$��/֝�����L=[o\��Av�#o�{������R>�U�8��x�XwqGB��ޑ����}�k���J�[z��p�@rj�4+w7!��4�z����
fۃ��x#J���B�&����s�[�w>,� ����%��o�cY�����
��ez�uԫ�2����+A�0�`�Oy���6YI�:�N�j�ϱٚ���y%|lV�1���;:rҋ��;�rI�����nA%z� �JA�ˍ�*�ݯ�g��k�3�9ʜ}�y��W��0���~�X�q�)��F�ת͏�U�?�FH>��ˁ���+�u�������Z��gWiaR� /u�ִ��"β]khW�P,�6T]:^�'�;A�.I�;OY�D��2�m{_#��M��ZF�^�bQ���\��ͤc�N�@���l��$�.n@F �}Fĉ�:-����$�K;L7�xר�h�=GH�-A����Ju�}T6�1	sOW	D�_�R��ᓣ�2�p��~�NvF >��&�V�MH�Y3�0FyZZzO��x�l{�Q��)�\�T���c3��C�����9����Pk/Gf0��ׯ��+ q��c��Y�1h����ʨBg�I
^�|�s}�71�����mKk�",����}�IZ����ɏu��wr��":A�ѵy� <����?g#$W�{��ܗk���e�k�؃��/8v���%ޫ7}�52C��a���L���`�B9�P�m�cY�N�F�r�Z.Y+���a�L`30�-x�&$M<>��?�}B땹66����MM��\z�'�<QvW/O"R�b�u�r�M���*�/~��9�7��$�:��IkM�!�!�=ww�Ve��nC�}b�Eے�e�u�2�hG�g/N*K�X��?B!ut�D[s�X>����l��œ�iʤ����o���ha�}���`s��S5�!	����5�;Y�@�������#����������=Ȗ����
]�V�A/�����M/�t�w��Gf����6{_L����`%����dܷ���!�v�s_j��@����0:��P��Xn�D��l��IY`7���X��yʕ�K��Tv��i���QB� p]�ni3����+�5���������4�d���۵m�U�dҲ<����X�`���!�v�Q�s�Ǫ�����t��+ D����L�vUB�<1�6;l~ Im�J�L�S^�$�_�a-9�=�w�<lq8K�w�-�bKqM�>��M9��m&D���Er�f�.o��u{��D�0_@�h�er���J�@���[�Y�YzI
�̭zDwb���;�4�?~�j�?��}�=YP4Pm��ŧ�;�ˠ7<�7��H�5K�a���@��Lȶ5�`/�i�n��U�WX�N߇i���.�1�AF{���_��1�o{�=<)�����4����;GQ�p��>��!���_ɣ8�M4v�O|-/�b�.Nw3����v�;r�'m/������PT���ʘq�W �_��ͺ?t�����StgCI��$�r�}��H��Du|1w�D�I8]����"(r��������Ʉln�G�<��\�+΢g�����A�,HyxFi��.f��`J���H.���	�S�ű�����*gEL�0��'�AiQF.�"xG5m�#ǲVTGo�=�k�8�-�����cx>}z�V�� .���81ZL#1`���!J�6J��_Z���������$����:���v���t�����,\A���B�bL�c�?l�1��)�h�����۳=�`��!Jq�_B�4h�[�jF���H�1�Ik�@+�pd["a�s[�&�����@�=�c��J������*F�c���	n�a 8@͞"��,i(z,6�<5�9��1{þ�4��"w`��[��I9|s���f"3P<B9���.b}Ũ��*u1�=^�FL��_CP��{4��@�eZXuQ��k���,�����`媫P*V�*	캷ʊ�Q<����A<�<�l��
OlӇ�t�#�:�!|�����WzN���\��:��g���h�r�~S�
l��oU<΂�ӫ���gOPu&{u����(-2��b@���f��E;oa�L{4�{8���| }���駧˫�	� �d(�|-Ƕj�;�ve�W�A7���:\琴��y��U�S��j�_7I	��5
�o`ͩ�����8#7��'K��Ɍ�)t���o�_��||��~�n��	����_���=r3_�+��=6���Xh�0���k"o&|���9���H���[�����p-���ѳ̈́�@ǌ=yz�3��VS���AQ�|\A֧թg�5g��to�ƿ;��֙.��窄����g�_��ٌǮ+�+ko�c���Eo���h ��PA�g�<������{�b��Q��	2��B��!����P�� �I�P�m3�ka���`�w?��<d��}��#b��˖BDDw2�"+2&�ڟ���|��c�bG����BQ�w�l�-�
�H��;<ض��w���\8����<�<�U��4���BX�vl��<�%� �u��Yr	�N�&� ��'�������|M���0;7�;�M&���v?�e�����0�ܟB�ٽ��^���q/�p&���j���Dͱ��P�9�] P9ï_����t4��h�J�	qR��
�%E�U��O
1�ho0���eޟ��ǺV�0Ҏ��[`��	�%J��^��Lt�K����L�{���
�L(��3���j�mE�,��ʦA�C_BC|�|2�h�OQ����d��נ�~�:$2���<�D9J�P{$�4�>����%;���׏d���bN�{�Mj9_�b�;���	��b�j8�~	^���8m4X��@�:�I�_���N�OJ:���`nGU��T����ӞO�R��	�*M�2,$F��1��G�u?���S��iҖ<>��3��6�a;�ȯ���Ի�o� ����?59�̐#�	_w?��Pl������z����QA����_��X��n�)X�fj�G��c�����~��k?�Tl�6�s��tG�l2���]f��_V�~�_��<�_,A�[�VTU<�����P�YV��ۧ@ux��5�aw�CtϸwO㕷��SW��w&ګT��.d?ٹ����F��C��	WɒS��y��0k����͵��?/�$0p6>^��ɂB��9fa3y�����$!�X��U(�1H�G.�I���J��4F�q�����u1%$�%�ÉD�{�J� �Y��ȕP�œ�_�����EB!�^�i�ɳ�|����l8��Εk��Ci���7�qH[���yY+�+��ړ�e,E%�Qz��j(O�b���c%9+)������{2cj1&PsO�=��;��IԎ����qPM<������a�R��}��N� �F�J[�0��d���Il�U��S�1n���v��cLtF��@��D��LN���@��H�h�5w}��q$B���S�)m�u@��m������ćI9�= �3y�,�L@>�l����\U�j���r�͙�/����Eɚ�B�ę���UZ9B\#Η Ye�@@{e��OǕ��G��@�,�:LdQ���~Z񫳠wxk�#����I�hdG~T%�1u���o�шU/8��YC�s����*���y\:?"�%�J쥿ꉢ��439~���N�ի.������}{�I_-G�������P��O�i�d��3T�Sω@�}^��o��l��~8�#;���}3b���'Z�����?I���Ͼ��#j��N-I�W���$�/(��E �e���8�TA���c�E�Ɇ��8�@F�ǌ�<Pᱮ�I����D>�x3{��g/N���k/�/,9�%*\�t��i@��V�q��ݝ��U�����������x[��9��H�˪� ޣ9��}��h�s��ں	͘7���h {��H+�n"v&ڹ��\��_�:�Cb����zO�*��]D��!��N�!茞%��<�h�L㹆W6�@�fϤ�wV[+��r�\4B0�%9���$TkmT����qR`b�:G�OO��>A��o�|�4q��9���|�u:�5�-Z띠{��<�;8��UG�G�8jr��U��E�����9�H�t9G�J���o�ޢ�v��.�7%�&%��tzPEr�T5��N]H�ib?zC�>d�X�?Rٔ*5�D��\���~ol�	F�f� =E��d��u����bG���<�	Z	ا��
!ג���.�m<��뜙����,۝7�VBt�<�s�wf��,l�����[�'����5j�J�� �	�@�m��Ĥߨ���������8�-����F�'�bg��
 �Z�7N]ߚM��]8�8mn�q�+!R*�5��b̃��	����k�҅I^�1�V���f�&11.���u>��i�!�Y�!��ծ��4�rKѽ��*�3�)�汰�5 �xZ�8�x������@��Y��~Z���/�־�X�J��A7 Q�W�n�����8��p|yU��� TPT*Ȑ�r�t�Zl�vW�/�(PԪ��K,$�,���:������U�E���Z"г��]~f�D���^i`����Az���z�z�t���l{����g	�H���L����p���!���%Ƣr��(j͇VY�˫���X�U��F�D���t�g��0`CO^��ǏFXnPې^���3�r�ӳ1y���w��Bu��Q�W��-��
���/y���K@X��4b��x"�M��R���G��9N�g$]�UG=�=E�RD7[�ID.��wn���D'�hn6��� �^OR{�g�I�<}�/�����a�g좿bo�!�?Ä�k��_a2#C�U��pw�{f ���א
!��2&��8�E7̟(���S��mAT���7�r�[�L�&�2%��z�R�f�V�8x���pv�/�,��@e�K��#��k�;9FS�A!6�4�#����.�T��c#��`�4ynԙzIֲ�9�Q9��R����Am��>^�uM�Z&�r�R�����f��e�:>hB�����P���M;~�:���Խ�+���6U��˿,��Я���#��U��c�|V2��[]�9r�!��۾W"O'�����"EЎ|fĚJ�S�EWa%��n�K�k�>�^SH�˒5��i�mlo� �s����V�EL��2��x��/��p���q2��z�>c���/d�(��K�a�j|=��߲��0� ���
K�8k�Kķ�H���ۤ�Z��sc���S���{ރ�1j�y�E��̺s�p$�с�﬎�p�6"�Z:���X�Nj��/��hj��I�Hf�3L��O�3�zj��m�d�.Z��Y߯�5��"��<��?��hE���ߖ�����"`�R�`�F��(��<��OI�^j<F��*@�raSR)=g�FҲ:�(�����f)��9Bt�̢��+��4O��]�p�8����H�+�W�w��
Vf)D�
�²�Q��aл6�?tT��ބ�)���c�h����=`5�E��8��'ݝ$�T$5�z��RE��c��W!���f��Gph��q�zڀ0�d�%�x�H�7�?Cq��HL��
�ٗ��~�1��2�=���4�?��2L��/@�V�4�c�`�a�9 �g�f#�[�"i�qqQ�{u�aU~��:���Դ	pav� p6�w����b�X�L��}��ԝ��z�c�j�1ù!b�lֻ
Ӭ�C��ۄl�-�`|pC�X9ځ�fD�^E�h��	G%E�����l��R�m��Y�#��W����^w6�;�V��� ��D�ǅO����Y�z�2`��k�hY��ګy!��W�0k�B�K��H����[ �P��$����ms��U�l5��Qt|�1�ޛ<�h����Qvx�ww�VW��V�@��SCְ��O��96�2�c���d'ز������r�o������AEԴ[�n����Pi-{(�)
�@��uX�K�X��=$M,�⠮Q���MqI}vv���`��4HH�x�&<��PE��2�rڵ@
�ʤ@y��:zd�x86=���?�5�J7�"'.�-�˭'�k�f��E�zR�F�@�j�x��@lX���w$Ϲ��х+0�!�9�2�����:��7`�}���_��ne&�F��.���RY�~Q�u܄��9���t͜�|���aF�u��|-�VtU��c�� ����\ѓ���D9��q����Ц!*�c�L�e�>&��޽���c�=ӄ�n�țT4,sA�$��9� �4�Aegh+�v����>�\�F1c�L:#� �/���7A�\��+�ʏ%d�}u��� ��X%�9��IO�ǵ�(?��~�$��$/�G�x r�1ڰ�,(�i e^�@S@�������W䗆V&���:f��d~ �Dʳ�({2]`8�����p������O	zĝX|u�������,H0���X<�{&/D0c�l�(V
�����Xw[����p�f���g;��F�L:�0�䧰=>�	�ւl2���s������?��4>��H��\�`�9[Ycr<�5���S�¿���S��&�0�/M�s�`��{�����o�[�4�G��y�k���	^M���4��І�9��p�l����^r`���؋u^�=8��m��ͭ��*��6��2X6�!�����:/�������,r��oZ�X�w(Y�x���aR��,-�%�J��k(�O!v�F��s�\Ň������N��I<*��{��<
e��� ٪�B��w�e�=Qvs����~�4/��ʓ��%���r�e���[s�R���� G)H1w����V�m.g�<<<�T�E$����=XW��r�bys60�8,�'����B�a�0�AS"�@�+k��v�5W�{@���u�s�s�"������ú�����ѿ8Ų?7&xbm7���RX��k*i��ǯ.�C�U�5���Q��U7`��Lb����"D"N��hZ�,��_�B�Q�<W�؊UU���2� Ɇ�� ��H�m�}͑n;�0aֻavh���B�Z+�whj�.8�����뜞**�`�Gl��=��%�&�ݢ�خm��X�?,�es�c�[n�%�L>Cd���/'�$�?X+�N~�lH���*��d�g��IA7*g<<=6�֡ ��Fj�z����	�
>��ﭔ8Rx��t��~���;n�T"1|8��6dL`���2����W�X5�rl<�i�H�%/D�Q�RU(�YlPO��B,O�3�����(a�B��D�7_{�c�{��˂�Ԝ ����`�d>.��ޅI8�oº�6܆)6C��pǘi5��A����U\��$�h�Уw�D�#q=�'s��� Ɛp%�ZUJcG"q<Ja�?|����s���pj������j����ى4�G���F�I��^���8Z��[�
H
�ː��B�_�г�!����Y�آ0k���62t�L��jn���.� Ϳ�A>ێ���ϱ�/[��Zl-���_+q1�zB;���w��P��@9IU-O<[7Gt��6�^�d328��c'�Ɣ�w��2!�"�����}n�c�D8;�	@?5�
�����-�X@6�^�EL�;�zf?c�fz�ү������ob�s�m�( -���&c�7e�/
�R����m�P��,6O���=�׿D�|V�
*�~y�>���k��ф0�� V�΋zn(�}z� #���{����_�R|���/�~;/���x�Or:4�M-Ƨ�hɻkY�����$)��
m�J��c�ўW����E�ꋀk��Z�|�E��q-�=��ΰ�/��B�f,(��og-zׂ�yQ������QLeۍ�&����eE�\+Z��d��}����a>Yz=F���_ I�m��.n�vBs�d0�w��I8(j`���^z��\K��?,"ݮ7q��4�!0���gHU�|Ï���]JroX�ڧ �"7|7��w��b?ޫ�����u=���ZE�p]��G5f��ΰ҉#��}�j���?1̝���{��R�d#N�.`9.ǩ��G�a����yH�}.��d��p��e����ک�P����$j���EJR�n�1�#"�U1)����I�j�].Z�6�O���O���d�u\0щ*�߷藜("E*��m�3<�w9����)a�WTSBS��-��1gc��A�DR^�u��n ?6G"(v;ǆk&O��C����a(p<ur
���~+H�D�$����[��
�6f{�+�9�9x2�=���Aq+����{�mT�������>iAd����?��z��kz�)�|o���mԗi�*�Sc�
W�W��d�J� ��;��i�iu��J/mO��5�.�aI�ɄŦt��Ŝ��K�c�]��*���3&yd�v ���"�_�)9�׶�b�</�������g�|�j6��-mϝ6���zd���F�h�`���(,xĢ_Smω�+��I\p�b3�����2���=f��+T}��s-+{��׊�|�O�eiVB�֖����@����*��c0�9�ϼ�q��+R��˔����2`�tbyt������K�["�O�b�������Aq�Y���/���g�-����?9r���֏R��D�Z�p����՞�A||�%��;=S���ǔ(k�( =]� /���)�wA�����%���<I��TBD�|���:c�'�5ߺ��\8���o����Ӱ�;?���/���u���*��6Ƹz(�~{�)n��z��2�R=[�E�$E��0x����P�!�'�y#���F驄-W����b�pz��m���N{
�V��Ϧ�B�i�q��������v�� ��ʣ�� ε�޺��;cۄ�����OW��5��46�s�!�K�T�<�%ޜK���IS*XV`V���@�Z��ա�aUbz����H���a���>����r�uS�zS�q�M��ȗ���\N�FM�!��Ǝ�[���UY�3<*��:z�퓤�DB^��_)���\��uY�����OV|6`��Ad��ܑ�_�sC|��;�����y�&tyS9A:���+��,_4���T���d����$�
#
S�Q)%ӎz��M���sT!�؇��B�����65�;OZ�]ߊU52 1Y�kdR� �,vCeLBl�q�)ب Җ|4s�Z^��
�)b:���Fo ��/�5�~C �s��9}�V�����ӌ�Y�21�j;����#" I�y���ש�N�C���D�O��%�3�_A����I]��z5�s+��Ӟml���O�;�\!r�#6�~u��{��������l�dm�b���R���J���\X:��i*�?��,"�$~�S�������xš��P'`����若х�ќ��8��ԥ���>�T[�x�HGE�G�������E�prڄ"MǴ:{��p���#h,T�̩�Fg���!݀��
eŴl�a�����B��'�����R���h�Ѻ}���9c�y��C<
��\�@r5���#�H5�&Q9� ��{�Sa/c�F��f���T3�=󻢐P�7��Gb�
]��m�� lW�4z��U�N�;$�RG���J8����B�y2�,U��Ĵ�Z�QK�K:���/e#��>)��[��YGg�U��@�`-���"�7p��~�� �o�q��57;VW���%yRƢ���h��������D�^�V���Ҝ���Xt(M����q=yN?��"���f�=d���T��M�/Su|�h��eM����jEh��e����|=����t �&D�yv��/�@��J�r��4oF�+w�����]����B�d�dንsT�H�	�}j�橡�e�F1���k.�c�M���l�|С{>y[I'&��8�N�,i��n��!�&2[��s�ز伕���¨&�Rk%�~h�+��$� k봃�S��"ae�c@K���gq�K�8
'�(;���'4�١�Ѓ���K+��j��"G���N�	��\_vx���Y�c�(��eO��j�$�X>UV���.7���>=����'��Y�R]*�Zbw��'m�h_v1�\׊V�Y�p�B
� œm�q<���mV����z��H�5���h&�b�;I��mThT&VdT�A������؆�j�UW.ۇ5�.�1� �U���a�	׊�]�Y���+�k%b�n_�9G'�l�`B�~�Y�����3�z
	�1dYٷ�mܢ���\��7�[� +�!��Iz��� M�i�g�iw,����1e-׈�hJ�����e�5�����l�Ź��a��O�����q0NQ����P��o���ߝQ.C�؈�N	�<�U:�H!'U��Ş�F����(��Z�(�����MT����6�︂r�~\[�Pʓ_r0(ȊF����Y�b2[v
���/��;o΃n��}u��d�9�����}N}�d?�C����S��i�:C����|�ҷS㈴On����C������C'>
��O[�Zlh�m��'�:�O�!�����9�t�=�`r�p{_����&0b�t���f�i�P@�L�ct#�/��M ��{ h@���C���>G��}�D F��,���	z���H��<L��K%�[��������%���c'-e{�9���Nv qă�"�cg|�{�`�cZ�y�����y#L�HN����1s�>��3�goo�ڻ_/�F��$Vw�3���j�����R�fd���x�I�az�@- �We�lA���Nt�Q�s�l �5�Щ��(���"i]�҂ϔ��cw��\�.�	[<u�%�KY��y�s���>)�P�G?{d�!�^k����%��c	g���Nl��EG�{~@Hc���Fld�v#�t���/��I�0���z0���k���W�]��z�dRJ�G��ߋ�^L_`ķ�L4gR��s��'Ȋ�����U#?��}S���BRc����#��ї6+�q�X8���i�_/"���)��q4��,�rT$=�q�r8��CM
�RD�hQ4�Q�K�����|	����o��UB����Nw�f����k�K�صAoJ'�#;���z�ۧ�_8�FX�#nL��Ʀ��jK�-�G�R��62�*54PV�E�ܔ�hS���s�L�t���b!@8mV?��������[z����h=��s$G<v���Q/ջ�<��|�u̥���I<~����G�D"'��(�UD���ŝ�
�Y��0J
e'���������M�$�_4����a�15����F����zq>����qpֻ�=Ĵ5ܣo��B�_�d)N)�3�"`V�q��"�;$��n���͇8��I@�i2��e�S��d�A}�JP�ͺ�j�/5�Ϥ�C�E�%*�Xh�*uHc�j$����ǳ�g�����be��� ghh�,l�g���K$��.�}mX���⫂X"���af��R�n���#bl��n
J`[��Q��x�2s�|q<N\�w.���7�t������}xb:��,0�Z��'$��_c�(F�|��*����aE��~�zKn�d �M�VOMW?eq��%�v9����H"�T��Qv�,��3���\���z�݆��D�*+=r��T>^wIS��7�0W���ʣ�
~i�;�n^���(��A�r}S����*�3����'��@s)J[��&e�A�rg�JO��r��rhyE��nR�%�H�i-n[�����r�]��j��W�9�א��;���Q���El��"�s����zɽ��ҁ��ӏ���~yӟn��R�	�uZ(]R��gY`^�s��M�?g�6σ
��"��d�6�����H�}aT'{���0�e^�5�d��$	����;V"��S��1_�"jG;������"C�h���x��Sa��qH�4\���:�DQRa��쑌3|^�YB��
�W?�7��U	��fN�_�Q+�|��zvm��z�p��sn�"L2�n5���enp:n��ܤ���;�a,iyq�A��ll�^�����9<���jU%�����|��ۿQ����<��  ��2$;R�=��kq�m
lg��L�?�3�yPt}�N,(���g��s��N�b��ᐸ�bk��U���*K��������d.]��sUS�H�s�Ƞ���2�\4����1 =OW�~q���W�*V?�)W�~̤�ܽC��Ѧm��fxN��T�yi.��/D��&DDeX&=�g3A,Β�B4	�h���S�Y����yрd��_y�yL%{�̷�Ϡ>q�Fd���^�6��[șD[�V�KZ&�rY��W����_B���0�|ֶ�M�C.i1�NU�HN}���;�1}�7V���T�����<76�A4f27G<�}o��f��`;ǋ�I�݃���f����ҳ�jd.S���a� ��d=�{ڔ�F�v㣐Rm"�U�������t�v_듰��Z%X�K̳���/~p��ƚ�(y?$��&&���T�3`��*���~ E��i���hD����/��g+C�Dĵ�U)�N�1+���:.K���{�s��s�T�E�C������Ҩ��}�����`��{mJ���OS���5�0D\��_�DLT��n��k'Ls�Y0��Ӛt�cǴ^5��1�fE��h��E瞴�͸+M��&0[�6�m�#�'z�~��E#wdA��I�w
u��\vsT
�kJF�R;*�e.�I�"����(م��"���l���M���@(K��9zt�< �H��cK[Y����Qf=Vq۫�j�4�tWn1��pߘA���iX��p�,4N�R�ªSd8쿒�%��̖-����G*;����w�
�\��A�8��������ʱ��5j���͘�4�Xо�#�af9�-a|�4ۂ�w���у��j}#υ�6�\�B�#`�@Eg���8�j�g��=u�����i/��48���'�����$�c��u&0�}�9�x�����J"�[*R���f�<��/�'��HO��t�2"���1��ߋ��8�:�>d) #��|�l���z��p��B��+	���BɃ|��zN>gqu�W��ر�@���C��\��e�>�]��'��NH����e��l��Ŋ�� ��Dm���i�r,��w�'[�E|�-����vײco�|c�:l��<�z�,��e~ '�kROQ@�5�}ϱ��ZX��s��Mj���������8��U(τ\3�qm���'u�(�#�/����%�'F�\���CŔ<7`�'4�U �0/z�����#�3�@>��Sk�5��Ȁ�9�n/���I�X�xa�v��8��՝�`h�$��؟µT2���n�6q�JZ N/��ٞ��O��4G����t��_�9k�l���iT�٭��fqBe��ǎ6��g��N7��*�p1W1��z� �O�f{��}E� v��_���Is�7���C;��H�c���r'�����={���w�+&5��B�8!m8O��G
EY�XZ���5ڹ����	���x��_�~P���J�J���V_]��zzj�B(�?Q槝�m����3�ipG�r@�u��.����Q�3A��g0=�4�B��5v=gYh��6�
����K�MC�w��S)�v7���	��0/�|%Lp���9�I���p�v��_Xi���=���Kɺ����̑�m'��]�	:�i��!�q�6���:��[