// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
3K3hBz7ydp2lEzzuBJPM/9VI6Zb+j/sfEncVkG5t6pP+u+tbSs3XLc7CnNlByPU3
eQjQaY6y6GWh1GNKDVmqMZtzJqmiPtO2GfqwQAV3pdNOLMGn1Nuh8xXeQeha2P4D
ANGmAwPpag73UPAXm7rly41JHQKdRkCkCrRZMhEZkQI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1280 )
`pragma protect data_block
9vWJvLakfOAzH7pROdw58sN/7xgAKfb4nl3SYMLCJCX5DOVJmT33iiemvCKaLxik
ek7v6P/qby2OOz20+3siS4itVSKVkrR70zcAlzQk6Ui22Y7BALxoOHUzC28rVoT2
2CGgjCJR0rNyYBNnLuIWzUUh6vVjhKTE3M1TGtEDX+8lCIkk/gauLkHQ++F2hD9A
naDmgvCkR0OQN+oTBIQDlruEdzmemz6vErM2s4ufdfJJdRGHhjDZ9M3bK4skqDuQ
EgBLtcBbnpTwP5jOmnVyPPlB4fy+gUX39RulpK6GAVRQPcEIV9c1BlxyTL9x9t6R
SAlVhMkhC7Y+VglhjA5EerWPY8QOZhwKBObEUynsBb57zXlPM1nHEP1dK4I9KkDk
+cYCs0PwQl/4ud1fe2xwJOpoagu3woqansTjDato0y5v9Dcsdg6QmmCu+Fvx3Dtf
7D/NaBL9s8NE1ME5foivLJ3pFIN9TJSoPl2YGqcVZLY3IDz9/WHqBIxhYtikqxk3
vyXZWkPB73pdvWSWw0Y1OaiZPTufEpiC9MSImnlyNaHNwvagTHCm0SEPAYAh5itK
rhMtxGXM5ShCWT1dp9Vg5PWh4835DtDjzB5m70K54AmzDR6pI4RPo9ezOgGt/3GU
cwOBmKs7I5aWTvsg+S8Eagg/TOpJg28im6b3LBax0I998i7FCPat1skDWv1aokoX
xxlA9712g86hZBhcjPGvXwiTg/blFFjYT7n2zRErOLEIoCH+00Fw/ElY5S9OPx5K
UWHSQgejhGkdcLQUHkuMzMmWWca3JtAVrKqsDEcMqjoTJ2+MUlFVfr6KC9BGcrRT
tdNVaTkOEYiV5nyYo+jj5OYwPN5CTls4/Lntw4ZfdYafuvB6+xT+y+bTKJa01JjO
ZsHSn23RpFX73qt+ayFEl9CBRwxf9T1y+bKvT3EwYy+e/hYejr7XDv331OsVV3Kr
NRveD1BavdU1SpRYFnLLilmC568ch2ZXx5bb3zKfbdXXvn0wyIDkupWF1kUbeFNB
itgABxbaufpYROBr4/ZmQvzx4tfqs96g0tXMARTk48owx9rUaiW2euTyvXHOrJ3p
Ia1SgvuPR7E/gfN5ZirplWJFj7BeomdiN24BFKHo2UY/h7UFZA7yZvX9Ej37MvJZ
9OvPuZmyiYni+IMZJnYkB4uDPg5NDCO7g56w3xf52es2iXtrLcpLU6LiFB+6aAaA
lLXTCPTXHoPT4YAgVVKQ0rfROmQBxJSZYOn9t0/qA8DT4TeeZro/aQYIlwVyTrcQ
3pa9R9j/pZ9WUmovI8jLcq934I4Dr/xqIFt8ZDNXNh3oPnh4Sevnge6nzn/HlkgI
osJU59ntMTP+EmpeRYQqgi++RrbBrSVp7fRhlorBG9dV/WFxQyuWD/P0tkLa2Q2N
jkimZB5dXbQIbzo+ArDcXKHnLGUvQkW+ItNW6P6CQDqoocfHr3HOFhYOrJ/m+I7r
q1ZTd2rr94ea25yhXogjcCpGojdTG/DQsPGoCMJnEHlDkGlVvCEumCdTXKlN0ysd
xkgtBANMxUsLqMdx8Dv04IVkWrN9tVdZjjlDPM42jEr0xyZfRW8e5faRrr2w+mdE
+hha4Zl3S6Spq1bz9im+pKp3sGroUYiw79eQabucyIeCbmR7PiZLco2MXHcvsEXp
KKCaeErzjMkpPaAU9tj4TNezedieBrDTKFoCCiHubF8=

`pragma protect end_protected
