// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GyyJ+tZY19RMyoNKkm1t0VeT46U4JMMybYQVRw6wuIZlpDzLJJXtmyN0d1ks77R4
veEm6qsEnXdLdXKaZZpo9/i7EcuEFQ4pXp+oJ2Y85J9uc+lbmAp6WLjfFFz2lPA3
w7seFszDnRWCU21Ix0Vp3xrfaLksKlIUTksgwnauUjjwijO7YGBkiw==
//pragma protect end_key_block
//pragma protect digest_block
AnQUZMrj8XitoqtxKwyKUoZdvek=
//pragma protect end_digest_block
//pragma protect data_block
+RwNKarDSMdYq0Hl78sX+2IqHmJwbiShnGBUe0ixThcUD7Jvm5Wcz0Idzt2Ar3fG
RqYChBlw+2QDrf2PLY1aiibBaYjOcSKDGN/XnOCzdEZsF6mrsmCuX8kFLQdyIcMR
Ff4jU57UMCsB4S6A1AxOHGx2aEof1yYjPiTdxV1w9GG8zJARWf+25uBxY429yC60
WgRiOb3ZnjAtwP6E8v0BqKbCeg34F/eG/8PwxOGp4tmQh0YaLMSFMYgAqxKrGFQ6
bbRv6sex2AOjvopHBTNJwOYE2Wbe6nUDqkC4XRV9ZX5tD/3fwvmVeVTbG/lkH50n
BCr/eKNcAPfuUf+MZ3zeR2vSIaEMAU+gyGHG5mbN7AzXYDJxvDuM4/6RV4ds9YpT
6hmsATifnP5fDJnR8Amkq/BpAaaXaWjespwNKHDYEeFnfMHl8Dre1tYt1KBP8hoK
I4xLwZy5y/WmzukNcYnqqVNtnaCJta4kx9zammzjeLgNiyM97koK6KIIMSrsRI5l
oci0mbzXwGKkhfjCJwSiydNami5RXZzBwJwZDDsZ8CBRePaDIxGm1gdt1UIFcS2o
F4myN9sBAodSarnbuBJTmTxAZkrbrQfAsfIDTn3mmYthVpwwUzeQ6VUySO45vThM
2m9zqes7fVCzXV7OPOlmoIxUMmXS5b4PkFTs2aGZp1mZoPabrGrlM7igZbPLp+h6
BHtj5z92WnoN2zrBcOlFnZ6Xuu5wIu7b6MHlYq7GE/jxJJdZj41SUlWbDxZ/sAXR
zAwPCwlEelvMKniSI4CNcQJK4rzqlnAk6R0Z/JP/CoY44ODBHXOJ1xTBHMlc24/U
5ACqeViSJSsbRO/upMXeCPqWOUqzx2aAa1x+MEp3reK0mOTRDwK13yHd9TBvg4EE
yv4JR8KkL0ceS7hj3DW1VARMZ/gElwmjZFkuje03JaUtTKv7w3OkcCYB5kQol8V4
GVnX+66fdMDmde8CMl1ncUUxnK5VqO+7RRicmDGl7wg1K1raNzhwPewhMsS/v4Ec
Azpe88rSc32CljvtjNQmhsAwPHBeqbO9T40VSefKwGdl3mMsG2lEFci0dqvvOfpY
IDzaiIORQ94EKOoBrEXnPCHFCTTKN5HYLImx3Fzae3u9okDe28BLZx/eKgiJDjHf
5weozOh+8ge5va078MglPA88cMHVwxJlnM02MiRU5XrgLJq0ghZzX5nqPM8kUydD
CloC7stPYy+OhcjeVrOkZQvYFcO2PF96XRDkeU04kRqTZX2IMmzFY9Ze2vPZf+Pq
Ub/UhMC7b1rbe3nr3uG0THXJd7fJoQ6r2Ipw40c/kBp/MjYi5wY5CdBdYvNbijjf
LrmLQ7UodgVkJLdHivXWMXv+/H1MoMXIRbPCEQqC6mZ1aoGpT6OUmsVuIyI+Bqto
IMPpd7NwLU+RnIJo7D15PIpO31z8t8ERLOZcL2Ak0A9xd99GuKHbHzkmQuplJuJc
33n31qdSH5B5wFKuPnPyVJEtuqxsGPPlz3IQ+wh8SIVGSwqqxqUWPDGl5uWK3832
v6XJkcqOzoxqsRGjr07WyEHK0kwiNZ3QsyR1GDHurq8MZd0jX51YRmyQDckquEnL
mcl92hcjrtz7v6hsGHcuc9AQpZhK9kbSfs0Yn3aj2LmDobB0c1ZjY5taJ1/qIEDK
H9VwPHPhPVTA5FyrhV98IQpdElscg5uGQMCatuEBEDkWobtuPA+jN9nHNhBSn4PA
tYftGhLMCI+jACXYjrVu2HhDIJE6xLCo2weS3AeT88MIFPOsgyVfZUIg0Fj6LJJp
lS3I9f2CbP3T6JPncEtjfvU3rSlV0OogZrD2FwNoyYKAwWFhTWi7tZSO2vHI8pVS
lktHnzQ9QCkAZSwkDw3Y4Daqv7VXQOgR7c5W9ckZ8rsuXBb8qGkPz3qNgCMg6/PE
SsL3P5RfGQS6iSF7t7+u6MWo/i8heIa/pWxfvftihXqJdxQhy4SocQTqwqfBgo0Z
EIDOQnYDgFqGL7KbjlTdt+6Yigon/AE2e7yZShjIjKJzkQ3ZKcTiNxZNomi6pVJd
RREQXlw2GQQKNw1B/yQzTcSUx4jyV1oMeuAy/KjWGLP6gp3hdLVijHOrIA7g1BA7
0ts7Sj2DEoBnfoNMMkNRUHpPEInXZ9KKbQImXZeBPtK9ozGi1OGxQKaV9HlERp0f
AGu8JyBHwdNqyqwHH/K5iMu0FyJuDkL82RqLPZ39zNx642YlzpQSDhwJUc9uS7nc
qqFvM21YUq51zHgJhb1EEDkiJt3pbVSoZG51i2f8yqgfgXFKtgce2rT4dKZFkgmC
msO+lZh9FDFFCh56v6W9gK1YBl38/Kv7HsPLkbFfAKAV77CsuqqywMvD1rwlyF6P
iQb745NzTOp0GHsP4RleGhTdD42308W20NxLqDHoD2WPTNYXFDq7fS2vrSClpmbL
Wi+K1O0Z1Vjf/ixgJHgkoWF4cP0yWq6exh/7kEgw0H41BbDG4vvdhLkJCuQ/n//e
m+xz2ouaCP1+tzgNgsQFJj0po1EV42U+w+eqgTNHmIAX089xk8FVN4QSPd4bP0BW
Hv8+AFWPj0HwJsTmju8LjVTs7HzjmwzyrvtR2uv59WbyA6J5qluvWzIcoDUcVuPs
L9vKS4CI1qDCyw8W4r/79wtdxo1sEgJsoHjK8H2Hu20svm4d0il5TtaRb+p7a252
fv5foDbD1mhtdzTImVogBd3TFlkftAmX8Qk9vL69Dcgvh8SGStAFtHtdb8TQEreo
y7V2C4ozW1LCEhwp9dTlOiz2GSCMYLwwe8ViIwcOMLOrfKxIqxgUoVsakIgCWcjT
woLDs3LsY0YEmT6OH5arJtksveQprrrXj+eVcknnO7QAKxRxtVenI46fAJCvMjVa
/xQHjK2zM3hdlBbQOlQS8AYMGl3G++ae/ZN7TUGj5/ORH7fqJE8RAt1u8jWVwcTr
BuW0yFt0SiOr/MmSuRxms04RKycwS/wrnklBKnGcaiZe9EyfVdpWQtiPLAR69SyJ
4juHdH8KRpqmCKVxCG/0Y6yZ4kKOFtiKtmDfXLg077RG1mPnDuUWji3hlpG3jqzt
nAD/U60XKmdJEXZMxqmVrDLZ6Q+M74lvk8rqbTP/e5liQoFzdj3eBO++xIJT0UP7
JiDU3jtIVeWYhfYA1K/AYd9J5ZV6ePquxMJNgjl8pAYEZzU7YpXvVI8wK8M9M+7E
mUxd5G5QMHt+V5s7oBWuTdqWT66iQkeOVazXgfOatP8EllJIwSNuwKWlAh8E6u6D
W/yU7IPFQu6/NhvV4wlm1JkUap+OKwCJOEyKIk6tc9cysKSL8J3x6ug3BfsOiFuZ
QCq0o30LMbcEwclayef5px0hnbnFwoBlCCoAPCzcILVmTDTR+BAHc722JQqt1d2P
049isTKbHriJT9C7ptzc0P9bkcc2+O/pdHgOxc823nM5NEx/6MjlY5T37Q1HhpzM
1ckCKHDj8AitsG9/WOpJfDnkT8AJr+/wCBJTwSQQjhM93UzY8P6+7yQAeaYTusoR
fRLuOVpJdDXUFA1CdE9E53JhO5T94+QTtx//5IWAlYubzgq7XgR9ooN+21PsDOvv
G3A43ty39FkswSCL18clJOiUjx0QUvTAfU38X7G0l9AMVD5cjPRmfo0EovZP+bXL
aUvc9KxoOv20Tx7DZBs6R/f/Wz0yAtULBxajgdGHowt7IehaubpwmvC7ywPWpqJS
qV6MYvVj42GfZfgsyqL/qGdJ2Q/oRccY+zBo4gsHLxEe2Nck7Hx2Fj+wUMeofxAB
9OPOIJJ6AhaP3Hx7gg1DvqIhs3W90U7WE5BzBs33jbzqejs2XsN37DOdC0sQUmHI
6jN0iHOa7Ze9C4cT/8qoX5of2GLIGkINIuRI1QTuwIee0SvU+x3h3G91goy1ClHO
zycNhg2cnJv4F2iWsWwFYvY1r0GinZu0LV6Y92yTnKbeFXYzcU1GcyxLEhDq4Cox
CGZdwnHZibUWDY+wV2X+Fk8GrhqFcOp9woWkq7YRHGqQ95v02WO/dRjps+gkPTk+
YxthoyPUGnLqih9YNkmn2n19Cns+JkBEjoGlHOLiu2ZYEgM/s+ehNQOrXAu4DQFv
HGC7HInr3QgzwbtjWPEbHUrntGGTRJg1OGdzWzKz5fenbGlvdfDyLVzI510snO43
afrepCTh24merBS4BjplHaTKsuIoEZDx6yt5e3q18pneJXooknS5VoVSSmwSxjnh
hbEJb6GyIqutJicAK934f3lZ1gNUkKHXTz4dcTtF7IORSg/09Vzm40i7YdOfcNxS
ziRhp77PzG5ri85Qpxz/6XiGqtlE7UMT/mEBHTKgNUPAy4aKBTtSlVpAhuNT3QQp
9f3mdsICI2f7GnbERnArm/gwxoI3gICdLK3/Sdk1ZgVaKFQAPIFfXDp0vVPZukpF
MROfYQmstVUWf1z3D4KOTjS8cqkUlpjbt12klVNtz55m2h3NixI6yVh7q18TuckC
UaF1fsLniijI3+DE/Xb788nwAQhJ2mWVEtwmRcwFCeFRR/i4ku+kPyBgjEjq9EER
rHjCsvjAkxHuP6Ve03afgV93Emafw8OJEzM2vGWxlmm3QV8UuxRAnieZYqOxtXqF
F2MLReQscglwBF65RNYnAJNROBg84EV9BDPOD6w8ps04RhX/Mu4Yx3VwccfW50kG
NJ9dOxYjKcfRsqG/gU+9AE2IqVQHLBWM3Ine73LjzRP3Fao7ypeKJgXVmt3U9a5o
nalCNUV2ppoStOuh+4u34vIqKKwylPqmbrjg6meNNtEzoZyUGOPd+RDB1axVPINr
tpk9Dt+bQPP/NlmxkOnhCTTMw7Noth3kOtw0CJvdqVs6I9K0CfHYqQVgZZpCeINY
N0dZY9Fg0XYfK2xvCmA58oOp7g18lpLEv2M3+lpDBrrStpbKWOAD608o7SuNOQHe
KwXpANhU290dduRqYqQ6AQ1B/dQYpfT5qzRo4Dzyc3I5ry9ANKuuiQ2cp8k7XSJs
exZcR5MjuqORetBvkyzKrvZr4hpG5ZVGb0lvTB4jIVoKrWCfZPl3t7dnRNIcRvzM
2OKVq1plGl2TcAOHTCvZ9JcWbIE+B8Yj+2K/P9dCL0zOw251gpVydawlYM+55iXZ
zfZGclRtDiQqHu8tfPxCu2nVocg6QFEJjOCh9wFdb3pmsysEC1yKHexjpdI9gxY7
3DU1yYoNu5z7Dt0Bts6Rkf1U8zy4Zqr5n1C1ITN4gjEwZSAW3fXop91iuE/x4VvK
/WDhO6uF6SJ5pw6f+4d9B0nz4tLv4OkXkHN5/yrtUBmHYZ35KUP1LMgYJC/VJbkx
zfUw570GvVqHjS50cZHzQxLwTJe79iOrZ4LIlPIws/XweP67XU2ujgogn75bqcUz
G23X5KOjWaXlPf2oWsX9AKacpxsscHIPvpzNkVQ52u4r+mZIpC3idjPlplm3otT/
ySRP3c5jdTWDqGDrOlON944NWubI882lEz3jApDZHoEB/EoDP2VpR/HOndKHQc0v
6S6W0OKq2RRnx3mPcd48QciNNuYWPDfmGmEe09nDlvj1eFDWjY2AMC00rN685CYX
xfpdmVEtlzkhRmWsSpPSau5lqnSRN/rjnAkzm/yf/PffskfLXi+1NoJiZFesADFs
+FHXib/n6Gh+WDsaIeRHm2/ei4rA5KZB3ZrkiqgXlXUu9+FCTdMrnC4m0UiUvpu1
7odtlTJ4Jk1E1w6Y7pXxy/Oq3VvQYiTEZvWu3SM46vw0pg8E/b0KBN2NcaXQYPZa
+FjJC5GnGeD+cmuWBWnRWtSfzsDIrG5gA1+ZiuCUhfTOUsvXMEAWFaehyJBrU1Y9
ehIpQy5/HzOZonpsdaPF+JED+wnVGnDDWwgvWpXiSOt5XhD6aicIjSutQHV/Ztbe
OGkrs6jymniIF3Bw3cq+EetJ1qZd5UyQ7p3/6pWxFvm78ilpZCk7mKlg0yGB8D6r
YkdP4mNYUlyDnyskKMasqhwEVQHv1KxVacFk0T5k0Tuehae2Lj9zNrTUNVXU0z3S
5ljHEUWhpBYGCUwsQDePcs6DwBky7tPEpyrau6MsPkcJUPggRQw954GZzWmYcrsX
gBTj/XhOkVku1sNnlInpT03C8MSXl+/hlqxscly2B5ciWI9E82Zj9aYmTeqZ/8sw
/p8bE549LwenUOChoTmcgWFaWaaWo73J/gE8NAS1POXEyPX6wui+xKCccy0q0l/h
vTw8Hj7qxH/dfkZl1KP+RhJUxBB3dmVyOG5+GwQ9BKOkSHffB4YatkgVxMrlKK16
Pk3lslib0RTUpGnsO9D0yn0gQDEhrn6nl6xeUwz+rcKkRDtB43LtT3xpLQGrJ3Ck
pGidadRjn/NC1+CkJO3x5IycFGTEMWMz1Yz/2FMiUN3XdLruDS+8rKIPah5tgn53
0V2XakZSXlpSBlkAkH0SgkD0Kw3unjL/Hcx8ClIv2DDNepKEKcrSJcP9y2v8e3F7
IPupDMp7A+Pf9D0QMiysn2O9JanmOMrE0KiQVuNMCsNuu4Cg4zm1FwV6fYHocZOl
EpjHWb75fjRwg/N2AsLm5fQsSDxWe3BCONynAbHwbx9JMfT0vuFpKS03o1faT4EN
QA+GS6uf5SDWrEwLv46XovJpHh1ZyelkHXHOa7D/fMBwxXoBLoy1YJ9os0naER4B
uOJyGMHRivjgualMRSrSEFxHD13BU0OIUhO3F5x6tI9SFIDU4avtLe86CSnymVYC
HOfvI4ocjRKyrGIg7PwYzlVi/48TRSC7lTdPSnv6D3aj3O3iYfobrE1kJAfLY4Zw
Nz5BaoI7L8wE3pYJufDCuaCvAyIgvkW5+IRnZ/KbzJ/FY1p5HQ4FgcGi+nUvWi/E
IC+GamuqmD3W6ZLn3y0tF68S43Szlgm2k/TaQ9P9FI96t/U58DeW4TTCzryMpLRb
HtOPqt+QlMIKdbpksuEu7uEK8d2A5Bzm31FRm/MZLjIJwga/0ZiQeUWSUj5vPoo8
x1NWcjcqW3aGAZ4ELYV97EMdCQByZkVYhtmfxZfoj2w7AVNdIy3dB4e4ujPkQ1Hc
p1hLnfgbpokxxypfDJT3cHwsCL9OgI9MQ4L02qbZ5DvUc8lDTN3U+Rr3ppz5mLqy
el23tZWoBIbK+HsAo1cU0AeBujTgxmkCawPTE5KRd3rukKLA6T0W5IW9+lKQQ3NX
y6XnfZe5ALOWGZWD5FJ0qtf7JPI5xlW4GoKEcHrtEB6QFEm3W5gcRbJib3esH4G7
LIysj55yH6D3hkZQKrLJekqU1IxNGVfMz5lq8caRxkXTRR6gRGTM/YZ4sA333F+S
kZphPASUgTLWZfqIdzYK9UOp7s9HJ05qHUtEc1Ko+Hda12AYhsZh+QEN5sMG76Je
pE0BfgEmufHVSgN/JCd/uT7lb6Sv+feotghEvJ/qbsIL9t+BhL3NzBjBlKCYjb6m
wOe64UxzI0gNl8Z3rS33snHGEJvkucpyB8xkrVjIkgKmwiUNryygH5xh5eQN2P8F
qnlu1/Jth+YfFokybtn63KvcYCkc9yaJgCq38bLJyJH3aF99KjrrB5sWmdBHFx2d
zJhrYQU2Ekh9ti16DoUL9utLke1/YVNVnLaTyEdohqYyjKT5jXuWPCf/Ug2rn6Lw
nTX73ehrN5aLX3lIO2FSgBYneHZKy+to7zQUQ9z+t/QZCAvP1WktElFCkfEKlgQO
lXJYBknWWVfmn+XHz19F6vC7jtiTXu0Qf1ivxgEADEfoRPZOu9slBGrtQLJlCPWe
CBYxZ4Pjgo8m9Ndt+0xj5gNOGkKmyDtr+0TwQJWLQE/B/uq+iKccaY4AyF6pIPZT
UbkcHmbwdzmz13O1hctS5a28sXNjwiL5lHXwYtVSJtWhsz3DaBA1o0aKk/ei5HiT
Rvx4fzCC4jwocBMEKliNC052bIdy/DbSkAXN8cpkKuX7c1WoU70tD6qI+ML1LHn2
ZDprnQrxXU7chWOpOsWpWiMaViyx6K8Mn5LGepaCCizfs3PTBrYTlpRvh+j1U2yw
9Tg/blG2uHQOzK8PjrTykuqV1EgbQEjxZnafhzOtGqmF88ad3vK2mgskKJdOS6Yq
bY7j+IQDI6wF417hF/E9pMK2v+YhUxx+PNd3HorawuDbsWsBP/tvtLvu0HraTcUV
a/QlyDHdX/8vnZYiSHBYmUOPl+0lV3SS7nYugwb/iSTP0O0Wrzc/e3e/RPjge5jU
Kgt2PlZSBu58GbzkKrKjOYXWF5gMCV93LWZC45hihVb33m3r+ahT8py6W9kGxsjW
0dLVm3K2cQZP/sSg8WbI38y70eQpIFOSDT5Pcvg14RB8tgsDv/ImWsGxXqduza29
QHQDwXj0bqydcydzz1/z4f2UImJuTkhjiedoo1kFh9h3gpqwBLn1kiqOHtAiuOIt
X/h8UPjHttL9R6t9Sxi57VX/0kXQNKvFO9mWRuLRLPLdu6pjJlOI8B6XAgeGkcAb
Shm+g/YNZgQesp5Nt96PiH0FqPIl6Ea+MX+pMP32iGUnzO/oxPXPO9DjIZcAhTiQ
xfDUPWd+JOATA+atVooYq97OZBUzPV+tZdb5KoTCilJ/toMSLcCDbdVViNHEFSbh
zZHG+hgscFxyivtqfqwmOuAbloBQWD47/5XPt4Jz9QD0c8mfC1E9ZIJ6jGLKvikK
hcoVtw/bl4bLogvqDvAuqD8dPxtctDQNRhwAWkjhEJ2o93jj+h2bI0srVVjFMYYf
Z70GJYsOQU1PayPP6me3oSyvHcH03BZfdBCOtuSlTzSg5vSGCbTfWxbTSXn3kDRA
AZnM6Q2/FSdIIs1sKnV0zFIf9UK0kuZcIXFc0F+p6AxNpugriry/sUPBvMxUTqi7
fRR2JGyrIke/8nU0BO5mwEI5iq4NV2oRox9YP8BJekLoXkOAgwDK6wcMuq7CwXUv
sAoE9KtP79x9o+dAf/7GhsGrHg6ROuvW8WzIbjuOJb8dCtChP0gTgooAbJLh4oAx
mIwIgvGzzTOqfPVt1oFBJk9NT3VKp8npMT7o9mf4sNW5mgmZiXo21CGSG0UUsrcz
OdXeb1H93Or2jDlWx55Yk9d57aPUmr7YbnuSWFuddRd2jaAFrLDI+TGFUz8dNwyD
EUcJ7Zr/3ZY32BqFNEqhMcUr291sgfnvg7z85pgqUYNh5FpfgJVTPH8U3YQlPkWY
bwY3cmWB8a1Q9o1zapNqIyASYCJL5K79uka5e0LTkXM20YWidMqZbjajkCdlGqxu
5g09PCeQ0mmOpSsDfPOhXMqFxl0rkGvUbEasRwoit7pM4NZ7Vg7nAk59GLfCHQZS
WEWa83nLqvkhl22SqusCgKUThgzebqWRTn8MqqnUPGaufuiwORdblqNbhifgAmbo
Ib48y8I3gYq3egQ3WQ7USgRdnqd9bTg1+i8JvQyc1TpYYR0qIums8KEdruLAgalI
9Mv7kJJHq2P6C2DVHrguIlOaRofW+YeOfiVq7fnAnLKfgHAMWLW2JLywb+rLEM5L
UZApDKKphQUhSZ13rR8rhIwkN7X9BqVruSb6EnSfFwEpn7wTj7AWxJBsjHpRWVB2
Dl72WKCzwrxbpWFsO5e3f2Vo6LZIlxdXutz9N97EHtMyEQIUA6DjE0sCvDjG93nj
vDn3qE53JLT3d3Tbec8XvKA24wj2UzG7wEeLdfJttB6368wyyWNFb45eN9szQJ13
0PHAYzmlMATMnia6mBbxg9jpw3ihK6KuC6F6U6WVpz7IyhJI2NgmDVKHVq0Iyj20
RAT+L/daXW7pdXgQjyCb+J/BC4l+4FpXNB8x86zOHBbyGbQ0VSBLjygKqDQyG9U+
wk0d50Lv1lxk3vVA8iUXf9pxvMrZHhZqa7n8ZICxR2pmy5H0P12tLLVKUXtaDl3U
xuKcPYyltM3gO9HuU3buYyysDAiepTVIcoOYHGQaKMNea6Tf6mPj3oBFEO3vkVaE
P7HsRLxeyNxU5Db8ZJLScV8/0pERfMys9wV6CkijmxxAAD2v7xQIkaF/iF9zFu03
Wyc55JMrnf2PwThdcJeP4/PvEiVFN4oGUhJQrbaA4HmcZIwEDZnVsKEscsYjkkKC
Ql2brwoaVHba+8apNeVVpggIG6DowANMH8ddvau3SiQbhRNxarOYCydMPHUvKpd5
R27YqFGOPy5Tt/n5tC+rx4NwxnYPdyXofmq7c5UwYzrf6foYfrqUL2B7BqsATrBl
li7hug4/whOqlKQ6KzYExpkXAQULVAcbGnmYB9So4LBqHmyxkrHIjmELsG4NCq4o
y1XdHSMPwyqmi1EcqJ3FIdY5s/5o6qfWaalDnLNqEwVIVHBSTMrGNVUq0qkmjXUV
tOvHq7xZ9OZQvsVM34IWR+jrsTnYl5IVkeY4MkR/1Iu6lW4MxQqXFiWPxgb5ic7p
1CCIoOVgIHkhRLQDNJfIZCxgzMbSGFKRFSf2rZ5f6Vkn2BxpvNCY+f7/TJITRiCw
nBjktarwnPpplRDA9ys3aO51FOkiHPmW4hzEFQv6BCSjPLtAxJNq4UwkA4JSs4po
JYZN01ZOA7qPTIGd/mOcLqs6YBxSlIc9UbMSQjb1/lnFpctVwuKkQ5BKwwpxSj33
YG6NSwAf5mfufj/f0NE2Rw8f5LfZRDSrsIHJaYvSWL1tAr1fRi74PAaGLIL0UX0h
dwAgqpF4K4m5lDKrHqONfxKlS4xvDvdJH9sd1T/EnNqRRLyphcQXWDBmtp9MzW7c
LymSDZjN6oF/FJMsseGoOZEHF+5ws2QPzoVZNiHzxa66pfyTLbB2olc6T2sCF4pR
ZmeJsw8YX2vkBzRLMC82w9xx60tAD98siX2t6JO3Sa5DdngjyDZBqxJ+9SXjau8Q
nDU+HxojFoys7uzgP4DWKCXKPLcwmt8CeIExbNuUjsJ/+wczHD+iUavNEvuKfMbH
oEccJ2oIQHXvaueeY6TGdinIntDaC9H8RgXLNopPQUV1YCTZ69TICizvRHCQXuDL
l+bTjIH3hWx90ag6gcP4R6WN8a0Od3QnbPrHf/O1LRp4UDbqSdrOIXFEs+4I4fiL
N14hqLq0LHf+OmXFyZQWuCjxBfGjkBszRwYthyVxijxp/p15z27tYGDsHmUGUDF0
2IRVnirLFChMvVTYrT0sclS8mhysroVM7MGfj5QFNLp047nlKr0VaNlSKhViWST7
5fu40WayAc+2zZdZhTRWC7t6/4A4iN5jOFcP+AnP1XLexUFDKoFyjam21Ma/y1lh
BpyRavwm1Z4yLP3OT7x0GbPU44j8p8u7jKetVepKsviDlPLQfFi7ooLsfKwJqm07
ftZKw2GqDt6oqWnL5Dz2488niffMZhs7M+0Y/gDoLppOQ5qHopO8Yd6x/lQZCB40
6NaO9VCIluv9zt/jEbgXuziWpqxFMF7mY2+RHgcU6cPw2vpcF8zeCclcoWm/3s0M
7S3pdsyMyixyVBVZy9KsnbGxcJmmjJjsAGuZ4KpzZ1XxMuJQaZ5Y1zAN0KokFasF
ghOcGJiu9M3li/WQOMV+xaIm/8F2y9Z7AmZElPQoNlVhqDTWSNqQRz0VBjhW+pem
kJgR6ddyCLtxIJa7VrG2mMba7/F8GomCMAW9D32Rf1Urp4sGVOGnp49iEwCw8yv6
8v3Ct3idDnSOJ6DUwCqnKt2DfB6Y+hzgbO0sTwZSmlPfClAWkX8Z2hblCyupK+SO
3KitK+JBFRt9V5UprYvpE+bUOmO5EhPb7pF+yL/lQRuwuGAvacbQDZNH0+KmKlLr
wArIYBojmBzF073bkeUK+52Sp/HLXywn6jWrvwxjbotCDl43xMTy6KLPcETAre8R
oKVR+qWjqDhs1r5hSn3J7D+UPfJqkwRARM0NYIuikmGwQb4HcRzkcn7vuvAbZJK2
saYxMC7OeVXa0OVHx1avCqmFTj+Vzl6ZcsYZML71CNZqj+PlGubktQvxK3nV520Z
Hi6Rpqbm/zRRLW4UFoZuq+9PnBxSfRnofJzgbqgK+9Vw80vHpWr/1C1NL7UYfMRH
yrcZR3JJRCrgOq3O6xMg4rDc9Z/mpFhFNFEN5FTLaxX0Xk+eYtXFzYitmJKTobdk
311YwC/3mEXqvr/i8mqmecF+wxnamFdSiRkaXZxlp3AQ9T96a0eyW8V+qERmDf17
N7AzaLz1Lf2yCbCObGisgzNC3wDHkLeLCpoElp0Pk3Ozz2nmU/OKfl343ncxCGtk
cH8a3li3zjVxWgrKW5BvWwz13m/EcZLh9KG6I/vlua/uW+LZU1QY5H/NHvw6Gz/N
0P6W/7lNgI59BLudnZIzaE2svd+6v1SFlyl7EkbZDqfSrPK/wnZJdE91QW3Td4JA
MzjCYW7tZCmDcWPcJY3CV0uihd76+2r3C+EuZRpOicWA5B1C2W+3eNvP2Xozc/4z
tKeciA+uyFmoOD2ZYUO/lGxMXi9JRaltSMtadc1nt2bPlmZIp2XLzzRWXR1qD9Wn
3NoJeAhPJlZ9Qoh3j9gvQGvx9BKwtTnIsJtrFCOIdtGd8vd6dWNyvNRrhpn4paqO
H03+9UHRbJc4qZJTJvBuSj6w8NuO64kf8U2EZoFxbAeIjVXNehi2/z32IO9621O8
G7lK+DEcgjJuMIlKiFL6jBHyJnhvwxYpwNiDiDvp9rCkor77kca0peqJewAjzslB
Tw33rNYuAo04LxMxfgWQKE7oO2BTP7NyW3zXIGcTA13mJl8Y1sEnJhCOY8FEx6cz
MA51TIQufnwNdJY+8pdKdSVKUY/Zbm3JbRWZx6h1Yu3X0V//np96kwJg8U6+CRwj
Oh1a1VmosEpof3tj0BOvH+bfr7NnFlDP3B0Ca8pd/9v6hsoK4ri9fShB8V1EIN8w
hfPB2dJpe0SjkdbqCBw2bX7dMz2VSusxBGYNDDRB57qdgGMTORLKy/mS4N7hFa7R
7pz/4CUEM+PbPME/JOLTGApuJfO3iHefjCXIIbwyJHZNlpbRAm8sRi8r94ZwlD+I
RxtBlnCqB+KzVzr2O59EDODKVW3+dbvTvjuAHaAq7FZxLlZPpzEMXqptQj+s+cyA
U2omViHchlaJJk//9LTorg7Crz0GhjKO+KUfa1STlKAGzCGHxT1dT1BLvbNwcsov
XaUWePUV9/EY3p7F4ibSGPE4S03f/KlNNBo4WXGIEkvGq+vWqCwi8m932+YysI7d
vC/Ld5mXNZKQbQPRIsftyiva2ET4OPmqU8yLqOK1lsZBSQb5bG2UWKLvdIpEoAAA
viUu76nFE+9r2rIebUW1TbqwNCBRcZPccg58QpJmFaKgOElUA51/xF+5saimULrt
irL78pyt8kmyhtm/n1x7e6ZL5SmzF8XdynRQhmsyH9wLU8dOzzlYUCUGZFgdgLmp
6gxjNwL2GoLh2fI7zRYy5r8A0eqBF9lYYJtpigA1r9JPSoXN2LDFG8kjLl4ki/Mh
9xn+d8phdwgGXx4wfngXn1r13W1s2aKaFRmsvqkOe515Xc37nMg6LVEadlNSsEfd
ZH7MBuaGPYNNI0iTmhqGuMp58+7eNfvVlqYw9gqdw1EMwdoTcvoQlUUJDvJqYhOm
Lilyx7WZW6GKs5apsD0yID9Uo7YfiiqEB4ewqqA8LcvuVtXJFqGOLJVYgsblZ6TS
4ypoGN/IUZWYx1iIP2alFjH7ph71Ssrdgeq8rAVLJSKZ0b+YJs4zxqx1AAqIXDYT
YL09T8uJpWB3n+A2K8Ok5GO0i4x4zrC4GoQrJv/MVk3+Z1fenetP1T2y/PdJbcDL
aQHl+QHDdxdbW4fTkDCmm+k2BaJ3JLNLmVjPf3o3JKgbnd/sftOJzcUhynLzrHmP
9L8CqY6w6LleSzr4rxuna+j4Gviu2HggAyEnsNnrw1Lwmg33RhatuGcW2iHrfcO6
Fc+gl0d6N8gawQhNJb9NE7aF2a/nxD3xOpmsXpDCi6CUwX68907DtwXKLRg475NK
htanp6D4oVGWdueoH6vDy5Pt8ELvPukjra5IQJlrCtlmGTn1MQprWjRDyjb5P+kl
Res4rBsaW9xYAaWJPtABMWaMD7yE3fmK+myLWwi79JZErivjYfHTjY5FF3jRs2Mk
WD7oqEBykCWe73A/Xlz4PcyhpWoPIKfYkZMJOw4DkR7fndhqwg/lKaAdsgnVT5mI
p9aCGSbvB1sM+6NonYC5dp7WI6NA/yrQSvW+SCGS4UuNoj/nHXcP7MGs8l5MnAGu
pqk0M2EDue0+0mf3XleyzCw8qA+bYOCZz8BFQcLvZirlXBr9GXDjqwgxdfaItmYn
dRXQQqJwl4UwZCyVv2FjhM05tghVzDQuRbQIFMnNjK4qOeMsU/KsoKIZFUKfGupQ
AIMwZ3syO2SQ4/Wbw+KsCtWbw8ojeqXy00PpPpq3ozpUqR6efzHUw5lKSouLfxQl
b0qxg9gdqB2/ECSSzf4U72GU2VSVyteD90joRkvLupfOqSRe0p21NLPPMzokkQbo
eLhB3tO2KoTCYaurER3sRm/05XAaubcazecaztm2PPl/4Kwht9kI1ASwL/+cX1AK
zdMbuSUFY/xj72y3YDDWzk158FczXY7oQOby6SHgK1ufU3M+X31yd3Ahga1p1Crz
d4pd91/1S6zyy60FGzv0TEgfHgBmTOnaRCf1BTXN1jNCCD9Ri87GdU44QOrwhSR2
RDjnZwgudwPSNkmwZU2xR3Jlf6f82XEJ+Jc12nKlfzT62+1xzAQnxyOsUoCS8vtN
GFbMFt6oAIVcYx/9j8ufrEKuPrEf5jNqOiTu1yS/nfJEQ94CIpuFdGE20643/BHz
ZJnxJkvAEQeuH7yTvPiGUMoCCxR+u/YSCM/3c0E1vJvG7YMl6ouX+LZl3qxyuUI7
lYjtgOBcm65qPUX9VDuJG/LxrjWIeVumppklq+Tv3/qh7yfSndBaAXJM1U7ZpJ7T
pZfP1pGwoJJyHLZ9hrIwBZppevH9rgTfIb0NEoiZ8aYGl3S5iYuGaQMZGzu5l4dK
djG8GbaaJJuj73Tlw11V1Peljqex6U2kRWM+Zf1E+7U2zUhVSt7VzENnYC5h5sl6
lPQUB4JVZ41eweaL4acKYruJVDA47f2oUCJcqEdAPrDlvgewTU0JB42Mtqn8qjOW
bkMpyzGxYGOZPrLb4dnqdA/wV4PTwnhjI5uYE3hqVbHF67Y7BrLAbPHm/Cr8z70u
Y/d52JAa57/Y9pmVV06VAOrx0t6cxlkZvC6daMYZGN9b+ACRVxl8hYSkU2fQ2inn
3lkYo75AvWbhEXTGkREOrVqiMNjrAImCGoqhrmp6Q6KWtZ2pTP67LDnJAjCs9oBl
4KsZ/U8YgWHJZbkoFXPzxnK75hK6QciG8spqfYv+ZT2H8lKTgfPrS5f1o51br6Ae
sunTxOqqSKuzDq0KA6OAQB+fJt4smAsc0D9NsWJgObRzM8gv/Kn7XBjRvv01kWdY
MESfHkz9u+EbW+11PFv+YkwgLy3EbVGhFtHm4NnInJsdYk5TPXf8EW5ZCDdkVom2
Ri3QpxXRJrbQ9hQNH/ZHD2vQxVRCFmXcSWV7Um4ZOmgsgPg7fQMcd73CYIz0jtw8
eruGyXlXkEMFWOnbjb8x8SEvt8uDSLFCJdiqJr1obfjpgGvAWhYDdrR8DKwymtJG
JDNPEIGzKCtoVHdimSZ3ZHTHV5BAbvwq+KLwL1/LRY65EWj43SWwvURJXu1DIaMf
buHAMm3295xvTvrOww4rMDrw8lJUf1OgoI+SfcLGH/DEmNOS6/LDsIowJwUL+crY
MetTygykUmbwsv2ZtrD4XcoRhCCWWIWxKW7HIoS7s8yCPDRDdjZzJmlcfqmxofhG
ZZU3L04XsVUFMbTppKy53Z8mfMFtOMTrJZFt19uE8Npsf5xoOPRXE6PHwHV8zqo5
ZxOUlA7gRUBUj0W18p/CSJRV2Ku5UHjNootNlozraKIUOBsPx54XCHQLqtg0NCVN
nAoi1y4qMdhkHAaJX1hD6/CnhB5qSesfxzkgaYtBfO5+FMLBK+eQ2AjNT5uxIkiZ
w42JSkePelTZWqwfMzYU572+hAe06uj5Nj1KCef6Dw1wu/y7IRMDGPp3grV+aFtY
SawWJLCZQRvtpYLLwBufGIai4gc9vynzzALrl2e9Ih9UvY42jCmVJsI8MU4l0glA
0/wj0vprycVy8l75o9bHy/TDd1SeQCGoEw3WPzXO9zajT7e3hiEUSdExHecuHXks
D+7JiXrrS2GpHUpFoYRIwyvjQRqOc9Mc1IhsPj0LSQb0PqJcWDwn3QM7FBl6tsu6
nX+MlFmORj9e2pW5rYx+ACroLr9uxDYXO5y4ElWdEmh4xL7cnQDIWDTmYy0mA0wf
W0C4eXkv6dnjPfVwh8/BKqwywSzPzW+8A5dZ7hiPZgBfB89FxmLALkzXAr7s5+41
+zHggzImgRqujSk89MgWzBVxHRGpltaQvX46bLpN/LXFXLjrzgriyfdYeQnhQxXc
DTGiXqiExGlByK4FTlEUojMwzgYtnfjgG+9zdo8WeqABKF08wa+uwugWMlGO9pAy
3C1xruqdFELuWuD2MUiltzohO/bBlXE6C/dbWSy15ecvtErXGGD3mlE5yOeJ4dJ/
4/ksMLML0T056RxkbEgzHPWiTNpRs2ov28GALDaEq4IbD3qXVmJCZXf6Xderi+Ag
iDtonwcWaCovwrTYfwLgBHkPDHh0FfUzIwsHRDepxnHnN50bOIEEx1xDaVLtI/1Y
G68q1wxd1JEBxVQ/FeqACfRg2WtzmKi8s0XLmumLj9j2BKmXykRS7mb9vI8bsGE+
GIS8Ukuuu9hu9V3TXKFJmtg9WU70yZlWt5/sKD7X0bAYqawbl7ICKXmfS8E+nhB7
zRCSqiN40a0Hb4xH/mLxTVa3kLJ4uFcDQBRauFo8tLdspf7G3DuLSH83TnxJfdcS
PblWLLz8l33mhY4EfpoIwJIeWmR6BPmG7tL4HYme8w89QxknW5f78C03IY/nlzDn
5SblGwTsHdGtGsmH74QAUl3jJNDgvxXr/LXdoQOOZQHXkIC8MQ1fOmTZfht/w0Ap
Rw1wpXCWnnXtg9i8TCY+htd8Pk1pIg/Xs1kRS7xUumsniCs4needjn9bQk/WB6Ul
5Xua9BLDmecGTMJ5oW2qv6NB4w8TiyFc1WeDAB07gTXcMs3j6h6yEkyytMyhYWXX
hHdqRB0G6q9HVUR7g3AnqTmDHDYGDrrpysDk0FP1TJVvSjcP9QXYLwGDiM0RpAOF
IRks+amr4erSuZMx1qj3Bs8MCTRz4S5pgW3iZLJPlNf+AuAKx5OvsNnnR+LFIFXE
QP0qnePzDcP9C9/OOd34Sj5qKHdp8I1+WacKgfF6wObXjKreZ1dAp1DimeRjVupg
OFYPzQ9U0k0gcyR6mjO1RMAnw5el7LQGo0snaYptMyebNXkosgRSSI2g4Glw8l4o
YunL5xoR5zJO+MJefUQuUKy0CHX2CuJduV+g2XJXhWMPh2emCW8cvI0EVvfGPlIG
UC2W3E4QaRsgqpW/gn3hkPzXcHqHA5ON0NiRVGfyWmgAuThu0py2WC5DdBc+UU7b
dffBN+/bOTj0bacp65tQVzIqe3sBxTOP8qGiErafa2SvT3GN1001iMZbn9afv1uf
wQtVD0no5qN2zirporcjv4eqJ0VzW6aaSERcxtMj84rn4CPksXN35HpBrXVsAz6A
e1QPN3G47jzoYgN1DkQJ9uTCNc5fPvHF/2yRN6rf8QrB6NK3LV9Dldp55MtlkOLP
rYba78ac6wP9vsbPgNaTPLIdpZq689D6kZP3vBIXz94i/TPg+YP3xyoAuLgL6mC2
j1aF1fw7VezXuOSg33HOEWeGqeDGIv5GgE+ix7Cio6w1JkxJRKwQZ3AqHoRQxlgZ
/hRXObgluy7IZUn8O4feUHtPtAqULdyaEffYqW+eAS7cMtdxnOPEIvKnH918I31l
sY4GM2/6Mmj2f1xQNHRWe7ywd2W4M9+1wHM95VS3FXtXGVAkq2VA3e1ng06N8lJE
HxbG8THCUfZLxJfjGXkqy6Jrn/zw8oJhWTZBqnYDSwujA0qggkgHxCnkQAzvNBwS
QWKxBbBiD7j4FEj3qHPXXX43M0NSjJYajCWwi07EUz+1r1YeG/e0wv0YqXArDDEj
aZKlSp1qhF9pznJTR6oGSlggZM0nUP4c+DYVRdul5/qVc8AwJrMXI5UaivLqZE0O
c7DCNm3qe1WVUfT7tndDIL/YpCSBobliVNRcuKqMv2zDWYK0my8wBvmMxmXX5BNm
cTQavh0jMPxg5wCRnN3MofKmTel7vdsLS1d9Pm2cz7cHlFFE3h/UzZxhouMqCeIq
tLwsqzM4w3BXLct9eFJpJQP4vOEq3Dj5dT1kqGAMU/rcIGIZFYFFffG8rpjh/ICb
RmKL3jiUdqLSTSXrXHwkz15G7KhT9dbfJDWBPiXUgFoQbhYHBb56QFSjymbaS2M+
qRse+wDLWYfVdF8f/dvS2kxQ8tQHrOsnVE9b+ndxNA09QAKd73+we8Qn5NXV+2Br
3lURNaUX3BBGlksfB/b1Wd+/0QWX/71YM+bkD31RCntlxtFhVZZWqX+0LSknge+7
FDDchNEfnnql0vYlv7CBOmGbV0CRMSg364IjDIk6G2haN4Urn+epNzmeBGM7q+ON
UOLCzdPxCfonM3B3Ce40h/jkxLBdUt8aLqJx9/iUU8Ys5YjpMS+vGJYXPVQf2ObD
VtyGIAHtsKWevdzcZ38Ck34RIAk8FL9OVPvW5MO5bVyiVLZy/aS8K4GCW1WsiWKM
d5rUgzhmWjOqSr0GGUnpKR1owapVp7G5Eewv/AuLGM+sGdW5PlbYAvZrI+3sk09D
YnQPIeVYFNMrBGHtShzUAgTy0bpCkqJQ8Npq+1j88TmLLENU9pqV+ykOKAcKao5r
gFExRKr2MwobuceDu0GyHwb54S061efvljm0tF1zdIt0pI1DmCd5dHWWbMV1/Mq+
1iZPB1q0GDApPve4dyEMWf7uB1PM0IWMVzBL5HzzcMzMVbmnppYrldGC6WSB90dZ
XuPSjI8NUgVv2Co1Iq8GohHNb2/QrIsm/QJUxUCmRxsRnEL+8MekqJOVAxqRZL3w
LLeBb6FI/Wqm+4isj7lQpYFPSVNpyBBuFwZ0bFu2roATINhl7+vAJu4Dl1RRP9Wu
/7iDedoF0voIBskedb8+8poC98PkvG0+aH5RRSRbBEN2piMNQ0crruyscffjSNAJ
W7NMJXMyOIpTGM3Qv2t5Sp2ohWRKPSfbTQA/RyRXeW6n46l/vgjPrM8VujmKfXd4
yyqChspltG6qrHciNUh9yf2bRdefqiyFnKNWaDHjq2Lly9U5T/+PLkzbIvFXXAJs
qDzwRUSyAOhvRHjlQ0rkPHqi6PQWgUdFkyPT9MSMnCaLZcIPwPVj3OZY44H6jlOz
HDw9oQK9nAcDvQqZRRv4XnEzENyI1zeSBZ19+upoob7lpsYG6toN94MlYASzPO0U
A8QjDeMf5tIQzYtaL+MPzi00FI3FyxuXfDxeuGCg3jOeJVmKC/pk5MOvojYevoIQ
yFxCJp8PcqiXIFNh/5rlWc5MwxLwj5Vd4mp8gsEYdD6IM4tvaC8lNLc0GyGGS2BU
yot+7dNhE1OJYen4MWSuVWhiFK/YmuwD5I9a3gtuymYN6lLgRAMO3gadVhNfGF4g
QgR5u0uj5+F/73RFR1FAF4ReAxhisoM9xxtNt81hkGX7GMQgDDUMEvzwVGVeoe9y
/IcjAlg1YmRloGu9t00hs3aO06OjhJM9PtUWkbfEAsC8OXsUUyNnP7vg3s4t4u28
h22FmIlVnyfzUeOu01bBjPLQoBDnn2oKMRDj8n/BKvZLO5hlg+3Y461J1jt6fjno
DKrzyA3Zr08ipObF9Y6BB5/1cmYrhWu0UEpBJxsjTlWb/rcwXwlzvuIYoiPhdOE9
Rqtn0qTsV3wViY7kaWn8Ptmw8lWk54PK15t/GCJtEkBimFIuC46pTIX1Cct1zShU
kAGgTgRxYA/1JV+hNckQhqQeG8YLHsJCPxu/iKRtYSeS5xZtOGrhB8Z3lZ+nWeJx
zQSs156tTuWxTWhH8DS4ikInVhYntxaoqqvhd0MKsRul6seSXLIMvsfSU5x1o1qb
EFBSt83hZfsOAezW1sBX58jU2jF3q2KE6mjrFKyWIDJBb2hGSoXL8/2sXXDTMrQS
NBGdmDN4ialfLbssiiW4hZGzl9srbwDiCVZiq0w1NGB8e2br8avwUIkrBvkW3sut
1Xx4gJ+DksoP5hIL7rAkfuzJiMgUlXcpPHdgS+m5NGs8sSHuKki5owivrnCRWQhS
7UY3HoKW0be0Uu5bLrSTBB49An3mv2t5RmsR0YIxFC0DrCROKS6wi3Kd0bWEEhUk
IIFDs0CvILObplgXf5z20m5JQ7A1nL5f+2+r8FMWYx1vQrsPppwXIHQiQ9trBagT
MtTjVJgbYOi7ZlGYuvT2j9mHuVlBNCUE19ZgoxpmxRnDGBskvc5H0vrSSiPzmabX
4qUEc8xu/uyWxQ/yHhZJINSPS0T7nyAolO3YIsy0DVwgWld/1HPsY+AljInLVPOs
/Nar+7Nd53TFtTwAaOYmwEM+GFoqcB8xrUF6eGez2kkapnWxXNoEiknAJR/m1K8i
qQXEK2ll8ah+JH0Q+X6KD+y+bO1cGz8zkrKS58iHtrAxqQDsMIyQiwDqDVweNTns
JMD3ltrhfpPU6VRWmIuv08n1VpS6uidKzhjZpQ32wXnxPa+FISPajVJRrOl+C/G/
6cwPDLQfwAQDChd/6WCF27xoJCOEzCb5CJ89taviEoY48MnFv3pEofp/DqMuFAd6
CSoI0eDltZ//DGJG/100w2sSEdGr2Vdq1fDFxwYkIzd6znwzB0pYc8sXBc/D2cou
U11DDQS0NQENOLhpbQHRxuq6BAQ/QmPfczS2He4ZGAaU9V4e/TomVAxjyKEXKgkj
iDjrkJeyODw35jgrK+2Ceh4SvKbKXJYnHRahlgaqKHAo9XqVdeY4hNJRJtAB7R0t
Gn58SDxQ8pOVfqVcswmU9nprqwwyaqkJI3/xt26+MYT1Ixm9R42mOyNocsn0F2ik
JWLrz8f0ekU8yOueJPswUzVxSe+bXG6bVar+31717lyhbVsqnaSuHjk4r0QLb1zo
YmMvqDcF6AwM/gKmN51isr8TLLI6Z44TP70q1BsQ2EaXWeChIAsa1bKTQ35I3t8e
ujP5GSGReF18om1lHBu0U2McH/6rKV0i7khpF0OHt3NGtvBeL7k62ntvX5i1hzTt
Z0V0ferDMdo2QWgIJssjC2qEEQhGCM6HPkQBd7+aAIkuj9/N1/A/gQEF9VYjyg2P
7dlEu66GIPw9u1gcfPLJwQnbcJPR1CfFLpqc36o7xaYZZHN5mvgbYlHDoVk22AYM
p9SgjphAQ442wvBx7XjHJ1Aye+95uX6KSDsuwF6gv3eZk6YUdFB9ZjmAlYicBrCD
+Rc3/FXmvGofYLQRjRVJTFUdQIkDYx2HatrbIEcsaBywhawwWkIaKnPsBtbDqBcf
oNXVImHfgUT+y2H9CcoBovT6jfZIuzKTmAcoIGjwUlA4JAbySzZhE3FL5QENiyHu
vwvNyHP26aNhWryK6RtSF2R2NLbZ7C3QfW+rmbtPauvaaXydqUo/ZKACWEQbu4i5
ntkBcT0EERtOP+7R7R/ZuHkbk0K+PRfC9t48cK6xmiPOcKbBOb1TJQ7/p0lVcts8
RXG/P0boMysLjvrRg6Y0XObngfSw5+v8RtiPnzIMSZbPVzgIbabTt3aAjcEUVokg
lzfLxZqqNIsM1+fKvZHBlsmWi776TrUBJg/EjfbTklEIjwQjFrqV+yG/0QIVevrm
fXTBOj+KtDhMdReESN3JuFL3KWr3og5PqL/wcH38degHKTJ1Li1IJGw0iZYTubQE
ber4uMnf60RIHZ9KRGQavTQR0zsiWp0Hj8NcL2vRjSRKyKv8m6Jr8HCy4mb9emSf
rEBeDhzPHk0wcE2JAM5LoWRo5i2Y1AOBuieAu7n4T75eC/OJ744GAzxovVm0PLHZ
TRfXt0AElezj4kIBjrjo8MDHTl5wMiW6qd7EIG+NupR/i9kZlVDbnuuLbh70mE/X
bdtALIiyWQnayr07GxyvsulLKG+soXn4yjN13US7IHlUIRlKgEZbk/km+HCQcjWK
Bu91/DQGoJQ01ha8aZiwHVo4/fpYDiZOA5SKpxLdF+ThGxPbELgUU59n1OQPgGdB
yfL/YN3t2J4jOKDvljsFvXFhtcLyXENKaeFBKkpugZwyBi8pHqQSS9LjY1oTMpMe
SEMUjIhJKOxSxhe0muGxF+WNMN31d1AbRc887i9rR04S2ZbzDCaN/JEW6bLVZ5cu
rq6//UD5H01G20hE4edqRuRtLZuG6E8G/+UtvqAHQmUq60C8xAlvBHt/wgNHqwEx
2i1MtogLkPwPrJy3evfkdqkVMuVo0RYCBNMXfj1oUg5SkofZVTNt3MfM/y6tLLAO
DXAVVcefUCP3xaBA7ZX4J6r1Pn6ff1E6ZYbYnPyHxX/dJRasGPTxbo/EcYvqfoYm
OdPm/v8GulCctAs6RvE5/wwxuwnwcdhDmyzojzgrSiOR4ACnuKPXOZmfU8DbA7Ab
jmqIJ3awk3NnRt7Zs+HNIlqqiY2lxH5F5A9xmVAytXX6zd8O/z/VCj6ng0Ewy31X
z54HaVwbgfDgWC/hwMrDZeXUd8hi31cMHr/MmLChxCt+Nh8hUlotSIyM3Wvr+J4V
noDCfN2G5UV/CcM/o3wRfz1l4CT5F8Br/dVAFAvbPjhg/LkzRO4m6g8FcFbIps0O
aqsT04gpd3qNmEZYwh0j8DyaUmp1bh7q36oByH5Vx9CfwZddspoRCv2wppad+0Yb
IusrJlJ9pxxC+CV8tIY2+pgW/H62sHtFqa/kesxuZPC/sRMLSIpAZzMA+CzDba5t
3mfbHbAb00Y366yryNlqVnyh+XtKbzDlGTDOBEBvH/tWMbxcuPob+SKsMHkvJUgM
NU1Azik/0FS1im5sD4Cxt12fQhrAksdeslhvl8cxmQRDT0y+R0LdlgtA92q2kw91
vpV7EO9ZDzXu02K323RDR87jy5oG/oN1Wf8y5wcSwnCl01Jp9lCeSk9GBGlifTAP
OC2hv7mUkW4tGbg9iAlP8OcTHaq8pbo0j/l2u6Lfw8FRa3T5YmiwpYCtNSYElhSo
CxeQ6dCLuRrzBCXHt6x+KF3MheS0ImwEFN1m8c0OAqyIG+QD503E69wdXaZLGaQ5
6k4NGRbDK77+RmvNjeqfszuGjWyq0c+/rGQMzc2XfAzMZSJfi+T1vWOotrX+joFx
WkbHkrX671dVD8hWuo5NrfBl2/xz5yHu702h83ARH7+95JFksJNEo7U60g50aZ7q
TsrBKGYnbE0JVNDDrCs/KKhaiesofxWx+pCBJV5atwCNuqiPJMA7yzD0qHPpU2if
ufT1PmnNV4kUhcoXbQUzdu6+HuScqKbrYV7f1Y3x2zonzCfIrNDPZVzXmuJd/At1
2xjt28ST/9FE01xwmDDc4D3DrKlYMp4rE1+VHnVvb+6Z/tGiA4+JRmcLeMezIvmn
XBtjtWwD6cd+Ya9Gde6K8Pp1zMn9EkxXnELdLGFSSeLTvp7EVVEHT73eP2GrGvX2
8zYy5EjgW5TNSLx1E52FFO7QtJ4Gz4M2OpQTQNgBR521rS5YIRU54kpgSrOUVq7r
i7X610IGC87WAqTw8Zg74CbMRd2y9aInBUMLHIrIDxCKdPE7eq5tIQg3QcYPnxr/
BrLmPLsP5LS9xh5cbz8kCkXEkCbvdcmWlOFMagIjOt0wlgJTwDbcOEkE7uHnnLbo
GfxPmBcvu8S1AQ1eeGiT3WwuLx1SyHhFZ/yh773xi2GvBC3X5CpKy0qjU3LAQgAh
Z6MJIbuZPzHVjbUlHGdi3iWguTEK8XMeAJV1GxEYTzjc8VpV1r8rebdcNz3hX7Lj
AQhvtB08XIPULO5ksv4xmm47YMLSqJ1LRIWLoCkk/plkY2dCFBxHqQsn1NiWTADT
cj5WoPb69KxTeI68oC4C3ATURH/O8AucO6fAgoovJnjBJIYOWCPPnvX7Jsl3zShK
dLomigoDqO9L6F7g8GClMjpBiD/k5w8mazJXhjatxnpl1EWINt+RL0lFNcG/tiD9
2vVYJ43+GhihTs40yQwIj7R+KGXKsc5VYsDoVsjLmQZVK7qz8RxEiKt7zeocVvmm
GRqsUA+RCEz+HgBSlOugL3i+K5MnXpQcrPTwE96YGsjAK6q8P+igBF+VOZSSD5z/
XcpEmojIldJ1GlDXVN7+0r2LGYUVhu3EvzENu2XHsbOiv3KX1mdUmbVMS5cGMvI5
GvikonXa3wWsvTthK56Ucd5pMkqBtaQSTPQ6SRJnJSoPlMq9Yi3P2mmVl8mARkBo
LDpqMLeRreiPCpL4v+arxIuYXt/dqhxTvJO4LgZPBD2qw8ijA8Ky2eqIcgwx8iQM
w53qwRaO73ERsa5iXgVxri3gpTeWmxtABeRtjJGUweEm0Kpqox2+Y3dbP3u7Kw+f
u0m/hXkarolo+avBiukSJW6zxQ8gn36G/dGdlPKm2ZyMcDzLiiDBpqqjTbn0xWO8
J1HM7KchKi98dR6io3EqoiZJ608xeW4D+wg8+LBrQ6EecymkRmamT3zEp1ZT+3Zh
PPcKoHShSJItXpF1wX5AKjwgOEFqu6ldKFvYqQLBxPsYhq8Pe+cH1u1E8AdQ/lP0
XJeQem0wby3zBD5Ca3LEjft6VIaNreKH36Z5S7xoO1Ol3geBD8K/mwOG5JWjl/aR
m4upiaAS+MCE/Vo52JNzPmRn+UBCNO96Z7ZZ6IZA8L6gtrUqp0m2zsMu2T57Crb9
wqlc90MGCMeN78cK9fwlYs9EUQ5e3LNUOwihP+xs3g22NEH+nZyna3oIWUx1v2fz
orkUNjSitBBwCQaONlfUiP+eixkyYbqDEXuvKAFTZKaf6TAQ4B9s7gzjn6K7hvvi
UUFDAoaUpScLQlriheuFv1Gr/lDx7RxJrNeFlhjR9NhcnPjzH/LDc5rifbY8UBzV
x/IUmzqRC020yxDTVr+9nzecdrsDhjzd5IwV0XjWYF2ghLEKMkzPkZmTuLccXmVt
MeMmQYPGR6DYvdKzm6QkadvlezQpoVZBCdavERWSlfup8AQKsKMeuagvB1yx8woT
2xIfDzn/3vYCYor/s5ipU5nfIqOVwP9OrUiAYmSoWBQn6xo+demZsbaZM+YSQ/Rq
miZU0GV3AYoV16YuCLm6rDuHlyVTxdA+n3m0XBuMQVEZrUOAAmarjTAOrW93X4G3
dRcrKCkPdM3xJlb8570eWN3i8oO28U+YOmDFKuEE/vQgw2IiiqdayGuNTpPX3ABU
L1lknFvQZblb0PQxd1a/A15uBy3NkexV5B2xhKpV9zwrCRxOTQTA4hodg3gUItdE
Tka6/uDZNlqAxgRX40WiBk8KBStHoeQe6fOF+fA0GLshR7s3Vlc4jlfEvREJeJ+B
P1VPDLzykiC8dF0q1FxBaQ6WMA1RgVp5pj0R2lDhRn328BM1X0zMWsCpQpV0cPZd
ZPmFwlpVrwKt2fyChjn3yN94HfnWmODSLY6FiotaQnZYIm5gdBGzvS19Q5xJbLqR
8gXP1yqO9XO4totnKCtuHTZF9zMCFSeOQrrMoOkVbbgxTOHr2TEJJF5uFGs/RwwX
TvmnXmQ9IvkB973i2i2paccg6xSRJJkCkb204ML5yjkhuut7TxKCQLHEDZIT/BIe
dnt7t4eSdZOO/scYK7bDvsUWa6UGHwh+gPDkstjdV4AMnk5L3AtnLUmL/+vxFjL/
kBjuR9HCJRuHy7bDYIN4TRl78VAkSKIXkGzRf37jDdAGHbt3HcRChwf6k6AvtN0p
EvYAiJ0bJToM9ch3TkqQFx2CpMa92s/SrXJijm9osIiRROxE8rLpzJpyT3QxisTO
EXLTbPetqHlfLg9oWzVuOkS7slXb4mRD9b0mqSLI8nm/yGy64BlCuQX/USDySrLj
rBLchpvJSoLiXAcz5vVV+FIZeQGeif/dbo323sbQfX7jY3PJmHoTCFmofG4VGiIh
7o3C9bDoTBC4GrohiT05GTDODrsb/DmovuJsyID0GWO5j090amJokOshYeHyR/Yn
kvbs9N8BtyVs+VRfzD9SfxHR53BoxBr0lJpnfos+Wc9EUsGebQrbqbptyrxa/hBZ
NKUyxkXY/em5LfA4HVtb+jc+Pqou1aSH4JBj5+V1biDyGv2OreCTVDbV9ODG8gj1
DeLo89eBNn2Zo0GEXLwLxY4Vh3UJPVPJotftTYxsEEqPmwRKmW7Af79GaAEd7P0X
YczRAOUyQj/4vlLVndL2pmiz0QEXJYZ8lzo0TRBG77DR0vuBYsl+M1boxDT9MaFE
OBqJPTOPukegXpnpdwhB5TTaRjgrXt6RaPOku8y2FxnvXL4dkWjR2EiQIMsmcSgO
LhbQC1Ml3lu1kCIOncCzgGQgxnScRwgjHa7yleGW1tamz5SmBuAuJG0qPI+hSac+
jSjN4jeuyMw1pXDu/4xRPo6oJ5i+Yh98i7VzY9mkoQdDHlfcG44F+V7zEvHSuyuZ
gVe5O7cXhcP+ZajiMXBjz0nflSKkIo1jEXk/GAWtcs16awPh6ogBYXRUS9H4lES9
94KdGAxGJrVh+b57W5VEqoNpZVqf6o+iqVA9jIV0uP8x4ZcqMV82nZVGuEgN0p1m
maEC8EsRxctmC9UqpnMex/5qhddIV4WBVTXErmnES37ZACNScJezZ3KdVlQbUNud
MYxgRXlOLGCfKfpxPVSs6p8cN++aHcCOL/yOTbO2h5kWVM4Rjn36BbvWwQMvpogR
qZQ//zLE9uzImzUmSh+3dzB5dPkApWoM3SOHKY1hZuy9jFwXMkSuCwFl3dVk4fao
EV1pQUCk8zJoafBFfUj6Yk8o6JJY86Jlu8YPKI036CmU1hKKFiPOdNVmnqq/f8YL
oXQZ8WSYj9yqIcwKMXe2dggz57uDhzYgBiRj4/R5AF0zuCU9W+RwgJkSSSQlex+z
pp54t3en0lodN9wQs7tto9joSEnk3rGVKzZ5c5YxK4gRBjXug/BN8DTPTV2jfggy
V+x0Pi+0gQm2uKRFK49i7O/X64lDV9M+usuBAg2NO7GeApjok20QQWbuF5epMB4f
2J0vpCAqDGC++5EEKDh1zXQaBZakQby7bPXNKSJY+NJsHzQJwC86i/l+oZLLABOS
2y5Ggk6PdNmxX7HV9qJMbeLMFXJEWBg4rMkui55ogypyDszJZ/EduX7EZdRsJ2bV
ArIgxdZr2H2CXon1/2RjwFuiruR5hO4hpo9c3sh9WyQpyIKGFUi6v6moKQSi1Y/V
H2v7CwKXKVPuTDNez6BGkDICo8o8ud4V9sxwMz5iktyC6gQ+1BZAZoQAHoo0GzFO
uZskK2dq4J+uj04a6T5g9e9BWTTkKcue9cRso8uuyOlcG4zghcA6hTcby6p7cOhv
34vWx4NBK/dUGUdTvbkUkOjZUYwrf02l6FlN6eK7+lLYjRBnFRsDYqEjNh5vbstv
g6onpGfVxMLSjLj8NNwcbRup4We69U17Q5nUpBeOBnTbqj2qRNjzm6H/lfvmKOJM
Z6zGVyFMVMKumereAgV3OfHGEiNemMerpb+rtesQoT1mRFoRK7wVJzKOtbDf4U1C
Cl3YejoDIsr1ykbX3CkapRFsVIwj9w66uf2LUcFk2Y8fU0XkfH0M0eyrtapASGdT
MNphZIZCXC9hUh7DCgUYCNOumcVzu6IiTa0qiOTu2xqwqd58r0JkOmwoqw4Wlq9v
ci0McY6zYF/mYtBgPMA2HcuBiCCrtVqvkCTzeksxMXeiTTVpq6Xr4hgkx2N6lizc
JGS2mw2y/ZX/dq40gBgT+d42j7FR7UWq1TJq0GmJsvmAT2d0cU4ps0w+h5Ff5UQS
wiuXMvok3VE+SDDphu+pba5CF28PG3Xh95/+9G9FUqFnelI9SGrG6HyZacMK9i5y
KNv2f82Z2sQNHnav+6o6Gn61UEfHtoYA+CPcy0N5573qvEy9Y+dCZ0L6+Z9VxG2d
uix7/LWOf9q8Nh/s/tpVQbLN6sivwDEBJGjw7LWU90unVnuOQVAkx7zgSNo6Q5Np
/Snx6hBA8jTwldj6m09a6CZ0r4Slfz/mulnUtW5iJVlleR2mdLGMYvDyEAmisSl7
kWDWx7i40mZYNd+C2SEvKM0DUjEHbgOrgiFqKQ60mrFqLUChdiMoa83eaAXfbN34
UBcwrNdbf71Bf2hQK7jEF+9xbP4gO+rGnz3NXtOYObT5dW9d8EGJkcOsRMgbRST9
nVjlMgh/SSi+j13MA3cY7zNd8Km0VEcpY/g/pt3YkJ1gfQuW0rarkbZyYwQI45NP
EKY+dOnM1dx+QUErr3wtCc79xGroForkzasbJd3EYP15JA7g4X9biaBtQuBf+NWu
CfWHJvivq0yVjnKOCnqjtm5QBFhUZg6En0ccsqfxDBT0jyT8s0MXAMN0hZG5QQoc
S5MefTuiDq694kFrYJaZtEGF4vOFvlMkUggBwLFMDG8r8i8CXOOHmnpVI9VTgV03
y0O7X6AFrp4YxLHiSDQzNUv4+rKchpHlwmxt3RqhroqkH0UwynbJx0VI4sO7s0s4
UJjrNbQpb1Ql8raIgMevSLsGQqwmvQy2D2ZQCUJOcqDh3mzRPbs02s9jVMVo5cDg
8N3GWfg488+ArrrLdj3WxIP/3o9z47WMM6lcYE5BcxrirOB6BMQkYftybjeC/nTf
2pTd2XMF3cAxn3VE8K0yGzR1SqNQudn1zsSe+CNxpcrtmnn9R/hJQXli2mOYY8i3
P9y2yoc+cqaj+VPflAy0bW81t1OmcNK3tahSvLJpg24bJc6BGTJoRrbOLNjdwdO7
Wds7TG4vh199qJxhkJifIb3XlLo8Z4ElZvkNzlBJ9C6nq1uUFfqy7Of2g5qTd0KW
QVz4C1CU+SmVwJMXi1ESwuPmoS4GR6Qqf24cHIbXfzxAY4FpNVbMudERSskHX2gG
wGzfauCo2NplGgLI1fHRufLlfPw7f4k8knrmbwY3addBh9JjWMSmhf7LG8hwyjQN
xn20PDs67cK0eN3eNriAPBiB36b7lRvjg5v7/+5gMTmyWQQEkn/Oz4ZcQyDFzzxY
PaSUSKDlrIUGfyPbBu+ILosrX42u5euqJm6y1WfLtdmFWZ7nqU+rnL4NjCwflel0
SSoLENUjqKNJwxVRVHFjnSwIYJDXKzvIO9Ec6JDxYCuWn3qG0cZKswFBlOklUnxp
O5acqZW+mQWV6yYEWt6rerDJ11r0tjQJs0I2m74ReYwJxIsv6DXzyvctH92tGVP4
Geof9PAFnimQ+oglhHxLbYyZZTv6m0Hkal4E52lOABLUk3DGi7IbI+4GPWz8PZwP
nU0cJPAc6kcDjYgHjHPhojEETbX5F+zv7dLBYgixx+m7D5OrRQ/nzlq8uaN+LxHD
I6Jeg2PNXGioPQBDXXlrLt4CYXgF7OZ4XtI8JtcXvsBfZZgm0j8HjMSkfrEoybvl
ie3wjb8fTurlDjlcNbRmQx+kx6gaAUgbHy8a1aJtuiFfwv0kXpZINJya2RV8FiGY
5L1PYaxAsVjunXre83GzyWacBdwCmqDiBbCghXhLrrOQhdGVYqKKm57XQaKhVJEJ
KH0aWHoeLSZNQjGthl/yasf0qszkkPpwV3R55QkkmTu+2b44DEPnml+5HOCi3v9L
sMBFW6JzC0a/DwQC63uvV5DRtzJdX9d+W0iwYvcANQHLlOzHPMHMP18Zd7Avgfy2
K8wdi4QIOZRi0NJTvM+1cDugVdU8ivAcGBdRt/L92YVkmSHrHevB/m4iVzTOggPX
Z8vpOHNyaECUVGWPxpMHN3WApRzw9q8xTR/zWGoLNOOG5ufMXRx2Dvp4zUZDWnnP
mGHT4WTtXiduoi1iImFQX6Zuc3mupwO7Dw5Gvqmt3DHRRYT94X1QlN/jOrZjXYJs
hF0IeSwt4ZARlIsXRcruhR6BkxqadywiGAbQdjvRPEKBXJUZLOyzOfeFnlIdcGBZ
v6az3Rchdm8SJExusIsmWIwdKZDXwRjf1khKgVrU2TaveViL5EOvZ2BYUqBNKa/P
QVTZeNB4Rrqq/cA049QZUO1808zQrDYR+PeXqlP+z+B3FG1Nrl+RB83LfCFMB+eE
4w0k4Rys3orDkXcpHkY7WQ6Q0KfPQgtO/vhvO2WqHvV6g20QltOz5OF5Kw43mNn+
AvFvDGgU50KsyhUuwxU2a6P0ITev7lbysRQ2BHPrOpbjMbzklvG07RK8rvaeDSFk
Pd2qHszJYRFVazV6UQ3GD6aK39qXL1G8OoRFgu3uqBmuh43qX7ys1JweFpcpe5k4
8Dmh8D1RWbd7Lw73RutvgqKzFl9LGrLYl3hiqWAUBUIDBTJnM/9enm9CEzUsLW6/
Nh1NpJ78PfDmS6Fc1UOTPEfdy+qzD4D1DiQUTYBaCgWMe6YFfgiRUox/r7Zczetn
DLGFLWlqvmCUoak6r/qQIB6pJRAHN379/ozTmz2sB5+h5TrLj+n64NYNbvK/kp1h
+wzM+qtd60yJ4XoppX7eTfDStVjmBpmNXybe6DHIwYdINQYaTaqdowpWMSa21/hB
ecRTpA9XPUkacWlIc8VwYEHYvktIASYW9xfHV1+hPfO6PzkOSTyde8FG7ld4qApJ
s7HWJn+6PzODsPITJ44re2fOZID+HjOsmzqCDTgsHfHImfpXcAi0iP9pPmbsDMnI
r6NkMxjYdyz8xx150P+zKuYp3anug+nIh50idV0LHcl2LcZAGY7nVbkHfmHYUW9N
w7l+bJQbeH6qhwlnUrldygE8RR6F6Y04KBsmr49CGknJoBVJlL+Zfm0ulceieGld
6kqjC3uu0X53pswuCScLc2Fwrie+SZYQpNsideAmI1Iq5FKJxcFTNfWCHMwkHhFy
y9P04W2mb75Si0gywk4HWI2eBnbC6MuKVPUQmfn2nXLCV7+t/m22bbJpy/4YXt9E
sDMlgG9NPN8O6Si7RRqe2BGbPotwo38AqQ9oyt+GveivYBJr4WopPbh0Aa13hAAT
1BKZ7V7Wn6mVWjv5wqjb/MyhYuj/dUVb3ikJmCmBkLs7aKzmPBM8w5cqNsiNrzSz
776o6ryTu6qaAMH3tuOilVXziQAGusmNZ+jgaq9MvR9PVSKibiaSdzdoDM7sXVsB
rALP8FI6lBA5z9HdiLHy2POBUuFrWhn0FbBayf4eKZO9WM16M4YHr+jcepnaZP7M
nx8Kr5UhHUHIBlRwi96TcCKMYTbVakC5sbArlSU3FbINPnwrHiinoj7CIWBSrTZc
tyMH4lB0ZWamN0ksTozCAkbNU/Wi/otxgtaOlN7w1NVEvIuov7dQsi06Wthy/jrU
IyyITWRVQLw+uONVWR3JwC5bMGQ+8uTu4u0pYiKpOJus9J0EaqBpAYLdOsarbI1x
jsI9oFEFgwqadowQfT6j5tpUZNlc/+8usqxk/IyJNM/le8RqRQRW303WsgIStgwC
aH78jIyvv3K0K6R28lfBChxjLJJjs6nq03/3p4nWbEAc+dqVPwEMBCRRuM4w/k7y
tGSEhrZCYIYelmoVphze2GYCtoQ2+U1TUxn7pPEK8jloDnvCwtQxZ2cRFNfpUMYQ
2LVpUX+bC7y2/UD5zYzsMTmJGBQUG/kNNr90FSsnZ80I85Ux6uJsATueQvvuyrUP
/Qo2oQQJGDFXzb968khUXyijlUvOEcrYL5oh1PtL7bsYdZ7jj6y4vs2YguVzEX8q
O5JtLleRHLJpZXTtYmMss049VhCR4syZFOVIoFCI+nWcIJXwWVhE+wfqcpr6CsqA
zVqKtU1RlnCjUa4jk6drT3/Bo7tQzcGQ3JK71oqpuJ4+RkwgRXYSeA7gewMW0jsc
Sp0h27SPqYWotXXdcedfr2nXJWOrischQEXx1lZlPQx/WXu8RYcsLP2Qx+UDSbWA
zcQPOUkpJE0zXfbavSZY8V4yJ7aHG2JhD/HL8eeCXlaP250PaAXBMH85AgiVsftq
O1mm1AgTA2EYFl00o4JniP99fpoENqY6tF1DcLT2GNZCjKtZHFbEs8e3BaLsZej7
jJvlx1zRnmneUjEt/SD+/WvVLJVArWrBi3REMuNGFOK+gKouxorGSJMJRJXMhHAa
ZAmUkx0BY9ZfwOM/Yq0G8MdL6VvQ4UldtkDTIGCsA+EqoBxc5eQfjIh0MbXGK2bT
/U9I49IGrmbgdkJP6OdOLiFZdHYoZN9xf+CSgpjm8iMpIvw4c/6hokONkxc1D9+R
ixNekc6Be5d+DiDjeyi7GPSI1IBuM6QfNxYPiGdiGY7TzILhLfEflI+GLAPjoS7e
ua7XemhOjlAvajtGzrHFmEytAXAtglZ7/GaAVuVSgPFI6SN7gFZvYM6J5kQ1Z82k
sJoe4O1s/0nlmKbrnKUtFMS0Vnj0lrlVh6lHdlRwF4ygcpXQpj/EF6AexYia5xk8
XsIuiOrZ1io1BytT8gcGcm+tsxqRJ86DwrgqOF69OxTFcyB3ls5dZj/7pxKBi4C6
RQm/kIdbKuYFNp60J4D4y09z6u8A2OsngV8KJYti9Tb5RGQ3zhcDCmzp2Al/xVaa
kWpeBfE212uTxsrzswl8YlgqC3PaFaQ6/eEgEV8E/i0TZOd8KbziPQXDge7U89GY
rgF6f+pBCMLOXDsGmP40COt1VlSMBcd5FGugWtER4sqCr92Y4oHmncVT0yjEeD6x
Mm7BgzhMJnqcG9/miaPYpMSojU5BIAqtwxBrpN/ATzS0P++WdNaCaGYc6Rkb7Xnu
xoJCJqqjvxDPfxvPEVqpC7CcyEubOIas8hpihPuDsGhdDxW4jW+fuYk3Y8GiCIso
NlnwYvUXWp5KAgwYTaAxzC+W/6gPmSlcQzNdiBvxdi2b6ebidA0++Nw8hLqfUFH5
2E6xhpI6CGe+/RXuP4+g3t0njlMFCVe3N9Jhue6gumLOlWtQXK3y2mMOcpX5V32A
T0GPoH9vDZzWWgS8J2Kkgj6khyPnEla9wZ4uSUwJaVro9GiAEyo92ICTp/SOEiM6
G7SyiVRdi2sSolUjfNR8uGyXsoEATTt5uWiwkps8qKJ4qLSUNdqprm9H0aHE8ZvD
ubB+rZLLNHA4lFU5BRaDIFyREuoEgzqjOBu8Dsbx75kCb5aDdXgUUbDrl4DTP7OT
6yvvz1pCVsDkimiQlc5I3ixEJ2FBz/qgZ9UuF+cqbeEh+vgBWClUVjxxI5lSYTwL
9hvRx3coEQPLQFqoYF2aDqOFIED69MP4pf+/We9QMh+BNCnPLXQSpndOO0U7JnH4
Q4BftSY+T5nlY+Lp3FRc+bgBXnTweJwx+WX6bqaB6rsPmo35xE49eYZTQchkN9yE
OxPKo+aSROZkkcSkWqoiUcCEC1Xu3d2wGNdXaO60SKLAEEh27C3aejO9RGzPp/8s
t6iylSNsxfp+sSGxCZnDU2gpuql9Mp/immcID3T4kprBawMhVwpbuJy7QvKRLqrV
WBWeLsgpr9Kbs+c94jk90Z6n2EOt1uRgTGBEQ9vbijjAWQ74a/fEFe7F7YIzimFp
lBKM4M9UkTKuqmKB0wKy/81Qn1RvJKCj6Ubf3WZXnItmU0LkC2Vk3UM60pDlktVN
mTm4tCnr3FhOVtbzAEq9r94ghxep+bJTfaD0eju1aqDRdIM1p9Zw+ZUHK4I0PXS9
qgjqVZ5dQG14OCpt3Ufw1egLFrzhzQxc1W8skckdiJooY7XLV7ZFaE3mSBCXB9OZ
thPRbQcegtwh2wN6sKRPSzzTPA16K7BSgq7GRQOsmCC0CsrYRiryjVmfWWy45qf1
GAG9vJ8Yw7qwBrdYiNyPRq+v3E5yoUabQVUsvTKWG0oDFbHKgOPHHQ6ze29qndBr
D7fjxiO2CJ7w6l3Z7e1XwUe88z7r4pEck+3LzP9O6q1nCM80NOsU+63ZuJfd5FkJ
aT+eRZdBMGFJ1dhmujMr39O0pzwJi3dZ41I7u+ZE9+AasqbOwJE0uEK8UbxoJFwn
/8KJcd1MQTmqDCwl6D0aVezYcLEUsxF20PSao0FHUdBUNa3ypCdqkaXRuYpKCje1
8PvN9noFRaqUQ9xu2m4JI7e6YpsVehPohGgbbfag4CRusHYYoq20jFY1iIX/j2YG
71TxgozQahxcxm+77PiyrdG4wV9+CGik8uxUDukqP3xHKA42jODmuQ26JzenABzp
DmDpiQ/D2U/iXs0j0tpGI8urrc4ItXEgl8kIGwEd3Nnq8Pr68scd4GJD9gEaIvcB
VyIsuWik4pRMO0wokvTCyaUq0YZzyZO3U6QONhMG7LFStmxKXoWpWBkzuSw6llGu
gS0TSL3m5AS8FXsmNUN+n2FaNuglIK2ybo5f/Df5LjdogtqK2E/1/N5OqYYQtMA8
M0bII6ciGDufFrylYK6hQUWJ66vdipYEHqhN1aWiJUnLOWnWpU13oO7mfFr9IiVT
eIu6bfj5t+zKmCuyxye/nz57LzTZUkqxGKigrIL6+9++UdhRYp51h1J4tOifyCh8
Xi0ZIm/bDMg4ee7p6TP3m+fK+wNft+wr3M/Fo6gIVz/kXjjyiU/I9yFLqgeLOK+8
o03mtUU/taYUvDdyzh/eeHnIDIZyEFe08qAqHSRtgP7a9Y7YXRuwizMGIKFC9evK
wkVvTGOW1H5/4Nfjabnbo8DwDSEUShQzz90mT/V5MC/drbkJ2ktJJZKOZfawTjEA
QeOQLsoFPJq9yVkc34BQXQXmKECwqeE7w8MrWFvOlrGzupuXXg6SiqqU3INsFReK
MYkmVuQEOZy3KxcfJGZZE6jbnXwaFTwuHhJT/oeYSJGTG7sb4vTp3MszGNKy5hU9
M8dE5OCRR75gX1j+OMVl3aMnkvM/XK0gMBpPl2XhUenmEVaHu9AIPNAYnAgOYt8C
byxCAg9URbC1XJH/XiNKIBiaa2dbIkqpOm27lSaVGy+D+/20gdwStJsz2bJ3k6jg
DPFlxTA+8hGYmaSSCI4kXzK3HLtXetdsGJpBf+meGTIbJ7727mf+1f1AsX9N8dKF
jVWDPLcU42xkHDq+1t5TjVoZ/fNxpagQCKE1L2WsRujWuqInGQFGRL6JfSh17Nld
B7A7X5cHFpLPFpm9Q4aHXt6MvTb90XG+M2sP/VPKz8upM3+kxZDeEpBGwUeBLrsV
4I+KX0TWcsOhC+Qm2m06cL+1QrQP0AyNwj8urn/pcGmQ3OHIwUMDjWu5lXAMh3dv
3TwWBaRfi2cXHbS05M+a5d9XCDc7m6/ASBci5fxNIyblgm7NMUsvibIm4g+SAFwq
N6tuvcwPpd9rY55dMgi93jrLQYmJu2adhl61+2uxNUd0gJ0f8cMhf6/gVrx9+7Aa
mPn2/0koBGy+7wn8WWqq1EUPy7Sy2gH8I6NKY62cvzqoBRCwiW5CB/BmM99IfMSA
ieWJR7u/Du0G2P2osAlftwj1YykgSvzHVhcCyCqcHxvC+qQ0L1tEuShysCex/vky
XKiIt0Kqxq/fV1vcA2kxklspn1XbAocJUm8kZjXIMjoRBngpHp8k0vSCkwGPZCQc
nOpsGzJN4uuJWHGyPq92G9vSidut0Hs15i+ueKHu3NN+KlwhFN8YL4YddcZ8wsEf
zQdqLmmxDSXT7TBOPq1SeD2q4dcQx8s0arn+Pmfv8V8fOTvYNioy0VokE+2yBOqz
JZ5gax3IMEMbf6LKjM7kUUmLGoNLNTSXit3rhq3sqIyql1hunMu4gsnoRLi5Pwvh
UJDJmlimLr2ptSafAWmktEaD1xKVDSf0WAQrGumtvPHJXkRzYm5KlkMmd4qrscth
nB+cVgiKpxl6DDteHtzDzK267nRq+IpevaEZsFHAc6e43uMwSD9+4v8Cy0kPZpbK
FKJznKv0cZuBehxItkOjGDA55hQHyG/npQmWOXm8RHgLloQ0hCOww3Hwx17145zC
SubLdzFM9gq/t+c157Tcdhnide48b4Bh51PsB+HB29gUULXhhabLtR/o9SymuFZd
uPOzaZ8fsirr5X/Sljlc6HWVBNbjoWlQrCxM9Jum6pSP8D0XOGKveqL9kIyT2r+q
Qfqjln6TnrzLxzoVfDN/W94zqud3QMfLCOCPjAd8qvYeMohrpJy8h+HigkjkmzEN
hPulTMOVTaeDTEkbKVlqjMWQ0uPLdqYlvxRljeYKYmdeHHbTx0egLOAhNnxTKxZL
S+F1jzjwLnS1wBLTQlHt9sAsf0C9qQC5ZEZ6Vz6Pc4Qn71SxXZa8mYBxF9nXijmq
A3+W0jDeV/x5PaRIq+/br8KfYJb9Tr3N2YLFN9ScvJE7zXP6OPWQPA573tpb1Znr
hLPXDw0Pxt2zXbcL0Kob0gXIlS0XoJigOLJIriYtzbLdm7IfAynyix2OXnpDO8oP
hq6do2aKKujZVEQzO+8d0AH5Zx/QrhqpegG5iMXRhEZjzJRhGumtpbPWhHdW6cqK
3YyxgSg++LhFD8m1tKzDC6vUADn/a2lfO4aaw519DAokgPqYKMf2+M+fOYtioH4c
Pe6XgMHbp/UPqIio2CojTYk2qaAIo+wHLPtqHv7HEvPAj1hKGqFfgjs1bZTiz+mW
W2ZhQf6KZ2sFPHI3PMCfXf2gvw32ZQzdxg4MqLL8oYQW56LS3VMRAdB3CzvyvKOh
j0dbaiDcWSfOtJmtSi5kVBz5IUXoPj7FKM48tMSHw+zrwmgY8GK1QoiBr0ad4c3w
pSf3p7H3w+HUpORTTYmk5kQ6eb4WvUg2HI9PbTTZyC/OlejWbYm5JGKsvWzCLmJV
Ym21WzTHIMjJfPnNesWMsLPKoquTiHkXKtBdvKHNi7lJDr+POlxzW4n0SsU13y5s
bGeW1nLwuQQaSBZ9DaQLm48nZm9nYQC/E2WwYJuvlh2ZmahfF1CjF44G4Wr1ZDqR
C2ssNDFMOg37uQSwAJ1tfpwDvPF90EmnmtQ9hzVctKKXdjG5idBPLTB+vesSU8gd
othzB+3g5MwdlvxuNoupOGoVm6UcCMblDI+xGO3E3f+lO9nFgawL8VYqFa9ydq3U
BsJm3XZ93bHAEBBwdAIenkBA2aGAWTw0vmNjofs2reTp+/ki8QoK8ZQv8Px8MQJo
jfHGl5cROwpjEE3NgayUD4MOVeawBZgi2XEBxclHfwqIruujQ8tkNFTqY/gm3Kjh
6ZOiYDYe9u9BY4b0HOKmgTEcHgfNTAarXsZGQDKMOD5MUg6wWJdllF3xaAE0nEwr
k1tsZsKJLGQKNlXTQnfSdhukkuU+NmCrqcuzJ7QaOdh3awLfHbx0zKay/Mg1NbE6
rKuGs3l5mYOSprekTMCDEL83VpDRRuH1ul97X4RGexhu+HRb2WUOOZTzU7Cxg6c+
dJTReIwxCWWS8FX26M5ovUwvP+1mPUiugU2wbFPn6/wTgVz6TcP1Li25oyWA/Xvw
BXqtKOxIzQt2Q4g7SNshqjsPBkcoDzs5rda2s4SW1R08n0yje2G40PO5exthdNqu
WlkY/5kv/iVl0MzZSrBkxXyjQ/zZs3lgDbBEjZL8IzcXhizsvI1e3rfw5Xg3Yf/f
rtWrDXgnCS0bcrB42X7SmPumUrqd+czEj9C3ugk+DJuU7YnMj3HZp8Pm6nehWSo8
VlDW2d5og1BF53zvqaWHZDAGCAnL74fqPmG7wO0fdsmC2koSwly9Ynze3rssN2qB
h1jy8CJ/DynTBhEDEHwbdNlKR4cDchsrLOKyqsnEhZ+sdfg3xLo6JkFSutEyzG6H
73qSYDGxV9i6+L3GvwDCY+v2f96uNwqYgqfuzW2ONv2c5xulZPl4krhDY488elj+
OG84qfqLLxKdXmUVdD/XShqqqJPAd8D+GmborZ5gzB1erDldzZ1/I6ZVbroVEOhc
rntmQ7QOh2jCO7F2FQsRahdHdAZN4BDAiYuK8ssD+WwSoN/sHTiRdtScw7+bsOGz
Uv6hdansjMKbyZxllXhmPFbrDu7A2cwxgL1YnE40i24S7eHl/qtFuAIJpzVnXkij
NcDRPcmmbJKKb+F/BFLsAVOZ5v3duc8S/FBZLFLwwye1/n+6kg23ji6e2Sp/wl7q
Z8Dh6EYcLeIN8r5rj2lZdk+un4R6jP6/4bc9nRqI9m+nfTLQJ7lGnNFi8ByUtKnA
bk/hUykd+9cnBY3g0/9oP2+pCIVM7LOA8e0DTDeYjVsiU4c4mdTgfJdATX5twTYz
mv+PgnJXo//pvbWcEeeE8iXwihLKEuM5lgKzzWBwwZlyJDmytp7HTSQsMciuomeC
viZ+wfCX3ppURpUk2+/BQ6eR1PPG1JDLt9lIfsLalBexqNzIhJ/o9YoU8s6cDMGE
5KsdzCT8poWE9f903+F+CaNm+F4Z/wLNL+zoTaW6A1ydtSbbfulZKKnmtRF44sE7
1oVE5cs3ativqMgDsBcmhkvjUxfs91JR/lb8xt8UF3fkmFF21oecoV7m1pxLbrG4
aAy4rAFb+zuq9cg3ZYkH9WpFH9I1MyK/2kn1KUQRL4SKbd64X2YV3tksuAJ/4yBP
GT+knmz+sxrybHYfxnYbhlUpBbQscSiZXZEMbXBpeTgdGqa/vlLB2F9IWN4QBaMH
MBBdNofZprffqRegXDmwjp8Ss/GqOQ9vS32ebZGnrIQZWbX/o+T3VpV4T6u7XLGK
dKrHhk1vHJw3Pd3mE8Io+z/lmdrP0VYLVBr+Uc63/dp6UajFrdNscAE54967B8Ql
ONwUvheDgUe1xTLHgAy1/5xR+eCE0m9UElqLyHpKvCWhaBvEy9mTSeUoLqNykPCk
sD5Ckd6m4pmvrs3gvCiiJCNAAoYo3mxrTipXF/MCn/BBJyTmtyoAvilcA57G7dvn
h3pr79Hsm0Oh2n8Kux6PMiN4TVQLRWiJcTpiabLfKY8q6WA7zleE781PqUtc3mvD
OmDo487zwlrTNsc20e6HRiunr+WRm5cLeJBJljqbuTHdOniNzPEtSqtTDjC1g0Iq
F5leKnKsxgOWUeTmcARfMFLHNa8TE/8DDV1ohTsQjmsu5SbXv/VUk15dTUcUXH8c
Ff4zg/QC/ZYZNfuXQRIzr7ECEmbK3n40ITqH8cdzmnLwjnBKWQNdt8NVjYGISbSs
xA9pj/YsB5J6/YDFy6Sb1gilWidhV69vh5GpDk+3V5DXuaP4Gq9oW7vMtCy55uhC
vAOm0HxcpW5L7svbgCPJ76+abiBtZQ4qpT0/UQtC386ejOv4xOabl1gzVdgQhiu9
dHgGXsh+zE8EdKcyUWWJgaOPycrq8R2e0kv+LEkvsnmgVcpswTfHj+7lS9kpegsk
QDxE7nrBhU16h4hi/qcf6xJL6zN9B8Zgc0OndKSkOQE9BPZY/FJsQUifivbWtAv3
DpW1sZSkPyFUDSBP67J10x2WJlKIgl9SoBvGabx/wEQ09Sr+aDeCR0U6WfAYMueA
xCULM9qMuj9IAinCOMlchJ5UAg6eYkKOjVI4Zu4QTi7UX9TylYon8WD13CQ+m9Qt
c0R1y8WEuKHVq2xvqW7GqXhCZqGj/vkP8SmMdKbWNSIZfjfwe+NRhD0HqVoH30Bn
r6/sgh5PRfJQtHo4BZLX6/V2wvls7PFKV96g/eh4n6KDoZycxUxP5PrZcxOsyirA
GH3rs/DN0bfnX8/bTrxp8Ete3JVPWr81XE5npHt1lgR4DY3VVRYfv8hhvh39nkib
KLdCjnTADKMWkMV1IKgYUavE4lZPziTsbV7MbYZ6LMkEJWBGL2RBQ1NunBse0mTn
3PEcWWBeMSdwGhz9ZGz+veiRA0hn0ZTlGcxxqGF5o7DVvopOFwXIXr912ZMP+ZKp
alIOQ+tENzLDvbAlySjniOxcJImZB+BeOqbBxEIcocofmrOyuTsd4jXvoo6qx0dm
J9EMpgXM1baMVhEGVgcWMl1WTEoPV3DS0Q/iIJ7lII+smyTO+Knns3GJU/8IiEfP
TtMmeEcaNw2mL60rEcZlqFOGD8LY31Omw78GqClUok4Iyd2VR1BE4w6nXjWEK9g3
UkjQKoRamVMrSwaq4PdVf/x5LXESA0O3tAGz/GkeXmFRk0NrkdN5gmBdZ2N81HUm
vtZNzlW8EESySvaI5+FtHYLv5/DAI//hiNkC+4kbd9FRBsPaxD3sm2eqk3rIVjmy
ftoBLPc4KInRdcx7yD/itKKPQpHX5iratHCDDcDxQH0Q7zm2MbVZoQHuuK5sDqrs
jiv7q152hhaBOJac8cNe1NiWls5kCIwEQq9VWDM02eW+OhU4PDq2sh64bVymtjUf
nMDes+p51luZsJu4xRKUQMvbNh87iWBKnTNAyfEIfNN95qe00gMoI4KDzuio1R8v
hN76U3R1vkq/gMaHw7zLUxB/7t41xN/DKYHVOJRCVzOgsx0A9Qy1mts+rQwq3NjC
eyfGRAHcoO1KfyzyjMBBnEOXpFq8TjBLuVt3AQpiV22/K43IKUuyIM5E1ayija7H
Ye3cNm7kbO88BKR58vYSzAAnjJHBdmlJMkQbatEh9BIPv/ARBguXWJT3axLMxPs1
QQUzqNsCzwdEpQIoDDdGspcdIp7PO88n3AFVGoYZ3e8OaJ6gHcYLGZQDHOxg5hlE
rblramy65qu/Xb10Hlabx9G6CBfOmUVluwoJrHfXrfbIivs6yIIDThvzDvM4shEU
os52VrJSN8QRLmxFZgqsNTw3uH9cP90dSRetR1ULyqsaWKfTplJHQx4Ek+aeNDhD
N05YZDmlI75mnDP7bzaOV6tIIcAJAo0Rjyl3zPkOXvZcPkyROZcnAdrGSPLS8buN
OO+i2OelP+dTaGxsiLCpHv+RKY4NibgwfnVMmkBuy0lU7Rn2GO8ONxsOBqPY0zvD
d5oFjVCRfiNLP8PpujnSJNRiUqXWy7fgiMWSUKB3o8RCZ5SqchtiH34OtWcis6ck
cRgtv3d9oKweGTuVQYIFz2TUuqfyA5/mGxaBqpf6ureI7l0t2BNzQ4qtsyE0bTx6
Mh5cwfAiTwcbTtGcpSbzPYPmn7riCGhc5Bm5B/63JSb2aZEDdgcbDcuhFBFbhej+
qQADxLue5EZF4HvaogQvHD5+z+t5Sy7NcAVVwHi4A1rdT0ws9NsXoEvTZz//KswE
w63umTBwOM+VvrkgcizpQBpRSjJu3eomPjDp/Bc+mMtDQNAS//6alDy3qHXQfB8p
rLPhJWK1xQ2V8mHwi9qlm+zYRFbjK4FjuM1fa5F+1BKvZs8SLoZjNxX4PF2Bh0eX
aDtAw/xk7XfpEWm1gvrUDcwgT6bGsig1NnxfmU5ysmJPaCiVwth7QFbmPUM86LR8
tiKdStI7leR5H5x1DWTyYeWpK30H3CDC1j92gXpxor3M/ct776nFls8C1C7WK7/z
2t/ZlAeLIUhvKTuUFwkqRxPMQ5vZdLksz4Ch63H2ZA+HJTWmcoCbPtJG2U3L0jc2
nFe7Rx2lwwOWVOAefcwqfAsqoCCjat40iR43BWrw/ojBa13ewrSRDFTl++/FFpIl
ABaS/rE/gS3oR2FRvqhPRY5TbfrThdjG6+Z+ccEiqLSGNFwrc6ymqkMIuxguv6vk
KxbBt+Dv4Qqh2rFo1+zQJFteWRhRKkYtvcpwTw3vyfI4Sfhie6V2+ncpXpGKgvVv
h6rAMnF1tp8RJ41gqz9zTyn98neEJF1twem0ezjmWkor8FY1n3Uw3AkaULiPiZM/
y9B+xRxslCyWe9WSXaCWm3PGrbfRwAFkOpAWgOff4kHYruTna3nvwIBsVUVBfdCu
sZO0XVeV3TtGTjAUaDULG52x+rxNTlMoSiZ7gRscFegD8mHVSxMdf1/MNwo31DuS
4EhatW3/1ydRbLmmHiAdiZuU9+Sv69qDt157ho7MNfg4h8ODBxna5EKKkGmk60MO
Mhlv/rwMYU09PxgqgI83Dg6/KFCUHWE1ng7FBukVIOH97Vn4hCon4sUBbC/zJMQI
EtcgLDSD7eOGP91VFrkXM7V/zNZmX6qif507QuPukGxqy5GFJlTvmIiSjo2dU3Hn
leLI73RBaxMVRR9MbO6qX3vrVa2Xf9UFkz9WiWD1fVKwVIXX9AFrQY1eHwsuxfWe
hXCRLAlHUJQm9fzK54G8PMLK4/aPy+iC+ziD2S80Hft46SVSdbdVd4GWwQwXBKrs
1EZ4cNaTz60qIpUq4sBe3/sNO5bLmNYLJ7nvzZ5RgBP7QcmOdI5uiVaj7mfoibhL
rdLULJh4UABL8hAWJfrsBETiNTI2xsXWQUOocX9YaWkOYsjvaRU5tvUi8Q+y44qX
VTTVUc21ilsn9k0Icom1GTr8w0dAg18mUG0Y+u00tCICvCxLl0UV5hVCohlmI5EK
C/QnVhFplYIWFIrzvOTO/98PtduJPsKkAHGhgBhmXBKP9j/Erbq4aOmcgba5MLYy
dCPrsS3tqUK9RYdRDh2BS4rHDoFmqIn/y5o/52D3qEVJ4qG+TtL954vmajMpxmuU
UeE6xmq8jJ1KuVYJmTy5Z3my8obGNJRuPZpgsezKJi0sTvAMbQV0uvAAzU13BDI6
0vMEt8qDiyjJCcLuaTdD577b842vW4pC40eSzJnRXI0T74oY7rOvQsdfO79U1i5v
wNeW3B0kWG6nv3RDPpeEMf2edSEHCqAela4JrItLrrpBe5WoTxgg2GkwRBXXagWR
iG3Njfk5cTIwl583LcUWHSQcO/40P/iVZw0NCz6pznNQtaU0nfbCvSQVHD/LeWJ/
nouP/b/2Z4TWdTfKs4q38nPq47A5xdxYe0BTRYUNXK8Z+zKL0dfQm/aRq7BvyfSI
WEaVXchUUi76E7BmtLjp4ivSISxJ+uQWyrRHD/+2fEkt/so06aHkZ7DKcPOWseRZ
HR2jA1PhVcSohZlB3QThhDIFuIxCvRpflNgSlXuBJk/5GM/BFq6haSaQ+PepjQ+K
UqnOQutBxqZ2m2OOjiRBlC1KrCaYYViWtFESelRdbl78djdxY6gyyENysOUW5iFH
ClPIg5a9+DhmXfgM9fQxE9c+TZtQzw7rh5yqPfPg789wnm6E/2YK2xX57tR8PX1f
tAW6h5n5QXFKZCJHmQTKQkPLnmsSk850TS72tjOsYBwbiGSOoSP1gubhlwFNWw+i
fboF5m/iSLnHOKQfz1PRNf2NImbJoMNowg4vpzPjIU3jKbZr7Ak1HuQfKlfl8Ptg
5NW5LcAvg+rkpoiHgLNxXCRez1byD/8/Z7rx8+5uvWmHjwWUAY63gzWUlBg0FLas
LBR4ml8gG/lKsfmwphKVGVPc8Wuy2R/zk0pC1eboLtJeA+HJz2Oz93edTQXiTjE8
dGhGMBl2xUhwaYbbKe38Sli8gUii/oEJFY3fnRyNOR6elO3vOR/bwMGaoRsuF9HM
RZU28tAsPdZ0bbFfWDU+aImLWk9sZ8HmbKmocnGFymJBuRCXCJUqCk8Vqv7eVJWf
hjniCzNQ5rkbysLERtVxF3Y+2yJYqu1fUWRzWjGJzkEdrtSgDmkkBdBtrM1GmetE
VrSeFIVwg63mEVeGg0xlDgbTESbVGZ2g7AQJ1LETqfw/ZKWzVuPV0sgmHbrryWAA
bIHF1uueteWrDtij8HflrKQJHOClRvnVE63WKxGVlN6lrdQb92t2ByYTJ7cdl7Ck
Mr+SFC4aK4G3PkoSfyf4CuQ2aXpq2nNfQEwipZN76UxgZTMmkNeamtswJxpoHpZD
Z+iC24jeTVvZCZ90VaaChAh6a1SZGCzRYNZ8o3jsZzT1TyLsRbTMRx/3NhJ8dX0n
avEeU6u7DcY6j76F/yz+4RJ8uT0WuJ1xJl36W/iVihRo0s/ShpVjLpcBLqfeSeB5
nubDdXoiY9SyENn3YBvXZwVS6cnYGNOzcGPLaZBGdXufqQfjpadX11itAfYArCuA
zvLdYys0qGMbXh4m3z7kI8QRhZElk+7A5vbhCwACBD+SPzirXdYQ8VX/Vk20ZMem
qBm6tcaFOQbyoiOaOocFewkegyy/gSONGhEKmwNKVQ73jsDmyoxWeMCjBfFF9fM2
Ac80WytWkz+O/ubVzThq17O6AQsFBcFcwgvoOjjJVlrazfWhUysYb6d0o3E231/M
KCxDnligXjExR9KDW/JbbDsbtBTZpdKS8lA9qXp/sxTMOOFmzaO1HJY+HhQtXEE6
PstHCrCZVtJkOt0AbeaTOsfI9Rm8v1PNNZwP1RCTsZuBqmwSgruujf4O5FPjCpjq
07qt+o9xRGJebn0ULo4J7D51EF74TaBO+wQy64hPzFbcfLonm1vd58eE91rBVONe
jY8qu71OdRIfkdMvW3BAhWty3g2lpVbx+pUuvWk1df3ACYCmAsXVtoZkhO6lejr3
D1W5uSsz88yXwSSW/gaZz6APW4AGfsHj95WYwBVLrYr8uLakvRSnWUwUzRGVffUo
6++gJ4ZYIPfrF6K+1tf3z7fsrAo5TGhETzbdM7KJhIuFRVl38Wu3IMg2J+fTdiLI
o5SwSOYUvnLBLtF4V7T5f2kkJSPzlGoUmbrSGHt9SwnXcqn1zfhZSPZzXD6qy/27
b7+2AP8cWESL4o28XtnWaImhfJMelAHW+ORNlpthahRWYU2P9a8tJ+Wk3IHobgRx
uqCDMAcGwqXlEr8D9f+R72jgcm07BmXeLP97f5PHkDrmPB5HolMsDYPbnPYZXDYI
QSPcHn0/GXdw/fulz0mpATC4LaLrlAbzsa8OmNPA4E9woEi4QnIH6soSmz9jLo4g
nBWGALxwki5nT+O4N6vxprXBoXz3q5qhnyeF5XaGnBp3g07EUEVuh6zn59XAiytK
7PqCfRh4M6lGC1NGEHEO+0fAvtuvzi9P+kW8ZQ8IXYkFvCPnaEGAL67/5f1d6rIz
O+QMAv/95AR/XYOyl3mhiF1auwKT9hzsR4vA6wwaGg7hDSDrJlK1yHYzkDdgGY/I
9tcRUPXsQZqKb4rkn+i4CWQuiPWiXrLgbBN/VorEDQEK0iqoyj+y6pJ9YjmG2yLB
ZDytGrw5xQo3hI8fxVz6OvO26ZUpk2mbljs0+DthU7WGqOLFzfaJDXMJaPRMD4vC
5KsGNFB6jxGhYp+BaxSK3emxKG9h2e+ICgVY0cCE5oA6tslA8h9+x2td+gvyxWx6
PFncNRzRzoECHXW55h0iuQ8dLg1MLVsGi/O8QPtGmKKt4ji6bFDIQ3aTljGIZMYO
sNOhalwiN2/kHch+Aay6YM7vdw7V/YUD8n9Ub9cQnapyl7OUZiB55fVGbuVc2mPx
ILijzzPb67mE2GgqXnq6lqoCF5dMg+37W/51Ic90V8an3CAeBA6dNv+s7Y4ARU7b
FAT1gcihgXVELE/M6QLLJprQ5muw9wYjWiVg9qYp82eHOLeXDTmoXnoWwk6Gx4qT
G9N8eC0yORvQ7B01nl8ioPpPUMASryaIh3ZeDpJ6a4HjDFCOAyG7DlW3Q6O97Qsu
5n15tm2LMAzoD14mMPLmFvIcGmpVmVWikug8lihkM4UzbuR/6jjpJ+1yOx0lc+Cz
0I2mrV7uD8wP3g3GvPZKMOKOmXNuWN/7+ta3ILbDNMLVXJNHa7qA9UNkOA2Mb7Sj
Ox0TPfULYdEVcoI+cr/sjL+5MPfdFRN8zSIyDLRs0jCkza0NMgm/dt+H+8KRVd2m
IuAxjnpXVm7t3WfK0WJ4v2BLpggUfS5MV2H+jQHIifRMXir9bGs1N6ooRviv+Br5
vx17l3LipO7ZulxhTY3vrqShGFEpaYoBR4jLf6U8r+rhC+aBJkFitbhL8YIAxcEk
99rhaROzA3xLDQWe4ZiVnXHZW4TjAsr65L8c83qBDaRyTvcRyupPykwAz1lfCZRi
Lf4p6yYbLQXuiTz6cBIBvEWId9ZfgaM5U5w+AiNkHqiBsi/zbw+BvDd7I5KgCJR0
xnDp8SpW5HoNJ1KEmB9Ncx7szpVsSG+kcTnIR8gyO50vLxMivnyLyrgVxhcXuFwI
QFgEhA/Xmyact2Xa4x/ppRzZ9M9up3Au/9exCNQnzhRNunrP9/uUzCHjXXJMia6e
jhZQomWlDUsmXY5oAz9Ff6zdTagXpzk2vicBPBUeAQ4mxRt0NVKChUoTmnOWeFhk
u3OKe6lM3d2RQfMwyiabtOu6J9aGNQkThX0pZOTu4wiaw6BQYA5kUmYe/94sDM7B
H+fq+ltm6jhULrQqy/nuyusRGn5rMeT/Il7lOhRDeD27X6ZCGyokJoGGjkfMcCD8
A5buWIs4182Yz1QW6GFCSGp1fyNAa3MNy1uZ1TbCRR0ceHI4oILh2+h6Lgma3hc7
TH9N0h8wLzxGDlKXhj6OzD4D5b4PD7Nv5A6Bq+pcrtY9AyYL2SSpAJC522v/Gi97
GieE1bBZNgSFfRLoJ5ms+gnVSHX1JoQ9x0iNPkiu0M9JBuIyw0P0xLvqQJJcmF+W
Er/yY0qymwUQs7uiLUhA6BZTKWker3n2wt7W8TbQrhE6XcxbI2vl+gABOxaj26o8
qNdLlc2J2iPw/EJIsZun/HWdVkFcr7Wd9dCQDpMxyyMy2qKtZQYV0kzPUC1Pj+TW
4omWhi/h5OdsnBMT2KcmH0HLogeNbFNjm4FX3roHgXiRcP1jDL+fsKTDHVrg3RMX
cN4aurDAcw1pVb3mK1tbKEcj78owJ1GAF+VIr5Y67PBgQJJmy5G9d5BWhew/f88F
qgl3WBCB5j+o5Hj70jeM4Dqdae9ShnG4VdKkGhERoduB9v5m8AvC3jXIlVLI9u1B
j9elhSXOsyVoj7BCqENv6q49xpXgf8PWbs3NtXd4kSn1yzNqM/E9XS8BXWCgl80k
otr7F5F+UMR0PY7P0eVbw9h2rN0eLJsab+Uc6VfrJw7zOBjEqRQYAGELM7rF74HT
tx3CdC2fpElC/h9JAMRfXkEmFDl8c0fLRg305CdKu7Z/JuyR+XkbFWNMl7b0eNcM
JrzPknCmiZjWhQicwEmMMN2XAD4QzggGHajbHi/uImC9eJWknnTn+Emib47YSitc
5grlq+qZGXQFmIZ2Jz3qjPm7QRhXVGo4jYKeuuC7LwnCR/6X1RbbflHLq2HjIeed
2dVXcfVok1ctovdchJZ4V0ZI9X6aaZxFY/nFy1vFZz7lDobzoV3HtKr3OpOcb1qN
khde9u2ZwQzR07+PGv4BhN0Hq5furh0UeuX5balo7/69ivwYltt77/wKDFAiTpTk
9w16DixSifdgwi1t+2567R2o4M8uv6Lt292BTXXusbCc1V/8Y+HD3P39IMN05kgx
yj4Ohcsudh64qQCQdslXHRKl7R1vvH6ZkflUx+4HEApbG1xwpa/dyoif0iHuTXU9
mcD5rxYOQ/VgaJOUbWVoJtD8Ikutwv8Ud4JEFWT8x6Nv0acocCWsKKoPmgYwwZ7J
ML2bzL7LA9YMRrktLQT/gJJTgA9SA77/j2MgW2/Evm2O1vIKFdgbr/rzzY73ncvI
2I6jPkvzpyRKjLotw9oHW60M57Mlre+ZhQUN4tYXlZcePF2ZjVYPWH8ggUcOg5vE
PBojG2M1KJXuUbB7SUqMd2qGM1moIliytInl1z3y5YYuk6Z2yd5eJr7U60FWjCVI
2Wn9h0GZF7za7RTVF5+3vUI+snFhV72QDMrriASJyAJDgT/xwkioMSQYtS2qfn5q
D0Ner4VV5TcXwlJbigPhhX2UC3ZDNPFMLJzPJ8dVGlNIHBxGOu8DCDWVRYDNqEGJ
HRvKiJqMN6ApRQFG2/09VdwlD2eBl7UAkawSe63h780=
//pragma protect end_data_block
//pragma protect digest_block
txUHnzg6nDL0zSMVvCbJqF5DLag=
//pragma protect end_digest_block
//pragma protect end_protected
