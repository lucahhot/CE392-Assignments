// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
cvVNFM34KfGokCI8jVNmeUc1BDMAC/Yv3VrS+OEMYR2yLMDd636hSzyDL4YmxjMO
xE52JiW2FiAdV/pdpNC9GkDmlYaEjOvfN/0oYKbqLJu3JQw5fy6G5OyfkG25O6pd
GTbduXj0xvV4FkeOx8K447jrxyUvMuCzXh92AbKQyxc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6016 )
`pragma protect data_block
0HXwuB6kXWl46g7ioq5WwFB2faEBvprSPLSTge8DJGoVtf5tIwhZMd4qeY3f7tWB
NxHy7wh3tpCL/OUIaAguKCEVrXas24KPX8zjjIpBOkadIUmBbFeKBWXKLNDKOxlM
fjCc+6B6bjyHPSMGUsNck4iLJ86pJmcxB2OaNfSIdXGcDy6S14/+a+Dtnr8EpxSm
lP+MgFs0JZZip3hQ7/nnEWZh+FommXVwXwC1wv9O1mYayrM9BBVQtko3nIXMoaTA
NYMbgAN+eImbRrAyCbqjMJk8bbH0nTgz/Ta4E0X4Q2BzWslqnQVgvpeBi+jVre5r
Rbc2tdR0u+hbH/KsGm/Bygj3PS8w/mQQCg4XvPQpge580WP+jLX3nKyigh0OqEXI
ilxguCKgXJKOcIlH8E6cIGOJJFamQ4ce/vxnUSTdMrN2vriNdu24zXaAkL/1YbLe
fajEyVjAxHN2PUJn1b+TLJa4CtXKO7UUvCBIBLny/SOjBcI63aT432wll04T8QIv
NDq8h1YnAj4zrzbM33omogejaXIY9Crbi2wElQZ0JIuy3eiIq9pHLAbr0KE1iEO3
KhEq7ckX8NinWvTi7mct3OrOT5w/lHHLl3W2pTrIUFeXJ0sFUIHzTOqxPNCPsJn3
2Mz1/AxTNRxMz9rGfjTWbmaldP5gBm9iLm/6G7TLPI+sw7OMKDj7buE8ncY30Rpo
1Zhn0xA1/NJiouZWXsj7xK2ErnvmoQeT9/M/rc2PrApMhVsXDjSNo4ek/hSgm1TD
ZXzFfUNNCLBy/cjKXEyyaypQXOh+DfIpcedq5iPpIH48OHWAF9VwOUS1pSr2sFDX
B3C/W/yYx4MFp6jxYXr+lnv//fra2QcU0Go5Dq3TbNoJTFPHM+AqLeEooVj6U2tK
3xuZ/1K5ekRZVNYtnQrKJzFFA6syUPxmCoN5Pwwlsi62pMGSo13FXqEgRAuzKVuH
uwvk5olH2iakXYvJe9Y20Cc4hJy8LxipsGNpfMOfpMvAd6kGjvrMDzP2M7OfmACJ
4SXQ2NnNcZR7XiV1A6kuq9hA88RLCa+EEFc5wTh5wx5gr+hMhgYv2/JrAom2PP7N
eDd39Y1ZY1H4TIShFTM+NRt3x5c067p3GbxZzLG2EC6C2vJmlQtidVO8Nm+OfO6c
bGTPnTLAqsun5CAC9KNfGYjjCc/zdgFR5k5FjvmsmBQJ6ddPmckDeROo2VjrYIy1
kKUgWoXgkw4KRJveagV5cjYMbpm7pZQlMPrRZj4mIMpco3m/242M9EZsJtjsitG4
Kg/NGSl/ZpDiNEhYb9xvcTA0oF3ryZZxDrywT5dwbqp+AGQfakDFRGW1m1iGrcOa
Q2IqwxsGgh9gJuhCp+UQPJTvtUQWFgPHTBfLzSwuAVzIf6j3Ucz5O945NbT2FqLx
iIzoGZ9C98VJLTlUlAPr79eG+KW9eKqJjn9VuRd7uenl+R3RT7oOg6ZF4tPVqMrg
TNxCEI7GyBlHGUT2gWnjJlkSpnVHM+amhCJgMw+BpsIpGDNoSOc0gfecWVrKopZ+
UB1vpGmc8CLgNvI4XzacQYQZ/40SaPUVuH2L3at1Jsche83IfkXPt9HHTqjMqn8d
RbAfE0YH2uHiJmqsF0Eq/Ddei6v+jM8a2/BfglFLjtKOvT+eSLwgq1m7c4UDGqGT
EHtana94qhdNKwWIwwxIiNbYwlagJVuepLKqasaSUuypZMq3i+0//8k7z8B8Heul
xMldJoQkwkwKef/rR3NqpMqXQEI2G79zd2ZIQ/RrDM4uyxkJctZbFZe5XFUo/Rer
kcE/PqqBbI9TeiT/HXUBEbgwLG2JPXupJhK0xUfWPP3GngV6of/EeePC1ZIfpwQ8
/lA8P4Wc0pqjPtn8VlVuVZqVAcGmps+Emxv1QoHtyBntWzFOCbygiXSK9DpcS8oF
tuaoqBhOvQ3x9jKD+D1jM3W3clG4wIiA4+1m3fGWioPDxigzdjj+O5FDa4zI/cmU
dxqK+dRbgqrLNe9u07rGRFDLqOGEsqCqcpbUNIt/PyEQkZFCB1f3vA6RZvsbQayU
c+rEhWvInXe8N9fQpyKIeNdymdlDBuNNtjbIbRfzmH/IYpB5QSuAeDelU48YTR7Q
GeiWmKuCoAf7gb0xYtOG3zhisksheOZYVnuWXWo7k0GHuNqlfqa86MxG9CLJab6G
JAQXk95ViW3zU32RY1hJybdSBRigYz2Q3RyPfndETC0mC6HT790oCPnYYPoJ9+x4
hdOQQd/4nbYzJqGQiHeZrtNNeFL/9N4pA1rRfKB2htnf1PIcOh5h5uSb8SVklR5y
jsQKgUxdh/MhVCZXn9rEmFwhHJ9+BzKFE6uBWJ5pLNgn1PeiIUxV3omDvt+1IKf5
Dzg66ujUYejwq4IHdy2WSfqO0gCoIs9l/SdFcQ7jwGa7QYAHpcCBR7EeTbhOYcTh
SSyGJRDjhr58Ts2fbI/J4+adc1VPdmCxqLfpDVREgS2CJSwGSj06yZmrjc+97ncK
BeH4FkHt0D/B7Ez3U3SoYAaD1un29yIvENlJL6joAgNQNnH8iSA1TJjDPpa4l1lE
xvmaaRbrAzQUhr1J6Qh56Jg+PXq0javBgRDSlBTbRuSnMDAkMrWgvqsOqEPmGlwb
aP4ZVonAyYfPWdFoYgGhlT4ZXv9k3uxecmMdle0kk/wKSBRnYg1lrIoTkALYA/uC
70rBYfrnSiQYdg8oCXTH2xtruDs8FcSIj7lVDRqgZqs6B2jsh0A/ad41nvfs7x7i
yoAOvUgJMctRAOV/aMfW/xkeFVrTiswx5C6PuuiuxEHKBvGxeadKTTbaphSbJnaY
ClnfK28jb91/+/FCnGqtos2ChsQzXX9v9JkIta+Zq26QzeTQTHezZcsDyLeZvv7m
fuEgy7KCXwEVEPXCmUzSEgpuRHBwoFD98Td5bYRnMr50bSjmTBOGjZTUFbMmUn/Y
A0lCM5mrl7XzwRGpfssdNXk/bWLjrA5tRjHv2K6y5MPXznwgDMmcxD8/T3CJYZO+
DWP1fOFUEi6nH1D7kwx7U4evdDDsuQvAdeX5QoT2f6oEMP2Nmyy1nR7aS1c2UR7b
cw6ngrc1qYcZTEZlGohhyvZwEdqkRRtb5K7HnWflV2Yyl0ADqRKrjUPa1RuxeNxh
Wo1ONhP4u79GqKitflLXon/pnqYfBFrYP1UHLgbj6oYLaN2uu8xQWMejQMMQWlTj
DqbyDwOPkufVpubxng9tKw4Or7kf/m9PjcaZS1ufzomYF7KkaN/ImnApDL7xqosW
gsMH3GCLxUMnFHnjnlPtFs4bcjx+d+iUaQR1EGkqYIRw/1kX6Tz00E1QXdLMqLNx
3cAPNFB5hQpcYl4xbj15dK8aDq8zq32oMgdPzGVQmcliGyYUvlIv0LVrG3tN4D7M
YZyg92hojyozNHsO9ROPNXcfpkXnurYdpHsY4BHSyL2Sz1u/hxSRyFxphV5+J/3g
13Qtq+fdUXNEXGRx3IPav0CsBQTrY3u2bk/RxhaH74KYCayE1cGQnZgVyeUBAsOb
CvMMMZ4r56+brvt1Othev+DiHSZb2xTKJX8zz0x1u0mxl1bV7H8tmVwdjH2EnJF/
cUXUgUZYlsmu7b9A/M9fU++uRm555CRo8veZNmA4GYwZbevwjFYNKfGpyxPJh87m
JFpJXUuCHJJeoC9Z0Al97lHKeLqK91+4lXSU8MHlGlIAUSsm6XwL58QVUZWvjpgj
vK7uvJjRl0H5grHqjPPKRLWIgTAU+gmtKz3C9S/y7Z7a1kXdeDuAZTEmZK42EiDQ
MU64jNEw/a1Uv6kdlaV+bx1+TRJ985z2+UJ4Q7MHf7B1bCJrgPNQ0y2r/PLC9HYu
+D+TYYOi+gaxBHUuEG1PM9Zj4kiYWbhytmTpBUhKGCfvWvMDcqa+9XWWD9RaDa/Y
dTiM/LTpYtDg+FD0GYvBi34Lj7tPLE4IYIiWHvVIcg4Yzqr7KWeVJAPEt1DGObOo
7O+Pnll+gBIOhzmiMwUsCeeTLtuwqHbR4p9Je70f06ihpRFot00JAVeyogWIspW1
1CfALxBs/ZzXhD7Ok5BpWnDEvL5HBu9XEDIzuNM8n9alhfh4mY9Y8WVpE/Wbadcw
hl7S0Rh7ysg8eqCcWSWzl1+gq1mmuYdfKC/fcS52iQkgRreoPrYFSP1Y9JwzLf+L
T3hToBj4DtWurEIxir6yui2o/yRAcU8WQ8FyJ/wa9pow83bU0HRZiz9EO2SUMOgI
dXyuMWk47QJ9JoNlBp88htX/65tZU308nskEuZzwsQxtYp7zQPhzrKfMKg5VQD3u
4Qumuo0aMGtQMGOCypafxejx83BnHYoyxCBqWGVb6AiOcqCOmprYGucQ6KjC7X8v
XTKMpvo9SSRJeBU9M+G9+R2Q7LMOjv/tdLqR2j92kHaGM/7eoRe4iAkcHyJv9tfM
7eTlbN9JzZZtJx7Mt46XwxY2Oue9H5/lHN1q9xAtKVWGve9VXz6nQz5JnCMVGChs
6+Ik7ySBIQx32peLv6IT4+tVtWiSrAEEu2q/Kdo0CqoO3C5bwqW2dZJwcQQotPA+
HFQnqwEKwwc827DIheRPrX0BfuBUh+6TQr9rOM9GfAffkPRMOc1TeFyKe7zffq2x
7TQ2GG1TTSXUVabQ/4MW+QvBmteoiRrpLHpSrNlqOiNV1ztAQC41h6F7pP8LocMg
nAY16K423K+bK4eEIff4Kd0uAjMVUM8nYDcKEtaM5tmT1KOrUOtXbqUDPj/DLgE4
sW/cIKh8K6WwqRwRl6yWOl6pTiXzCw/FPmB6SSC/EoK4wk1SFmb1W/y3yT6hje6K
opNiJACt2Gt3nbdQwGSZ79LTuMGci++T6GJRFhwjLKTwCMsgyTjEVX7mMBHB5267
s/Y1K9d5z1tF0eVmvaRmrHB0dQjnAqnGUGcr7cYD7i5oMhZCCEir5wXR7mrDZt2L
56xlbPhR/RiZPXuGjBMh9ixj1BaZtp2FUP8Xba6QAa3LagkwLq/EZEW5CQmeiYlL
+4FDZTO+VdEL//TMKuOEYjWeTerPj6nkeAVjjK7x+BdCwAq166V91Sragt4kD2pU
aNHaCBZFWNx+G98r4iLa0YjE/32j+YEeaTSV4d/FPJDTxV1afevK6NFqWTY7K4we
epkozEbrHG8jaaslNZvj0cILrz7ae7jWPzNImdTfsL54rTtXAK75ROsYL0h7rt2z
m6rM9zCij8GXIKsnNIj5M0Mpa9h6RA6a7Zhyq87uxteRjhwCPprHx9zUOit70TmS
mkkdLreOjFzhZBLj+GxQymVSJjkMarNjn9L0/IpDa15CkbIl53H8B8vILYWUQhgv
bXFyeawiamjLgRe5k5kX8LC6rIKpvhPkAYHN2dXkHQnsJ88K6SsM54omSY+F1TTR
QXmPpTtb6t/C3ZHLHYl2w0tTZR86G4j2kDIHj9cK6DuiH8OIxsfQHyYO9Dm14O18
VjuehHWqzCSvVScbzr9iS4HFlO0MziAVw3iCjeHTzczIyPgEv2oQahsdeOIwHV3c
Edgso/gg/slxS4TTSUmTbTq3VnHUSmV5PJQLvHeoQn4eUyaZz224qVmAIb2l7ouz
AzO1seXH9ooRIKpUFRqymmVDGTg3Ff0+eghZgdslEj57aEG/9Hbd62f/MU0VoYI/
nYIleVfsh8COBc0TdbAqQsVdaCTfVKyfQcYGAVDH6d0PvpvGBjTpVwVH0ox5Dqix
WX0zwF718snwP5Z23BBbrjcWhrYZzWCoULyFCF8r1uYrwgF1rOOQX+S59g9A7Y+Y
J1dgozppTJwbwY3JIicp9aqoozR8tuwIFZA/F4j7/xcKeAxKVOhlYhvju00Zslol
AiijLQeqA/V0cccqpvL/gmnOvatg3+qpgfH9z1KOaAY5oNTU5PQbHgpKCMCU+06I
kj0OgvxoR+f4YWzxrtmCdcaNmPutACuMTA+8otp9myjJd57vGxJlROYXBwUTSsIm
l8agp8ITZhFTm1VVbFz2PI+DNQX+KaBE1YOGItJlBhrfvp96wHZNn6kHhsRTCVND
PNjrbFnxgys3pq6QnYPqXzqoR9yzVp00tEQzZ+ilRHabL8VA0CuGrapS9mwCL/M0
HKsW+7TZYSBbY2w49e5On/naoWfybrVTMfnYerxSG9Ufb+ECiB8a/5/VxGXvSOCN
hNhinrgzLkA8yXnub6CxsuBjtD+00qO2RjI4yWpytIKhQGmqyObsaKiLLAkchCiH
jZap+7JM3N8yWtbDIq+l9kIAbRndNuq/SZpVQp/JhqRT8SOQsip7oWU039SE6Zoj
Q8FRl8SrsJaTP1dfMf1naoMIyQCnzKGHFbZH7hGG8u7qsvNA2gyIwR/JgiCJ7Vw6
v2O+zlbVGicmV42jZAQjbA0/oWge7rKtcub5fc2ZMYRxlSy4b2nUgTU+PWa+Dsj6
1BZTY/1Uymv+o/tAs1BdQwEF84z1S24/LIfIHhz3fvlk+8GDNCiePuGcUk16Heh1
e2cwDBv0Wxs5emb9WDJyH6Bg7odk4XF7T7onKzkVPHq3+4anDhgNgdV92AZRYuUV
x3LWd3EKJNP+uE49wP5Gdi5QJSItNb68PaeaJzuoY7JNgBtqy1OChyeoLh9HkGJq
y5ks7590/OYnxWdZ9fg/lFKp/QpxyKvGunMQDWNqZm9vmN2MNIbsuW5YMhwQCbRR
2XYFMs0sU4W4B2UFGAJyw+Q4LtLOWER5OqmykJyqJCThmwHDQlAJhvo7pZMfiXON
HnvzhrYhlXRLY78nsV0YJy9cD2wkoXxfJyr5GZSgbXtwUjEL4wuTK9TjLxZ5aJs6
C9PpMvbqfjooUs+CqYQ9xboUY48EhZFi8t+RzjL5zmrXv5QEAGp08gT7+GfJnlRt
UTZuQCNNErJEs5MD/mUvZ+BxMOH5YRXJpu6SYusipZtrUbJ1YxsuWJ0/ByTCFPqF
DvIMTvscroYrDvDwr4zLjjjquDF/uJXgLcOZ2hlSnk830g2dLZSAgSye0za/umAI
EVL6UjMzi9zb3DJZmX+7+FyFL0kSwuHz6OEl8F9l5mHYlHaZc84stEuGlaTyJya7
h+fVQCnd1fEtZJt8oH8dNTRtG695jjBfkp3n7Y+M8jtV7eC8tu3Eu/DgN2AkdlI1
QEc0v5vwUhE8unkLejyYyDxqmcKdZRGJGu50rRvfAwCdlji3yrzxDkNAa2qY6+/Q
LEuiPNSgDkRWecVzBVdK4jJXNyJUiAlGwq38tifL1a3WYHRFmg3PwiYQsqpAec/y
PD6NMc5fye8uJNMlAWyFHIkLoF4E8ta4a7bKVmpS9E+irYmXc+gUsk0r/SdYMjtf
TO/2vi2eUyPvGIbqheVvzwYcrXJSE1BBxOmMkPZZn0n4VbCNy5QYJfoUXPAz86D3
7tAk9ztOr4QCJJ1JTpFogPF13zkRnhJff1Nf42T+uK9YGN6NOKDHyCbFefCd4Bxf
cWfazVjikzYYWZhzRKKsqTJ8qQ7eEmfcPNERl5H+E13o2FiE6S7ayrR6j66AM6HR
Sd7E/tlxJKbml4qxhG7WgWv9gLz9l7ng9MA+TJCgRBTaET+Qw763CJgRCRjmLGIY
NnpJa86/Cuc7YGzfFGK+AV7dFhiz+yqcu4/RLpOR4qgD9trFMCJqZbTUaSc/2NRo
MDgYUOvr2/PjDAQJVX1SgkwgaAujYQvxxP+l6ojKUSWd8JjJUYUAv7QFRFiCdaTn
2NJDTl5Rrz85op7mjlwgYApCctlhS48x0sXaAIXoUc0YPnc3pOZ4lu04v0xpyJ4m
MCN8vesFNM0VDe7qVNHnUTNKT0VI/jt+rNK4frx4KsKIy2B+8DAJvQ+d4izMj10K
18A5aNdzn/+HGY65B/IaBqyLiS8ecVTox1oYe22j2pbWmpKGZAuBfdlfuy259cgB
J97GBKHS1m+kobTCuvBayNAga1kWDzqlgZBUi48jWC71AVfHyvDRbKs2Hm0aw/at
t104W17pU8Ce+Gv2hiOsOe/lh3tSJohdhwmtHziG9glFpSOT51Ep3gVP9PzFsFLe
MJbAiB7sPfEQbxri2bVn8w==

`pragma protect end_protected
