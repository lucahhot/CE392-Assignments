��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�a�ȝ���,��p4���x��-&�)g��J���V�5�ֻM|3�|��1���v]�a=|����O�t�HI��Xv��W�Ԝ����hAi��6._�����+�����Aw�� �G�'p���K��KM�M�jL��#���O�k��%�f`wX�vx?hD�����P����;�p�b.;�a+�p[�S�h;��F]T]�!�ѧr�^��!�+�Jw�:��q���61��3>m�����Zy
�|�hj/e����z���\����wsJc�ִ&���RvzB���4�ad�f��裦_.����Q��8/�RQd��/�s2�7�3��;�dL�e^���b����1qofQy�� �3��|~����7���ڐg!Mh�ϮC�v���m���7B�)�q�
cI1Iܐ	lO�.�����M��qzrZ�H0�t�)	1*N��Ϟ��6E�)����݂W(eX�1ei�K���K&_��`U׮_���8'��$J���=�@Ŗ3���rT���8��_V�p�p�`�vF]R�8]#��ZYvD3_��<5�٧%�  qBy�?�b�F��6����nحϱ��>L�x�Ij�&�Ҏɉ$��Y.�V�d���d��ϣ D��tE�5c�9T�*G܉q�b(��c�f�����2��X;nB�����y��Vlp�4��f��U��!hm��]&<r�)�?��i����6��~Q��DKnxR{�k���C�3��_�����b��%RIX[�_���e�Aa�V_�6�1�1U�5o΄�/���_2ap���>�8C,%}�o� }�����Mtm��DgF�1cjw�m�9}��t-=YT���;c�2�,W�]D��'� ���|�/�����
�o���^���"F��'K48~b�Q����F��Y,�	��|S��`�i))�xCX�[��*���o�W���nS�n.�Hu�]�C =�A\$�n\g��P����+�;�M �Rѓ1�H��B�q$��l��÷W��*KOq
�e!����ꨤ��J0_��?+B	P��h��P��[�����'���{U�1�*(I	C�|���W�FvʑK�=��2h�Z)��U��J�g�l6���z�+���/3��梃2�F9���9�}�Dz�{u֚"3�@����A"9Y�8�]5��pL׏L��z����۫u��6^s���D��9O'}�+�a�&UYT1�B}��G��gIDO�8Uir@�eP}O6����M�Z|�r��8���/���'�\�t�᭑tl4�DJ
Z��������F$�F_n�Xxx<�54lcK"��ƀ_�M3x��2̣stױF"��Es�3{X<��&w��s�����s����z�����-���;	ʗ@̔&�&���w�O�Ws�:]ي7�
���'ǡ ���!�W�KʏaS�eĵ&d��eynD�o��ˤ�S���P���FD��8����u̹v֕�� �JF&�̬��P]�5�4|�Vu���/}�Le	s���X�8Z��W��yGB�E*��.M1r�"�"ء�d�)��e:�'YФ���Z?Q |�8n@�L�Y/�n
�&�]�8�4"���`-��_c/���!��#;�U�>�D"�[/�TphV�j�&/,V���/\��-l�`&��
d*o�DYu�c���Bz6m4��pXi#�9H8@��� ���3i��ZA�W}�/�J|fS�3�;�#��aҁH�	��eڟX-��	�sǦ5�1��Hc����rxh��8f����R�2��R!D<�y���5��8����*�5��rR�Fh�W����m�m�Gw�m�> ~JG��%;���HbZ\��S#�9�zK�ů��c̑��s([��|3�����'dj��w.[)��մ�Y�-Q��z��5� d���f�����d\�i��p��vS�j�[.lX���R�"I���i��_!�g�p ����}Pb�SV�k��%��H�:�N��?��!���@����&��c�� ��ϖBU����]��2�Ç�D�%�?� ���;� N��Ư�r�M�4x�s1�A }�!�������54]���<- :��7�6Zn�p�}�I�/��ՠ�~p]�5u�ώ�����G��C/��� ��/Q&9%���.�������X�3C�C����0A""��Fb��Oc�!D}b��f[����4��#��h���b�{pU���Q4홦>�s�?a"�X���J�g����X�N�.*�a�+g��j��`�����9m���q:���/���_�Zc̮��C(���:*��OV �P9�Ǐu�u�>[`����>0Gbh��B���n�~%Ai���u}`]��Lng�w �큖l��dp�Y��,�ʢ�D�D�� �_4O����6�B:v��j�Y���a%F9]<�������z�8߲�C.m؎�;�k�Or�y5�B��5B��l�Ke8��5dٽ�����fL�����ӡe��!A�EA��3�\	��x��8)��'� ���Ƶ������]l��l��\Ի� ����{]�9����V)N����22e�|�$��_s�b��Շ�Ö�A���J�����]������#�$�W	�'�(�B����z�SSz��k:��5���`��ظL��52���[A/�@�BhF�ge��Ʋ@���y���PZ�B3��Q���H	�%q/�*+��@��ӽo����&Dn6���3�U!�` �o�\a���mP�FǴl��]���53|�c��^� s���IS�Lɸ���/���,t����RI_��4���=��-�w�s�uj�\[A#