// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
sQvXigTAwo2TLy4P1px1Ho73IFdW71nLCWE91Xw5m+3jh26mLsXGxIMOcJAIrvfj
rQhI2deEHXft4cSJS54pHZoqxDMNkMdA0UxDeOFdXFUIrB4FnFN7IHjuXuGNRzVG
5VAbGiIbj0oG9m6IqdK9Zvejn6t/53lWX7pyyfZju0PxCkTS4lmeCg==
//pragma protect end_key_block
//pragma protect digest_block
M/Ahu2BqhnCf47u+avaZ7BlP6jE=
//pragma protect end_digest_block
//pragma protect data_block
dVfPTdSA1+p5ef9MHNAetURFb4HLOw8ACrul1nQoWNx2TedXkFYkIhieBggrKR40
0p0OGeAaSRThTUB7cr+gRv6xcqHKRR8pAR2AZg2zE9xceDn8Sh2svQZXqXhu2sIQ
I9EQKMvruxhgBfR62Dfu0BARAmBInzYXRd5pF1mgzaNmv9PMV5vtRwGK9rOZbk2r
5pCF+l/zQ7z4qMDQL5cLVgPZ5bad/V1GXTSGXQ3ne8gaDoQQw9j6DiV+2ku9Hwpa
w50yVJqH8h2ImjLO2jE9Xpxzu/OXMMRZKrN4BnHa6CypOvK8nEnemExtL+lJ82Ir
1EcaKBt6sC9lOGHbHDwlbswRrNT4UE4z1gJ3GX831PSfJ+zfy5gzIjlb+925loA6
awB8MeLNlvG2ymzUj95CmGOEnuSbKp8NQMrb1oDi9nUu+2cDJ2tttDx90joloSZD
nIdqBCrnHFY813Gp0U0bLwrowFd3dkEBQ5bG7kumI7NAfHLsm359MWcRC4INBDYK
v6XC0Dofop5/1Cr4WZqtCiVtTya42zZQ7hMmi+aPxWs7CJHDgAcVZu8jH0oreXGQ
G0sAApZHpRCSfs2IT2oYmAXNcW+FX451axamuWuKZbxYSIXp1Af0vxjq1JKvyt0K
qXhtzlLq/u8IyHaKQKjg6WXi+j/KsXVAx67e1T9hSEyVli4zZm6ImpDh370Tvcju
OFE6GjLBJVSgFQ2ouU2s/7ZrPIaZ4CHr4tSUW2ZukpfmDbG1XI2wteZQFcUwe/E6
hHvVSKkcEzojozIzoc4VvxS7x5CuYyxWkaXaUYdfDs341OkPmMOdjxlxT0ad8bB7
wNxKSpVVGBONjrF4atRiS7ANButsWu0tZ1o3NQjQJ8K+iaX74sOJeHJvUP7AD7Ni
Vi171+sGg7SwnuoUHglSxDHHZrcO1FcbGoWj1jQ/H98RijwhfCHGSyM/IB0HLccj
WO2OczYrpZ1Og9PV2VHkOkeMffPAVurQx1VF7Th+WoBQW8I0gefAeaxCxSUxguk0
bM2qw902UQinqTPjwHoyqix6aIQH/vJPr7KIRkJNjJGrRpULuN5NxzeNb3MLGGdZ
AhIGhi9WRMWHBlArsdG27S67aA8UqfyKycEcaAZqD6YEPIAKFFCs6LgfsnirpVaC
yZ+ucEXiCowwEa9gfjx5kSx+fa4X4KC8UjSbgnAsvJkmuJGtr1ToqVrV3oWJr5u3
mii1PpFiZT0B2bwxU3GT2r3w00+ub/cXxVkChbNSQ38xRJ8I+N8MPey7PFtHCy8z
p0/36p0wzgpoWIntM2KbEbeNfBuejzl6N4BdCX4ZLKBvEogENH8sKU9MUhUEWBor
bvC1JW/rHzuKc+FeL5xwfYn0U3VurY+zWLDJKNRplwBsE3SpW/iM76jm/7MvFe30
AVqzFO3bwygPQNdke5QbpW6eh3gJcg8Nd3oNtT+OKwHgGcb1pGhJnq9W0lHK0th0
3VdQllr51wiI9VSoZ+ZQiHN1smaaNflRBzrjAwK+dMcadLNAQHbPxzEtR2TlNiZc
qccn3W1j1zSJuBUeFLlw1Cy1hVHJ1P/2ucLntPTC7X5U3hEFRS+mmLZmNwhhFViR
V6+0D7BBnOrCK7Gj6fJs6W75lhMaNW2tH3m8oAgMePsEGXNxtqWI63xDSXDHIVfL
qbfTentWcQKLCYx6ULSYUVIqFofENlKH5ySt/qd2NrEEni0H17CjIAMGzNOxwL/i
5ZVmr1g4j7brfHyQ9G37MKokhMZW/qp5sBeFucStX2pQFj5ySx5QtJK4M20nIaFc
16ZGBBR2zw86WiN6IiIpUepVRzbrmHcZlJwPzdxFoMy1d+QCXwXc+HIpjnO7hq6Z
R15sS24k+veGHUdH/k6fzn7JlsO28dOCPRNDTWTHOOw1J9UPInmSaa4fvGMVNeG7
ck66pYoIa8uRIyUfNmKtH2c9C+LNlmgGllRmlANrYNYsbYzmgd2ocRXF3xNiVc2I
ozoPxyyF21lm5G8dfCx1lUr09+43Y3aaU229PPtBDjgwrhn9Eip0WqGPewUT067M
YsnF+M8d0XoAIlDSRFDDi9sEpSyBTh1uqjHrH7Ooh7a4heU7l6I2g3xqlGS0fDgW
cArzzrXCv/I8RXR6atGJgifrK6EgWHObDAbIzlqqzZ9taClNJAWVSD5r3w6f/2I0
NavvLOV568UWT3OvW/+3Axq4yIyGcnI92zDvbmG0vuF1yXYPn28eGmQ0Ro43UKF1
jc4hltpEmiHwYZqGKqWv2T+3jGeB6vDBxxF/Voo5zrId73CjjD88Foj7eyLEBLgo
PcDYg+ebzehAleATFW6ApgFAn82dnDHsmGd+otrPSV+5Di0bmqZuwd9My4PzVXCe
xk1s/cNR8eLwOQVY+O5uNDWioLL4Rvp0UvjQX0Bbso4SD+dCWUR9sjCtdKVAXhzn
cO7pEuuL8mI7/Gioul0cePYGl+MTLO4MdCzzjL1LmVDB+d8tSrEfHbozN5c1J2vU
OmOwoWMMXXuXT/Tzc+mh5MejMfxMPXX5CcLi53ca+/BxuX88aH4qH7MdgCzXyVmZ
55QoNXxdp/BI2+AyFUzJczI95vEMXbkU55ozkZtQ8VqZfy9SjlKzdgfjnGKXCfGh
RDCtbkqjCB4E8f7l+z4GpBIzBy0fl6qSxbyGenYBpO0pGuOmcheyvyd2KWVFxnz2
w36+EC9oiakklT2DLK6ElUAbpazeYBCikdUX/RcZ5g6SSRvTYMcxbTPuMOqYkPN0
Jcw/f5fNKbVPDCrDC6g//ZMdB73kQRDqTmv0EtDsbRR5+PvvbcdU8LgE33YygfRP
isiITFAWa8i6dOPGF8uoKEkROkTWYmYJEAZkIXKFAWkwO/LhOZwpBV6uAEEknYwj
kctRhMuriggtD3wPqHbTYkkvxktLu3XD39ulKH6DLwpSRiybnvE0xby5j1VoCzmK
KiaKCd919jrRcS9qWJJPNdxN6QQ3D7ddUiyhpQYSZ+GtcJk0PXQvLhjGwIJz4HgB
1ZXHpImBYGHeh/pfA+jgx8zaxbLOXCeJnfMf+O0HopcvKnhauDKX7KQRjtX/sFxP
ZUyz8j/a32rfO/80B/W6C+4ZWBMMpmf5fxj+l7dFqFhw0peXqhXtxFCZbvVXmKch
hlBk444yDRbISn6lhcWJslb46jtAJcH3Bb/SHshTg4AC8sRLzd0G08P/4uci7SFY
qN+/Cyq9r5PDSXgCo4BymDQ8EF7oNukNGLpE4aObFMQMW+cgWc15CsqcYwxEnWeZ
Cl/R+0nXWu9ghqLIUXi1z+h9nhaIXvcoD2kujtJf6UHLZ+n4S6Ar40OjHYysbJVe
lKu0jIiAmN7Z+/COq4iITrJ+qJLoYGcOp5rxtaJJ7bGlKKk8FujCNqTBIYBNYHRl
/sbiocWANNwF7LekECgwhsc/myQFIf2HpKdkyrXwUFvQuBDuklhMuUk/Qoxq0+5Q
u0lhTx7RtqI6tHjbT0p/kC2uGm0CfxXTmzkkj3n1fsLJFTj8363DiXu+KlslRSJT
TdHZACxIG2B/gF8z301S7wFrYQyRzqZ3EcGlcszyWeRccYjpSdnezCmk+QDbjOjf
HN8g/PChHql/tsChFgMPLGqWBmpcop4JrmTbWKyCEgstER29GCMfMq1HpYuSLLOW
GY2rg7yddkxaFB/i3a9welsQPPZzIWXXVaYEOxy7gmnazrTC6vQ/+LhoWMQF4Ayf
6hd17i9ae6N64x4mOqabl6FzpKwR85C3/2z9pkuTHboEd/R4PvGuVgT/7AmmyIB+
OsAREQ+Ge0qQjD7MQw+KW2jbNExgLVimI9Gpva7/iwaayPLNAf/kZDbwtydicS2r
n1lMCt85k2kcJSIkzGwM3mPmIthggSU1nYfQj3VBA59W7VNj0LeBhsJzJuCIP/nf
I6ZHyuVvFNoZdYExtRoixhYCsvHn7elLIsUwMne+wpKrQkdJzLld8ja+7HxQVefv
/wKjQB33uBuYMjteg7xaSxGWtNiKkP248eauS+LwY1KXoA/hBDvQ6wJFCU6PkOdc
TQh7aAIIXIctl7zeevEsEdFKmMr0dpSbhUHTD7nYGZwWt3jptL5zHTgNpY/r9EGY
RoFb3r+SaZQXRXIvWa1J1gTMcsi1jFbcO9EBgqWYtDQdD2K0OVReuZJDZRj0pbK9
5M0p0KPFp5isXYKw+yGm2GLA+HUZ7V/AfmDAkSCAmUO9tXlnobJz9uzm+eUmrtQk
54rIdmuBse13kVoTtvWPt0AkMHYxNii1l4C74TQSYf418rU2duTDO5DAMVhElr+a
/Mj45Os+5pqsXkLEWi1WaJebkO5ZKS1zOBcdlrXUoBD0WNc/PDk2hNasM0stmTnT
qmjf6RTlAzsiYzGOlnPS7Un7fK9P9bW4PbeBYZAKALuqU6Kd21Cg3yvtWETa6Ed+
wtN98v+eBeuiD+bUcgrKFXko4L8utW5pochf+T9TTOR3t1H5JP2sjJL2Q60/Ge7M
dvPSHY9pnjzgrSFA4jAnxUYYks5aneFnaktiqxQADEUk6g5lUF97MJUDQs7WpFzr
SomeLgDx2Ege9lA+78oCfZ3HoIf7x7T0STfzoniMywn9wunqob1Lju3giP3t88qi
y2R45yKMY06qXKz17Kzkr5UQJYzrjZHORJgm9Y1U83BV9nGVd+GT6QYeZCNZWIwG
uqvDWhE/KDBbR8rPkAJG27ToAeaWBM3hWOsjCliDWaDbsbofhgORV8aWwzGHNjBy
RGl5EzMw8myar1JfCpKYiAMX9sX5TcE8wy0KvQDRpbqtxvT2LhXEcoWRxlURMr70
qH6miBtY3AnSF19fdVSLoftDwf3u/x1FFIY2wpRGOnSacc6rTCsSRO/w99wyQXVq
NVs8UaeVrPI6Hnk5lN6M9E10VYfv8+ZVYLcmtFPZdZdguuUrhexcA8PKzEfxScV6
DdWZcs4FWVxRjD5ecRoN6LopGx2PEvCCkk0vj/czxM1rO+FH507mpLwEcWNirS3Y
4sJMfp4f7GJoSHz3JleiIeBoJIYEYMQyxaxFbpVIFervWfX0bBEevYxMCLbJtqtG
uY0KU3rUw7qQuFRlRnd11kl4CTuhgCxZeXGJMYF9zZ2Z9eRJWLfi/kvAOBPud1gM
ExaVhU0BcfOedcKkuUHuM5yQx5Bup02bXg2huWX92Nem62aU3/zPK2SCeaBaJfw2
imi8JLASvWALW5NQO8M/0CzrnP33vY6AIlnyxVxga68OLR8yQtaOAAhV4l6cEYx7
4GoWn6lukYfuqKxucyNcPP4JCDvkKac8AZngXx2twj5w5vH5h50ma4N0bZWzhahz
iq67YgYlOVSeZDj6JyR9DVjRjaW27ItycCv2qFDDTS2yNj8NYK5bmwS/7qvwnUtu
Z9DszgEUq8Fkjw3Tl8D+MsJrG3IfINpQRr8nr04LmmPLJQ3tNlPy0dtG2B/nrbFe
a6AWFJCy4balPmPH0YEs+pbesXwrzTF0dG6gsxo9lpZ/IV3lGktPkxS0k25+SmNh
y5h5XIjxUj7P/V9nHvjv2DI8ZuOnGEXHM6S6hJAP4+1hwt0XAqK0VXvt6zlrFdE1
pJYk+ps6xwwWbF/2kIfUMX+nJHNabeB0arh25ckNL+Qfjn4nlMBFUHTK8GgETdFL
pvgYmwn7l1YVW+QM9rswb/+sq8T4qsdVQ2lB0eru3ZCx7LwhQ9ei/cbOpNggHH8H
H3s/VT7dLA8WxinLtWFhIPN8uCh8+iFEzy4nERAodt++8p5R2JrBH7u7kBReT5u8
B9kJ+CrZ9JTi4aVvfcf+eFZKMxPU6azkAzNwgCoubkW/O0XgkwFFrlB5ALaOArs8
Xtf11T6uNno4Yz0kUUo89dy47VO1pnwB/69/pCLS7BpSLWUjcbUJbQYB/TxgQpCb
g+zy+Hl26SChQtAzUcFP/r1mEzXO7AmugZX9kohkK6R0l+6AKTjfBomgyHqd2XoK
tq0u6ZzpjilwzNx7vFXHHrAkFx21/cnoWvDmcAJp8S/AP8ezMRCaOEToZWYdWuV4
q0HTujh627bj6+duHJzoPVLJFSBG6BGJqKvD6LFQ50vTjQX1G58QvNvX7wEpEwx5
IkcBHlz7XwvteC4u1USN4Hxme0hQS1P78Tce7lnVmD5xrvh8t8c0c84CPYfHPWQP
pKVgFhkE5lpHcKKc5K/KPgmbJzy/H5zw/KUip6JTnSuO1N02fP39CPomjCz2DvtT
uw1OQuj4b5CTEP067PHhyxb976U+HdkfNaFKfgCx3qesXAzqxxZ0J5MWQe3sTQJY
DxmbHdhtHXxrxTY587BDBYHCriu/2Fvx8kEzBvADLgpLOZsbIBdcLtqSntuZ2+ch
kGXKE6qEnBtr8z4mXQFTwKTdERs2lrLjgGXf53+SbFCY0h2DzyWTAe5KnFpXmSEV
tIt/U7y7+NhTdBjQPT9JW1YCFSYkdYdqUhKNV4Eq8PX61WGO53T3J744Xn2m/Wgf
mreLIDQa6y0yL0YNf3pUH2MKGzt72O0paI5orYrdq1PCnQJ0WN+Sh6/a2hm59Lf+
8vzNXO0gaB9rfDwsNqZsxeD2GMQdzUsd3qMtWGf8UQQFYNfAL/6/c+g+Fq7ZOl4I
KFFPzRZSSrGVzh83mEarVllKJ4cD7sw+9XpksTYmWE39OVirnVvqQeGmal2TwkRP
VQhV5KNzxLVFGf0uZVqSqYJAJVVQp+jYa/YucGdryt62d2wO5tSTteS8/URe1i9W
LKzZfLjaRBtJ7C5J5oTNnHldTy5/rAr415SiEfO4VZGMqmymaWbnWRvhuvIkJEVv
TCbPATIF40nWwEwhBsRM1IkVg1Dv21uBihDaRo/0AkuuNbmYKJyMK6nJzCqzdynk
0KkEzbMj9kb7ttC9tfUw7w2Hh9s8vKymFQPvzMmChuKuO82hETq2Odf1N8nPVTLJ
T30v+z5zFI0ddf7T/6BmCxWbX7EVFsVRLsmy3sGIoTYwPHIULUoLVzTAFo4l5BG5
5JhBkFcPXizWiKnjsvLfslNJ0LOZHb0b1nWmUP9tpWep9ou6eBYjgW5An/OgnKjz
pVq65zvJQjOmMg5wengbRBZmSg/Or9tqUDKg7NP0tetxexbgvjhoxKRXMfMSt8zs
sQ4I+Ssd+Q+64Nv5dJB7To0WL0I/RZeBigoEvRkx/bD/0rP0SF3vGweClke9MsgT
nOi+67ig9hHaLjgGoMwOGV6LFSxTdzedgouTY2bWWTpEBODSFLiN9w5vzlTKm2lf
eMpL5o/hLst886BkLx09/N94Ub7M1qRnDTTmszkoE+PilW2HvLmYGmcz1EoB9SGy
pczAeOV0K7+ZeZKfxEc3Km5EJaY0ihqtTSkXlBNxf3CTM7FIcVOXJeDtap8RNEFD
a1zEtxLZCZ3lWhDJs8r+TcLBKHSTjXy5HQjhc5bNfTOpUJmYS0U47vow11/q6Mp1
cinBPRu2h/pJal4u3jbhmy39PkwsgHCydN8ZNb2SLrQnvjpKYEQ18sbIj6v1uVV5
Bg4GUCXLe3VvNC0dpbBkhi4yNiaUqYEqgD9/V7ma70GfkOsS/ZVIVx/vFBT6Kfmx
F30H6QjmNPNXn0yudsw6Y73qythYr6diJt41yMXHWAs+HWENvNcnj0n7Th7jLimH
Oj9wbPwVz1qunLbMxfY/6nsGsU4jCPD0n0E5etufNwETx1fPGoiKTMrpeTTm/Shp
rc2Ih3lW1R4PnEsIysS2x/E9RkElntjgfbSoh2cbbL5Cvxjfazng27SlhDRaCqff
Nk2TpCFfV50ggpmCsD3P3DdMDvnLhnfViXter5kNUO7KyScJsnKz8kJqZcdxuDV0
HC+xZJNjE72V/yrJm9RaG6bMEfDH52R7ZMjMCpcLudl6urr5gy7aj/ArF8IaTUIg
SPC7kYXBayNGLBpH+6TmozTb9ahjHM6eA6FL80I2cVBkyNYlGYoOa/X4X+h3QNKq
GJnW7c8j2KwrwlIvTIcTJi/ot4vFlb8JtKDGtOxxuuv+AKd28Hl3nZCSs1lj/Imu
bC5cM7y2XXhh+l0zl0Tnqzzhi7ZIZgQkFRlBLuSdlLPwqVX95YuEkhnS6dpXG9OU
gCBgGPs693/2XQnohR1PMrG2SbBYGAxtz3q4DMYg1JWtRyByaf7LCyNveuvkcbXT
ZjCV+fRyTP/pstNaxDNEnAqwXdOLGuulORqY4vFhhW5PHBlMCJECVFSJnwnGNut2
bMLM4JZq486ED/7pBrwoGIfDyPgz3fyVYrCoJk8MoX/siRGkE31hEF10yHVnpX0J
UrcCcpZ4B9lLYTmVVYUzun71wAPMhv37ysdA092ZGm1UyK1ySVWofV3kguRfHF9B
4arhsYO6yM+Jv/1+0aB3HP2qICE7tOi0F9JaAKhAlI7gjWM5wJcRFq6lCVKkeKGI
y6TH3MP2B6wWHm6n0MHnncDB3evb1iNvlQrGGO3eVnayWxPgRHjMahcuyk0XI388
h5PX0GPiUQkz7rYKsq79K3EjGdwMIHztwMzoyJ44Yrnk5kYBejmdCl9dLK7ISqUk
aMPBZsOIxU6VfePjYxQm6BorqBJgdRZ7YTesN5fKPyadQb6ogCOgItAveapciZX9
amBaJq4Z26BN3jUNgzgTYR0Sue1iTJA6ZxzKHGGgopgWkS5t8Yp8N3rb2TP28Q/I
wAb6bHDSfP3lWqVSO8ljtSkhHbEFWN2OoYxJfwADeUk0Of8YlkVBeUHkpGhnEv50
cVgyD36ONZhV0mqXIIXp/ULukblmdJ5TKymTH/EbowP8FVj9LChSPwBV63D6yGwI
naEEFy2wr73euiNYhl8CfA9WGEQ5fQbN7do2GWZsuJEwTehc91949YGCa3Z5ke1i
2XlO9Fn5DLknTUc1oOiy6Yc22B+EHvO4zj4r54oC3tfZb4EdfexSZchOUhs0/ShU
GWa2YNPKH7+VhC9N9eHleV6iv6yKxoLO6H4ubPKXvOnGXVWYmEzRxePEqGI+jmac
Zve5B2v/fEfYcaBQxKgrchmb3SDB36BsPdEI4+urRg7ef6P9vFPExyxaKVqvGD0q
CrzsRgkBq7ExkEDkDSlDDcUx6CciNjlInMyLAc1xZDV3flJ3AXZOqS06bF2V1AA3
E0ma2ZliWy83Pz3NOuRI06C5Vs2jkP+y9HkBYXNAu2Y4Et4LhiDIpvkMjN8AGc9F
zZS4jP/+DJ8ZCl9c/QCf/D4Lm3U5IsHJ/FU5ZmSRBstaofxczOUxT3/2oyk8GRyM
xaz+RyXzwkKA3C9p1Nruj9EVMDMPTA6nmIeLEt3Utd2LTdAegvJlNli5ZrfUb4uf
7gFNrgXCgsA90M2/ODqYwzau7QYcjpBqFTz0B15IFGnjLqDi9RFIUTCB4D5gfZBl
JYXOrPAtWe6aRvNtKoJuqQZlwHtY4f7dht9t8+FT8SjI1L0StqAxj1k53hsU/u74
5kIA+KqVmlBeOoMr6pgyXXfZLV7J/RKCVn0xxyD3+1TuzcxkavBis/OKPahApxUo
nYwP9LmGgAUahLXg3R3whBCQIH4L0j2JS8IL2L78cGAmhpMQdKuFZMlMlGi82LTN
cNseb9SSKoXaSgKHSvKz6VCkBXT0SIoSEYtrqhPq7QS0VEz/4rYcvSWdABI1M6zz
rjMAAAJEBcyhuaa+0ihgOqaNFM0MmvqSlRAL966EH87wqgztxefcjzrG8TsVV5K6
OtQKNu8ltqju7fd/eO8RNp9tDwnROrAR8w/8jpe+v8xJkQv/OMyQI+/+wlQ7IAjQ
BIEWxstH/8L9qvtnGZ7HEQhCgZZZysZpbVpAzo3Bz+4TwuDLqpIL9/ltp446Js73
KbETqkQPBKc07rN0wn+dsWO5QvCdytNk0Y+WTXTckg4XcN6VDwTKsq1ZprQQia7n
6u53Im1Ofvxbb1Rwb6z/h1kT3ZERrHkH4T/mfoQ9vRi+x9/RnCt3dp4fgEVbMPdE
h9cMgicFSSQw43JzBIyrb6N27KIGNkJ9vfuwQtH1rWqqVx75eT4DAMA+lgJgkjT6
Ce9w84qnhl7Qerne2HmRH+0zVsSsVBD5bKRSynejWrkVzF3p1cEm3k9ZWTD8spi5
9585AWaa7iFKhblfK6pHEYLR6iuWBUpB1I6wEi8S3LaosgZ5YAghLPeV3jXqJpt0
W/btAXQUhagchtuM8xk5QNUXinUPB3u2hfedlEqYN7PZ6E87pH7fd/YeZoAc0OFP
OsFPg98qkn3LAx8Gfh+av3DEmIyU+ObJlIaHYa2f2RJQQbuKjon9bHyVrZM2f73p
quIgNhGw+7oGR3Z6CpamN6QKzXUykvF6IR1XgNKtic9IaVV5FKLZhSG/z+VSluh9
J4V1bTUAqfJxGm4oAzHnlj4ND60gegIx6evA6ZHvlXO/qV9W4ALD7tnrcoXOlGZo
Sw6DNEuN4C6K/97cWxBiC/vNqM+stD8HqVEyFwoiEvE3BqZahPUnaFpYnaPr8F4Z
k7j9iOE1jK6Y54661UUzAp4T4NPsAbRe6gTwNVwDVdeASwxqTcg/qSAUOmwpWLO2
pli5cOzHQq6foo2WgdILJINbWGMMns0ikdxXC8YdMKDZ9QumK0JkNU++PnbJXtaC
EXNAHIQ6pKbM9dPo13qcPBb5lKgF120V8DK3pD17zouVGejEmzfHlzhftCxVU3PX
U7FSvxdu5O2oShL+ODiGXOTOCgeDAa2r9JlrZRSLyr3f7jXou1fGQx1w6sfk3Kv2
7cUAi0NKh727cqujko351RSgy5WMlTC8TFL83EkDUvu7pUfhP/KDedSDsbTQPmql
VQFsotQTUSIEXf8UCme2ltD5hYRihKyAQxsuaOhN2It0Zbna4v1ictPw6Q+9il3O
ypx34dlDnuxzBjAy7kqiXWMF7AamdNNkkEQ3yA2UokP3/CL8P0OuAlaSIpdzjyzO
aJhnoPDvpz6CNEUf/aO6rRuxgz1FGoYL23oGWZ5y2UFYjMVYt8jRHDHeP0b2zXEu
wPIarrurMdOID//0LxdIXmRyVmpFRfjeJAbma4Ag5pq5LqcCU1hfLoxyVUTWAgcQ
jhiWv/PEXpcfQTfNrfo64siUflLgD2AyU5GIrOKusC0OMz2ILBEoM2xCGYi4uhAX
RSucqbEWE6Lefkpty9VSE7oPbHBKUCUeIH/e1jzH/Fbrr/ioAL8qFqvPI8uDmvIP
ky6S1FSDOcbQIa06UdvM1RVb2ydgAqwJewtRXUZZwlILKlnRrDpCqqre9OAWx009
P1NMI10Iw4wopMhC/g54hAiUNl5Vgirrjk5TxBmpoz0RP9RO7lnJoiRf2CBJ5THj
8LJBSQO1Ilk4AFn2m1V72U13ByFbYfpqJ3//ShVW6gEybggsQslW25ccISVPi6Rt
p5GtaLwXdEk5oQrWX/kjVxxtCYSoEmhYh4SSoHGpLuEykstIm2UJmxyXmchhlhyB
cMX21xUk0FcNcLj4V6a+diljbz6H3eiscotgSq+pQ43Wkk5gAJ32JtgnovvMgbKE
AyuPLe7I5xrq6WYOSBeQ/mqRFwkTmhkO7LqY+IN7Rn12W1wlyTX4KgBMBSBFovBj
vBtwcTIXRPJxoYwr8NyHNAxRQaj19k3HgMQHQkkPYyaoMD9VZgYfggE7u71VoZb9
GI0xHtCvmmk1h9vCxlKhjmq1ivFpLG/BAq0PUkkXAUzI7KxspaaePA0BwcI0LtyY
YF63u3tvljI/W5nsM7IgZb3bEY0rqTMxhzdpu/DVwkQPFe525YJv3o+W+ZxrHbqA
yWuK/kUsUxsYC2GipidcEK+EAO/sxZaN+JFwXsWjRinuKX84Ce+8XorR8hLYPudR
pPS6uJwP379zxVChm1AfQ2Ek90zvP70LISLbSLy1n031+opM5IghImgBSM7sbKxs
r0rw1owD2pYdaExWoCLZSdBiXjXjiOyJQ2UxNVOZfHbfyl37Civ+22DF0qXGI1/U
+otBvbuCA6s6TrP3XuPkCD/kTQ9QYARWw/4acFUVIM7z6JUSOZn10790IonpzO9a
3QimCEYXU9h9FeNQWuGwDXgChz/sVtDXINjOehi8PT3/oG+R3xqzY3lN12HXbeXo
PZY4vKCdItIz4Eh+dhIrcL8kUHzTxr4I5kPbU653003lslKHITDzrJZcacJHE5bk
cK3oRw1urjhgQ6kh39CrQR0t8T1NHpnout6OWkC4Mlur75KOL+iVmTY0H9zKMOJL
kO8YliiGue5p8ed+HCg0cmhUbDTuOfsxQEh6Pd2mm3RMYxJOhsc+/JiUE0M+GQw4
vJW8C42DEs6T5O8AdvLevmMn3u4Ezq/6EhujA47PNr0p1fIf5D7YK3PmUnLPyeyV
z1hUbaOz7QXqY7fFEgy1ni+uj2x7WfwO0cxQr2jlFZ1TUa/5H+8SLM22V8E4VvqM
1Lj+1Qhe0w8zcg+GlZmVUjx5KWhjyVXOufHexMPLBHTmqo6+wutaMz6p0X3n2K5B
6ZtEotQKxv1eTjY+mbBx4Hv/LIAMP9p1G+uBR5A/YCtrZdzRgshEOWLIEN+YLEI+
QIxqb+NwY+Y0Zl1jMNsZBrebUjkL08vB/u5DOSYQFLKL916YpgTUCJo07W4Btl4l
DN78yIBR1ZNXwkyWx+FkaNioIX3jqIIqfzllqu2e7cymTlS52/JCqKI2p+Z9ur8e
NXZ5Shgyb9a01pj/LWHUvAovXprO0X8bA9F702OycCvIzJVXqPoGvLJpZFD9XwcK
azh1eVAdIzgeJXtMAAk6kk/L72Y0zLN9Td/4CBw64RHMspiKjv8kxmdz+bi+miwd
iyJJQV0cLmUcVS6kevmCUv6n/EmuVYcwMolrebw6EAS/hllpdpIbxjS+PKTa+KLx
66PuDOxs5J0KnqpTbxsWnURySGw6m/TIGytjc9L82bQX2qLlzlFhHWRxAkd55Y5n
sZdsePHab5n7wxm1foOpi798T2pwrX0DxtXiatFhuVcBfn4j2RbFqE7M5iR+69y0
zFZo7BONZs1L0LYE9x1BGQoUESyzFk2ErhzmTkMWntchgOXaWzdWKw1N67sd2IF5
4zzJojfIeL8u1PQRcx3euclT7uQRPw0lj1HmSAczJQRYkc+ordjKm/4pLBD5ZMT/
ei8v0xU5QsV7TseVzLQscFIDYDm0jzNaIyG3a3KlaMwKtSNhpzZxZ51iRUeV4XGT
NIPS0sGS6w/lOpigiRR7IDiGSZR8Tk6H/22Y1v3ukxHM1qa03CgBXopW34OF1Ko/
IC0tZNYn/3hsAzM3c4NN7wOfSB8UQhN4jtu31x5zMCIj4RWns7D1K5mQCoKrzapk
q2VYhCtdoBzaUb50Ki9/XRdt1kbULfId65f9IvLdFZwVlMmv2AgvLfZtQ1v6dcHR
l2w8STvlOzxtWJru8y+LT+ZjgvSv/8Azk95irJ/1GAbd5LxIWw2HhKVz2YiDiCBB
uBmkJ0ukFfjGBBsYdgi74WUJAyqiNr1lCpPUe5jw73qQj0Z3xOZROxAhO9YEt0rV
3oFuI/I3vyAKzEVKpx3gXCCDnu58ruc4cBme7giojl9YgbAEUU7WNeSy+1Hoase3
AL2VmMjvHzjw+09YLAe49htnHd4qiUxwtOAukLvdLAAFabn+su0LAyBM/zKw/urC
cMzHCvgc5sOeJRfXqZEu9biYvP9BBLbXbkzJZprwO+eWRnOYgi0x6IVoRY5Uw+/I
0CEL7xy6pNnxrBnFa7c9kzZuZhA26lqiXZHs0uHrffzzGGbjJTqHJAxpUlsGT6mZ
pN775IHmxnpN22aGK+9cDtLkvb82zw6uNqW8oKVZTnjfemco1yPRkNjtJ9GKBep4
BqsQBwAg4tICtpgE0Rvjdak6CFlMDu4bDM8Xp34sagFM9eEC5JAWYp5U6oKpU2I+
mKmwV6VluDBb7XaEqrW9o+XUif/oWqawN2cDGHgeq0WvcxGQPidB34M+VkOs9OyO
mzn+/GJRtnZmc/+3nQ0szb/D05FvaAeClUwQCiV4OD/Oscqkv/Y0N1St8p9QriMd
TuItG/COPSXxK+PVG4JtvZMOY8+zro/VCK4DU/IQpDU1fYjhAFph76SGQtYYy+F3
hQ8jvhHTlYA7eRfMHI+vDaRLoMKyMNYih/2ASGz5Uu2ilL4B+Atb3BesFbTqqHj5
pNttpb0DCE8vWGCIy7CFF7AF9S1340MGmn8iOgUz+z0FELUsCOB3jF5XXwI2/w+Q
I7V0NM4V20EXhVmqthnoTD6VwHbgL8diqeY/FkevTsEDHk2R2B/80I/BxXvKdcpY
rAH95LwRIqcZwCHS8CKTN676ccDXHcwWd9VrsDCSP1oWP7qj2qjvkH01UAabovVY
Y27DjWJUIq3zrjqAVs0FgnlGaBxbORQZIuLpMEhzvRq63nP5roWYJQMd+gL6aUox
Wj0EYilZJPM2JdyuxKxDMPgBYVHtj8A9q3iZWqF2u/pxvPuYrTY2XvEDnPBf7FRU
CotxJz6Lvj8hzcrPfnXpm2Gz9nq1Yu1zAdMQ5/9CWbkDMJ6BHhFwBK41SDWYe4Sx
cX5Nxg+dBseQibXlE61RJG0Jn0jthrjr/c2SY3Ej+i6QJGCAG6VkLzCYMEk9qHoM
z5DgU3IqMYJR+63+ppzO6Fxa62EJlMtia+j4BsY5HDvyBSmUcubLyGBXCyEuRjhp
50GO/k3opyo7jmOVmS7zchQ6fGDfC5DLwf45pfUqCxTLHslK2x8S689SLQTMaGJx
DM7JF+dS5DX7P1Piuk04A5wRYUiPu0QDlxejamaIb0UIDQrHEQ2D5hShPIhOJUD4
TmP46Ioxa4anyFwgVrTqOwtWZfCMwU0940POAO8CbaJyXd0FzpEEzJK4V09qlJiR
F8VunyVzat1CSeU8AmN7aJa3fo/3vv4F/JhBfPvmBm3c56NVAZbnrvlElJUd2JBo
MWo05PmR4Eyb6AC0idSpCj2Tqb0+j9L5GHlTsVS2424eJqSP/iQ7F8A+EP8KyLfm
/LNnQT6SJs7igw0mikkZBD4JjfdqYBTsuZUU6S7ua5ikuHORPyDMCfbjhK4GyN9d
xDskg9JJIlmv/WQHYEEk+vEoSRDf/EX7Y+f0pznM7EfgWXcl47xfEdaLWNUx/SSG
R3rntWRh1Dz/KHhT9AcQS4523az3/b8ok3E/J1T7kMPyXeOBqdjf875HhBRYSdOP
uV76jctUjQCghDgdM4LXPRQKHRU+cSRfEYKFdz7EadLHdAjgokvSu4B+grb2gdHO
ep6q0Zs6DE5mYJ8ZCN3D+/7zi3J3aF7sJNtUU2DdW/O9hNCIL8GOoKUsIhPevoQn
jRJChosxVHQGRwT32loPwb+2umbr/eAbomMGZLyHijb/f3mUOYi43rQXo0qTMyBL
n175AhRDIQAwpANxjm1vMyIV2ttsxtKLHi4DyRSMq3YrqldSqj3Ns8vBWgz78hNp
kavpPObU0+RO3yL6T6zMAgrq+8dxEMNI8OK/brxc2Ip1lS1DVcIDxNo48o5olvac
yFe2uZ/P0wK0K43eF3Hdft6rR/gua36b9n6NdDQzhkujhJBJeAkYr/awDv6Kddw1
xHg6tbB6V6JCU4VPmCAh9UCN4L92HFku5fQ3l/GZ3WXz58bau7hqrb9xNpK9wg3B
k4BWb93wYnBAjRd3a2CM7sXqMBoxCzcO59h/NLS5WgYUvqwzOJn2QfaiBlKzoqzw
mFMAdiC9ABFQZSA7rzj7tvWFAAS+8nt5oexouWEFn+yPwNMNBJl6jMZE6OwNKrJQ
pgSwTHhNSu60ANyOO+HD72jQN8huGN96ZE5V1pOpQwC/8RcE4IeiK/Yg1MmweQx5
JNNBuFpb2Fl/6XxvszmHYeBfjE3sVCbQIoSwDKkungz9pquB/MQVbng6VF8trKt1
NoWmSv7pPuooBi3eUbZlJ/9/GT2idfQjXgrTzan1JzLddlehqveASDhgIsb+TTDw
bXI1IAnRQBuf8RerUMbVIOwB4ZGhTyCwfjQNcaKyUlXsrMaAr4wI9JvvGFXdBRhD
c1npAkhukhIBTp2lx/Bh1m2LNe0iyB8qBm7cbIX1f3PVCyPF5WYcB0bTtNHyqa7c
cOjrmbAi02ayn38S6UNgEC5KOZwKOS15bPJsDl/zI1V94t3Rq4SDoeAu5XPbdvKM
gyKPASGKjbIL4fga/xouWh+pFYM1Ohny6euAll2bUMNJpazyBQ87GH6AH6wm/mH4
cU5eT2tM2rbV/esF4ve1dRTatpocF5YFFeUS16n31Z01W1lVIjHSJsnFHHRsVXt+
wBlEngvGliWeG2WCjjP83NSJ8qGJS9SjSjz/+NZT9qniq18bjOqrkgcxyeFY+wc3
DrGzcopqRGGuYXywUOEDlWtpNpEk7M8zk8C/naMW/JirKlR06VPG/kYPx/qgFPM3
T99nRSGs/5WIG15K88u+AVdNpYgr1N7QOqTthD+P7EwvSNzGQGQDpK5gYG0NFkWO
/Q67pB3y3TZ9hYVW7lw7FkQ1yf0boWrDt+Kqj+k9MIl5gbTOTZ4qTXz1m/XO8EXp
oTp4BfLB0TotIYGOIfY+6rshaVmLrvvtM7s+pq5+uYAkJ4sUp28cc6QRt8Tzry3N
9x5Y7y74d3HTizZ/FmZcWT7gsEHrOtELw+i/VYWyfFenqxzlvxug6FAm4AJ8yqba
bkhQEjpO6cAmVUckRJurmOE+vuUDJNjJxz01gyRo01srVrC+jUnL2i/vHnN86MCG
zQKzXgsiWrwNFD0VrYhvbuY2mMn3iJNK8aTmqU0IXvIh66h2Q/EsKC2L0iOwmBcE
moN5pJqDg/yiWf0oZACvK5P6IOez+PF/QG7z9+BPREuOSRMYxmCe/dSFVVqoYoeZ
WXq3Oo/kEayMux/FfuJZHNgRWPBe56/5ZfCxN+E2oHs3fekgM8pFOh0880txJZSy
E1a4eaIv6q/oNyXWM7bVIpRKZmM+QhNuQ12bLGp26Wmqc7or4RrXH0yQ/9AeyZCz
swWy7oZlCbRoJoy4GMrtPDeDNoHstklgXSBC7c5lkXdg5OArF69/3bxj88xJch6K
EoJdW5HjAHkMD9GcH+kWog7Cc43KrHdvnlJas0z6CofMn3TUX5btAVX8R4L9P/sj
Bnle6hRJ5ClmoSUGEJ/g62n5TUBNn1nqSVVtqNPeJTFeZjecwEWDDXZ2fJWr8Q53
45igMyicPOSGqlL/9FkPcd0EyRucxkSlmfRd/zTs8D2/abXX7pgdFEVF7f/KQz3G
1Gd8Gii2F3oXNjnFbqCI848tBxRnkbR/oVsQwCfnfgzG7QUTR577vx6yShPe3ynJ
k65fEE1Rvbmh6Z6UXPpqs7RPT44n0OlUjPgyH82UdXFni1PTX1aZpoWz/N3s9oAA
SASvoJ51EkvfBsmgyx9VTCAWw3K3QI8OnuUx8toaxXeEd0wxiTOXkPa1IDyUkeWx
S+JdjXWQW/ksf+gGzl9beeitdazOElZ4EBsTdePfRiIOr6fp9R9MGGkhUM1+d47b
T92GfU2AEDZGWJZRvpdJxSFZ3pqY7XrAC/zMj4pXQfVkCr4mfWRePPedz25jMMM7
r9XsJNeHbCuk+omBDlYeJaz7jnkzNVcoKTO4YTrlxK3m/cmNxQzDMcB7uVqJxc0n
SBm0kDtjatFpyjtXsNVgPV+hR9yMzMzzT6g0hKcf3sh2D2obNoZl7dyATaF2DC6u
EiwB8Ddss1XDbGnW6vzl/7vyr8lZYqyNY+8NirlhFDyKbftvnN0okXtQqbRuxuWx
BPCqaKLX+uiFyQRLis9aJNMThjSzupYBa4dRH8Nd468gHXVHKdUbIT8rp54iMNsl
aWlRFcMR7j/5EzNM1kSBJ4/9kLpVwbVKZQVmL/3xkc8ZFU+FoMFxexXzJ9SZAwh8
B2lVy4ey10yMdmb9L/DE+saqKvaSh4gM2HSwNe0rPLJtScNgsjfN+hjgnoAcjnJk
MM0CBYul7u22XEDNxgeTJTIBV4DRbZzDPR1g9kkYXSrTt5i8RN0D+tYNtnRTVtia
GSe2Qs+aSzdeadLJswzjmDOBcAi9tHUc0IfHDe8cgOow2Qb2GjJko2aYdWfrDGmJ
Zbw196DWclgv3T+/an9hJBO774/QpOYYB/kg9HOTJwtKXhtpsMALg3VHVJoutRRH
YSNo3tVOqMstN59g0Bx+6CEI+Xn/mSDs2Cb6naFavc8TBlsFu+edlI9IwBk17s4h
ZxslnyhEuTIYFxZioAXoQXM0bf64Skp/lw760Z31Vii333WeMeXA5E3zQJ6YIp4A
w+rjugj9yCBSZ40xtYBMdZUGlsrc8NWaE32AeGRDOfURjCrwPpfpQK6hlUf2Ah3w
4AzeZz3ntW0Ek6XnlZrseAmiAaYtin1aFzPsAn0Rws82fHumkkxL4tIUlTCpIYxG
SxIkKWXQDhw7kvQSubGrx+tZoddGOhNGzWkq2B/BNa9RRdni6Wx4kKVCRadrlUTe
wcfHgqq0Mrrp7psMqGP6KspCQ18UTVUqOazU+3BSDyouGkeDf8LriKg21lHZV7qs
QJrIgc9LL1FTyNP+sGoQT7CuO7E365C1DTR+p2TGLru83zxrkD8fHDGn5EC8k3sM
vsOUN8tan6dekD9modc7Wpri/QBLtpqLVob0fXlT0HMcPyT13OFuwNW7cwRDhZac
hZ9OKmkk+QeAqizNz+NpBObK9eh8pF7AVROXup++FiK8mj680HnE/MCFQyUliq89
EmCLn36WakJwfz7HjbOl/687bhWCgrGHQ92SIQrJq+NInaS5uMI1QhTevhKssHqV
oqgupTq2+mnhLmevKniDKLPkT/C9jAF2fZu05dB2z0fVtSI4EOEB3LBVX4tzo6Cx
0K86ZCM3xdWWJHMB906mn16WZHh2c9gCHXow++RB60CfEWy6Ndv701Qrp0mi12aC
LtKyCohA9e9Fqj2VN5SJEqXQ/Vp95kpD8QMYbHlOYFXE4144d85Z9STuSI5gl4Vq
nuQFYuucO5wRLxZ88HEF4cL7G4wwtPxX1k0NF6x0G0Ay9/zao4waaKAaEXHB6u4d
pnNa0O7fALuS+HzCEi1N5YXX4Xynhlpqe7O+exncpdUI/VZicYrhActXZPXkt4x2
lR+ZKPBPH6nChF7YjXQ2xEnQLXSzYLAv4wbepVKd4VmEvTsBTCSg4OLfzJy1gjz/
9b53Ve7WjOgDtxFZA4JrnuxqmCp+TAolUBT+YNGbwLTlefSkEotUMTzmf2IiADCO
xx84l77UTqbW2avsuBsH1f7IQDH6EnqLsbRf9kVzfe7A0BqRYxNiEyOu0haa5CtG
9WcLsW41Z+CJC3u52TgObqe35pDCaNeN/JAPNAAlmEva1F2Aa4jKJXwqg3XW10gZ
YLyCIF4W6zLDepVByikvNzN3QT7rJuO90Xrc5V+3MBlodbpVaEoWuQvCtOyLfuY/
MqkXvEQPx3NMEdC1gi8YrkNlXUbb/rIGrkXzM3UEhzl8ZpdSyG82ktJ4kR1hPGHL
K2/7wAmOLVMKdYDynzpCw/gvq5L4hwyIxkTqbg4+juRfPH3yDg3Hy0jgjV5MkfXw
ScwZ2OwOXY3lZ8aOAyj2kZz5eYy86OW3HLOEqciuOBKWkl0TuZBzHtb99zerntHK
Pf0RvfYjyDOeOMKYFAukGsTBseVl6bM2rc6qRA1OXoaDMPQQUP5QX7i0NiTElzzd
3KY8ZbMg1HJtXELO3ymmWUGSyFL7JPGLbKBeg6cF6/9swQnSrL6Ju0zVceax6K4e
keKNAc4ljvDMl4tu9gJDRazHSenzS0cmBhpB/WpkTfJliDseIOcTYpijQFiHuEGL
sEtVPif2LFrSe4HxkeAzN/6YYtIQ0SWESFFNidit3oYY+gqWVn0aJ1G0wQrtgPH5
cAvcI14OsaNZ6DkoTCwSyuJe0b3hX9UxBVVr1SztR0g3cgLRgTQQjszOOtE1BQDX
bi9XP+k5zZuv8y24v5qCCxY7amsp8qK9NRPG5gA8MvEYWX3a5mnDjk+pMOLZs640
g3piYqgDrRi4ct6Eu1KJLaRH7uP3jI8HZlv0G+kcwUe7KSHXNy1KWjmoW4Hot1Q4
fO/nk63v9m1dcluW81w/xHF+p7onE+KzVYEjLdvxgHhpKEssr1LunUdfCn5U3uzM
5XPz8DoF6dCTZY6AU8jvGlR2Sr5Uj9jZJ2Z3Wh3gWYObmtiFO7+oYH33bGTFm2Bq
HThqtEiuwA6jha24Sz01wIL26P7vP8RnQjmZo13fBKq3qFaNvlt36rT76gAmyDiq
yxO2dwoCcIzDagHDU9xBlwEVuPLefr9TSiaHPB5yCZpyItY8SDdOatncCq+L5YYJ
VR1cXZXLd+a9NevO+tK7puN0TEo5MJMSp8nE0OmC+TpADpKn8cLnjTMrnRcCdwdY
wXbSefG3dk90yTIwDbXTJND9a5gn7MBoVMuQ/x1VAsIl+d7h8iC/6zTyJyVJcS92
MKpf9TkEk7AXihIAdEDy5Nk9Cz/RVCY2HwJONBHLvHa1Mbt2Jg/OziLXgrsBDsE/
Dssamv+ZsGsEUdsQR0Tjvs5sm2c6nfrqn/zwm1tum9osMJcnh5gd29qkwPyirBgW
h85NMnGp+bQPUKRkEKyPuZAqKRIC6oTWg1jt+UoLiBWeGxTybv5pTY4L6UvsxNo3
p09aT07IWZeKvRIhALG8IDdu6249I0zUZIzvaFSHYXQArSQ8VtsCMSuAmVB0a5LS
QZorl2dlVrQQ/N8rPIrYkSl7vKUHNurInFbCb3XPW+0hAWoo9dNwTDne004FN3mV
AzLwxAlrvTyB6V6vELgrIxzbpKGGrQyFXmYgeELe4A5LDgtj0IOG0p6q3d7T0909
rFEeM2mKmCBuCdpVb0Y4wiuH6e2bQkxle433aIDHNM2MhZK1SlLD2JSfSbU8w/XZ
9OyX6+a8AUtHb5k5FJt5c5STO6h/ZlE0UXOyd/P3dHKCDolnrfFGx7TroJICKUDs
RfUr7Lm+LRSwXiJuwkKbGuGvmC3MNy+aN4cSebEu2QFEXlnguKJ9KsRvmf17XUSX
9vRNekb9QW9W3LW0KgK/DDR/mtv1AeEIUr6v+Bd+EdK66k/wrLKiLkv9rEBGJApV
C+QTr8l/1f6wm4VUADoTToMtYjGIGALYoWOPeSaM/jdhRYMwF6JkpNOhJ2akN2Zt
McWZFM+SDzOGCGVmmfLZXF2BgUPlACWFJEhmvFpExbubE6zR4oRYq70vPk2y+3BB
1zRkaZoaiqby5LsBMtxQyKiGqddMxFuHAYvcoXE3bbVIa4wKemKG+9wPvLzl8vfk
WYkkBOVHC8zfSj107Ez1zVOp+M5Y8A3VOmWs/+R2Wu7Bj6U/rA/LSWbpN6NcZwQK
bhJEbnEAfG//Zp/6fcWcXT3fphYlXwBOH8VobSFX8BKRcMBpby5U+HqjrdDXdYhV
jfhNs8rkb+YW11x8dMuulG70s5wpFafoPL9HaVpIObcPipQWdjZ+ZWfIP5hD+dg+
+SltFy1euREEFA9HU2ww1Ns1kvhY2XllNkxwCvVAyuvKLngiRacj7YDkq+22DDYc
UbnHmYlrLp7uPq9R4n2uKw9CNREqLf+0BXVa/mN0GuFtqd6GOREV9QXvr6XpkAEp
GeWS0KXmi1/nc1W96EAxh7ceO0KS/zWlLcPpmEJ8HAiww2EI/qt2sVSlF+rTRsEl
IEh21pPRonvlzA/LDzne1Z+Og5DBZo6A+Eudye8FlttuoYByiOe5H417WFkK89YS
4Z1jgeCiS0yvXsiN7si6GnpuqI5GB7tyKBVQyPO7kBnEDgvnbPTx7MASi5nfzPmY
UCCRUIC4YjfXfmJtLU3MOkaxxBX3EbCYmQkatD95V6b2WAeZRRBb0XfXoA3vCD3K
a1EPMusKpUwTwwYOV3Vf3+6jPa/uN9DRPydc9NEbWHiUupDWocf7+vJIRQK9mnoY
NF3WxIRpbKEY9wMRKSDS7DbWVuAMlbj1vch4T9PqXW2tnIbcSmKWztPYe9Ch3ceq
CLZ9SazXB5j2FPEZEixUsfqRkjHPfioad79kxAGNLR218CN8kjesxrFhYZD2alRB
kD6sKOGoUSrPy1FePBZvfrNtEx/yAXuyHnXsPVfefVy3hekuGoocSSXgWSclnpd8

//pragma protect end_data_block
//pragma protect digest_block
SdF9wn3TktROpWSPiNzvevXToHg=
//pragma protect end_digest_block
//pragma protect end_protected
