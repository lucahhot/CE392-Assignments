��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_%�=��� ��}��v�����L P{u3��_�4�]�2(Z�kB�2�ׇ�T�fay�b�=n��p������1�w�L{+�+��b�8m�Xm�eذX�����Xǆ�_�VCYx�"w��Lȸ�f��:�h��^�3X�5F�|�����.F7E�ũkF�IA���&)�6�G��D��N�7V����Ou'�,�~�ݶiÃ�Hb��Q(�́�<;T�4��)~����ݣ���۫p�?/8.Fa���8�I�0�ߞ���q"�fDT:�[�S˵����U"R�g���<)M�hM�2�&�z�z���~��Z|����z:?�H�y�a=-��Uٮ{��[Ԓ���O0�������
��U�<�N���9x7u;�{g���ͻt�[7|\���6'�S�{k����d�qS���A�h]ݙG�#�ͷ��btaq��a��1 Q��4�'Gl-����)��߸ $��9C,qM{����L�m�9��D֧�!���,���v�-ޕ�Z��`���qaN<T(4����/Twl�����\��C����dC���`�1rv�I�w�,����%cn������_�T����d���^Y�s����H �J�Le	d��bփ��.�ע>" �q(��5�l�Q�bn�;�D�7��Q����"���	�mN�d*?�?|�>s��=Ǿ�tu�����ǁ07�ٹ��=Y���.����k��*OY�PҾ���T��US�?���l	��%.�)܁�x�E	�,1P�FO�W�4�T��F���Co�M*0{-�w��eE���	 �:�l�(#�Y�v*h���LO{��eSZxsXɬ�3�&���vj,!�dg�z\�䈔!�]
���n[ɣq2��3��,/�O�u�q�~�Cs1��,�h	�^{�]�ܜ]���Z#�������vXlz��R~��6)�jGA�f��=v=�]c�P������H�r8� �'��(�ml�5!��Ґ�Qw���XS�v|�aa��bt�;�&�)�I�SZ��L%=��F�������ۡ$>���E['�ˢ�4"�`Q���Z�d�]�t� &��v,b%J��_�ґ	����� s�A��i�!G�3�k7��H�����lc6XU�.�_���_��9?�fqF��=)ס�m�̱H*�v�/�����?Y�g�I6;tL�a����1ƪ��C�o�sEOF�`�@S�z x�/��a�I\(47±�{�x�%�M ��R=�@>�ߘ\NE�� �^[ρ�3c\�z�8�}ѭ ���>RB���c��+��%	N���L��,?N�e=M/���P��X��xw#۱G˞0���������g�C��h΂��ǋ�g�,<��g(�(�o2�Gj�`ݩ�_�a{� 0��=�������ub�nki���T�� �O�p�j�z	��r�nx�-��D"�b�FP�]���Qع���sC�T�%ԝ�P��0v����	ep"l�4V��g�8�A�·����}�LO�ײ,�wF��� !X	�9����mV�=jr��>K������ɧ@.
v��Κ�a#a���,dg��
�d��t�2��~dr�����o�H4�9�G(���0)#�.<[���Ho�̟nq�j�-�Vr�O�$<\#�Z���"(��B���8o=���eC�y$ �~�y������҇����� h#��j��hY4�?_zϰ�X����`&͗���qO^`��2�����&xq��4#7=±.�C�%|���U�	�����xirx�2�,"����H����[E���	��:L^��C_�v��AȖg\�l��|�0�79�rJ)���g�<h��5\#��=C�i��L�t�h��[VV�neѝ�g�]hl�@(U��S��ʸf�O�Q�Ә��]W�O��ε��z�]h.`z�;�d�3C���2#���ɥtѩ�KE���pJ���+�q�7������ul�ߋU {Lj,���ut���˫�:�)�8h<���k���;�b�+ҝ@���4��^���Dr"�슭���K�Ǥ��N6QArL֚$�ԡ�H�5�D),PW���ܴ�Qx��zIu�e�8���;e����R�^�R����X�K��i鄔�j��W+(%��?���ZVE���ѩ��*�V`�$��DA��r�a���-N�Қ�㈣_K��n�� ��Gk�)���<&:Ä^@EN��s���%FS�'�Vmr���4�ƫX����#9\�Y6.x�P����P������%�R�c?[p@4(��S�ݰj�Π�]9^̦7ш�F1w�&5^�7U{�/�3;��Ҵ8�
��)xr$�&����mk�%MR,���h�g!?i��Z+�i�YӮVT=G�`~��]��XT�����y�`Rf��IU��]F��{�倅Wx�BYE���|���%,%�k�o��l�֯:��)�r��J���
�\E�Ax q�'�(r ���w���7q�o\�DKx��ŗT>_2�poTj��?� a�$�=;��)����7=�W�U��O�p�n�OW�.�V�:���N�)��ٵ4�X�Bc]ωU[�*�P�O���}�HOl5��=�Pr�:����8P;U���5�aǮ�l2S3��P���Fa��A���1��0ˇS�J�D�e�Ƿ�<� 	�Q��.�:,9ڨ���0x�k����0��>���-'P�K�xkb�_��Uכ�sV���6�_��&��u!q��X諒�X$�����@9M >�������7,�UPI���Ppo����H�Sj�˛_p̡��k�&SI�<W��*�$�/�5�b��-��O#���E����|c��Sb���Ƣ]���c��l
��*EW�]n��w;&�AњŨ��8[� u�ŷ�=a�mƞwH{,D��� g%�Wi9�e�2͔ro�3nO����lh��V87CfS[���nQ�
u%g�
6:�cW��lH��[�:r��M]d��ӄX�,��>���N��s�ld�#� M~5O�8��)$��*Y�(����lİWu-�#):*X��=�nMeg���3WDSYÚc>B�G1F$������,�o�r
�� ��ӲZ�={"8�mi�Մnc�E��NLMpdZ�
�x9����$ub�������z��}�|+��GR����p�{����e��P&!�(bI��S���>>Ԫ��B=͞i������Պ���_{�n����?e��/�(q�G���
M�6}%t�]���_%GRG��uc]�c�ƶ���#����S�����1h��X�)��S uU�y�?����V�^�3� ���8n
A���W�e��*h�D��W�'�t^"� o�S��X`��QEg�k���q9��?���,,H#��B����H3�ila<W}�]Z�W�_PO���304u��������ۏ��~�|�۞ö��s@Y�������O$L�x�2+���C9���l�����/�ѩ�KE�
��X��e�_���мw���Q��
K���M���6t��/:�/�(�~D���^���e6�l�/�P2�l�����s�B �J����Dw�SU8`v`4s�MqYVcy�28����_��g�-\��	��OO���t�м�o%5�����3{�M{�)�n��������І �*#��dƚ]\�DwT�#�`$���ϧ �k��%���A~�̬`�S!�wQ^�p�*?���!s������������5�����7�H�Ň$��1�>���Y�a�D+�� v���3V����+��+ּs�%^�R	v�.�%�R��Pt�!�h�c���GS�AB�o�	S�\�k�]����9�8?w��|�ʸ�Qz�����h�,��e�[��}�ZQ4eZ#B V�w���X�/=C.�>��U^c��xy��V�Ʀ<�f�0\�v��
%[�3T�q8�&�J���$����8���J��ZQ��K	 0^8�-@̖d!�R���a.N��M����hސj���bS�3Y:�l����/x0�3~�:2L����QT���/��
����d�OJ��܄���3+8Fy�g~��1�ח*�Jd�Ҡ k�p��-�xy� e��h:}�ץ��)����GS�R$Ƽ}��)��Lrʺ-'��b�ԟa+��V� h��H�U���<�x���Ʊ=�����S��3�[Z����I��u��>z͓����� !����쨩�sWj9�C:���w�Rtܱݩ.VV�ʑ��-*)�+�.����lN]/������;uC�oM�z������H����!��J}�_b��ݽk�D�["��$�H����SH�M�^��K@���Ǽ_�dJ���.������Z���*a��"%����d��� W�<?A�h�e��r�}�"!���M�9�NVࠗ��<:ן��g�nܰ��)�A�<�\Z�$<(뵭���~�;7�mI]kv�Kbaz�i���1D�l�IoVݷ�r�:�5��s��g��gҮ �~�-�x���t�n�/5*�hs�r0�W�� ����ٝH���ԅPT�9�>j+�$���XH^~õ��{�re�J}�h��BI����rc2_�N�Y�����n��d2�͍�W(�y!��Y�t���<p)��7װ�/�u�$�J�	8{�з{��b�$�n�PHL� ��Z��B��#�%)cOo�[8I��C<�\~i��ƈ����ҝH�w��s�s~(��xՙ����y�l��H��9�-�R�e��Ŕ�		�955	co�s �?A<�/_�ܤ³�pq¸4�*�ܤ����qo�t�|"wϹ��gS��Ļ�1�Q�7ƕ�|�c��H������خ��s|e��ˢ�i8���n&�5�YT[G#�gn�
5� t�����ɑN����"��`������1�H���B w�z�`�Y&�0r�07s��Q�}�ì7�@�Èi[���W�h������22��hk���.Ur5���Ȁx��$Fϣ�C{?��ƾ�.j�ћ�����k��x?	�R8���o���V���GЗfi}�=�&�¦ɳ��WEc�ߩ����-�kj̄s�`��>�>��5)��yc`d�[0���^-��ZA�{b�g�ƛ��檍� s�\�W���Ou��Z�1Ѫ���2�eԽ�n�sצ���9�B4ϔ}��k��Tow\y��O�臵d�^�~���p�N�c��]���j�iͫ��%��B�:w��Jr��E��O��mk���i����o�
�#U���w�uNkC��ƹ�~�K��^�Uפs�a�7�3�(�VV"�{�.��a��ɾNgw���SwZ��Q/�7��)��u��#�*�+��{$/[�Hn4����U�ah��<���~���l_�yi�uW ����(�3��P6�'�S��߻`ڔ<�P�{gg �o��&�81q����̆�^n��l��2p�OYjL@ߜؖ�5 ϖ�g�[JXpW��)^��g'	_��r)�ykb�aA�e�0�5RY
h�:7f�K�o��lsU;�þUB�x�\�~�Y�|�2���8&�����ýI�|g=gr���iԟ6�1^O@G�X:��B�e�Â���E����\RO�NS��`|Z����ޏ~��$I  ��[�wQS)G���L�tf���
V��<�;b���H���kÕKZ귩���Jx?��ԙM�2$��g�8&�;<ce=ǣ��>i	����(
�y2�(���ڤ�!t�cQN�w�筠g���	�/½)��.T�G���I�������YB��I]x^��	5��"���T�x<P��|]�6�k�n��޸����[�s2*-����N�ZdqY� o�g�U��H������ ���G�y4�8Ќ��=��4�8R8b\�Q�7�`r�9YU1����r���?a�tiJ��=�F�5t�̡�R�k�o7Ł�*:0�h�����N) ��xs����^+i�ެ*,�a��}B�#"Oܼ2�c<�,���2h� ��L����j!�n�!�\�E�vpkc���|��HH�|�Z�&o_�!9k��Tt�[�<:�����)���q@d���c;1��tw̖kW.�N�1*��LmQ��}�ck��*�������tY�m_ZA,�n�[h�'냽���b�W��1�5Ф��%�O-ۭY>',lͪgu>����O�x�� �B�z��-�n��_Y�0P��A����zi��C�#ǘ#k�B����؉.��?�>���u�q���X�(�o��G�k�e��Ol/��Ꜣ�Վ��y{�@ɢ@h�%q�4�KƫP��O%c�x��~5C�(r<m��o+|�5�SQ�;��I⃆1<o�(#+AZK�_��"I��y��e)N���W���V��W=�*�����8l���>}M6��V%�:����J� $0�n~��F���&>��ԫ���Kgg�RJ�	F���Jr��Pn�|��� �t�م���2w.\��uR��0Em8"��f��A�x���%�����3Aя	�BA�-)�� �b���a����n_��������K�W�b��K��1��iK�Fn~
 <#!�3�0�����������;�A$�qf�O�O�.�Wख��M�����q�XT%����_o��Ȳ%w]D"hlńzN��<)�ڝ�/|C0'F�;�۰�6鿻Ym�&r�J�/�$�v(��>-�)����6=!L4��zt(��4c������,MaΓl5��"�?﯈A�OA%�u�g��l�??1"uD�p�G\P����K,�w{����slr�]>Y'��j�Tˢn�e�K�'# �x��
 '�l��T��Sۑ ��<Y�ݨ�����s�g��<�jiB3��ч��)��|�A�ϥ�>�C����DZ�vƐzfK�h����H��@�����#�H5+Z���d�G�b=ɗ�\������L�T0jɛ i�D�$�H�Q�Մ�dg�_P������Y$�P�oz��(�!F>u�S��i�Nl?w��M��(�"(�s�z���(��`�	\ n!�ѥ�؂���J6x3cu_,���5�"F�jFK:|��e{�gq;�V�����B�
��m�RgLP�a�V)��N��|�r��=�`U
���p�����0���:�B�ow[�~*riCZ�S���k�\��˘�Q~C�v���S�&���$��xi�+`�Z���N���F���_ɂ�F�t��еW�PV�;��B�Xb��ߺ�#m�;%�K����>T�6�d-�R���y��F1vӾX-W�}�6�le�,ݩ!%����X8!%���b��\�,/W����س�ё�#	�N�])��PZ�n�.���c{��д�Ͼ�x�Q�%L+^l!`AF��b��g1�7պ�8���\��-jM^�ͫ�եcU�;w`r�{�n�����կ0uo�O��<��_M�|�9��>Mmo���5�dsӧe]�� �lo6���6C�"B*N��<F�5�n��V]ڐe�K/J��=��7���J`�\��
C�����?��zQe���0}f�Be��Y臕��ˀ�y�uY3>���~�X�D���+3��/���9YsᲳ5W=̴Rc�:�2h�´7�ȗ�>!�6�F�0��+-̡8�0O��3�I)�Z68����)�*	����:,�����Z|�L��>�S�AN>�q3��jݰ��Q	�M?���{�1�䨞���*k�<Z.�����7�^���'�+r�P5-�}m��/[���*d�d�`�	�1d��z56�-`�,&�vw��Z��{@���TN��|�ƪ]�R��4+7��ֱ�Wٱ�E�E�+�:� j�B�CƷ�}�mF�l�c�S@R���� �yd'������.{�
��~������5�i�3�|�u x���5c�Lah��M
�]-�L�G>�aa���w�:UI��B���2rһq�^IY"z3K�i]z*Ѩ� & �6Gl����+H��W	�a8��p5{-��l�/���l[����F����}#�В��&ˈDI}��e u��;]ZU�k|�"��*A�+���{�k�Q0�H����՗W6��.%�H��x[��O�	������oa���	������хFߴr�kz���~���:�cԁ�e<I}�4�\y�E���������<��$�	�����'�`���dH�}pt�	�EK�.s�p��f��c��B�9W���h]q]y��*�.!�lw,��S_]5 7.��+A��m�$���tohj�#ۙ����s	>Ճ7؄-+�mL-g�ysq)��6�:����q��[�R��o�X�\	vfƸR`�>��x�7<:$ \�}��Nt��KS�^wOd��V^��wF�h�Q�ڿn�p�Xj@����1��J���ųM}ý�%��Ռ�z�������ۯƽ����ƶ����r��`�d3]=�K�e��[��d��NNe,ᒊ���	���ȉ`y�Q���R�l��i�Sٕ�$�6����i�<���I�/��\d,,��8(�vH���]nW�������u���eh[!�h����B�n1Nkb�<�`P��g�N����^��KOPx��ՠD_a�^�V�gR�)/���H����U�~Ւ9���/��?M�1�tE�Bf�o�}��I݆c�a�t��o���ke�6 =x��[ça�*�8���=�T��ɺ~`��P���z��,ɪP{'~�<
 я�\�����I����3mWK�u�u�}{9�ۭ��k��I��N\����*-���4�;����5���~N`�Zr^�֙���:Aq�K֛���(	�g�{������}_A}�Q@�-�M���_PE`�_���s-�I�ۮ6aYg��@��F��V���%s��zJ a/�\\���q��'��%�N+km<_}��cC��x(AO��Y [oK��z�,�8��Th�n=p�$�S������(� .M��5M�+��&�M����h�p鶊���Л��@ A`��,u�[�4��,���.��q[�]�����vnJJ"ޏEXR�E�Зm)�e����/�mL��x���|*7'�;{��F�O�k3Н��-��e��r9Q��xk1dm����H�O%5%f����v�㴢���x`�f��������B��q�("�-ή�Ҥ)��/�K/w�7����9��Y<w���֮=/WCJ>R������Pl0�:�a���蘚�;�i/j&�/�[$�dHd�aYF������B����[Jm���Bj)Yւ�jSS
Ҡ��)��3A6-��K1?�ܛ�-�$���\�A
����
aU\+�7��;��M2K�b�.7\J�l�Y��	#I`3�b�.7jW�]/
c�m��>�O���?�q��P��Z@�L߀3N%O���t��+���\��+��ԅ�ӴѸS��6�w���x���hR�����oА�c)��UcV�8�z��Q�1��`S�2Xo0���N�:V�5���_�l1�N��
r)w��_]	r���X]V��lo��G�S�O�H�o�I�,n����ì*k�D?)'��<�Q�����Q�_ӛ���{�]Xԫދ��cZ|�㝙&k�U��۷�e�Y� �ܲXo�9F���p��5>�fF��w���Lg��MC��S&�����L�	��

4���*����[]�'~�/��:/�Edߜ�lq�h7�l���Y��+����[n���p*�L�9�PT*���2ťsI{q�ju25��z�"���sI|h�����z��,h��&j��W�7&MM�Ε(�{!���/ts��~`!�ɥK�~�c�1�M��X�ZcW(n���G�=�V������5����ݖ��`2-�:.zU� +b2l
�@3�s�:�]Z�K����;r��@,�Z��y�)*��x"M����Լ�OR��������H����)��Q�Շ�����:���<�q:�W���(��+�+��;�C@_�'��/D&�a$$`��r���i�t�1�ڵa���A�:*�pF�������8T�3��2I-�U|#	��J]ޣ�1]�A�2�����4��I1�Ã������z��q^�Үd�^�'���,
oC�K	Ip�Ƃ*Q��w{�\�VпA��b��wj�m�5���n�����(����>�#VG����m�vR����Xe{탩��;W��kP��6�i��΃�R���ȋ��j*J{��Nleo$q�
�I���2+��X�d�Vu�ZK�N^D��6�}G\$&��j�F�	��0c�8�8Nz�~�|n����!W��	��n['�7�^3�����I��ѩ��]�������QvR�3��!z�*��]�:�X˨Fn�"�v�r��@]�Q"S����ɽ�-(��U-�V���;�
u�9<w~4Sk�$���K�r\�'��'�0�u�1��˶��O"_�ܹ����WX�r�W#�9��#o8љ�8�z[���@!n��	�G����˴�*8�A"�V�&U��݈��������j6/Vm��1_*����V��B\���X0w�4�S��~,I?��*K��.ڠ	蜷{����:�,�C�3�����wW%|��`9��l�vp�� �dL��%�9;t���rЫ�
�o�iO�J�D�y��{����A�*��p�m\�q�Z���!NO��M����P��%�أ�P�#�XzS�ko���T�y����>�+x�6��������݅�y��-Z�GB���9|�b�z����\��x��(�sF�J�� �}��n��n~�'k�@���L����)�ږ��EJ��FbH�\o� ����oJOaRۤ4�Dxb=G[!j�@�'�Mad������~ن�_�u���/<$cbp���,'F����'���Ƹ<x���Y�zow��:��
d�����Z�Ӱ����Є�����wұ�t�'0��(�b�ʸ����b��N�e��
12��)�Eҡg�`���oCD���s�Ԫ�{����3���@��&l���SY�i���Y��Ҍ��4��1Cbz*G��NE"�}I���|=c�����`/��y�@SI�v����R��P�EM� bᩖ:��D��z,�!��G�H��b�:��D�Z2V@��P�3��,.���J�����!lUm�Y��2�}�câ�1I���,Bٕ�4p�8�c�T�գ3��7���
H��;�:l<��5xA.Ig73W[*���W��˻���D1H���y�E�뭣9P-�ץ#�s��_3�!:����j��Q�t"XF���$��#��:X��hPDG�fj�Lpu���>�4����n�@p@��ǿ�>WX0)I�5܄�;�Z�@n�?� ʚyZ�����f����[ @޾�{���Ĕ��i�V࿰�U��������&�$��<v_���<#�ZA��y{+��\y�*�4O���̙~��ÇNsU��@���%��?� ��m�xȋcd %�?�ٔꦃ�`s~�4���|r�񏛛����>��ٝK���c��j�X��g��?Q�D$Tg��@n���=�\(I�
�h�.�Ԅ�$͊үz��OY�[Έ�O�����s�w|䯁0@m�#�S�9�Aٝ.�5%6�p���!�v����Ș.�/���Tr����Ъ����+J��9.���"]��;BQ?p�u�g�T�5p^n��A
���j��bI0g��Q�ʚ��\}�BK#�}�~�GG3>��sl���
�����N MW��U�,�k����Qv4;���E4<��MD���B��yR�	o�>�)+�:�A��SA>4p�K3�F�]�]"5B�@����\�C���e~�I�~Q��O�~�C������iP��p�:l���Y���!��4�҃�&���U�)��sU��}��?�oV|�g�
DM9����^ă^7ӕb\�oY���2��U���6v�]��u�j��x�n��)�F���^���㇓��
�Ly]��`�r���uB��8!�P�ps�%�,��� )��D����Ң�����g� �>��c
/�%���ϫU��?BT�j)�0㿰?�ق��lC����&�rv�7��P���Yn��|
$?V|��; �+o��M�I�н��T�=�aA�-��� �o�=��v+�˛s~S�Av���ƦS=E9��q\���N5u����`��Y�HN�BS�L&���@������+��f��+Qe��EŞ��x���brc� jӇp,��-�W�=U�,��ǸPU��(ެ� �� `Eh��<W�5�;EUI�T�=!C�TS:���A��D�������-��hZ�쳙E/��Έ~�A�\�fJ?�KG��l�5��RK����t���$�;u�v�&�&V���nbY�_D�"��&��z��=�Z;�@ZFE�pت���;���џ�I��'�Ij�D�
[M���>VP�:��9�I�ِ�LD\_ �^�i����&}=�6��8m� Y�"&���'���폛��}������!�)VH�R��;��I���gh�JsC=~~�dD]�cFc���;�i"ԏ��׿+��NȤK�¸�@��_X���M�Ь�!�C ��\����F���]�'}pO��щ����Is�^��&,��>T��Duv�X˱U���5�A�m��,�D�[�5��{g#�Ο`_�'�Je�pE�!�(�?��%��ڢ�����?p�@�ʘ?��Kx��~�������a �a9���F�6�&4�5Q����+��p!%�aȇXO��'�{�ykT#Xk���oO��( ��j}a&c����(��ei���8�I��l�>����M��q����k_��;�@z�����B�H��_X�= ��Bq�������$��&��d<q&���ًN�*�I���d�
�ö���/�OBKɎnLS��<E���]�lC�K�����g�7]�	�
��Az`ݪc� b��v������/�M��`!�����t�T�������Ĝm�R΢�ћ�9t�'������f��i2�������l#@ܐN��U:#Iēԃ��t3U+Fx���;��J����X1Py�F�����if`/��Td (�+�>B�����`)����+PVU��3����K��aT��R �T�K�����of������w�މ�����kE�ӂ4�dN��\B)_((�_?�x��F��a���MOf.�D�����9�֠6��~���W���dj������qH>���]�#L�Z�~�EL�`�^n�7Ք~,�1ۮ��o0�	�M�:	E��#�t�����7�x�5X�z@CB��!NDΌ7�d�i�0����~T e�~8^�T��o�S��K � �_K��������f����_$~��� ��617��%/��br��u��M|�eZ�QN2�)H,���^_��P=���(�I�<�ʩ�{�D�ya	�x�lJm� 	Vx|�ɡ����bIȿ"�F�* �'�[�'����m+5q�V��������k�P�(��ᵻ�t��6�BܦU��q��:�|�4��Wf�Hƍi��p�z��QD�%��۷��<;��������xd�i��Fi�����Ic����
%э��xAj���K�oqa��0&����;E���0����Þ����V�lp�u�߭,������y�';�b��Q��c�5���V���r�C���j&0�����S�U���꒪��@X�����7�Pාϟ)�$��#���̺G�QV�{����M6�u2�ՙ������\v<�9�V~{%���K�����.5��G��ݬ�kA�L�GXT{]DK>({��#����b�<cAk��@JA���۠�m��e�H��Կ֧�c��`����;{s�U�˝I�6��$o��&NC�H���wڋ5�#��Pӧ-�T�� ����?A�v�4��J�?�C#��@�@����l����h�~��ಟ�(�8ﮁ���O��i̘�g�R�j�?���cb|�U���l���������(��a�^F�+V�Ϲp�Ab�6�)O��SK�^��Mx���RyJaq��:c�O���0�	�B��������{��u�}��\����k̺T���=%tGQ��o��l��n��`!��c���5�8Py jz�f
�#&ƠN��@on�"�=S8���:���S��x\��c
�`����kc�\���i�C�S)bA,D��^�,Je�=,E���*�;���y�>`�� �? Q�� -1ڤ�=����瀈��,�{�]d�����r��ŶzZN�s��yU�$ }W7Ϙu�Z��ި�ڌ�\t���Dڟ�_�wђ��

�,�;�.�n�ߞ�T��{m�c�V��~=V>��y�ֿ��no�cɭ����5ЇT��<E�z��wNP8�+��=҄�U��{���yxz���Z���^�0dB`>U[c�h�r�����L��ƛOpX�������c�A���Kd/�|���
fp������p �!�X}Ms=�4׈�ʰ�p5,�`��$j5�j�9z��49埡Q����ї�*�̿�q��rPH�5
|'K��@�[Q�a ��E41�Q�dM�-#�H�L���9��M�c䜡��5��BC:���q9,��M'!�{��fn��\�o��f=|گtz�H��;�TO�p�Y�eۺZxq�?q܃���-�b�+��k��L��F:jگ��}�c2l�p�%X�o���V7�}=!�U����۞����L�{h����8�V�۫�x��~)X�˦�0�k��L�J�/�;��҉0z�.]P�u�EX>�|6u���q�τ]�ϫ�y�<B���c�Zg�D#D��G	���ɇB����ح$вK��K6���m��������t RNJd��@O$�o�RL�����f<`B����V����,�$�/���Ι�$qdeѡ��8�K�I���#c)$ E�|�Va�`�愪�@��ㅻv7~�S��Ur�T���`������j�p�w*������I�3}[��ݙ ��7�_'7I͒��?-���bq�Bn21��*�=��¦��V���/u�F�7˳a{��/H�P�(R׷d�8��mU���~p��t�N$ɉKp��R��keF���uv�����F��c娺ekǔ��&㾂`#"��*۷\�9��7�E�¬���Z\�|������0gx&q��{���=�s�`x�kq�ظq!�W�HCۋ��Aǐ�M�
�3�ݦ����:�y�� �ܯ���� Lˆ�V�oFq��dM ^�/��c�������U)R�*�Bh)�/�Ӣ�fm�W�C�Y�k4��f��E�O�2�-I�3#(�e�*�g �ن� �������}B|��ϊY�D�ѧݑV<0]ت6[��}��G�0�$a�P��A�����A�Æ����f��ܯg�.�=���<���D$�y�Mj���d��?߄ѹp��E8�x6ي�;�&����;���X�OA�i��9s��W�j��_l��q\��/�2M��s��vc:�f'�sp?{5D��ú<)�&c��T��M�$�J��%-�5ʈ��
��(o[Vy|�o�Gi&1���d�	��5�]� ��SUo�p.A:I�NB�beRA�0B��r����I2�A�:���(���?�'#mʬk����<�� �-m����P��3�Ƣӫ��&�\�,9�����ޜP�K8����w�՝G�qL��۩����F)�غ�W�7��A�Y,�8�7�D\u��uǬ�Qb��Ʊ~[��:��G'�'۟�O�\�n��Rߝ��46�qr���>;���!h�^(�QÉǷ9j`�e�'	X'p[���Z�[#�7 @��˂b��/(w;ݠM891������'�ʻ���A��%�y|���C�rsml��Z�񢓣�C  [x㻯r+g$K�Da�"Hnq�xXHA���b&�����h��Y@�We��$�U%�I���L�x�'γ��$��b=9AnO�=2���/l�'���fs�|�q�}E�S�p����]�`s�S� }�XP6��T����̈m�� ?u��W�o)�!эJ�,t����/�f�ӻ{}�5U=;�ق	�V��0�JB�N���	꨸@YB[�2f~YyGz�;�-�H�\�!�YC �
y�U `1wV�#��h,��2;G��éJs���S-4r-*%^l��]@�X�Ύ����*�*��c�����εo�U�!�4x���T�P�/4��Np��k0I��T�&�g&���[Βo+���e�������`���S�4"�_��4O%�?���_�n^DԿ���,_�c���8Q������Q�3�fIwJv;��5�0�DlT(���lg�R���0� �0��ү�Ʉf�IN/��?]�B��-M���(�"���x�%��z���B��6��'^�=�{��R���rKN	��d����c����� �P�+g�h�ӷ���f���݆�v�*O��\�Ie( B8Ft\�[y��a[�<�����;u}�38Yg/]���}p�*7�$ە���sQ����QH���c@�1'Z��^�|�§�>��W�ї.���(-��X��V�����RB��w��X��b��)t�:��>3@I����rR�.0�s�Gfp^���߯}��x���㛢�$��2����W��@���2�n�%`F��ݺ�q�:Ns�qo@��gգE�|���G3�%{�:�.�y�K�ӛ�?�&���]�Xx0�,�D�[V�p���+�o���P-��l��|%K��Fc����`�":��������O l��?N?��]���s�"K��lcW5Buupt�WV{��G��h
�8Y?���"�G8��h��u�7b��,�7łȪ���`�U{������L^�����;���}�Xc�u�3uGk/�?�r�M
���S�p�� ���T�h�@^y����{*6ʽN���a���=�kW�����n�o�����E��q�Ղ�z��JmpI�0'{�t�r�(2 �pjBȽY�g.ȰV\�hɞ>��<�v�b0~�@=o
�V����x:
?��\?kP�i������W�z{�.��k/KkK���#�1���kgݰ���ٝC�Y"[|�(�����Y ��)�fJ,�q7��-�]t����m��(D��7|���u�RY�����j�M�bKx7����!��:,~�^��/{���i�qnU;�ŵ����p;��# p�qq��Ws�H	&�9{B�G+[���k��n�r��l|+\$:BDIꭺ��(����Ϙ>�c�3@��>�<=P��,����G_Rw��NB1=��������8f0�X!��
�VCF�gm������j��`�8��y��0h��{#�L�5GŔ�sLp��.���@0ʻ��Xs�lAQ}�/�� �1t}�Cl�'^�
X��]S�����pN/�W�$����[�&�]���kmt{I+��=�s]ږ�o��h�k�Fy9@1:��}F~�{X�y���=����	��I1�Kx��2<3�i��$��`��+T@���y ���߳�ȅ��k�(�A��6L�$ ��jeOx�~W�|��E>�(�gY��n�
4��� {�#���6j�f�J�
�{P�z;	���k�A<�\h�5Wy�����|�d5�ٞq��z���C{��9X0m�L��p�s�Iı�	�F��&c�[m��"(�v��`�xY=�G�s� �F����&�7� �B..{r�Y�pF�*�y��\�h�$ff�ϑ��3T���KS��)�����X������oB&�50�`ML�����]֧F�v�����%�N>Ԡ��bRɶ��4.�v����� ��QN�ƃg,�J��ْ�'|����8��+m����M�ɀ�hpa���
kw�WӰ�K��VI�*����Ɍ/���3��D�	N1����z�)f�*�Oe��{w�I�֔X=��Y�cl�z�4U�m��pr�h��{�J7����ޖ� ��W���H����)gT�&|�k�0��ִ͚9ҧ�I�\��d�(9һ ~Ћ�SNh�X��(�7���K����c
1J/j��i��`�1U7$#j�Կh�đ{^:�pQ�Gj���-�7Θi�� [�����&�X��AF!&�t�;���ć̉q�il���w�_ڀ,RC0T��ݭ����t����#ԁ|ڂ�`?u���(�@�u��~U � �y�}�/�e�qV-��� �������
�zX�Fϝ{���x�GϷ���U*����g���zL���m��e}h�b�$L�c{G&�׃8��e�p�پ�MSF^����GV[�L���Q�t�hJ�:�p4�H]��§d����$Tr'2V�R���?
x6�p��2��b� ��6iD'ϻ�ȷ%m��l�����L�U��g�-�C�@4=�3�x�[0;�7��U?���c�P�Ta �+-�	{:~���4 �]�w�M�CG^*~td�L��}��L]ڇ5�S��l��q6��ࠡ8���7֞d'z^3��`�k`���p���#�YSN)�¾tk+�.�NG�.�$�T����}�����?�bЄ�=*`�~-�������С�GX*�$����D������@���S:�B����Q�B����{c�*v���\`y��J��������]9ᣥ-z��gd�K
�[3^
C�_��x$x�uH���DyE��t���[�[��	����v��G�����jO�~��f'Js��Sρ�V�gej�\�a��x��y��xS;5���,�R.����R���\0�:�ۭ�;P�^��(�	)�(5XT��JQ�T�'�(�P#��r��puqе�]<r�y69q�J��R!]tT�� ��e��e~���1���	������R�˪�mX`��D�K8Xf�;���-O�;(9��zb�W�:K��!�5�~ܧvǩڏ̨������g|��Xr�}UK
����Il��;R"R�	�LfaK+	��t ß��Nu��,�Q֨ܬj
)�:���i�d�Ada(ۓ�">3L��iT�{m�'��3B���_�>��#��;�}ͭv0n^�?�5â�F��m����ʭ	RP�%�a�ɸ~�j��!���,vk��f.nG��bZ>2��O�N��[���N��P�z[V8T���E�e:Z�^uc�U���i�>��C�A��ʕ���,o��ސ ��b���0��ڔCJ��+���o�Z��s�S[˃z��߅)�H�O�P��X�� ��Y�ܩƙ�3�8�st�X��ٓ���acu
���{�6l��_�w�9>�N�x����m4}�V���P_��+=��i)��Au��� �2�"9Y���cP��mxEe��>���dm�w�1���M��ajv�-���wT��,(�܏!��7�5^�b�j�Q�zr��`�u�����ť�r����~(m��t]�Zz ���aۥ�w�^�
���Bq��!Ϗ��k��1�y����M��A̢�e33�+�8模ۻ�d5�~G.d6j�UT�o���n�@���G �@?�O(noO+�k�_��f�a���,��v�r|�WC�]���S����s�%���&��츿�u� y�I6��!�W��=1�ͺ� �xvR��/v4����.��	�-�0,���y
y��[$ht��j?߁0�����]��Jhۚe6lj���� M���>֣�ʏ�Q�����&)��@p�Q��~�2�Ȏ��W��/u��ՠw"?t��ʄ��*n��p}/��m�bz;����!� �5m��1�n�R|���r|����I��'�i����`�iV��YTJ)\X�|�Ɨ!U+A,-�
?��ڜf;���E�U�2L6OD�rMI�Ay�a�j4�)1�������@<o��C��Qr>R���3,���!+iԦ���J��I�ʀ���-`<{A^�E�ag<�. w��7�uz�YQ�[��Ҭ������3�P寖Q�1"�P�	��Ã�6+�i��Dm�mcTz�ӻ�d�i`��E�����_����m��i{g<E4�����VT�.V.��%b�4���xY��4l9�~��k]�?���y���l���)4ڧ]3�s}���8�+�L֓"H�tT,ʼ�����7V��d�ҽ�8�A� ��<#>,7�"� �c�(	�^�z����R��"l`�+̼v��d�V�j��F������^pC�9���-�c�Bn-�2�e��:nz�t��$0�_��'��Qj�u$�Rma�E�!/��� BV�^~�g��	vSR*.�����[d=��Ð�����o���{@))o���5vCd�p_�!.���#$k
�4W,�s&���S�+y1�y,Z�"�د)���t��<T�aC�zL�md`�D�<�~f6��Lа��t��0����:#� "|b3萮�đwz�e�.��5�F�jP^�k`�c˫�]��y�r��G�a����X�l�~�1�C���P&�O�C��l@�,�xlCBhe�Ŏ�3�m���?�[d��	�0F �*�7`��<WEV;�J���H[ ��E��A�_�0MNy�.���fK7�z�vi�i��耄	jr�=��#�$.�YU��S��<� �����x��h�%����^aǝ�Vp��N��>lU��X��#�w��f�![�X�w�H��`ۦKb���X�8�	�y���cn��x@=�$����&�-�#��������K]n����X唭)�A��v#�mϯK@�-�=w 
̯���t�+���!�@\ج���z���0����SX��P�g7xM�P���i	# �5wBs�g��b �^Ƚ�2ļ���X�
��,{�i�.�$4����8�$��9���Q��%H	�����������k��_���v|��i3��:>u�kˋ|�C��j0�ȁK���v8r�
�΢cL�箖�9����[f��!K��P��S�p-U7d�%�?��e2{�Su�x	f`�'��f�Zo�U���J;v�	w7��J 	��3��ɓH���	sf����0?S��m�J���o|&���m0l�Jl!tb�I��e�+1)ս��#*����ee6�6�+��д�h~��dJqفq*����{4�G�%��a����|�F��� nX��pd�F��f4�:Z��ڔͩǑ_��.P��Z�\8�@�n�:i7Gae:c\�_����U��&�Hj�WQ2��!\�4觝Zi��B�	*px��
+��P3��.A�λ�
֢�B��r�� �6 �����c	
8��������!�7Қ��=[��./HX�.��/E7%4캞-��aZF�߼P{p�I��1�����!;�W%Y�X���AV�������Qy�
�Ї�x;-��m�r�n>�m#)g|^�L��&jm(�G���v ��nt&�9e0�vo�h�i��X����2خ�w����U�۞!5%xǩ��q+6Gc?S�gq�B9
���{����m��D#?}�m���ef���P@:�VWRw��fа>|"eNL��\���Wn�p�
�;E;��ŴoEJ�k �����������g�»�k��7.h?h.��,����
�5�=�>�?��)L��s��Rvr�Z��2��j���T��@ӻNk���O$�P��b>��r3�x5�\�y2IX��l ,%$�������jŐ�A�	�9�L�*��>r�j��4������"h0�w������ea�����kPrू݌e��u�/«��U�J��O��G%�m`��A�(i[O(�� e���Y6Z�t�}���dG:'�Ů�Z�D��j����4�_�УqhfEov��̘�UV��]���GjU!�i���a�����+[�Z3~q����:����i�E9:��Ս�B��o�t�$�µ�C5rl�ďEN>�b���d�_8zΡkN�WVS#���4��'UqUo5��}�
��Y��ė���"� �P�}�̲�O`]ϝ��1F�݀����S9��]�Ş{�O&�C�����'u�gݩe�?�Z��(x�'�Te(���.��s��Wa�D��t���I���F�F���x���4���a�#�|v�5�ˁjF��a=C��y�	N�aj���K��1��6�gr=ɟ����.��_ZT����&���G��diw-�%=�Ý��ҍ6Y:��\��n2/�9���_|�R{!�Q����
��.�@����(�i�e�3�N�Ah �<�m�@�}l~)���`f Ҳp��ϛ!�7i�I���)��}(P<�,~Ԏ���D �ȓ ۿs�+�lӉ�A	ĳ�S�ݼ�}��,�������9$����A�X#����3�_�<�BQ�3��jX�%��׻.�g_g�#A�Z-�ڠm��m���҉&���ə�i�~��AĎ�}�>�,�_xQୄH��u�B��a^-ᚪ#����S01ӂˀ���OJ�P׽�*�����)��.�o���׏����U�S��f�`�����e�IZ]t��js���h�.u�R�TP�`�1.�3��߰?_�%�W�2�$�T������{���e���ܷ� ��3��l��"z�ڞnc�*�%.���ru�3�E�f���Ldc	�)���g<�f�ꑞ��Td�`�0D v�;-��>Jޭw�<h%vI*	�Ƀ(gG���<����nB]<PO�P�R�9��RO��,H*�
��������M�Á.S���D�o�\ʋ{_:D>%���pN��*GY��{}/��4�P���SL���B��A����/2����O��B�^(h��B�/~�����Cɔ�q�Y*�� �m��C��Dv_���NLp��NQ%I�����*�e=�2���)2�]�i�w�e8ѫOA�e��fn���l-��JsVخ�h�.���,��}_jSi��L�<�ư�}&�]Y:^�#�Cճ�u����]�� �'���%��}��X��Kl'�������ej�٨��l�W�(�֡v����Xm�}��%���B�h�5�Ecޣ�fr��Y�ʣ�C����iP�Ոxt�����9@I�+>�נa��N7� ��'U��M�����0B�y�T��?���Mk�qm��b?r3a%C N`���D��fu���`��H�{(��p�O�]O�/Ͻ�w/�#���c�˖P��Z*�6l�@3�ᙙ����a�����e�&�7E}�!�x�Pɵps�d���iZ/m�8�����������k��2���Z�����|8��TH���?��=�4�By*����cc�G�3�ۻ���8��Z
ś���7�E�8��q�����D�(�\�����a�Ĩim�n�C�= ��1~OI���f�""R�� �Хj57��7�N.���Ď
*�0��,/�3O���PX9Aޝ.z!� �>�*���&�;�O��p�L��Gq0R%�Њ=�'�/$�+�ܭ���D��#*. VZ�b�[WH�b��d��v�E��W^��ß�S�r5�d���Y4�Hi���K7ܒ��:�`{0^<Y+oʳ���/�RX��pc��6T��W����v8Fp�ԁ�b_���r(���	S-˷;&g�y�����(�=��#⍡�
�b��$LH��3D6����m�6��V��R��N[�N�@�w_b���'!��e�z���� �
2���9ͦ�F"ڻ=\w_^�9"���gК�s�y~H�)ƅk�����t�]Y���.)VpR�.)u��!��b�3�f��>�\Oq��	d�r�3�@$ �������@��@;�d��2��"�}7(8��a79�(��G�Z��7��┢O��b'e�Ժn���A�O��9�	���-\��Ne�#d��
ܑ�Ϡ��Ku�K��ug��9ሎ���o�a��N���O�c� ���f�]��[8=n�T�u0��=;��J^�Q�6��|'�w�T��jK�RTa+�`9����0J�g�vN�m�t%D�q�L�����%_�0�Z_�Y�F'��n����#��5	��_l�� �t��Xg��/���?�W#�,ly0�y`�?
=\%f�Q�h"k���G�1�s&l���=�sw)���|0��<�f�,���@1J0�l�OE�����E��f�X��H��4�<�8�S�:Z@Ov��p��,pj\N���HN�D�ܞ�؏��'�<��mA(�-r�]	��r=c&VUv뚄�xê�,�c���łf���� ?�6�8��XO�+jQ�`�\Y�C�E�t�~6�x��HV�>3��ŏ䪈��*�����M�,P;��fd7�+��0i/�!����Y�r���ֻ��%<{#1�PG~�W<�.���I]������ֆ��
ä��|U��,�����Pm@`h�G��L��uX�7C��z��x���Qw:P��z�Gƛ2�!��Ƒ𚰳�tg���H�H.��0�.B ���R�j-��@8��n�nb��W�Y�$,2ю��r H2^�^=��@	�����zP���p��3�y~�,`��t9�	@���Й�\8"�2���bJ�?��5�}/���aB�n�|�D�]�'��,MW�UH���؍ܺ�]H��?A���N>�Ġ�B��NWI���|)������^�R_Ƽ������챻:��=jH�78��H[&��J%d�k��W�Vߔ��̋Ӧ����(�;!�l�K��ؐ��rJ:^)���R���B��4VFQ�D�}�x��vm#�1B��ȅb9ݰ|�5�I�Ȝt�(����cRt/�yr���+��^��/�,!��p�����c�>�V�NQ�����"S�����2n�z�g&G�%6��?��@ٛ�#Jb�!P��<���GX�+}Ӽ�93��� .�vD9� �ѵ^��ˑ�������G�c�
�O�J�6 E�w�Nq0� �> X����Ǎ�D:qh�8�/Tvn��9p�{��l����̚)W�S�Oy%*A_�ul�i�"�f���d��/�?v#���f�2S�|��*�(�D�k��"�	�♨��������*�Y�Z$��ο(	p��Og�H诠�1�%��N�x�V>r�ʪèڎ�U��v�RY9	}�֢G!!sw�E_Z(��~5ى��K���X9�l@��?���4۔h�ϳ����v�-��pX=mAۍ.�ّ���0�k���Dީ��u��oR&��9����f��"�O�N���T+�dͦ������)t,c.�~c�5r~z��^FN�M��C���MG=�_�Kft>a0΂�.2�����0�΍?�@��e�.���V�`{����V��|�5��5��}z�y2y�i �]b��U�Ɣ�H,1 ֢8�.V3˘�[]�6��T��^�쿓�SU]PVmFf *d�	��p�o��5
�	���"�KY1?m+�n��ռ��^h ݮKD�t�|��Ɔ
�}O�IV�GI��T�-��"6�s<Ep<F��8ۋ�����N�[`�/�X�L�É��  J��[R0�b�ZSu[���2AxB�m���m�M^��6����2U�KWg���D#�;��a7��cP_�M��Xы�߽N���{�!v��%R���}�
#"���95�x.*M�F8�����u�e��'�"�n-�ل���s�C�'������I���'��h�ͦ���?ݷ�3�q�[��c\�����t&&�����j��aj�CM����R�؁�:�P�
��|�\/��P��"��<K�\�k����-]k%�D	��X�rv��^᫜�JK^'�si��y�� +w?5y�?�r���H�'��`�%��l?ŧo\�am�a7wk� �X�גz��H"Ũ�;Xe��������X%d�b_��Q��3}�Eܢ�6L�q{�`W��}�~�S�>1/wM�n��ܳ+t��yv�Z37=+kb��cDi�S\��r��U&�RkeR�V�	�	�.�E�?��+���Ǔc�H�!�����pBM�ブ���0�~���5ev�F�f�~�&��
�Q����{�nW���y�9�%���-�j	�=M�љ4MCX;(Z u
�v�f����k�P�ؙ��Ŋ!��f����϶�Np×�2��k�0(Y��p\oUB��D�g��H]��g����궥�A�͝6��&\7��ړ-5�ΰ�1��Ӣd�д�N����)4�͇��ӈɴl����zLL�n>	��|��/M��a�-Sz�V?��ӰboGGv����ʳ��3@����ΐ����*F���n�U�Ǿ�Pw�Q��(�_����TPsQ�_Ъ}��� ek�����/�NM�0J��?�8q�G�za�R=���;?��w)�(�%9�.��)��("�˳��S�0\��.�s���h���W���?*�����.߰Ǜb$�3�&�R|E��S��DU���?/����J��C@�!��e�u���\~�b��w"lPq^��,�D��NK멝��y�-�zdc!m�f�9	/�����T¦��K��?<Xt~,�;ns,�z$1��H���'`U��0�n� ��;=�O��"��ʪ�����=T�<�\	�a�_�z��z�ՆIdu"*f�>����v�m�-K��N�Op�g��Ē�aV�\�B���&�`)O/���yB��o��ل����AA���ݚ�|�
ys��k1�o%-SN6��H��5�+��Ժ�I-s�M�v��z�@����zE�s8�8|p�F���I���1Jb�x���5�j~l���U���j(�X)	t�#�T\ނ��O	*��3�
^"#0�%�A����ݨ�Rɋ��ۥ����$w��;G�+�v6f�؄5�A�P���>�a��Æ �j�Gl�i	�:�1������͹�F���91���Yg�2]lXM��O�	�
^����)�t�}&
&e�%����K�F���` �
�$9ٴ�����������F��║�D�r�ڶ����g<�Ee��{Anz�C$5Ȟ9J���wP�:�<.{����@Bӓ��Rjޑf����F	h��\�n�am����������L�� ?)��:�g�!�J�Z@�J��_k �2�<1]@�扅����u@����;CQl�Oc,��rÁT´7cP�kʄ������h��Dd�nE5�����+J`��f\ϊ�k\�xdvA��\�k�c���a��*-oe0�dw��k`g��o�aӌr9�mP�q׷k��w[��x#k�i���0�����~�Fq�	�v��f�i��pԛI�(�/�P���J��X�o�8"��t&m�{�����1�b�M��Đ�eL*�+IHČ��4���e�;��R��G���.�7�׌c���t��\�֗�=�v0�j��Yð��B�#�彼�ԯ6�G.���'��P��w'�6	Eg-9��m�a�hE��U7���11x��r��A�G���m�F��*/5ͦa���Be�Z&`\1�5w3�w�����Z�n�����%��"yj��s�xrL�q��e%͠�YCSOt�2�QY����?<01��q]�⩽UrM���bO\Pm'S�6IjYr/�BY���'������d쪑�
; 	o�i�C���JOַ��s^��@ ޠb��RRC��խ�	(�B�x$�� �t���|�p��
X˫B��͕l8�^a��r�=ܱ@r���M2"5����Ȼ�f\}I��F��͝��4�a-�A  L��1Z�V��(�����6� �3�Ð�#�|�A�e�$���[SM���O�F����|<������	�}�r�Y�Z��Y�i�.�>)�4Ԏ:Ct�
 �#�6��l�.X�D��C#͇���J�}�P�AC�.���NN
��{|��?8�����j f�$���5m[R�
��5���ѿ6�?t�4$1��|A  �>����N6ϛ�����w�d�n{vf~	��ͩ�bS}�����_���bg��l�MiS? ����K��bB&պ4�
R�����H��XBe�"�fW%nf��)JA8��H���Yxz�9k����3��"#-D�=���68�#�������Ǉab8.�T�����M�4Ӛ?��r�8�R}G@���A_��3^�Qi0$��<mi�^e�S�����O�no�/E|C��T���"4��Q��IG��ǵh'�[�H�dz竑6�'&�t��a��x�����A���S�_��Dk�?'5 0{��]C�#�H�#�f@�߬uM6FKĳw<�vxʠ	�6��-�2=K�n��m
��
ȁ�`�ݲ��/�I�^��a}9�F�r�� ��le��oM׼�Դ��_ψIsщ�i0�{+�� ��-�R���&����qM�Id5�F?�^|(��T�[~C��U�
��E����h���$�'(��H�� "q6�S4���+�RZ���G����b���Eqs.pAK�F���U}2�k�i��E׬���Ih�o@�ƨ)I�>(!�� %�b9q��;-΃��똉"t��	a�{q�!zc�/�lN�V��
�uCDqZ=�)�k��5��E�3/6�}�L۠=7�#o����0��b4%�U��S+���Uˌ���g��4�v-I��]���	�"f�k��HMBۏ��|P���s"
E)9���S�	��o�h���Ln��jb���@��%eە�0Y�;�&���'��2��;`�����%��NkDOZ���l�>[���.�w�y53� �;{�ǒ0�w��,afɪ4?��
I�>M4~=�^��(�9S֒����fzZ�S��Q�w>w���a�=�\���K_s��Liw��L��U��/�
��K������W�!����l15]
�iC��j`�,�?;� ��2Ƅ�+������G 5�1����������5�34$7[�����=�`��Y����@*F�Ѕ/�i1�Uy� 㨧	�V9�`u
�58�6�`��6'E��m�.;�o:t��PB�~2�2a+�Uk��!���SDn�As/���uj��S���B���X��zK��&b����P�>����Զ]����8���ԧ�Qk�?=tLe��*�o0�Vh�<�mn��Sc�cJ���Bf�>��f�Fck?�DǄB� ��P�7��-)f룷#���<�D(��u*��6��:�ؙW��m��N���P�|ȷPKS�Ӎ�V,�]��L a��1�H6�w~a��8��]�h�iX+x���ʄ�R��C�K�t	����g�[�����:J9����O��R�%i�,�1 K��DrF�����K-��\o���i���k���?
��`��wԪ6d?��S��P-T#;zQ$��{l�tGǩ1!YB��Nų&>����T�xU//K����ۢ;�E�Sk��B����-moO�j����XX�k7J��x��Ƅ�{���I�/�$�<BX��i�R `U�����E{ƈ/�f��F̗��n��֤��@dV<�t�p�3���t@����������`���T׍�B��/���%�m�+ջ�$�۵0��Y? �Yvʤa�CG)򌺴_Mi��_�͢+E�ߢ�IE�$�,�dω�x��Ui;�d�M��қ��\a�a�`���Ϧ\���u^ˍֺ�t%Aѡ\u:Q��y�-���l�^�sI���%�w ��,��̦�7��Q�I߅�j_J��Uް0��28@���))%J>�Iv��bȎS;Q��袕�	����Z�Ŀ�|Oy#=,�o����w����ا8�2wv[׃���&��f��3RE���89$Q;�~��G��/v�o����Ml�緉r��؟Ǘ�kQ�;�G�s��O:��e��}����V����J3��-/A`� ���[�-�E{����S:dG��%y��sJK�Մ����w=ԃŅ�@>&��I݊-X;9ֹ����m������������AػQdÐ�f��V�E�8���Ic��i��s�%�u$ HaF�%�m�r��Y�J]�,�E+Ӈ��|��K#���|:3[��ԧ��FM��aD>���%�Q��(՚�.z��v�<�ث"P9��hc�8/�*Ǐ�,��m�i�kq����H�$��x�NF� C��j��s4�I�zA������PTCx
�2�:O��F)U `8�;}�:�%69��x�_���M��[9������?�q��$��Rۘ?08���P"{�H�!oa�|���PX �p����$_=mE7�r.�!rjx����Q]�,�V��I�bo�8f�����=D�\cP#m�Yy�w6
���ɡ�Eί�A"�쁉�Mv89r�4cću�������8+'Uh]�O��+^�G9�?�D��'&PO@�|u��p@q���߃Ek=p� w���o�P���f*�����8Xo"ބ � �.G9�Rς��c�*�e����`��!<(:�>�jO�?�2���A�>l	kWO	DŜI8Q���*��Kvq�[�����\���~C@�����s�m�A�d`��3�d�`�)V���`�]��v9L1�iu�����{c��T�,�Y��z�w���	qǑ]��S4�J䊄�w�#������p3���B��
��8���X�A١������|���ӹ�t-�1�m��P���K�����F�Q
�j����H��λI6 W%i�
�f�%oʿ.�Y�%��[���'���%w7-e��{�?EUŸ�'93���k�u}�L�Q�f�"E;J�i@�:^ʋb/�4�%��5���Sy�v�J����)�'�&rYw�C�c�I�T�������X��Ȼ~��q����hIY���$ W���� ��F���P]!�{`2k
�dSf
YoB�R侷��-���fl���ύ��jT��X�2��a���5�F�3#n��Xx�mɐ�2�jY�h����!�iM�����Jcݤ���Hy��u�KL�Ј���>�<�@@���g[Vx��+?<�r3��?̼�cp��Mu�+��PBge7	�X�����2n��d�T��F?�B���.��[�%�o
j��OJ�f3�i��9��97��q$3�W�a��M8���0�F�&��<���F?(B�v��k:�"�.}!��-/�2ep4\��.(e�oBF�}6@�d����钵\{5��6�fw��vd<8���s�.�?j�$�������U�GB��g`)S�Y6�7$)H%�@�n���U�E�X���SV;T��J~خ����IL&����)�!�y�&{�Q=���̽>d�^�wpc�*]�&�'�����x�E���橎��D��n��'�z6�<+���#�T�+=Ŝ���N׉ƨK����Ws]�xQ�Z���9�i�w��
�����c'�����x��+��0WJ�i\u�q �%)	�X!�l {6{�Vm�HՋq���/�X������݁�8Z��yp�
?���h��1��X���)
K�|�bi�x�!������NI{��0�u�cw)�_�C=~�d��@O�nڄ��)�c�"!^�'��m#8 �����^�/S3m�����Rm	e��ݎ���� ��+"lY�Y�v$�yX�u���0=��n� ���nZ�E�ϘJ\S�/�{&���5�m�137E^¿�ֺ�$��ܑ�J���cr��N�S�݅�sř����_������lK��Y2�q����4��֤NS���J&�c[�L����)cVU�Z�!� ����(U��E�Zǣ�I��V��#
}ޡ8/筎J�7���+�^rwL���ZD�>�ޫ4��	�a7*�'쌿����2�x���*a1�L�"���H�sc�*e6����D]�>���oP��C3��b9פ�&�D�]�	��ħ �#�Z��C�v.rU��W��!xI����p�t���7.q)z��8B���XުQz"Z�Ӱ�貼4к�)��*T��}�	T�|�P>���D����!K��fؒ|.��㰀n5fp:�d�թ ��)��|qX?�;v@!k�\$���7�X���1�iTY�mɌ�,HY��6U�ۡ��0�Ef�a�\�	���قL�m���F2��sO����q�+)\��p�r^Ǻ�[KV_L{2���E4D�.���"%QZI&�
:]�uM��&���E��w�8e#j�<�gF:���	~mMp��� x�� /��OL6-\1��;YTu!+W�GVN�O4:4ܡb|�M#ϔ�ל]fm����Ծ
O���]}L��4�/�e%W�X�,=<�{,e��l�W[�l���g�lp=�ƬG���������ˆ�+���(�a��45={���.y��FF&�����/b��2��*����8��W{zZ�a�v	Y	ϧb�O��� א��b�yC�1�!<Up:z�:Lo8fl;u/0��\��}�;��*�<y8Hۡbo!ׅbH�X�H"��u��_=�-Y81 ���Q�N��V��A�,�b%�#5�ֳ��MeC�km��3���t�U���se§)S�gj�q�I�1}@��\:7���k����N�I���M�`Ҋ �{��~«T�-$�SѪN=�xMS�gw~��*��&��hnZ���s�Y���je'p���������Z�r`��Dߢ���%#�=����U�iW���+�.?��bK�!�߻㸂15��y�,�`��@r�>�L�XGe@I-�"+�/?e��o*j�V���1�Ht��#�2C`���7w�y��l��H���צ�-?Kf<���8�,�5ȟ�hIP��#����J:�2���у��M����D��$�����*@_܃�a,Z���I[Қ���n��B4�b�r|zq� ��!DjR���4aB0����L�2?9�Ma����S~�,�ݧX�a�i�����Ui0��@2W񃮿��-���|L_�+G����&�؀`�}�c����:�=o3�bn"ca�oP�H[���in�7�	���|.^�(��۷7&���m�(zPi/E�P���OEa�߻3T�;��qXfZ�ݨ7t��8%%���RJ+�4�n��P�:u�P�ˁ\����Ot����7P� I�S����.���A��:~��1�A�+���
���`�z13�����٤i�����cv���=���*�t�C9W�լ�|	�e�^5B�>b��xi�.`�*e긯-}X*<��z�4� ��k��ER�������*TK�B}=�~J�����b�P��Y#��$+�p���Ȧ>�]��ο�L���ӨB�-�3r -���ñH���Iq/-�#^)9��G􍮔����� �c�؉p�B��|B���k�x����T��፰d�R�jhK.�5�N�U�j"W<ͅ^�c�+���\��G\��1<��羅�]��|O�2C��)x�Y��WsZ����U<�aw�ޱqJ��+Q��@%��?f�@��V.�>���Iq�w/��X� Ic0K\s}���xu; �Y�7�(�'h,��2Hb���݆�%!60�n(�q�^�ȱB�O~��\HW�p�t����yZ���m� ��T:�
.�Z������� S� �h�q�9�>�|�*pf�r��>�؏��JܺF�kA��_�Hk֥��	ig2n�{ے�a����`SHD��+*��CRbL�ң��W��.^|f�,�NGNOVo0W#��=���>jŬ'g`�P�o8�G�/�6j?*@�s�գ�%ј6nX�q��*.�с��3Z5U��Y�r�< 3���D�Z�����)�=����"� ��r�b�t�fs���U���c�p��v���Z���p�� ��Y{4�L�\"�(J����:l�s;�EK$`�����^б�2��r���E�A���7�4'��g����Z�f&u
��^2zb��MFLS�c�!,f�c������2^}�"���6�?a��2'�����Ȉm�!rJ��y���Msr�!ݾ3�mU�1��a8���>�z���؈���瑛)�\4ť�'!_	F��)�<?�?j�O�sP��;=���Dm>pѤ�<*������	�}����s[r�z]K~rV�K��Մ�
�Ր��CLa����c���ypV��UE)��Ԋj�+��.{	P��;��C|���q�2��W�D1��W>m��O�E���b���U��o�9>� �!^��aV-��^
��r���zNq�!Ke�$*y�@��m����
s�>D��o�ʠ��7���x��sKՠ�ͨ�7S?����ŧ�_�B!�M��oE
���n
��	�1J7UX�2S�B�:�T�
��u)�D�zW�r�����ɧ��!\�L�x#!T�ל ��:��>&�rq�&���۰�2�j��`�7IQ�R��7�U�i�yJ��fwP�U��b��|��_��fA�q��7xi�|ĈBr송�t��O͏Eh�B�i�SRWn';m�?KJ�V����7J���0m���%�Xv�����
�}��;�O�9Ɗ�w��4opG��i��������J��V�:��PW�o�[��
�'�I'<����H�����Ō����f�GT��3�L������4��|��f�d��ʼ�a��%IM��ߧ;	Kl���I��з��}�FL��, ���A���յ���Jo�gsuj���Bsݢy��w$=$B4��!0PIa+!�ɜ�y��b�h
�������A4p3���9�{����mE)1�3٪����i����{��;@?>L�����9���P�_vl�{�����L��֥D,I��4Qi�x�(ṴZ���X�6���A�U?Y�\�ZPu�6�7�|==>'`
��W,��x�F!�����&���s{go!$$wA`���z�\�7��SQ��xDd��yp���йk�Y0p�j&$W)�{\K�)+�6��%nvM.6;��b�>�����.���p���D�ش�w���#�������&��E)W>З!`�t�"ro��߰���z7��JZ�.���H{��*�',UM:=����b�rے���x1T��,�WUd���d;�n+@{Ta��C�M�_���?d��Ǎ�b��xR�٘�x����w�C5��������x��gt�6���|�a��v:ٛ���T�i�	nH�>�#���2]h�3�z���~��5�JWk;���E�T'������B����nf��=�$���Cu"�����SCV���I!$[��J��u��Ga�
�i����A�h�l�^<w�GWr���*�$	'��'g��*Zp:�����|0���k��X��b���^�"~Js�6$��=T��̬z��>��@����
�M�+Xb�0f6���0��fG&���4#��蕇^bj�P~8 �`� ��`�*��U�����?o�6�r�!��5�j�g�J����zQ�M���;�vwK�l��x#?ٕ͡��I��]�:�nv�t��T�h7�D`0*Y�\�@J�oz3Q�Qp#��`�B��»���ɹI�ۿn�����<u�ž��� ^�=��d��~I�� ����E��(���S��7�k�Sa'�{�Tx��@��	RI�N�%b�=1_�X�#���x��]W'ݲ�~p�2X�x�$�@��@aʨ�f;�,^��E�����iV��˛(�k|�I,iW�*�*s\dX�`�I���Ns���m���5�#�o	($p�,�Gf�iu���t�V�`�9�t��㞂$�=}��N3�Dh*ٍ5��j�W��=�o�-�-�g;��4��s��=��K�1i�I�XA�~j��ƺ�3-���cT51�R�u�w��>P�y�y�O��r6�W��r�FD�>KL	�����m��<@ٹ�6�e�b�6��Ug��W����	��CD��1��@�C(��,A�����^�����?O���%�jm�rm�1��3կ���bǠ��
D�^������V��	�~���,>`�͔�'0M��M�J�=�۠_��Pա�{�J
�9r��N�"�Ǟ˵�~x`yB�,À_�m���x�F�_�A��#jc��ZK�g''�O}9 �}���M,.�~ބ>�'�����pPə�S,>KvA�T5�a��A*�`³���x�m�����/j��]�L�Y�i�8�&�W�Z��R��FM�$t볎/��	O
{`3�DVN�(7&�����+ѯ�8��$/��Qy�^�Dh\�9�C�*1��mе�C*C�[c�1�X�5�k��M�/.p`7�`a
wg�=_3�ٜ #Kg���I�*�����\�v�A�l��vi&�_k����Oe�(	j����M)d�o"�N��~ۯz�9�N�!�U�ͱŸ:,a�Sg; ꖑe��=J��k�ׯ�7���X5]!���}5C��y��l�������k�Ҡ*�
�����`{�H^ﰸ\����+��^m�/� ���L�L��'S[�=�/$�&W=���5��{ZD�bSM,����(�֒���p���ʯ���`�_9��h�s�g5e�]W^	�>_>ΥN r�^\w��d�x(1d/��S�
���"�����E��!*��pE7K(�?|�6�5
�nHLmx�|���C�[N�mVLn��>��@��jK�
8�L�xu���9�[ť�����/�T�|��2D��s"Pشr�	Da�X����q�)�����h��3�f�!�)	@I�X՗�����@�f��!BH��= �#���2v�OՑ���T�෼�GF=�،F��?�uA��+2WI�o�f�̛�u�ӧt���K �g���!S�:GQ��[MY���D��,��F'F_~��k|��4"n��5ѠEYF�Eo�roFnKy ������PLBȎ�{����A+R|I��xâ(�)ۆ� q�C�:�g׈ic*���N���\�<{&�n�l%$C=�9����8��Y���nʭaΑ��ꑫ����G����|�z,��!eAT���"�Vns�"�����3�U
;���~)�qb�����I<E�N�dK�1%�~"O����B�ڼ4�{i��[�;��	�So���Q���ř��]l]lJw�����E���{�+$��TĄr�l�D�}�[�:ة�Z�o���������x��A���ZI�E��%�$ִ�5�-������t�񔭈h��tE��;h/����bb�e�<+���w��6�e�i�Q��	�hT��%Ih_��⸝�^�{��"�@��px��h�����}��R?~��6��� $�Jj�E1M�$���<z��%�ߣ-�OLj�h��eC�e���Q���>��$5�W�D�v����?D2|�pN2�R�ע��?`�N��7��4xI�ɄK���7����tk�&|n�����A���p=�T�0ib�� 2��)f�:w�O��V�K�� �����Iv��<��o�� ���9hc��~�����f��DZ�5���0h���<�O�rY]7[��[u�w��������2�w*w�*_mg}ԟ3���V_P�Ӭ���R�d�$Ma�r��lΘ��Nu,@�Y\R��b);��qW�~\�����"�ѓ���p/�b`���:.)�ѧ/�F�]%�f�u���܊D�t�q�e/�,���Ė���%\��&�%�[ܶ��F"��Zy��/~����P��Rα�^�+���O�K��qC�5���?k��y�+
���^�fNVc�ٮk ON�yX�$�����n��h�PD�����.�~9[�.'�m/��p�0v��\?`�aqA�A�ܓ  �E ����%q_4���Q/$���)�I�:Ǩ��������~+^�v�m����q�L-���'EX8�dQN��A�M�/�Z��o����f+ۧ�b�d�<a�Y	^e�)��C�k��5% ���#�bX S��F�Sx2Q�w����>l��X`��ҖaK�K��N|����~��3�4��'H��˙�ù�Q":;�}�D�w�����}��}p������z��EFŁ� b 0}�h% {��d��2��YRR���s�x�BZ�2�]�߿��[I�.zN����Tn�<l��Z�u�Fh/p���C��%�X�e��K?Xʠ]\�?��ث��#"�;O�.�(Xg��#����:��&��7��v�غ�Wc�;<u�i!���\� 澆t���"�5����=k�n���$���{)���1E�?���	��ԟ�l0�@Z;8� ��t}2��$�rp9䜟��O2��+h�p�Oӕ#��?����#�qd/zI`%1|~�F4�����'�\d��kP~xy��Hv�������Q�G�o��Ҥ�2R9�)]UH��é�+�P�d�P�	u��[�6��|�KJ7�kj���!��ԏ��h�Z��'�|�"g��+���eU9�}�,N[2_�7B�:Tf�d�}��oA�0v
��/�Ȅ�mH
��9-��/Ӵ�z�����8F���6����*5r��5a��(�.�eW�d1?Ld�aj{�!K	�b/w$�vXP�`b�=�&	�4s��[�qr�+6�X�%`�����MG_�8��Z�2�)ʓ��Q�`�Ȅ¬c�)���?�n*�,������﻾�0TNk����C�p�+�8@��v	����b�ib'P	�T
ǻ��Ѩp�䮵��8x�7,1����x_oX,�!ak�֟cl���O�/V�!g9����˦{DI`���<Gt?>���O<c~�*^�L�ԴX(�)�!�1�P���B��0�d��(;f�F�<�v�����_��,R������Kr��7h�F�����x���Sv�����<��@��� �݉	G�����& �G��9��A�ʦ*�;a�!��I��E&�����v\���o��t0z��Yi���-'�ʲ�`{1��&�TIQt�^M	؞����VS�]nUe��(ܮ�8U��xfIU;�h�t��q�Oxň��A�1���ok�E�΄&!��T�8�8���:K�B/e�e���_0g�٘��A�z:D�;E�����Ç��KsP4���>�����Yك:�C(�5��7��0�VҌ���nI*;b͡�,�8(To��kz���ʓS��>]�����BTS�(}W� &@NR3�_\FK�=R< ��* �ܮ|:I�Vbs�X�z�Ș���u��.��Q(�N ��!�TU�6��Zˆ�=%����E��(��J$���<'��;�@��	����`qp��.�]�G������lρ���k�� !�����4䎚ѐ�E��x����Dr��k�`78��s�;��hQ���2���(�7K����@��\i�T��n����R��H�嵹�*��(mhT�ЉN����qL��2i����C�h!)�`�ە2;A��M$�HUE�h������)�
"��Pe���y
�>xL/�|��������:�������D�\r+��do^J��ҏ��K��J�e[�]w�"d�}�a��a{*�d�?�H��^�Y(���xd���ׯ�%���ڛ��&��V5�-xbo�Q�Y�/�����L��"<�+��59������e���/�p�A��U��ђ�,���fݥ8�룙~���A�k�x����ݐt��KJ�=�;#�y=º�sJ���;�S�%3E���C�A��IW�/ݨ�[�ZJ��(��b�ԗ��7 
���VW�u]�����tu �m�4���-�S!!V�M����vCS	�e8}E}�1Q���n�ꔾ^����;�wK*�Y�؎s���2�tQ�ql���CR��澰8e����N�ޫ�,z�U=���ڡF����`t֕����.aw|��N�ۂm�2lӧ5x�n����ߣ�޹ހD����˹�N_pD�%�?f�4�ۥ���ޅ"�,�+��9eO����s���h�β�
��A�(�z��O�t�%�����_Ae��+u�:4���򿦃�c��<�J?11��t�!{�X��'�m�	��D�S�����;
��
/��9?h��~���|(aL���ץ q��n��u������<
�k�=� �K��^;�d�dt��s�z�dϑ�nީ���T�0�6��k��;e�6���³�WU��U�Q�B����=19�w�=�0ȝ�'/�bĨ^�Q�E�-���/b u�y��9�}�x�^�*��I9(*�=7^��j���Q�?�zyX����;״(N��tul�,���[_�$c��8ak�����7�1.�43����S$0	�.�jWs�5<ٔY��&E�E5/#f'A�ŋ:�%M_�K�n���Kx�oڅI0��R�{� �ʥ�CX���y˛F���f���������򓝾���X;�z����{����1�g���%�eXzÿ���sp��ǖ���w%��C���HF~��`��dVeA*|A;kr2[���Ɵ�8���A��Q���͠�ʿ3@��A����ⷛ~2��k��-�T���}��a�Vd�`{��p�)���ZښC{��s�����Il"r��n�$\�'>��Iu�\�jB��0��ޣPe��Mi����YuY��+ ���P�"�n5T�i�r)Cb2 ��5V�@�E��6��א�g��S��:5e I��\'�=��[�y���8>�&�:,Z���Ī����K�v���N�������4urbF��F�٭ۮs��%	��/����*�!doM���֎�}=X_�n#�۸ڐ̯���㉐��v��`��-�NΌ�g\�Ѱx��K��5[V�$)�*�� o�G���r,�ݫPz��rs�7X��F�ń�n;s�[����J����ve^��R�|���=�_���֧4�:0:ɋ���c�&j6������V6^���?�L�h�9K>��os������@�s@�3cͲ��p'p�a3��{jZʹ
} �1����I��[gWz\V����w���6�8��p�B��G��P�9D��a�|h�Pjg�+�o�J �z}ا�"鈉
�6����)Ю�/�;Z��y��߸Ɍ�h�����zųnA�`�U�]��m�=r9=F�J:4p=�N-l��O�hO}�FN�JL���S֮lӴI�mq�h�H��xP�*�' ���0sv�<�Q\��t�i0^���}VqT�ץ�������l�D�^��;X�xO���J ����Y4��Y���m)�F�^�npjw͔�0ܩH	L�5��?'���K��	e�9s��om�J�)�1�/�}�hq�Y�N��8_)%�Ҙ��NzA�qd�h�\#�I�d�ے%�kH��,�G	�_�y�}$d������ �f���\#1���\�B�J��!�_��-2�$�G�I�ڤܨӁ#�K0S�G\s0o]��$�N����.�	����P>��:�Qf}��_�JI�w!G������b�<�5�f�,L�D��Kj���"���7c+dN�����@B�~|��_v3Εn��ܐ>=⥱������?zE4� ?�ԥ^��|i[A���q$��/f�`�oߵ����e�C�<3�i��:��³�ӂ�=���tv�v�)ʘa!���%G&���-�����.e�l������$E�	��~���v̖�v�s�� fa6����t���3����|�1P����#���ݝ8.r�}�����B��yF�Ӵj>-e�1�x��\B�����EFբ_�6�ch�F����O�S�@v��^
Z�Y� �Z�Acڽ~M:��K����ӿ�57@��1_���]`��6b�PǶ���V�����`-v�$2�p诛%m����i]!>Q���͞�b1�\����#��?��������	:ɔ�?`o��x�Z5,}˨T��N�ʢpp�2������<
ɵ��NP\��h	O�뇵����I�o�bҪn�Ĉ��A����~I�\�;)����.谄�ǥ�\�VV�1'Ljū���Vb(rae�q�7�r�����EQ˹�q�w%/U t�j �R���N|I�+˿����=FIn.IUվ�르I1��D�o
�c�|��a�ud�X~�Y}�y�K9�Wn?dr��ƉN҆��p�|�B��U��e���^��ch��i����+�\a贈-��g����C�^�ekl��p�ć��fyڳ1y�.�=�tBD21��wr����<�#���@Ou����t���V�I!X�"����i������4|�;I����]~@�*�gg��~"a1o E(MB�2]��&8i��$q�5���L-�$K<r|�쾚���k��&��1��>�C~��%uC�\�\�l7i�@-$�ͪ.t�$��	��	�V=Ṽ�ns��b������5Jп|,�@���@� �^�|t%��F�z��{(3�Wc�,��x�/ �c{ �����l\^�Pl���R�7
���+}�l|�Qa"�i�0�.�:@��֍O�t��r�Тy���@��W�$&�'7e%nt��flb	NÁ��Q7k@b�^P<91�H'���3)Ltt��h�Q�[[
�-�C��)@�Ol��������oP89-7��d�I�"�Z�� 2b�va��{#�(2���H=�g^��u0�?{�����[�Zz�e��䲗	�}�d�:|��&�>~��=���H�;1F�����L{����+2�R��_C_r'���g��*�[\Ԃ�UD[h|θ��2^Y�x�0��+�C&f�Tǳ���eu< ���ѩ��=�/�;ݗ����x5���]j3�8�O�$�K�u ��8��7�9�|G�q˚p�:�vOZ3��I�<%� ��@�f����V�}��h&�=�?y��1������΃��S-8,��5}K��.�h1!@��W�!DƊƘX��UWD�v�س���^�����1Ȍ��E�� � �5���ץpD�9@�Vq0�IR˩��9 ��t �5����$�O����M�=�Ot��tW���a����K؄��ɳ��V�e����g� �OB�#:����@��b'G&]'C�k4�V���+��
&;Zc���v;`��*��0�D���< �I��R�����+��%��8�b���m���XT4h9�A;��>2e�n<���]�y:��T�y���:A����ɼ�:���\=-�}>� ��0WG�#=T��U,��Xp�f-E��	Ƹ���[�z+�����!��>(���_Qf�n���ܦ�H��BЩ�^4Onb�Rh��I�tЯ����VĪ!kP���������D��H���X��Mk�#"��hW��J(=՞�!�^�y�E�����)_r��,_eʳ6�M�0|cZ���ь�hZCo�>B��a\��q�
;���f��ZW����~�0�P؎�+?�d��'%�m�z����,3ͽ!��s��*���X$ɨ?��߸���C?�b��	j�#�\;�J+E<��5���5X�3�</7 VmL�Q�CM���4��J��A`]��㣻$�'�ȹ<I(���� �2 ��I)��|�d�a[W���6��5^
ޤ��We�5��T���o2�c��j%��4"�鼻�5�������b�L���B���x'�V%�q�N_��������x^=�5�P4د��[ys~�޲D��_�����؋�+ݸ棳�m������65�^S�r�*T���V#ޖ���d���@ْ?Z�f?���|�46!/��&��8@4���ly��`�T�"R��q��CM_�8`�0ŕ��{4;+0B�f8ډ^�I��l�jh�+�E�<��EjM	�&�K��o���֜w�\A|<�	�6a�!�/V��Fa�O}�aYtR�j�m�ڦ���ts�����4�9��R�zj%��z��`�k���:m�'⨰�<�`��ZP�bW�v��q�7��-U�(���%���g�����|]�-K`h�O�}Yw��Vw�X�,�
y��-��/G�6��>����������L��_�C�%�����w/0�DX�1[��]�!er|�Z�4Aܮ9����g�n9b�:8�DY �D�e��
��	��WqAy@G�g��ڮ��'�}�W��80v�Pk�(GR_�A}��F�PA2=0DM!�$+��q�ct�T2N�nn޹��6^\"y�~���ͱ�-q��઱�$�ʅ����������*���t2�߄ۃ#=i����x��/ߌ�Y�J�gf;{��'1�ӵa4fĐ'�ѭ�/cJ/3���}���s-oI?JI���](n�5cr��U �H�&��0?��
kh�J1K�;e��Y�B��W��w�Kp wF ߡzϜ�]�ks]ãJG$��F�6�i}ր���3�۲�[��d�t������5��p�rfc �I��i7���3�aE`M���%�o2�N�bG�'�:B�g�H�X8Bu{9�ٛO��m�Ն�pp|f�UK��&����5�*�tU�*�E0�
�a �G���
è�=k�\}��9�[\�9��<⯆'�������,�1������_��xN��wߌO�Lm�~n`�p0+��I�V�hK�,(����TIO���ح�H�41�o��+��O�Nk7�k|Xi�qri>��Ϗrk��9��(πIS�8N�3�%H��*/O�A�[MhS��&,㐲C�U7����Ee!)��	��j�����$2�9A�����m����q�)lok>u;T�bp��o��b�C�Lv��M��2�C�'��������>��\g��ld�.�H�t�P��\d/�jx�]y_c���W$�&��֝J���~��;�`Zo���$������4B�٨�
$��6V��3õ�K?�7�<ը��9�z�/"E�&h��w�	@����&�+�&G��|�� �'h�����-�[z^H���lW�Fkn���_���"�#g����2��w��[�f��g+�
y7�����<�1�٢>>��I���9� op{˦��>4ձ�C$?�V6�ɝBŇu��Y���Q�C~�֩���C�<��;�
L_�B�F2�1�Q�a���d+괰l�1.���RQ'�i�p^%z�m�)�����ה�?��+��!RT }*P�ֶ_(�����'A즸�Eˤ^��s
�>�T��;�������S��"�\�����j7�Y�۬'��8�}�ח�Y���i�5����_~*H6�\ka�^ۃGS��.�H?km���hݗ�i8��5ۊ:�,�?O2�gJA�q*�L5d�� �J���c)Y[�J���}�՞d��`��-;�-�6z�:��Y�L�dzV�؏d_PR��A�_��'v�X�
w�*>��M����k���y/��iמ������Vs�۟%*��w�9�����������tJ���8~�Df��U4�ޯ���+��
%��oY�t��滵�t��c��4�r'�l���;���^I��}P�&b�����э�1.�� ����~�y;հ��/F1���P�)~�gv]@�GX��R]�j`�l��~!���k��^�I�=��D�Nt��60��0܇�=��ֱ'��G���D[����MM��}?�s`���j��o}�[1S5m���4Y�B�./N�[j��&���A��y�+����r�(!��(��4}V?z�k�6�a�� 5x-�Ea!�5���).{|o�(�G�Bͱ�����+�s����gYTr���XW�����N�%�GF���}��йV2�x�;UĘ��a�e4%��3x*�L�
?J�K���Be���_E���nd�igC�����8Q�:q�~������`��6#���,䵻Á��Q8h�0��	��� ۟~GY����-`�$ �zFGg(�>�04�(Br�[�
U��A[ij7w��nx
��,\D�����F�T6:*MZ<|/���:�(�Q�����f�[%v⼞��a�6pMV)�(N+��E>?��f/V'�	{(b4g,OV[�%Jc���/mɹN��j\��4ˀ>�\�J�dM�pw��닅ϩpw�q�P��!���c����`Co�h�A��Yс�fO�?o�4=G2���_m�ݛJ���%�Ɓf9)҉Ŵ��\`9�@�2r*@n�xdOQޑ����J1�3 ˝�'��kx-��;'3qM����3�xM�(�v�����aRB?ҕ᜿=R�u'�KN��r	T��y1�`�����rU�Ŷ/�!�Vb�K��݆r�����2�����)���Ud�3n;
6wWΩO��*���7���FL�Qp�sk�C�9y�	Ab���Kb��P���e@J���䲶�_�}ygX�xhʺǍIRI'�P��`���4�O2:h%>S^���pj|盏��:���Cqnw��$>����*4�d��z[�P�ʹO':d�i�z�>V�|��z��q��ߎ�Pk�В�5��v/�80��4����I0�ڢyS%i4����L��`�n�wAV�k�9��\!��0Ɯ|��k8G�������u%����Ƕrǋ�Y�@hl��<�;�u�u��F΍Q����f`Q�8�ɱ��h�k~k8*��7�M⶞ӟ���1�W0s�wC�����A}	��7�7|5��.�*�c��*����c��w����n������-��K`Q���~yd`�$���-�T���ƀ�L����xp��BCBuf�p@#���L�Vz��F�߇$8=��'�=|CO���p@Z�1Ϻ ��ù�m)El�~v��������E.5�q��>8;��[Cd��'�P����c2e��m?u���-�+���ƪ��
�t6��n�@d�D�i�q�� @�_��/�����- ��ӻ7�r@I��G���,������O�KM�K������Ux� 0�)M��6�6z�ڟ��5=�7�.\�5V����.ٿ�P=a3��54��W���1��}	��s�;�u�t(|���G��p�͵ "*[)Q���������n��'I{,yj+Wl�`�!m������f�ݟ����!e3��3ޒֺQԘX���9٤�$��d>�,[PN�x���w	�w}�_Q�z�\�����7�[�Џ`��J=C?3�a�1%��z�]�SV #��W�^2���n!9e�N�}����7���GUnMp�3��+~(�Z�^zkL�����D��p�>+��L�jt"��TZ~Q��C+4��Y'Jqlu3�x������<��sq`�^�U�Q^�1�Y^�l� ^!�W>�<���J��K��6��r�6-�ʤ4'[�{t[�Hmm�J���y}�A��n7�I�	+�狖�6�K���(*k2��*�\��`�u
��������O>��YE�'m����y��j��1�|�G�~�_�,#O�ē�`���,���K��Rs?�@W"��;1LKQɾ��2�Zntz���˗�rL+��U�K����Q8o�\x��6��Yh�;+U����-���� �mPU]e���_x(g0������Y�e{��.Kj�O*�:�6�_O�`�}��(2�{G� ��Q!N9�=�:K����k!��͒xSv�1�_M	͙��.X�x�jE�=I�� %ܤ��Y	��Fp��%��H��S2��Di��"N;4$�R*�y��3��F!���W����r��I���B)���aE+�:r.��5��̈Lǣ�YmC1k�t�,ř�O�l2?[}q�'_�V�r��T���"����ƮdS��;��<u���Q`ӷu	����;����g��3�Ưc�_������ۀ�G?i��9Q`�q��a"��dE.��1�}G�.\�3�~gz�����3�7�v�4~�˵�v��E�{���Y�V09��ZzpJhS@�(�$7�"��b��ҝ���6���翹�2gx�Ϸ^��"�5J=;&�⭫�VQ����������u@.P۟T�3|m���S�)J81�%6��s2�@�����֥���2�ϝ���|靓��gs̬U�+�9kn�Y��+'Ε�1�A^V�e�(g�gg�V�P�TɿE����W����랧[���P�-��h���	��X>D�U�kc�j�+ ���k�&
t4V�����Ǹ��D&x�>����
�D�U���;����muS�'�y�kx��ɲX.����ώgo�T��m2���*�T͈�_p��qQD95�RBZ22�ޗo~^����IF(E�z��	)�h�7�N��>�ch>�b��'�l�+	ǒ"��y�6|��a*
���@%�C�c���6�-�W��)K��Յ��OK��.�e�q� �w�y���;E���dD#3H��#�^ɵz��l�U�eu`e
��<~� ;�A��Gd�,����~�{'L�������(�Zsk���q����h�x�9<�'e=�4�0�~9�Y�!���!����m�/�{@ק��Ye$j�$�n�X��&D ���!�E��|a[؅:�!%��G�4�+����;$��_��/0����8���|_X�.z �I7��,�Ķ&F�K���&�NƂ�_���{d����n��Q3Psm�0�̩D��/t��/��æ\�R�v�Z��R�Cs�� �4�A���7��]@'�H�<���b����x/���У��sNo+ʙ���vn��/�\+��?_;s�	����ƙ\�RU����.I^�U��#�S���m��r��t��V����Bo\O;�����S a�N�~���1��v�/�a�i4�����v��(;t�A-���D;�L̤Ta:�$����Ӂ��6-��C�+\��26�_t�e�T�EB@�[nR����hm��3���-�A�c���	��l`�6������<����we�Sӣ�Q
��y�M0Tx`�2W7Γ� Ґ�d׵Wuu�[ĐU8o���2�EQk�	?rK����*�	�������T�oK�N`x�}���Wuǻvb��@��@~�I�Yy��]I�d�j��'΄���W!:0�Э�,��t�E�KA�ot��Tm�����(3��e�#8o*T���ڶ�Y����&
]���E�@90������s��ذC6�v��J��p4&�~�$�3�"��\Dn�ga��Hp3�3�����
�6e����OLN9ˣ��-6��=����GM���%�C,NM������<f�����Sp����r��	�A.:Xw2,DĎ�Ww�F&⽬R���s�z�#�,�� �d*0o�?��ʬ4�������)�ǳć`�[�j�Q���`��t,D�)��O[�wx��X��u�Kl�L�ա�m"��P�L��ظM���ϩ����v|��LkX���� G��"�W��T�M�r�6
c	-WI�&�L�Bo��D��G�H��0��"�q���[� '��Fն� �@�,<��ߍ��V0$�B靧�	W9���s(?���	���bE�}��	�:��{O��6����/%��j�gշ�}E�UR�e�V~y�+E;IcY.k'���UM������$rU6؛����E:��d�0P�pD�^'��-���#��{\��-���(F�f��$��ѨF6$��*���F�aW��\�g�����W�pRD��o(2|�W>�8���׹%��[S!��lV�s��v�þ��*��*K�4O�g��t���~�������m���<��?h��d܊�p!���>ӧ-��7\�#�{5�{:|VA��d@�m�.E(�G�b�uӼ5�����Ww�Q�1�c�:VYd�Ì^��Ľ+�jT�(���\	x&��RϷT�N��L�>0UI��1)��^�47��~��7�Z�[�/�gte��?���¤[�g\�G����d��*�-m�p&MR��ØF�2���6��N4� ]
"��R=�v;�_��7P�2���v������Z�C�NEnx�UW�����(o2�`²��l�R��љ���0��Tp
k�!�s`��];~���#,�3�6˙00	�K��|��8���&��;8��!��A}���Ȟ�@X���K����J�������,2��2<�K ����@&.�p��Pk�^ ��Zd\�S'�x������Z.1�*�և%j`��]n�y5��Ku�@�x&qT�[�_�ǡ�%���� s%������?7ɝ^/�@I()���m����E,&2`t��F�/�E�G��]�6�U�_��oU6�l�6�����
^J�h�)w�����5��r8��".���ߥ�nc���cjC�����ej�&uP�ڕ4Ζ��{�n����0J�/��t@u!:��⨭*Z9����"?��$�ú۱�q�3l�8��r$�$Zg�*�̡�"څ�o���Jb�^��2��lȂ�E܁��+׳���$6��_�f��K'����n�ƙaS(ho��	�!�������L	��ƮzI���P35Tջ:al��D�d���T������nC��F{W57�!�-��ƹ]���z]i?���~�9GL.�_�j�Q��`�?D�$k�q2*��&z;��*���'�ss�=h�ٷ༈�q�
2
�,[- �ػdSP��=��r�W&����(nq���V_vd$��pF�ݞ�I&��}uJE���/1����h��J�	6.�<!x�G�3��L�a	h.�\L*�y�f������@�4��~��� дS�:���o�vA/�g�'�� �5�R�t%Z�������������L+��d\�.��dF��`�f�a�N&'
�R9�y������֑!g����4��%�	�t�DT��MȆ&L�����t2��t��xR��
Paq÷00F)1EJ>�`නQ�o^m�?�%��0�~�����x��R���Ķ��$N�"�2�_Xv���:o�2�-�;>&f�'�,é�h�G�z$4	��L�܏��w���DLn���'CJ�=�����X����X��ԫPd��DV��}w���'1��i5�[{F'�	�5 Fp���4��W/���+éyL�ޕdW��L�lo8��4�,)���?�Nb.n�U�1�9�~x:3��4U<�;TR���-(���� s}=�^��V��$���i���;c��ό�Sݠ��e̦��s�vۀJꡛ��0��x��c�,�\&L�����-N��zL�����Ȗ�XH	k<sqҙ�o�\����2����#C>Ћ�@��3[��6u�t��۶}�e�TG��ӈ�@th+zG�~�6�	F���@`�L���ҭ��_-��	���3����f�����u�,4g,O:J� <@0�\�m\�ʑr~��ƺIX�-���~@��������_����C�����	\o�K^��E����է�����AO

Qk�8 ��oj{v�{$ݳ���9�a�C܎琈��.��c���r �I�En,� g�c�$iGLŀ�v(m���bDB�J{��8д#�Fq���Qg���G-��Ԥ�er����o���h����`}s�?�L��s�hD���Rn���=��#�O?>�*�Ƶv�n�6���y��1U�gB�Ւ�{���|߂ޜ1e�v���
BX��Kde�P ������I�PC:�ʿK�e��T�oƨ�'�o\3}@��Ƀ7��c�C�љM9:��z�����3D)����lnF����H�j:3�������ߋD9�<��f��n0�x�-:s �;�4{17�Vt/P!ޟ{?��
j��@�Z�@�U�Z_��ه�y����D�r=vO���>�F�����ȫ��fc��|	R��U�rB�wu5ZM�������|ѯ�0Mx#0�}�w�k�꣸��L<���EX���lt��ƶ�uR��>lX��(K�D�׭��F�j�@dK`�rq(d;�MF��n����9�̨����l�~g}/������5\B���u��K��>�}ZA���_�r��̽Z�����Rv��˕MyLTp��B���)DsEΈu�xY�5`:�V6�)V8�B��R�^������N�[��u�o���;�����k��J���׭��?��I�i+��D�tP&!��
��!q)����
CRH����0����,��<��7Ͳ8�M$����2�6e�K_�$��c��8�ZZ�U߿���[�-uÐߗAG*�W/�^�ҭG���a�M�&ŒE
v�B�G�6��a�����=�'�{z�+֑h}��8Z9��� {#�_��.���5�%ȇ2��>pH�gK�A��(�T޻���{�*�������g5|}���	�sV,>��e6�h��T�_������"�[Ch��ώ �v��n��B�<���3����V~�|1?��)��4�8Y:a@���Z�ڐ�0��!Y9
��q����	�L��c��z�A��qǱ��k�&�B�W�A�gm�t���=���j0au����1�m�U��f'8,��lXJ\{�?.��#.�4>� Z��ڹC�"M�Z�ż�A(";�#3�t���d���hH2-\Gȸ$�h��{�b��F!B�LO��7Bi`
���~����t�+E�H%4�k�)!�G�i�ش~���Nf�B�h�x�^)��u�勡󠤙r��|�¡_2z���_|D������q#���ڳ��LEKD�"�ΕRjm!���d��JdoK��#&����4�P�hl��rM�w�m����JMFuHU������-����p�Y��U�>Vt:�{�_bw�� ���+�8�O�`������R������8m]y��Y+�%	��,���^cAg�t	븅�99�B�Nl��+�L�����l�|�/�,}ucv�Gz5[m�J���l����#�Ȋ��g���Օ�4��8���he�<!Y�%�Ȃ��C�E�WV��t&>���Quh�汸p:|�Bf�����]b�����:�<���[J%Ysh\� ryf_�J9Q>����_x�O�\�����?.p��d�X��-+� c�ǹ4^6'¸�	U&gW��k�}���/:��,�_գ�3IO4��O�䇰��q�Q��O#�N�oNR3�����ԑD�υ9����Y�#�	B6"O�0�W�;��g��~��<��7��������^EV�W�A[-�@���L�U�l�V'���R�X����s���]HKm�>�׹}�
���ߞ9�W��\+Q;�aLc�2�d�4��=��j���{95�7Ҁ�n�Dhf���מ|w�R���{��E@�P�S,`Q��7dp��oY��X��Ǐ�YB�	!�̥TS�]����IT��Z��s��7��^��h\��#�2Z�?1,�����<�~�� ?�^KH�u�Ɖ�V��H�W�?:�9l��
��۶p�Zu�&��SA!�Z�Qfψ���O1B摹��O��ugD�UF��Y��������Tk�8����	h	w_�j�����Lͻ:�ڞO�f�9:����B:��(�c���k���4ꭼ�A� p˜ڞWM�]��Gtך�P.��U �.[�"/�~��]���&��l���%o\�[t4��ԏ����b6�yi7o֓}S��FY�1EY��[#��}\>��U���a����P�Z01<}yB-f�=Ti!<!X5����\)>�rɃ-�	�(�-'!����+�Sw�q[ܖ���cЎ�\��,&;MްK�g\Oh�fE� �|�}���g�-ˁ�|T�z8WVpeT#>��(5}��c�g�ѳ�/��^��O_�F����8TJ�rט����HӤ�.���c1��L�)��N�d{�J
��")L�ك~3��9`\���N�363"*#-D���n�,xSOkrd�j����>A�����F;����r�OZP�O�|�Uq�9v��T��6���H�-3��Rk�HTRh�Q�o|cY�O]6B�Un�P�݃�G_��9���!��JLR^~d[�_�j��M�����e*��|*�9���oL��<@���F�{6෷���KE2�����Xߺu�g��°bL�H�F ��W�O��*�U��Q_��P�{X�ٯ��ݔ#�����B
X�.	A\�����R�h=�[%A��=�vV��Ն~�!� �����;���2o�{-E{��~s~e�ًVq�d;�՟�O�� �a��yWf/�s��~X h��h�4+�_����e'�=�섒ڤ²��;�/U�����NT��\;�P��RߒG�o��dg���8�G�t�z�����e�:r�C��	6h���bURf7��{W:�jY�!����(�w�A��AIī�=l���P�������,�%Y�n�%@\TƯ<�cy8�"�a�c���4��GC�;�o��kJO�&��L��GK�)54��"�Rk y�Lи�6������*1�b'*�#��6�!Wq�vdn*��:��g<�wտ�h���
�P��F�sQx^/ּ�3���7�@�����vI��+T#Z��@h盝�K,i^�Io���J��H��N|��^�cJ�~��a���3��iy�[�f��ؘ6�"�U	F�C[㤫ҍɔ��V��ɎAd^�")$���U_�w�������Nm�"�/a��M]�:/} ���N3����~䙣��m���Pq���H�����}uPP�6�m�|К�^\S,L�E�X �N��Ўn��-��U�7�S |�/d�&h Ix�&d��y��bS)U�<�����s����y�h��bn$V��=�6���M���{þF��E�d��/J����%��l�	�tM7������TT�j5,4</
����n!��G��s�aQ����`OS��3^k��+���G?ܥ_E|��+�:Bʹ^ɳ�h#���M��;���R)A�.؎���x���hj�����3��?~0ea�Z*~����I���/٦�,���:q�Z|�[�����}b��	+\�5c2�v�v�Jס`��SDr׵���R����Y�l�HԽl�-.����^	�:[.!�Ӵ��g�bk�f���{}�ur4v@�6���0͗�R���ӀP���?�7&�an�߮�V��N��`R'b	��	m��z��/JCnf�@�1���r�:*e.Y6����m�p{+�_͓�̟C�R�z�zJ�.Ζ#3�X�6����T��d�p=:��>��qٴ�X���C^skq�qZt��\�rH�q�����I h���dn�]�v����H�Y7�k�Sݚ0�;��#���g$*�//J#M&8,��+�,ZJ�NI�����\���nkڋ{E���mQKDd�n�|�@�`_�|���fQm������d���W2�Jږ��Al=򑇨Y�-t�!�_6��.!K3�?�k!կ��
��|?i��$�z��,c ȍJ��<QK�!�?�.G����c促?�}E�Ѳ���=	�C�FE6��<���Ew�~&��V���V��w�#1O�*����[��C��?��h�/)L~z�KR��e';��7I��s"c�l��R��i�l�5�c��:|AΖ���T}^��;J>t����q�G�A���&�S�/�֦�r[���7�����s��S�9	�ύ,�!���s�]!��AyK�}㹸���u��o��ݍ��oU<[1�T�HOi�1!&��C��w@3π�3J�A!�H�0|z�M1�Zj�	�+��kW�pd�	� Ll��]�04s�1�MSWK���VoA��F�mg3o��p��U
��GK�{�E2{N�S�q`J����_��1l<�5p#����(�l92GP��~o=`�E>�|���n*��K���V�^6Q�����x(a������~�B� pP@���zW�|I���[0��#)>:6<����C����ǹ�ةt���5Po��R�i�|�FNYP|���OͰ�4��z2k���#~�D�S�]N�4��C�������Q��a��;bX�3���r��?���uwgm�^p���%s+��t�!ݚ��f~������26KҵEC�؇-
�pܧ���d�U��]{�rq�ƈ#н��A�r�S)9�-p��<�64�#[95r;WP��J
����n*b�Լ�xx�(�{�m�`����@���7�.�(h��Cod
�ذ�V`Y������D�W�L�s�/B�i�n�#��/Pz(�;<�_r$˭h��8,�'7v�1b%P�g�r��0ǅ^���V��Ռ���~V�Ģ�i1�R5f"�9�76/mV$6ͮ�<_�����3�Xr})y�@�:�r6��`n�^�%��ꃽSԀ���|�ƨj*��Ae �Z�O;��S/`QC�T�hvD\�r�1��ԛ߄MĮ��ռ׺��#̛s���0Ӥf���#R�MM����#N�%nqn��0��p�J�;��GG��W%+r�N�{SRH��"�U�!�:m�������}�׸*�À�r�r��DQ�"��п��6��
/ϜP]y�9�a�`W�z�qi�8�E`�a�Kx�ПC�w'ە��r�����cjCl�x��E�/��Q��]Z1l]�(��scp��[��X�x����
xAsk�w|��T��Kk�*�R�ā��|� ct6�ӈ�9h;�S9:�wSI&��4�!�����w2�J�j��?\\�4ݙ�B�k���F.쌀�(Sb-�Yur$Rfb5�3E|��GlOu��v�m�{U��ԙ��`/�8�m��3�v�M�	~<�K�o,���X�o������E?iC/�{j����Ń�%2i�9�����94�ז'�n߫���j2�S��޶��By-�Y`	��k���6�=�_�ĵ�Υ�@��2�׼���_�J ��΢W¾�v�.,Ѡ��:Ee���>&����T��W������d�%��I���tc����#���͂a=���t�O�(&*�?t��`ie�0�K�,GOM�ԙ6"8LR�P$��d���� ���G ���^2*!��q2�X�"hV|B��Bx�GU�_z�#����M@}����%�oy���s2�_Zs�- ~D�����-P'HN_�S�[3�7��xu�0��q���\v��K��0���l�sٚ��������Ea��nB��P���v;��i�l6�Gc�W�g����# ��ظP ��m?���Ou-(�3���r ���)C�n��GM��Βe�s�#�r+�Wp�n�p�p���ٌ3>�Iy{�0�@ /M�V��Fj��R����
��[_�`�;&SY?lR_'�������6��dZ���*�oG~ra�RJH��5�3����x�}H�+y	P�R���ty�g�g���mH.�hh��<2�j�X��Q���f�du�@1��ئ���Wv�l�̥�.��t�-G��Bi4؟�[`�Gt&���0g[�>���7�_��ݘ�a�� �$��X,���(6g�1�"o��y����3Y�p9������Ve]Kt݇�S����s阬�d��p
�/@Dl�24"Q�{kFV�tZ��x1��9Ě�rA�	�.��w�b���!�փ���
��?}Z}~����Hu8��R���m=������4��8�����H����jII9_KB$0����n/3�Ν�,��,��eת_��hh���%�ӈ�"�w��&���F~J�<�~���F�"���+\�*�!�^��r�BX�P/y�����ށ��-�䢒&���#�}�n�xC�No��ƞ�,�.i;]e�p�/(p|xt>����/���G-]OB���p��kA%?�������:�	�H땰�g�@�E�ď��4������ǲ�R��H 8Ze:��:7Oj�	?�V"�Mo2�r�Al���C���I���2]K�5�Z\-,�F�R^4����iAQ���i�<��ܜ���A>��m����.�b�е=�\4��݇����X.{�?f6���T��cY�C�=��๭���ǥltv�;���ϷZyz5�
�3J�>�'R��D��ي�EA�����Fuk�QX��yUg�㥙���X�xU���(O���r�ii��a9��gǌ �ځe���"������C��+�:��YB�x,Y���k�
oc�	VC�(����&9e���T�:���æ$�ޠ�~�|���M��M]>Ⱟ�=�O
�A]�c]�cG�q&0a���W���M���_n�b��Yԟ�f���+"�'H%��ƻWh��ҭ8к�D����Q����J$�uCg��&�vm�t%�x�ՙPzgO����d����!r(
RlS�dҪ�U�9�ar���R�r��j�x~7=�}=�,-��gU�������O������#4�t�yL� �bD�6y�����5����GH�#$���ݗ��rȦF00�/i��ӌ5i�9�+!ܝyi���������-Փ�Q����t6R&�ʣa�f�#B��1�ؔo���z&���V8�qi���o�ۑ���#6�3`*/��+�w���V����J�3B-����p��k�O.Lyi z-d��{����A��$I�wm𯭕�ߎ�� .^�K��%Ԥ��w��a�ct%�
$�[��$��F���.�dc�$�\��l��8v�
����7��9�ky��V[}V0ӛ���G��w5ۖuy�ZV���~lo]�������;�G��� 2,��,��-7�f��k5&q��=4�-h-�>iSYex8�^+US�Z�u��|�������ۏ_��6$��͆|�aaME�Mr�g�����mۿ+ꝺ��&�$����+hL� �$S���\����R�!T��>ﬕj�W�=������G�WR�&�c�G���8�w��2�czB����:�;]-;�O��P�+�pw���O|��E׿ƴNd-L����Ԋ��g��j���*Y5s���1iw#��Tږ�����
�W"[ev��6�y�^�yc~���/��>e_�HU�I��� ��D�4u�w��q�~��>�_�[�����mMט�jA��jK�_5
���U=��Z{S��׳]W:^�g��)���ǉ�4�9w7ˑ���)�v�Z��y�R��J�E+%��m��:�`{9ue'/�6�"�WT\E��Q��k����m�)O	X��ּxʒu&Dw�j�T���eԭ�|���w�D�N2�"�<2�����5mGĀ;�hh/ҡ��2���y��xБ�����z�����hȼ[q�'�����'&�[�����)#H��)��l�A�}x_�\�P���Z�îs����/�%�o\*�N�=G�Db�C�馄T"�g��(��+_�RRD��sZ��g�T��kr:!s��b�.O@�{c7@��&����<˦��=������z�yϻ,�˲cl�d�w,쩄p�p
�����C�<Θ���6d���N�����[��55q�;Z�SKY�ĭ(��Q�\&J3�'���JRK�+y�Gi��&�H��t���]����`q��?�Rp��a���PQNC����i.���Ǵ@�I��ɲ#�5��s_���^6�s���yV�&[�6��`�Aq�Y�����9���$XeǑx^��3y����%2����9T�q�Ɂ�l?��������V/v�������d?&��a>�9��C���+�x�2$q#�Y��'S�I ��
n�o
�"��\���eb����+��2Nl$����>jc�&AS�X�q��Tz����K:N��������?�X���ë.L#���s2Gɾ�� ��RKY���1�7��i#�N ��t.�s����p��C������[�
�'�9�_��uY�;�������L�ͩ�������aM��rf�#a�RK��s�XCf����F�@!(m��T��*n>���;�"�t�.�^Ԫ��Ӡ�����i�����Iq��mL ��}e��h"�}���fO�?:�:��f˽OѤ~��S���S���9�"Є��C��#�U�k�G=�� ��������*Jk���� 1ȨR^�U� Fl��.d+�̶��3�^�
��y����V.����.�3�H2�\$�܁��*�zΔ�
ظHxR4��x�+U=���.�.K;u3���=;�)�dV~���7��� ʪ��L�r�Ć��5=m$��T˺��
��E ��)��b���x�bpN~�? "������A�ѕR���V�MMd��ٵ�IO�`I�2Lq[:�!;AEM��Ft�^*o?���xp�/��Y�~�#j/�'e�/0,���_�}
�S�� V5ۋ���5U�Ҕd�����BeХ5dDԓ�pqq'�3N��d��q]��ԚA٦m�u�y2���ީ���,�o(u���>J�t� ̷z��],Ҹ� ��_l%a{�L��{���yu(�p�%%{&PDT�P���7�?�P[1w�my���r�Xiv���h�7���������$̓+7i�5!t.rFt�7���p�<ݔ�p��|�������Z�K��-���w��ʫwV8��9��_���lnJ�q�.?Ӭ �����Ï��ՠ��!l6���&��̐�TT}��<�ͼʶ\}h�hm����͏�Pd�Z� 7/�0�ƨ��&�"^�N�^\>a�j���O����C|^2��7�}�l��9�qC�j���I�y���Ë�د�c��~dCj�>.�N�4��\���'	��`����045����u7��SڑY&��D�n�ߪ�Ä:*]a���R�Q��}[CS�\5��P��!��#��B[1{����Kn�t�u<�:��u�#�L�EQ�X�⴬��ռЍn�>"=�Ӽ�Dˡ?A$�2�Uw?��j&�~���Ɩ��g�R5;>8S{�Ԩ��c<A$B,�y�\_�t��(g`!�XQWkQD�^m=�0!!@�����pZ�f�|B`�$�X�zŶ7ܿ
�D��։a&1�N��X��މ"R�"fK�H$��6���1	�Q�5��Ԧ=�)Vν���ׅF�ixC�}xv��2|�:����� �3�N؀�5�P�2��<s��,Hʞ�h�W�z�����lͰ�7h'�z�\���gd)�v<��'MJ{��}A5Oo��<�S��`�	��:��Rp�{�M���22�0��#�D�]��tw2��E��|����@�l/���y���/�I�#F�S |����8s'(�Z�i�?�[�@�(�ώGq��4��h��������!#(0z)LPX3���]�-}�Z"R���`l_�N-��d�#Gdq0g�Ň�T~�B�%G�r"��h�KD-��~���{7�q��[��*��% `mL"�L�\�q#2<D ���}�֋��
��NL�����!��Ӥ7��c���6�Tj ��%�Ѽ�r��F��J�'���g��r_l�2���d�,/��c�zG�f�NtC1�d#!���	�f��K�g��!�@���Ԑ��q�_�(c�@b#{{�#$�٦�z�q�q��R���R_��C�Ɂ�w9HLYFn�����ܩBϛ���J ;�����\��)��Il^�3����P��S�j��.�H6�C����. \����F�h�t�!�]6FX
�*��Wsx��ﱗ����a!��cX��5�9D�z��>���aW�?��Մ�VUaY���Nq���^.��U���?�f����K4�����Mؕ-��.�_ك��'��5�� UY��<c@�����4�y���$&k��6�4"@B:)3�%��!��|�M�'�pƝ5��غ�����Z0�ޘ��<�3���h��ϭ�ED�Xk$�G�Tİ�}���\�Ѭ��#��#�E�K�D�D9�<G]�g���H8O���S=OШ��;#�r]|9ߚ�T�&����?}�?Q������Ee3��Й�{������D*�]��΁�9����\��)n��Fk=e��6Ѭx#�?��_�(��z�	7�jx��;�HvXn؍f)$��۷�o�ڿ�Ў���=�`{�E̊���RywgI���`����X�/7���Y(��q<~�;�"�s= ��jd)�m+���^��(̍	&2|�\|}D��ݯ<�G�@�]�}�92���^sBܘ�ԯ6A�>����0'�����R�	������k�f���?
Fu��W���&�!f�-��.�2��7<B�)@@` ����æ��!�qJ�~���7�X��z�A�r��_!Z�43�B�P �.�k����V��/Φ|i?����gҵ��S�y���GC�{�y'�/Ö��������'W\9��h@T�s��I��泑>�[����-[{q.�L2��L���9gG+Q��п���S�[5\S��1��He��R������w��o�qbe�w}�������룧J?&��?�Yzis7���ѷ�9d�[�d���B�b��h�pob(ѷV0|�{o�[��@����YZ��	���h��i��HW��QzXv1L�S����P�ё�?E:	9�>K7@@�1�E藏�U����ުZp�p��>��M>�Tsh��Q�ߦ��<m~�%
`�ج�����?��,"�L���M\�����9�-Y�l�3$+Cq�퐛TYUz����d�u d��m�/H�3�۱L[m8�q�����E�q� Z��Xii����� ���q��6��p��{�)���\���ed��[_qRd,ms�56�Ӽm�%�����_�c�|���?F�ѷ��.�K���������%�#��N�0��]]�%�݆���d�&"�@,��߬���� ���O`�h�:u
󋫥G\0u!h����_�Vw���Mf ,�_(���(�kc�+ag!l�N0�<�뺮�L�����$��b�E��O��Gj� [^�w�|�s�#TvܺSԸ�ܱ���a�d���c桻bdh0��9�̾�G��\h3�3��j��}��63ё�a���j8ũ˯���J.,l�`ٙ��3����7]N� �ױ���`�w5}Z���O�~���d��/e��}Q��p�2Xno�h/�.A���������+����>�����B�=}���,q*%���;'�߁�� �K��0����!t��V0����=��%�V��?�6�M4E�{Y���묇���a�mc���H.WN�'��r~w'6¢�����)�/
�md��e�pm�
����1�(T�{T=;��X�����s8�;_�))����}J�~�H����3�)Ni�0��C9�Q���b)y���8�+�

��3x�~����5�V�>�1n>|}�@-֭)�VNC��2�r����S$Or��)�脢)
[�@w_x4}���S�`|E���SN�K*��ֽ����3UܗO?� ��s*�����7�v�}�#尻ޫd"j�ܛkU��՞�����Ϲrc���c��۩>�[�� �$�%W�]U՘��Ay��6�3�߫�QDC���TP�4s���d�
1W������c�yõއ~l�B�"I�?ҝ�z�����ȑ,k��y�ĥ?�����Q$1���4��LOY�/���s nl�>�r�d����\��:l�f���xw��H%�j/q�%�S��C"�Y�(�ښ��pP�ܠ���r`��N��z}�^���L�1�P�d>�a���Z�æ�1������[b���C+��w�����;��h���UgY�A��'�ԞH�Iڑ���#[Q�N�9����P8|�'~܁�pV�%!w�-_�geXf��E$�j|�c��]#`=H���[�u�O����!~,�=�y��s������>H+�x��7X��%�v@�OA %�(�x���_u�A'VНY~�f���lvƨ=��Bf�9��]3�C�A��Ω2ր
E��ٱ��P�q=<��$�d��X<Xs�EC�	�(�L�%��ܶ��jH}�i��<e�o8���>��3?J�`��([��W��L�,������7 �^��H$�L����R���.�L�/i�?M�N�>��	���Y����ОG-�Q�kY@�ߴ�F+�nxzL������Ud�`}��֋. 
ḝll��}��r�|r'�����
I湺�U\$YxL��� W��vh9��CL�TĲ$��u�l�6��M�S�<��!��ڐV��Mh�}u"��Ƚ��b��ap��G�,;>�K0��'׀מ�I��x��4��\�%g�;I�J"ߌ9g�ظg�3��J��/oX�F��C����+�s �Io&�i��e�l�,/[2<��Bh8��4o±�vB�8��	�"�0��$R�9����	���ݺ�O � �k���f�?R����d�b@��/�G�@N��)�<.�_oC{%�R �Z��O*��y�cE9l�ҫxs��@uw�pC�^ũO�'���P� ֩�./U?X?,.I�c=J�l��J��JA	��R$�x�6m`��Mz��M���j��e�����ͥF(��5ƘWP��F���_ �0�_��̶�$�E�ﷁU
z���K��J���A�f؇�^���x��Cl�,y�R�C�t�ڶ(\�Tx7ҝE��_V�>��u����	ls82 ��d�T-O�W(�vkc��UA/E���Nw����fj��%��:Ǒ��"S���m�a)e4^)�,,Ƒ�d�ust$�e$-�\���A�^�����O��4�+���؋������tU�����W,��vC<�Ti�cE��d�C�w
ߩ�>�َs����X�CB��gh�u�"�W�`18}>|`r�98���hP��7O��)�{���������~�v��P���\�E8K��&�܄'q �T*��#����(��v���W|��������k��~�K<���=�)}"G9)gL�RIC*g�`(3c���#A��I�J�ө�K���z�r$��WvU)nPp����� �Y��Q��$|^���Ϯ�U"�����-�����~�hh.�j:͡���3w�"M�+Ir��z��#�mrT�v��;F)�*&7��������|jf��!�Ӯ���Ȧu��j����M�9i��t��#�Iv��̕�%��?���R-����}z5�a��w�����8��a]�-�V\��)4�Bƈy'2Zw��4goډ�b�D�	�٣m���y�&���b�@�*�yF�N�C�{��-���z��b�*���D�	X0`�{n�h�6~�5�EU��(Z	G1*Y*�K_���Խ�h#}ț�'��wz6lʠ���!�M%�Tw�,o�=�k��"7���=���l���C2&�~h�=�zC�J�i&�I�.)J��2ڨ;�j#&���O�n�N>/�`9�->I�cBB����xY��r�����3���/���R.�6C�*�?t��ݵ�W���Z�\f�6���:c��Oe�LK[OIE1��}��Z4��WH	���!�P���#m M�b�̦ ��k��(�'ŋ�u���HG�	<H�Ӽz �0�ދb̡z��//z��u5�P�|�	���ګ�bV���8�������������$^� �0t����9~�El��J��̹��r������,��õ}�A�Z:m�6`0-��o�,}ot1[��5�o�dT|R'Zx^���f&�,�kޅ��iB��lpkj峖�s�����r��_�B����g8J��g�S��V_��ޢL-�-�<=�:4T��iX�˟�0���pT�16>ڎS��t(»�K?�^Iw�$a\f'p��b��5��,X ���p�����}y3����/P�V�&|:hi��J�Lz/��1"�-=ʿ�؅�����/�Æ3V�F��|�Y��� ��64�4/��]����C��#�#�}�;��~�޸�Vc3��=5��L\��ccUT��H���X�J'�;E�;��xɳ���^�S�cnbV{c��^-wL���a�?��Q<ȤOg�ҿ�@N�����WI�B����j���7��,8 &�����'�Y�U�[`V@�)(�(�0��a����ϒqc����vb�9�ѫ�q�"�g�hW6��?�gҮ�v��y�O^�Z�D����Tq�~�i��''W�i)�b)< �W����˩G�4;�dlk��J����<��҂>�vP�2���&Ǩ�e�UɊ�_�G�V$#�>��Wx�������=���l"�'&"´DT��r��&��C�.�m�.�@�X��;�A`��p���A���Ο�p+s%��b�T��65�g�lm�/	r,P�r��G�:��~�$�	��c&�~��ҥ^�~'m��κp	hNiu�$3����B��~�F�UO�Os��B��M�Sڮ]�=N{9}�KV��cȦ����$�8@b�%e�v�tI5)��� �"1j��Q��.d�r\�[cM�FLz�.~d�6���ۭM�Ĳ2h0q��X&����̃����s�'�l�{5bAkn��P�*�77n�����4�mHM؍�PGcj���\7��%�e��Lhi�� �S��L�ո��ǆzz������,UeQ�ۉ@��6��b����@)���B�A��u������ځ�+������5��0�b$�!�n3��F꾲NVi�;�E�d�!^�9�a	'�ӑ�֤�`�)��O�&z��<勲��Tn��C��>��F�j��"�/ר����NU�$=r!t��?��P��x��"�P?.��ې����:!�*
��@C��՘׷9�[D)���UY�����f��]S��e7q�l[l��c��ai�r7��z�<�df��2��a���S�V��&o�j�V�CKm��0^X`M߰˙;���9���?��]Gv����>��|�#���P� �\�z �&^�����9xvfc2W���;8���X��,�ƍe�j(S�m$��R^�CVn�j�$�9���8�|�7�N�F���F�N��7����1]��J���(i{�:Yk^]�:ƎzHl����b2a����C7���(a��7\��H�D���z��\�h��l��c�ߥ:)Q�����b���zY����ĺ�wA3�`Do��x���t.p��,(c�6��&�o��*�{ܸ�l�*X\d��J���h%���{CO��X�J������3�rG�*_ANT����ݍ�X���Xq���S���h�����u�pN&��o epfw�hb^���� ����3�_wfIS���KIz���}i��ƫZ�'^T�}1�K��O�[Y�-GъŖ���pp",���/˔�#����)��`A��Z�y��"�"�ﴷ���dp����Q
>*���x-(�Ʈ�Z���x�������n���R��8�h9�r��s������pĲ�C�J���p��ڏD�����#��d���(+�_�`����1�0������ܓ�%w'@��R�����\{j�����7.�'���>@JU���_[���m[�j
$�+�� yo�&���ݘ2�_����|�"��S8���M����.Kt��6M��U��l�u�ht�u@,=`3��q5���HX�x�.d�"M���Ќ\V����p�W���z*�l�Vk~��W��*FshA�,_2�������J�v���q��
X<�������+��c��N�4��D�5�n؈U���Q�I1�l�)7�8#"���6�Q���A(Dm+m��2��(rf�f�iN������������aݵ����{sU�A-ʼ:��{��\�z����Q]9�{_L��m����&��$7��*G�>2B���ʎmU�R ���g��c8VT\{z����؛�)�Z�(z(� \��7���<:�!�$ֻ)��"�Ѿ�a����ic���M��6/oɑ�D)��1��i�sx���H���G��g��w���	�;�KC������xA\V�Ɋ���d�m��u��l�y�C���Q�M:��X��>����������l�j*Y��0������[`��u���@w���;��S����]Z/EDbQ���GBQ���-lw}?�5�[@TD���`���ꚨ���}V{�ռ�Q{�T�����u���)�D��jid��$θ���A<��Ji%��յ�At򡹳����L%9��jR@�dr)<HF�����Ұ�!(�&hU�l�H�V);E������Q�@��XVNJMܹl,tYӇ��Ga�qѯq,(�	PKpysn�Y#���5���^�zv��1�:�������O
���L!���)�+	���8 BqD?��,AH|UPb�e$��&�f�Q�V	���mݵ,��4��b�\|����}d>8�o��r����u�����:$��f��^oo��5�O>I�C!`��6n-�$�Aj�d�^�Y���425�:.!Y]��/�i������ 5�	=�I%>�I�%��cu������8E�Hңϋ13�.�؜�>��*:s��lQ�V�y�}�=H����U�R�Kw���D���50m/&>qWX�&��Ə�p��6�<�C�|CX��JXh�.�@����H༻���� [��:�E���ί�T�.�5����>�E��p�U��h��1:��\��4�&@�'�s��-4b�	p1�0hR�R����'�I>-"��x�b�GJʝJ��j��C;[�8�퍴`���A�G��_���D ڞ���}8$k�)��@]��/��u�U��I	��D��؍�������*K��J�Y%�����ݲB�p�D�o�����{o��(/�
���w���7viU�Q����'/](`}O���Ӓk�q�"�Iؔ�?��j�i�a�9ـ��IL��E\l�����I� [�_+ ���G`�0GOS�>��3�
3��V�m��4ESv���u�h!�J���)��
n$�J(���Z6�E�@j�����\�,�e0�oLIA�j��md!�����lw��sv�b�����.2��m�l�r��ps�ϠGP�8�]�A\��#Xj����DGى�ˊLF>$x�m�YFTnR�I���2�`7����^��52��&hK��v��Zkn��
�鼰�䑀��)��qJJ/��Xk����,�*� k�/������u!�s�Y�c�6�KLI�+�$*����O�N/A����d�3́�jw���狹�I�k�jF��y�h@x�H��%����d��W(Q�;6+W\Ը`W�q��|`�뫧p��*���B�^��:_/��a+���.�ٟ�jrh��
��G��̑�Px��S
b
�Py�؂��i������|��g�{$�|ߑ���F8j����<�[)�*N�X�ݾ^��D���R�r�s'�z�2�r�k�T�0�I��p"}UR?�����w26<���Y\�/���������
�����;��L$ *�ޫ�a���)�ÞNz�:��G��	�E^��
��}l"8�+
^�!/"�q}�.��B�S�J��F�h���ϧO��`�߼\��4 =g;"��yC)�O�m�Ym ���GmA�nT窯�4XRhM�U�k�!c͘����.�싟E��$�z[�k���C��O�N��I���6�Y	l�L�/��W9XJJuFL�d��W��ҹ�47�Z���H ��U����Q��T(Y�� \��L[�_�����G0�>ޫ�w������i���p2~��]�{ H�*�"�;�/�J�-\v�m6T`�VS�˦x�>v��Ʋi\���_
<	�y�$�n�m4��O�ȋD��3��.R17:G�<q�Ҽ^.�h���h`g/��R�# ��6�A�| ȓ�?-��ᚳ�я=N?V�w����=��l��s��s�|@�3���)*�)o��[�2�$�FȳN}J�T�7�	��B^�U����>���TL?���������L���?��5Џ��I?\�� �Q ٞp��-]K ��7�;���x��&�o��<�ea>96�$w�?�VǦ�5�S��K����H;��Y�U�YYA'�ȭ�}WhD����E��P�����U�+�8���h:UX
�y�#�/��?��̥�v&HR�<�]Ny�x��f�܁<_�KuV�0ͪFlT$�̀����+2���p~ƝGpUBbݔ��hm�2|�9�XRBV��x�}a��d[ ����WF�����l�h���;�X8�0���F|3�܄��JϼĹ�|�f0q����L��KrEkg�3�Q{7�G)�`����;���~U�t��1�(7�*`N�Ds?o�M�i�?�?�v��Rn�)��t��݅N��ޭfjU��?�8"��g�7����оv˥K�X���7��
�8�?�ܾ�̰�H?j���P+�',�s�|%g��~�;R5�:�2�*g��ވ�D����X6s}�gb16Չ�
P$�j�/{�'��}�0=�ͿF_��?j������Z��a��ʻ��x�<Lfi��n�&覚�
yL��T��;?*T�}堋���0�[���ԗ��'TB�NA�y��r^2�"�����|���C������EY5��V�	����'�%�ǡ�J#]A�JP�3�=��	����K5r4�d����n��XvG���3ޓ�IαZܠE>���y ��`T�y��� x�,IŃ�Q��O'1BV=2z/@},�ŸoL�ӑu�[�ڋ��U��s8�zM������#{��$z���0!�|����V�(d�.�5��k��f���2� ���ux�1;De���v�bZ��2q�7���K����1B���A_�7�$|6�EH
)�M�@*�.7g�VfYDN��:�}��N���	a�&w/��=܆��� �"1$�R1vRp��˪%����� uM��K~}F���Y��|4ݐ�`,�,��F�D��JO)v�nt��ʲ�\:N��^��X�.�|,"�^�� F��B7���ہOʖWg-���i"�m����}lc�a4�T�TL�i݉���/GK),�E�
����GJ_�o鋶{8��E�XH�7�\�6`Ǐ��w�N[F��"�{ֵg���#iL�5
�č=��"[Kޏ��
�[���M���9�쭪���MIO7�h������nXU��Ptru~���c���\,���zFYM�qo�rO%,p�א��"��n�`����B�2��Z���6��>[{@
�c0���uvG�O^`�{G�/���������bޞ��"��
Ýq(4R�^��.����E���~b�q�tI�������5������ں�#څ�Ԑéu*���)mpۏk�`Ұ��7���b%D��u�ʺ2H@�*T8�o���(����H�廢�L�?��MR�1:L��LxO[	GtI��GGWvbc�Y�:����qۧNd('N86���c���no		(�g�_[���N��N*��}�Ŝ����,�֧������?·H��������X��/��3:�gUaUiQx8�?�$�V]!r�&���hDi�=�^���ǂ���/�#B0/]�vu�-�^�phۥm�:J��ݣ�(�*��fRu*`V/7~�ԏO�w�"��مqh}�����֕���HdLҰ}l�~�����p�RZ��,��b*Bh�[���a6�4���d�C2n=ax�ퟛj���{�J��L(���ˢ�l�|Tz4�	�_��D����H���\�ćС�U��C�q���W7�Q��5��]nh��;�8=[����t��丐0�U�;�s�;EH��ON���[iV># ���� c�R�	��
foVw���d�����%�[G	�%���U[�KA]�	P�u[���}�M1Ӯ�e�ڍ��E	��0!�3��h:�O ��w��I��qǩ����\Q�۴[+;����u�y��Z۝�Tӭ�����釐�*�_�W���x �c"8�H��%T��Ҍ�r��Z�)�%��P�xt-�ӃZ.o��'�8L( �k�)>�]������WKT+)&?�c/牼GR �(���Y&�:��Nep���'S��!$P/��xX:�?��D\�nWt��p���#l���A�/��Yɱ=�q%Ro�V�(n���A�}���W޾����;�������Ζ0]\��с�#���{/����^� F�����OQ�d
����6�#
��t(�U���_&W�>���i>į�G�r֖�����,�ycGe3.#��.(,�{��ĵ����䜒����)0Я�#g`�L^�[�"�y��}X��d
ɔ��˼�j��f���K���HOD�V�J�<Y/̖�h�im3�i� *��H��d���O''�l�i�����?�V�@�h��In��Q�XmuiY(�̊G�g1��i�S���>����On�Ia��L%H����O��<��~H(.+�fF���L܍u-`����� ���,н�C^m]��kH���&�d��4����¬�K�؄=���}�c��.>:������(�[2�I/�D�S8�7��|zΈ�u{���A�%nė:����\�Q2Hђ��.(+�y;���NJZ-i�������j�\֣�{���""e���юZi �\R�u�|�T�v�R�J0�Ƨ|���Y�5.|l��xr�b�CK�u\����91�̖;dl'�b�F�)���6��z�i
��_+Ύ��ۨz��H]�!E2�� �w ��ʰl(h&x���ڪ�hBz�YK�J��l}�����6�Wv|w�3�,i�&�s"�$���|~@M?Bi���|�I�X}��`�ް�g�]�R�6֑���q���0������+؍��}�`���A���,P�Mo��ɬ�Uqy���PFE!���� z��7y��	�Ϝ��;�jX���(�֮�<���-\8�^�"��*��9!�2��z�?e�o��56��mfɳ`��� r-����k0���]y����ꂗ:�E�_5	�l#���N&�Hy�vQw��̀��p�d�+��\ƙ�Jt�L#����ǎ���p?	%���Uo�2���'+!��1�ܘ+�@��L�6�цHE��6]�:��g}/z�ɭ�f�CI�ͬ2�|�2��MBPF.6��' K-�k�i�E��*�������o��,(��?@�0:��O� �tf�? z��Nt���G���~�L�
� ��w�U�^�-t��'N��k��m<�J-��;G	*�)�`��s���#~�/xn��OW7<�f�����������{�58��3ۊ-F�ΠT)���3�!ƫ4��()<�(��Ͻg�Ƅ�;�h�4ʟvK9�@��Y�E+�j��Sjb�hw��Ȏ��L�� ?,��#h��v�����(S3&�\��e ��Y$\���rZ�F��m���`(�|IǼGD��H���c����β�	��%��A�7O�;(S-����OY�?��vG�ޘ�
Gp�\f��*lԍ[lM\��o�ހb%���R�C�$i��<��>ES��@}���ƪ�yM��f�l��d`���!���P�߿Z�W2��+m����R|���$����ػ��Z������ϰAuM���L�pU40��0/3�	���HY�՝b�T[S�>�q"n{{�Qd�M��-1����y:q��h�i�3�rPȃ��e�/$���� ���`8S�m��r��*6�iֲF�ک�ji�{g�~F*�����?HآlR�[���Cb��(�L�����dA��ҡ���?����`;�|�a�֎kw�	���{�z��ww��G �1���@BW�+tXx� jhq�L3�7YK`�.C��oD�c��|c�|���M����~FB?����<ml�.������8��̳)p1*�b�Დ5P)ח�Ӽ`ػ,�E�~~gI8��D��>X��>��^���>�:�[-��p�<����Z7���5`~�oJ���t��w�.�@�I���+�)�&�~�b������p��mЌ@_��T�����Y%��A���d}� �����a�b�H]69�W'Wf�2;����/��%�P�\�aH�����2�$�i��=�i��
G)���r ��x�y[��و?R+ND؄���j�n�Z�������j�>�̪���2\;�6�B�F@�.���X��M 3A��h[)8[��Z�J��\��D���W��������o�	�dO7�V���8kq@���B(~�_���e�i��M�f�X��c,��%
%�E|(��[��ե���?
�����Q��:1����ȫ�_ϔͮ�Aȧ,Ci�|�b\ͻ/���:�Ό���ㅨ�Hc�K11ŗ����>,�%��l�M��Xx�7����z�l��x�!΂�z(9�V�^��9��3	����=�Y�o�~yu �?ÕP���BGf^��Һhrw�U$W����!/�C��5�Ԋ����~a1ɭY��Yb�Z�U9�6�9��\m`�_t:W˿��U�FuP�V�A��Xj[\R���g�9�b������ b�3�A�R�G7K�043�!0_�C�Oٯ��Ņ4%���]þW�$��	̙Z��W���Wy��xꠁs�ICt�S��QH�0������4@�]`��/������#�"�u-�ꋬs�Pde��c�hL�ݘ#ڊ��� �k�fF��|�,̮� �ٹO�<�D���O��
���P��ޤ��mau�}iS��٥�����]��4wLʮ�^���Cִz[�B>���^Mi��Px<v�my�d��\��⏢t�,{yS�M\Z�w�4�0���ي���EU��u�rp�	]I���(�N��{��CӰP��]S�5V��j�M¥q�)�- )�n$������M� I��Aq�d���IG�W~-�&�2���-@OO�=�u���w����V���/\g����J3�֬���gE@>	X����-��o����i_�ͯ2������\Ů�7���$�K%���Z$w�nȞN�~X�X�7���T\���h�4k�=�.}݊2�#��x�ՌǠ�)Y^�
2p�"xb @�QY��Xv;]������x���m%QF;���:;��	R9�kZ��Lʘ��r/������
rKi)+��k�Vz@��V��1�#4�ۻ��?XR�f0�-��:2b��Tg�'��3�#���;�k�@�Gl*!6���-���4 G�fa@
[*��Z����G o@g��v�P���ݘ��#�u�҈���E�4J����UDihwN�V���H��Lpt��&�Ux���Ƚ���ϔ{�#Y6��ߠu�C�0��+|�2E���nᖧ3d$�P��Vq ��2ݴVf=cj�\I�|*>�w� m*�Vq)+Vr%IEzZ騥���<P/�����A�]#�����F06K�oL�t:��8a|�{��E����b��E]5J��T�}IQ�Q�w_J-A�����=�d��R��;,�#�g�(���4ψE�����^4�o��d�\�Գ�{9��`7\�U�x��#�h�L��S���2�-��CR0�mlȕ�I��J�g^�Xκ;�٠x�'���%��R����
Vf��d���&�k��y�ƒ2b5.�͘�'a,�����gILKWewA=ԴB珹�*�QHmb�������Jj�Zl�{�2?��c���k����P"���^b�g�����c|�4g��a�R�h�s��%�ʷ;,)�>��\�ծ��__����RWx��A�*z|���C�O�RԊc�
] ����{~pɐ1�.��\<���_�<W��Pz�������!��&�l�Y�W~��?��{���X0��J���&�`Џ���v�q������S�5�6gZx�p��Ω&�h�8��7c_����>Zf�A� �kt��5}MB�N3@�@�_8�j�S��J���E7�.�s���t��t.����a��=�(������B��z��+&�;U��ڷ��GNX�H���v�3ȼ� W>qP�x9OinR�/?�GֱNԟ��2��QJ�
Zv�͝(ka�.��k1��~�|d�(��Ʉ~���@�͜Y]nEmm�(�Gj�Ngt��v�N;���uY�J�$9�E����+4����˳-���6���Ήɸk�=S:4��-Q+�fBH�D�ˎ-����?�ZߓE��@a�V��oo���)9W��p�o��|�h\쵺'#�}��Ӄ���mm�P��g�ߟ��vA���٬����F.��οQଉb>���!�0|�&d��@O};�'����w|.�A<D9Iv�՞'"��;��M5�l8%/���}�]��<�o�UM̠/.<._�X�� �-���<'���ԯ�9㤘�Z�FE~O�R�����:���/�O����$��n��9���|�ճa�gi?Us�xp�;��6؃�|��,�mi��ꁳ;�e֟O�Y���f<QtK�^��ng�-����
N�.�2`��w���;.���;��;1�D���p���2:p.ޒ�8i�V[�s�E���yI�6�F�"g�H��U��XWMC�?�__#Ď���sx)������ؖ�o�DT�����x$��sI�B��J�S��н��������"AD���w�e�]���ALߨ��ql�R����ъ�Z��LF�(�KH﬐�o�O��P2���O�x�@�&V��O�Dq(㑑*�˲�\cڅz�����w��l[�N����� ܦ���8�w�)%ڜřA"����7{�`nr<%e�͞���
S���%3�t
�~�5��Ǵ�!��"i ��m�V {�s`l5δW;v1]5v���^�GY�(���Нy�47����K�%�`U����ԭx4{Ǜ%�0�D��-�:
���Ŷ\����A���K��mk�>����
Кb���,�b��L�L;�?݁��Wrh4o��o��pc�L�L-�D<��~,ڿ���`�
?���5�?�4/�
������Ӌԕ)t��1�p��S~�ķ��Y��3��Zv8Dǐ�"^7s���)�v��2� 杞�3�p�6�$�d�����"O����G������&x�,�l�N�ޔ�6��Vj�y�K;vC��{>ԟ=W�{�eK<o������3C��;xDߴx$�]v�ٔQ/����k��(��,W�V���
����X�S��eg��]]��M�B�?ePb������Y�[�F��0�����t�����-b� ��ّ*�d+[�.�^�$�Mw}aP�����.�?j�7��J�F���*t�J�g6?'[������ye�)LǞX�Q-&�ҝ����%�EFuWn�q2���]�<�
��#�^�iʪ��caZ��&i��#�b
ܬ���ax�~M��1�˓l�yBb�x�!�3L+特��e����}���Ͻ~Ԏ=���|�vޝ����#���������ì�� �͐�ic��&C,]*�ͅ�gՑ��ӛ��-F�jc.6��2Siik��3��Ww��F���{���r�g�?�f(~l��#N����M�k�;q��+�F�u�J!�Yă� ~`.�"�/�W�g����v����\-�4�NS>��Y���OL��6���*ܬ�`Ć��8i���䢜"]�*)Ty����R����<���c�x}r��g��i��^�kЦq嗜MED@��kj0ꗀٳ�*�����h��.��m�Ħ�L���G�,�}�6���-��
�� ����5,��C�u;Wr���~��(�w�lR�O�/-tÎbwXH��X[���C�
X��T�̫�N0��"VK����Z0FM7A=�}�6u�Z��Z�P���������hv���;���s���K�������(�8B|S���OO��� ����F���jHŦ�.�PM4�^I�b^6���$�' �U�Z��ʻ83�B�������3lB�˸�'�����F��nn߆��[�j�j�h�0Y}���������{,���8�̚?N��Q�&z�R�P����[�z'9Pس>H,��2�g��qt�	`�{w)|N_9h���$�s��"l��"ӈ�]WB��	BG��P4|�؏Q�%�˚����m�8� Ω2&C�)9���&6+�&�%S �j�_[�<o�1��a�`���jw�;�yޠ$�JI1�"RMm��l:�6QZ�x���O~o�]�˨9�����6k1|4��bÓ���+t�'�xõF��R 9[E�E~*����i�>�5`P�Ӹ����A�Oݸ��z�.����{)�a�5�&E���9���[Գ�F�����Z�0�Ɯ��vn}P�����&3�&��3�����I������L�X�L��T(Ȥ9������j<������Z-����@y�b�[f5��^d+��`@ v���,�Zd�F-�L����rj׷G���4�+����&߄��$��Z��"<��@�Q�g�4�c�;�ʃV��"��f�R��?�)�O��X�
�T���tTJ���+�o���9��|�Qrz؆�g�EK�w��I'3_w�+�]5#��]�6 �f����#1z=<u���h��,�N=t�h� Ƌs!Q��2Y�����B��P/z�$�6���"�Wm��Cz���LInh_�Z�u�|��#����<j�pQ;_ab�Y��旍U��܇���֞!�`��@^sg\{�����+�/��ײ����<a���f�T��jB]e�ɫ�#;ԙ�I*��������{��\�@��O��qb�P���Mk���s �#=��
y��XS����8�\��a��������J�ԗG��[S{P�lX��~3�#�6ǖ�o�k�ٶQ$N� ��i`Q��C��8���r��t�9�!�l[,ޥ)C��_M�m�;O�W<����HͿҬML��3�v��"�����k���l��و.���ؚ/�'�Xg�6�g����Q��78eMsq�%Q�9f��� D���I_-3�<���YHU�ψ�OU���D�6�^�q��CB~��p"YSk"���
��#I�t+e
cۜ�XC������q�TNC`�?W+ȓ�J-��}�_�=v�����X-WC��^��!8ɜ3�s��n#��m�0��O�Si�Z�j\��4�����*߻1&?�����V}��
B����->>&֞hT<���h���{ё����l$��E|��s�ﳔ]������ ��|LL�ȰlȊ���hr^�#ϓ8x��	wI��(^:�1��V4�#.����
�v�Q~�-��_2��G���_�͐���[v�XGBbAX=�|�拕����T/��=�|��d]��e�2?|�qIn?�����GM/��\�W*����_��Z��UƇH�z���I�P�P���^nHD���bg��+JO��k�U�tn��/3� �"T��Zp3�g�c `~���ӗs�_�Bi��*���Ha�ػ@��Z@X����ˍ|h!��H �S����fL�l�s!��_#<�������������y���{߄R�Q�6C# �.v��Ono���˗��*o�^(4J��E�� �䷳�.^��̤��cj*��p4��`K6��2�7���fl���9p�*�}}#���čST�ZC�D'ى��2'���ƛh����o!:��co��.٘�V,K�6|��E�,��/��r��F0Gtm&B��D3�R�3у��N�ɰ�Z�L7mҞ��y���������N���i�	^��
b�z[�3�)���!g�O!���:��.���_ P��C@{7�p�����/�L����H�h)׃_��/kJ�WJRl@�@�r���*<=Ȓ�'�DQp����AX�[T6W��S���Ir�!���#��x��-�����Q8������`�pü�=�MXoNCCrڕ2��+�������0��	Sr:?u̯��+1E�A8�l4�c쭘������Y?���9��f�E��x����6�Ax�i�V��� ��p܀(�R�_<2���&��K��{��h�*�6��~(և΁�ȗ8��	=����o�9<��$ړ�53M�S�����5�d{�Zf���O�<8q�Hh�v	���M+m�T+�xK�����LYo�o�nCP� �!졇�>�DX vE^~*W�Eß7������a�~��RZ�xy7TK<�U����)�W�太��X�x(/���0�Ԙ���O i˥:��]���%��w����
�Ay7}{��~v�">����4CXiY���s<�qo��X��%��|�(>���Q��+2�����Jw�#��h�.K��2���~���y��5��/��L1�����Y	s�T�s�G����Q�S c�}�cM~��JЙŁ���\v�Fb��c<c�~k%���5�Z��!�^�ơ��;E0U��n��qCa�\
�QOsH'Fbi��^7\������,�΍���
vx���������ߕ��5 :Z���r�ܒ���ȸ��JT���;��&��؞j8Y����#~�⃼��_�VX�H^��}X$������@X���Q#^��C�YfԡTmq$��Eñ�!vp��X�����9�Ǫ�\�P(�� SR.�b�����9D�@+��k5��&WƑ>
/�.�b�����ꠚk�t.p��Y�� �t���!�����G�4�<w?4�E|әDa#!�e��lFj��\z2��[�	:1+�k���>�ۆ;���4��C���5��TWLX2���>�1ؼ�jB��ruB��2J@<z�R
��.�E����G�,K	��C����R�A4�W��{����~}�(�k��k��Ă�rm}力"�������C�+M���d�^�Ru�r"�끳^��=r.e]:�Ct��c��˯j�d�o�h��RC��&Ð�Ҹ��h����A�z�R���hڅ����4m���iL�s;�;��d�۵�e�b��+8-%pD����5�-���XKQ�"�~��̸�
�Z�}�Э�q�/�W��߷*L��`V�&	�ti��	����͆B	�}g�R`�I�j>���B��u�]����*��V&g;]�hy����k\|���9(pȄe9y8 (n Tg@�]�:/V�s�UZ���Qؗu��9�)�H8�Db�ֵ��5z"9ۮ8@��(	��ȷ݆���z��H(�bx�5�Ġ�!q����D����/yR���11�L��'{yb��Z=f��N�x� �R�b�?�o'K��V��|��LuX�o��³�9w'@^�7Z�G�� �5@�Y��챍�q�@�giQ��Rnl9r@��2å�9q�uO�Ə�O�w%��
�q�t� =c�e�ޚy��Ȯe�~�}��B�?\�Qw��-�W��p=��/����P"��AQko<n��PS�ԓl�)K��)�)�J_�ӕ��L�Y^:��8���Q���%N�ϤM0\�d���J V1����o�H�W���rH���'��t��z'.��;��`��Y\D����$� �7@5Ɵ��������T�3�PN���f*�h�YC�xŭ�d���W���%!��͠�-�64��p��C��;t����u��i�'��xhF��
����s�|�f�/����!���[A��g�+��
*V����S�Ph˴ņ�t�\��@w��r�Un�a���T
Ѯq�&�%�^|E�km��%�X�D����//_�2�����8&�-�0,2�;�O���>�'u^hu�P�x)*�$����Rb�����_[ռ���	�0�H��Rw��jɞ�^�$�
Um�%��A�����|�s� �ճړ6B��ӊ)^X���>�Q��NF_{�1��G�ôm^�M#D1��dW�-j�2��$|�������,0&����2 ��p��U'~��IG	+P��ƻ�R�{Ğ��

Ў�u ȇ=��l�^o���o����U�)�]�5��^b�Ä�u�
�����#���R�1y!W(�%.7h�K�* ��}+G��`�U<�ZL&�Z���1V���F������ٝ�����غ�vU�Q���^bh��X��C8�޴�l'�EE�]�N$��v�l8�w�S���������1��QME�n��}1rd���^��@����[G�Y��������s��������3G�H�x>]��E���8���9&�29� ��%�`/_#��QW絉��r���_��6��h\��44�&�.��/~�0O=I�/�"������a�2��ݣ�Eֽң}yn���rC{��'`D��'�$	s�98k��pi��*D��~�j�B ne޺-�@WY'Oav���;�KƓ-g�}$���;��PO�#%|d�1���o�U;��;2J@���+���{w�{5-a�}��Q���o����Ż���i�8h=�C�Q�?�D`�����x��t�{��uػi�����ғt�(��6�Ȭ�5�2 �z@tYB�c�q�:�ew�9o��	��[�zӛ^�L9A��f�ؾ�r`�������D�bc�q�N$���G%vb�0&�K�vSܡ��SQ�,�K@���q�0�����U:� G��le��a^zߪ��K��D������9@[^����
+kE\�&���MA�2^���v	�VwQ0�ĘY�{���=ξ-����3�ñ�A�1�<
��_�"��^�
�U���ѓ����ϲ�a�#�PI>>b�w���(e'􍺫tf���|��Hb{Vt�hc�t�UZ׆�[�d��X���?� ����r�odAr+)�u��&,�9'�9U��9�q��5�fC_�	�Pvmt^�-�=�ܒ�>E�$F"��٣h���f�m&l �g9.ք�#�P_q�>�1��'�L@V�3�ʶ�� Y?F�m�'�U�K�a`��z4�߅*�/��`Xk.����a?����ew�����{���/����s2����ċX����ԏ��~��>(��LןPr�m��+Bi�I���`9�]!���}�?W���kT�*���]D!�n�[F��/�{�K���q�j����V�R��zp_�xr�����>G�=3o�J!���l7��(�L�0K&bVry����h�rU�+�M4��O�$	נ�Hy�a�]�z!�������T���ͽho�p
��
��H;+����,�s�y���͑قq&����s��Z ���s�G9�B����V�=��!�q�;b�I��=�NJCYH���a�!�p6����ʥ�1^'��_�Z�:�?�ǹ��nf�Rt¦@�|W�'���P�>��Q�c�*l��5�Yq�/�����������ÔR�N�8P(B�6�+.��,u�Ӓ�B<�XhĲQ�nw^���3�*.���d#��z����o僠p��u�I����~T	j��v��̳r5t��n���n�S-���;C�P�Ԇ���ӳ;�:�T�Jb��\����i;�bf\��I2�j\A�,����	�>��GZf��]��dK`���%w����b
 ���q�pj�CW�N�l�ܺ�ݨ���Z�ar��_�����2<8TȆ�������1|"�8����:�?b��8��ә�|�8P���?��K�h�NY�t��f=��&խ8�I�ċj���4.R�Y��$������Z(���V�|9�i�{��P@Oc�ԥ雐��W��5�Vħ;0x�Ŀ����s�yx�[����`I�F�r6&�U$$�yƺ�澥o&O%�o��}��;�4@��?΁������:���7���v��:xNkCZ����ҿ:[#/��}�73y��'�͕�F'�6��g�q�t�>��d��x�#��4n��E�F�L���c��C6-�� �^�z����qy4��P5 g��p�r���V��&����D�O����;(����KC�u��������J �B��v�OL����*�lB���0?�w��/�3�,�Ss8�s����6�%6�=��?�@��vaK���\�=�S��]%�%S��)˞�Z�M�N��HM-2M\��9������~Y6?��mӵ��Kv��i�x���}M0�!��Oug�m�@Q~�'�_׋�'� ��Op�z�w�	�y�0.���'?+n%@�d:&A�yY����Q>q���q����|�3��Bl�l���=5�N���*#z�N%��g�LW�*��ٶd�\� {������MC�X��d�U<�gp�>T��b����o%���C5q{v��L�
�����w5$�~�� �������KO�p&����b�'z��#NH� DR��E�"�S,���CB�H���hs	o�#o��`<�3�,�!Ǵ]<e&7�c`_[���5O�5y4b>'�>	׈X83���Z"���҄j��JE��p���cg(�b������x�ꖢ��q#`~)[]�zEx�u�4����?�-=N#�y��>�]&���(CIa��Ng��-hg����n5����$='�n)�^Ί�}/���'�Iǉ���*2�؏'�+;x���܇)�?!�[��!�6�V��m�
�p�>!H�Hl��/�4#9W���ʬ4�r����[�F��83�v"�@FZ�����'�1�-�r��pzy`2���"�M�φ�&;�w>W z.�#����9����ٍ�{�X����yғ����s��ڗ���u�L�G`ɡ��q���:�'�y��F��X� �<\P
�⢅�����o������|��1[���p��W�%O�����v�q;i!�����S�!4*]���;�پU�y�(E�"��i�|��$�4:��\�VR� �~�q��Ǜ!N��4�R!����8�"G�[E�~'hw��Z�1;�Mp!~�o?wƨY~�N~�[~���e�ΏN������.i�yn<��s�.;( ��F3�c�s�%;�;������,Eϼ�;��'O����V��K])��c�f�*'������Ȕ랶�pM�)��՞8�����)ǛNr�(��ї(MV�\WP����!�����Q�M��~�ƈLV�L�*, �4��/n�,��]�^L�FH*S�r�}�>����LJ�B�$�����Mjv谟h����ʹ8� dFd+́M^�h@x��|��$9�^a��t��JW=x���1Ĥ�.��/h�"ͭ�D��p�z��)���~��MY
|m�gJ GUn'a��!;U�Ґ��A���5�.����:���@�C��&�YrݾH��MD �%�h��	)�zj�'�i\,4K�-��vH4� �a�U�������ӂ-{Өr���ME�]k0��P�k�zc����i����]���/A2�����/jP���b��y�Q�N �KOUv�BׁYkt�c�H��1�;�k��]+�p��F01��3ê��Srck��u��#�{�F!a��Ѥ	n��������9�75p�f
J�7[�L~�����c*Lz��Ș���A��l�Wc�6Xb���TpԵ�H!)�W+��$2��ێ��	<-#�b��� hh�k?�[|߯!�%�.��.y7��t�i?���`����o�����>�K��f�a�T{�W�Z�������0�^��R�(7��;�?��^+x��5m��F��.*��K�C��Q2s��8��t��H�ٞ�{f{���	n�P�k��=�V((���Y��]����,Ktx;����jt��B���R�APL�Nھ������5n��k&��*���-~Nb��p���'��L�6��S��#�,͍s����8��+��������
�7�sQ�ڍ|�z�H}h*��ٵz���8��E���-HZY60��p��Y\̂x���{O�ES�^�\���h�柱�h+O�V�-ث=H����Ѝ�z����ŰwT���"�gǺ �ck	�Oa,{.�NX���`�����KN)���V� u��<�x6m��(Os��"��2JK���0{R��H�A9�$�-n��#U\׾/�ȷr��M��,eP�%=5�pQ��'G��l�>c2�Q�Y�,���p�Z�~D(��~�nl]t9B��(uL�T!R��½wέ5��|0�
��]�!N*�D�B �1b�.p��ou3���^^=��y�VMѬ��Cy��Uh^��y��t�҈U��g�g�j�.p�v:�ǳv%Q�~_���P�r"��π�`y����\������H����{�kt��,n^�Q��(gy���
�.����������!�8�����`�*��9="��P�%�֔4OU'�]�t�@n�{):DE�x��q�>Owu��F���N5�60Z��h�n�?�*��
� �%sis>}>�9���8�PH֎Tk�����u
������׍����ra�QN�A�?��3�����9ݶ��P���0�T��:�ȫ	��pq�H�]Ʌ�F~\������4���@�"x�iE���TH��|<n��B�`��9l/��xcZp^'NXDr6�W~w��&-x���ژ	��Ew���Ƅz#Z���$Y��Li�:K�_�#gu����i��������/꛴��/�!��5ԠXLq�W|�q+��).��.�D@TSP\؜Vb).�Ch[��J�C{�DCϧ&M�_��B0<��H�d�@�z ��[�c�`۹#��9	���f��GN ��A�fֶ�a�Ȩ��c����-��8R�WTm��Y�[�ܴ�S�M��-$�%�R��p�2L�Wi����y�<F�yPS��݁�A]M�޵&-
:B�i8 r�R	7��r�)*��Wc!F��;LGݖ_����䩻Qx/�N&܋	ݽ&=��2ҡ�gh�������Lc���`�?�n=SP+�� .}���4�VU�����q��qo?�ƭ��-+����%#�^0�H�,1��w'�����EPG5�&k��E��Ii��z�fj��k�(=_@���M3d��|�2��᯿�t�U3�</dz�_�Iz��I���*o�(Р�;_{��į��m����7V��;-Id��c�䯺ۈ�<ơ
�n���'�Eԗ�F´]�s9�,��a`Yo��9JvΜ�
��D��2^��ԓ�w��hVځ�d��d�qq�H�N1#͌���dv>�U#l d[���ޗ��u�xmo��Hf>��-��iE䉴؃s#f�
��)G_��(��é�Ó�)������~���.����*;�t��6ۦ�_R�Ýn+Y��+�cH��5�:�Z��V���Xt����Ӎ'l��Y���{�77�����	 
1RR���硐C�hJ�7�.��w�ƐM���'H��9D��� h��'��>G��5�c�c����X�.��@Ԩ �q�I�f/\FT�v������:�~���Zy��oG��Mk��8�d���=g���8Uq�w�zB����]�d�AV(W^ȹ@3��O��=�.�3��#l�~���`.RY̦v���"$Hd����9�N�|3X���\�H4�CK��s5����JX[�k�s�H��,3,�z=P�py�vGIv�_t�
]-^B�J]����M�a���3jb��e�Cު~��P�1�D,�x����2oL}���F6jƍ ��B�{������v����"vV����\�x��-�H���� xj܇�H3��P��& ��w �H_��;$��\/h]cc�&-��'c�^Ps�SeVf���T�_Q�!�*�@��c� �V=P2$���3���_��Lt�ߜ�,��	PC[�FHA|�>r���Q��K���F�ϓ1���v�1�I{��^2�ՈD.��ާ�
���x�ÕnZN>����7ܝOt� �C���k*B�?�%3�h#�����A$8B� �b?U$��'�8��/W Ȏl�X��$$�~�_�wSݟ���Bpu& �Q��c�4su��j
8�����B�ۥ/`-�zLąl�s禩과��p��#��f�o�F���
_���I����OU"�i�+�BZ:�����?�J�Q�W�$d�\��x&�� �+��d�m*g�؋��cނ-~�t�n�A�겊�r�=�8?1���R�(i�k)��e@��@��E��'�U�KU��B'������&��"����1�4y.����d��� 6���+,;����ᚱ)��d��"��NE~�n�Þ�o�s;�u�"^�Fc�Y�p�|�df
&�W�4��i�F���e�m���l�� aҎ)�(
�/ ړ�1�U8�#�O3%��u`=��4��09����}���o׬'�w9eE��F���񟔺������5���Uu-����+��SA�&����F�� Oю�!���8�[�T:&�禛v�W�� ^sc�z�����������O �n�E����l[��
!���{1,8��Z���v,Kr�5cW1�^���G�.uU�P�$�Y��|��dA��%��t�q%��)r���4�*�`A�u��u�Ֆ�P��dF��P��%h\x�@N��X�퓇��P�v�Z�͐�)���bx69J�"���[�M�VB��m�Miˀ�����X��Hl}?���ū�B���|�1ߡ$~����!ha�l���i]qN���B������z�5Kɟ���tג���%]�1>��h�|+:�#���$��FuP�5ת%˔�D�ΪtYy9f�Xّ��K�`�t(C�@̪;�簵\}��A�s�.t�ģ��Z������ �%s�(;u���.}	���T�D�v��#B�S��z �7P����hC��ׯ(���E�	:m��4OIÂ��LzX6� &�G�5��O�ށ�u7n�:�+�R�,�h�=��̥CC�/�yP�r8���a-���1T�ɱ^�#9ߪݞ�P��E��| ��#Тf�=�BU�hAc���.�\�Nq��c�R_U�GW�טX�C��-+hԬ����2�$`��(ݸ�Ȕ��C�ʪ�r�d�Oh�s�<��D���d��L�h^������Ш�������܁�NPA�	~S��JeO��y�=�@2��wm�$�FporX'��g��"�jS��W�!B A=ޜoc-�Շr�o`p8FߍŝůE*��M���	zWxpI��*�թ�i>���|�M�!��X+?�˧�w�AR��q�\��I�8l#���'C;��n���ܝ٤!�_I*@k[�5inޞ����NLU:��"��H��J /&����<c�d��$)�j�d�E�0�������eg�*���>]�(�<��6�� ����Nv���nFs�C��w]��h���J.{��;C�7߇B2�١�hA�?����-��܍���r��S��?��~ �Dg��aut`-���[o���u���&�AI2A��I��mCwh��m%DJ�^�
�y����k�rZ��$q<0�֕Q��;��%��i�e��=X؟@q�n�̩���<~�㷪����WY��m�弪E���b@1q��OV#�H�n��@��(/�Ȣ�������QԷp�����攋PʿQPT������wX�@J��~x��~Є%VgtD)�oIc��Y�z�FN����q �-}g&�i�p閹jQ��D�~ì�F2_J<2�GM)R�u۞�P�2oxp��`�-
�c��ꗴ��2@�ȍ���u?�}�� ̏�O��]jf@�	�s�G�S1'n���{p�H��C���y�w��-ܑe&bs�J~s������cz�*MD��tQ�'��޻58#�]����fj>�U!�иU��r�8Ӛ�MG�Ϯ�N3���@/��^7�7C�AV�0�f�c.Q�j ���Z���Z/��:bJZ�� �|��Ԟ�u��*"EӀS]o����ᐞ�SCp�k��э�]8O�� ��A
K�p����]�Px�[+���(�DU �tY)��s�p��V�͔7V�6,��<_MWI�$��cR����k�a����{U��C� �~<����m�ݳ���av�:��>�F�{���}6͟���Z>ٺ6Ds�Ր�'d-� 9܂v�!�c'-�q�n� �u=.�/�/����nϻ� �}��t����~�Byϔ,Jo���X��簽�����}Ƚ�	l��V�]������[D��j���̷�l�oD!D���&?�ϕ[���AOy�y�����#E�Q�jm�~F��os J\�0�ƻ���O2��Dv�������^��@S���ű0�1���u��2����էF���0��4�@X���.u�Bn�]��'���G�@���Z��	JUW��1��<6���2��C�T�ݎ�2J�2egK���RNޟRD��s�B��=�E�d;��I����K��wH5l��6���3�f� 83�R��
��4v*@���G�����\zxI¦9�8�z˺t��ǜz�2�=��zjE뱈ah�^�ɀ������y��cAP�Df�জ��B�6R��l�� �H~o�L��*A���T3	���1mc����%�*Q��n����<Q�[����Z�b����"�mcLg�݂�W�O�}���P�"���뢨� F~���Ny�LPw�<Ԣ��������k`���)f���� �Rq�O�R|1�c�P�89���W��U�G]�N����9��IvEF��E\R^�a�Tl1�0d��J�vR��l�NxUmW�k��߻�]��2������gq8+T0K֜=������)�Aa���u-����m+�æ����I����� w�d*/����7�nZP���� �r���HUЄ7s��&A��16��XߥL�h7�S�]gf��F�d��R.T���'�ù���n�����PC��_ٷe�=7+x{�k�!��etA9K�
ܕŞ��g�r�B���$r(�����<	x+J�9�J� �@V��.l�+��#\�_�;�q�>�)Ϫc�:�ð�I�>���	2�Ԇ�e޳����E�@�ӑg��W:�S�m'��k��@�yZ�츄����'�cr�&?���旸Lu�,����63U# ,��25�sF]Z黓O�%VJ.?�Ȯ	�5�k~��0�Uͨ�M?ׅk���[�OJ�	nO���S9qX�gFxLt,j�s�����8��6$�����!	��L�"z��gw-Tހ��g�gf ��Ne^�F͹ZdĤ� Z��=�~a�%�e*�;)F���Fߟ߇�eF!|�sD1��8����8�*�UE���n�9Ϩ-M�vub��&"�ퟪxR���â�54I�c���!9I5P������g��%)�sEgs��j�b��*�������nj�=��d�H����m�?^��C��$�=�X~�p/�}�#
��$0�K򰙗X�3��^�+t��_�S;��?��51�"��Q<ٷP��7z�F�3;r�qkه��'�DDJ��͂�<������.J{x�y��N�.��_s��|!&�X/�ث4v���ݯDp=L,��ϊ8�g줵�(�i����m�pI�9����x�B��;Ԩ����A%�O���S9F��E�K�<��n�N����YU2?�2�֟u�����վ�����Z�d����/�O�t�L�L�$�p��O��b˙���|�^CO�`-�5�@�}R W�a��m�&��\�1/%�|��O�����F�ߎJ+��-������4�4��q�I��1�'�S���#�
�1���>�#ҡKJ2h
^�^����Ydɲ�Y$Z���j�āz������y[�����Ķ���M���{1�?&Ĭ�� ���D@*�<�1�=�� �}*��2�b�������f@�F�4	���E�6�X��?�M?���a2kc��72�����SR�=l�4
��)�;�j�+�d�Pj�T��0ס{��'p��P�kv%���	�y��7�`�R�j��[� H���w��a�Ij~���<�|�=$���_s�s]D�s��!��b6%n�J# �#�󫸲?�l��R��h���Bap��^��D�ipwNFB��vA����W��Lj�}�ų�xd?vP����n;�'/V,��^+��n ��e@�H�3AJ��>�� ��[#��@��=.��2X��ǝ���$[���w�$&(�-���=���6AN����@�]��>�3v���D�MI�n{*x@H��N�SJ��bh;,�δ��w�'gp(��$�괸�F�['�� f�7����%kQ{f���Nn��q�O���P|̵��&�
���cy�ր������"��}i��e���I꿷p,�P\��օ^J�0kL1�!�ջ�6i�5 ���Y3�*|����g���̷���}�~)W���v�[h$�&!��l�ܿ���Xe���n5X���߮��d�~9�G_�n��L�_��g$�X]|�x���^����9oY{�c����j��,g�T,,�\�p.^����7�eA��,Z�p!��gB�㏊�66���(,݋���>Ԙj�~�0�/I#V� +�L�[���wK���%%K:_b�=G<�[L�l���@Ãi����ԟ~���+g�5�譅��>�J`r�s��	�Qڸ�[��}{�3�V'gwh�,��]c�`��D�
Zvb,,z��:��5ˌHh�v��8���/?T9�,��bM�NzE��pv�VT�p�Ӹ�� �u�+���4Qs<yv�MF�Q���p�l�<!r���Ɯ�]vL�.���o5�1�����6Ԩ�c�k/5���C����g��Nᤏ,!�đ3L'$VPhQA�:��V�kkkB�����䀭e��o���Ɔ���C���츺!��ݵ� �r�}�R�eK0<��3������f�b��ANU(D��A-�[
�U�J?�:����\SJ�)U�4)S������L�U>�I�ፋ���o2t,aշ�_6�Dd)'ve�e������9e�(a��F�����W����+�`O���-��n� O���^����:��L^_���&f#�E��?�����+�Н̳�u!�dp���s�r�����X%ԉ��wQ��=ͅ0=��7P�8]PFq�cWk�aP J�W8�;�yP#=
YQ����@���,l���(]Q����Rm#��F�-ƭ��.�(58�U�X6%[;3�B}}���m���Rm �ap<{B���O��o~�A�}�ہF;1���d���aƏ��6���x�y�Ck�9�D��x��.�Ϝ1�%�E�o���$��gұ}�-�O��X��}VM�a�$��n��]��Q,f��Hﬤ��6�m�����4���ү��}��R�b�᡻1���J��e�p�m�����;�k�`O�s�U��=��c6�^[��{w%,Fօ�%k�Ǯ+��Z��V���p$�N&M	��6��C���%>���}�s���sn��jPF�OY^\�=�(Y�cd+�
m ��=������.�\�$*g��	��l������ �lM7�c��O4�^���#~e�^:��8�_d����ڬ�T�c�Oa�"�oK�����e;]4n�	R�N,�w���Y��C�w".�I�/d�����#4 ~�S�^�p��f}u��,5)g���5�{��X1Q�v23�����<��&=+<�)�pJ����Qv�Je�0a�^O맹3Qs������Hݱu�[~F���5�H&�\��c-A}e�,o�޳p��
��HL�E4&!Z�2�'lB-%lO0J*�~����!���R��A�����l�6/��2Og�O�4�W
A�^Q��m�6�iM��	����+���e�Ss(g��!T~�4h��6g��/�V�y��t6즳��(��{�R���,ťJ��q�Y&[�� �*I�Wa��U轵Ol�hqؼ`����XZ{d��S^�����}��7Wx���$���_Qw8@��(.�����Y;���hmTM����$~w�� c�U��d-$l��D��ImƜ"h�7��+
�mr�bumbd�S k泰q����r�s�@��\�D5
Ϯؑo���ى�U�d[�e��_.pt���K����jd�F3S'��q*{ƶI���Yx ����F
���1TN�����֟������N���\ꔜ�ݵ���r���
v��oRw�&�d�a2�G!� ���]�gJӈp�݋YCLD����g�Jx�v+zD,�~z�Ƒ�����H{0t�h��2�9�����^A��������-��s޳
f)���k�¶ш^�(��@���X�
l3.�s�}���s��w�ˈEs!H���<���f�$C�p�9�:���򴇻��E�u	������K�bt��}J�h�T�)ܛӅ�%�L5�4���#*tٰ�I��ϳx�o�װ��YW;uz��W���rx�Bu*>�J~N�a�����o���A��
���C�c�cUY]��.(��һ��OD�NCX��-������g���u��HM8!���	�x�'{)ٹ1�<��}�����<����Y�U���8�+G>��\,�1��3�ځ�̺�\
sA�Dtc�+��,.	:��x�����q	��:ˆ�����n��Y���W�m0���	��>%@mY��x�N��,�]r�` TP�3l��v�2(o��<vo-��K,��6���g_h�?7��m���� J'Ng�ۡ$�16F������p�ۗX<�Z�I�y��˖�}\�Zb��]�QB9jz��1A?�{�A��ڎ������_���w:-�>J̿L�V�E�ȨPy��G�P7k�Ǽ�e���Yf����"�P�\�W#T�>�v��T�e#`Ʈ���Fc��#h@�mԡWq�!˛��Xm!;ۨ���H�4�Y%dN�����z��ȁ%+T��˼�C=D,���bE��|����om�F�섯yQ!.�?��z���z�s�8U+m�B�0�W�o�w�����-@`m��#�!'��ʞ�Kqq̠�Eu{5Z����!�����R���(�4Ms����
��x=���_LT2��V{�ʔ��?.}��@��:O$��;(��$�͒�L7|�_.��g[Cex�L%�R��0�"zi�ESS�44H���C��eG�r�XW���܌ � ������o	$Na&�0T��Z�,�"���i
:�Mk��+x7�ɠ�Ұ �ѷn.7��{j��a�f�P�{���	2k�1�Sj-�9�ҁ[U���V�AG�Ӳ]��<��W[G=�ĕX���l�u�g�H\��D
j���Lx���ԁ1������XB�=N$
;���O�UB����:� e�������P;Ӟt��J�,=��'tE� ak�:W�e~>��y����5n�`,B��GV��d
B�Kf����; �����v:�\�K��oĬK:x̀��*H�tj���yT?1(�w��a�fe,A�0a��_�P#�Z��b9�d��L�0�`C˙t�r�4�7�ġ�m<�h�!hZ9kd��	���.�X9�6^�����+�Qf�O�0U	1��/X�&�
��U/
�R�����:5ǍF/�&�X��Z�QRm�2�k8���C��G0tI�;��{qu�_�x���:����y�.�ds�  ��Ի
�m#�+���U�d^+�<ԉ�6-@�8��׉�i����^�7J^�x�G΃9�郒)FnJ8���maY��.�7=��.�g�i��}y�~��fx0[��� ✞��		��fE}B8�{xy@_t=�J��c��;�n~���,���i�1�ݦ��˄�ػ�X_u�����/dY��W�y�B"��Q�թ��é-�	��r�0�!�̽찡,Z�Rm�EG�SW���	j����H9}�{�B�|&����N>����AHW����U�8����8���biw#����Rd��`�5{�Gnq8Tގ[�̀^n�^�; �Q&ۘ �,@�In�,R�rPt���ei�3A��: ��W��Cd�Ҽa��&���M>|e@�r�B��n?�R�ʥ���򆪟m�a�����Dz*Qș"�1"�nVR'��X�\��s��(��E�����h��A��1d