// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Tjio7eW6SnBRL0+M7XaegX8NL4gQcLqyVQvMOQmnr+pugdKy0Ncsk4xib6Hi6di4
zRCaUFR2D/q/11Svb/gaIkuXVpVepr7fz2h2dBzG7lkzt2Fgfaj0Jj825gkkuo7u
ATEjWVgpeWAcsNJHYV7uVhs7PV4WKKU4kLmnz39/+O1v2DExoB/kcg==
//pragma protect end_key_block
//pragma protect digest_block
AWBUU6AatRew554BJOGCUxADL7Q=
//pragma protect end_digest_block
//pragma protect data_block
GEiT9/JGOhAKgW/fxY8PI0i28ST69XQUZ6M3rRTDm7Mi62+TOui8b3EkklWLcOHZ
0q7yTbuCXxUZP/amHQcESD06LGNt1ath7uHSABS6Ua1FYF7mvykrlEJyaV8utPmk
y31BpQllYSF6IrQ4NzXXeXcwHUEiSIPBjCvqKw7Oksn+x1yuA3XiHTbZ2IgABXnX
uXgwHGjYhUczfc5nySSRoy2EJKUDeCr4QR0KJ+B90242+02axblsWisoUg29syYy
vJPHinT+bBZTP4hfieIT4+X7VMTHuhkMWR9A6ZMK3DXmuE7nWCY1GeZ/1QntNxpi
m+1x2HSr6qIE5hUTfrjgeFcLpMMA3kq7DH9ZW+mxMb94f1ktn724Z95vDTpiO6g8
960h40Z4jzbt5Es1FOb/xlxjDQXr6Fu/RNNjewOjYF1frzlVCqAkqQtbtpR/RU15
iQpXMtwKbAbNFD8qNpZOJE6d8UhJmnhu1weW/Dx2+WkfMhLehIpssY1JsFcCsbkS
aLShLbdKS4hwWoSACXdtgM8EEQQC+A7qF57ZOtXhYon/2QspOfsz5uUhUH3YK5QQ
1LtuFPqACwyZ9CiHWnA3B8LQ5hFQSQnDlRlEiZZzQiU3Y+7sd6odh3Gb86s1lBxt
blsbMzKohAls5uqzLI0bU1iIJ1jtP/DTeMGxixYcad8EzGCHNYdV4UezCgvTnmmj
wDMC+qjYq4lzWJ/OpnAwoYj+AOezWG4fGCXF6Mts+xBG0GeUC8gwc4eCTpuNSMKW
Vg4RkU2gP9V+VK8o1pgBUkqNIkzuTXVVVO3OskFMOKmmnwQpDS7W8rVFL1PZDTnb
j6M56dMQ7z2nyrhzYP3u2nEBkpDVWlB1oZuJwIRfsmxSstwEqvQpdxLQwp6Uz94j
4p7KsI3urROdk32PCqCsq1Dnj6ZWCBJ2B4fQDXufxM/xdFXXqVstfOgNSvT0uVlw
VjDiRrhpGB/AIbOiJLF5FC3vr5u/I5TTi/Y95aAEyG9ej+wogiK0M76vheYF15nY
SzZI0lhV7BhjUzpxm7tlEAIuYwNVCOnLzLBswLFakpovuoVv7jVOC7NdnzGVDz8z
t8HkpqcowXpgz4Sulz2GYBw4LK3aitvufTpCzNXV8lmBdkxKu8JbeahvXtG/SBW8
q681a9/ZPS/BaygoYuEtPBdhCTs0lphaGCMjesWWgaX4KgY7v+y7vxKLb/DiR8bA
9FTqABfQWxbzZdlXVNhNU61wHf8WuJ5J9oVwusUV26kaJxmgF5sMGafpP5mz4Ekl
qa6PTZjztQHWZ0CaCohXMHz+bh/dOvSkwwIM5sHBRXd1NgkvB4uzu2DDVyCAcShC
2HgZA0Y03Ct2Auxq4EOlAwPOkOMh2FOKeTMSNq963CVfbP2Bn0cmdBdS5HhrrO4/
b1DEDqmFzsriUcP48gYnAUU2RfqU1BvPFN45fbhk5WL8jOEqYek+sCSrlP3GMocr
HVNS5c/GeHr/IKTmdhFv6OXPRyhSGSkMg/7RHiYFPzCiPw1eArucm9K7/y5U4vw7
zWkA8JDxVBTZbXIOG14XCj+aTW50bXbLCeV8nRiKj+UJZIkzOQSVD4AeGBNblsUe
VseiaQxC5G658mpzpwo3KrisawYXDIMxsqq3oKQAaJn8X7Gly1BN8fr+B/5IHani
fO1JlcfoYQxQCR54hhSpJVuAEOmSMpVR88oEsja5KeTyC06lPvPZaDkXbG9F7cMu
RVCyLGyqRpGnUuz+1IGMokbBC0TTjgy7liexGfOghCs3ueaKLNQdIoowUpBPHkvW
E4Qd606i0Q0T2kTM0rZHZVoBA9mU1ECOUGVwuPYvFNcsXIZgGksVNuYJMv7BBTiY
fuVmVKCQQLE3INeqxYC+PdvgrgrehI7XIu+lPGw+qGFe8re8QHWnhnqvJ80QWXZp
xGpNPUeFVxXfrIVmDi2SvMuQ4ZuKycUbwYT1bPb5uC+Z2ao/YKnG7cfH0m8HVIK7
+piVhFf1yZ3lYr5oSqNLXwI2f004vVRyD4Ee1ABnCQU+rmEQ+qDdRNUmSBzQxMjn
wcH+CogyKspDHiQxAk4aSPCBxldiPCw5NCue6dhANG2hx83ly3cTOaU/32knVwfv
Zz+NHCrhzlFAw8/07Nt6Eje0pj5xHyVkRkTi1XIkNxnfUNl/w2a/Nuo9hsfJiI/k
1WTe+6xX0pqWlkB8X06tlC9XAIip87HyRCVGWbt9VixZZW0WpwDcVbJcgUPHAEGN
aiKBDyypQVkYhuzwhYFn4UToXPZcI6b/LtEZU9tc0RQu2QzwKhkzc2Spjndj7JHS
T1ZIQodUIE9AfMAZBlMbwiOHixFjBdxa/kAXFScKXIxPl+ik8Tmt1NuCeoR347Rv
9LUEosblzmEiiUPeDS1RiJt8+RiGNAvSI73pRWU9Pvwo0JP6Mz8YwLUzx7JScnKf
5d8a1fuu7atjTNnsVWl2qsm8AJb3l0FmwLJ/1wxl3teVRV5VMqFI9kOcBXH+/ncg
473tiHZnbLKxRoL52nMtuWkKg1pBEZA1+jMOgbEo6fu9yBwfvfGr9/t5HOauNGSl
59/ukIhMttFtxM1c6rpF38kFFhG6h/OdV5f+0aexGGCNkg8TV8IqKeneGt6BypVT
6wRg+amsySmJqz6Lp1bYZlMfdhOr7m0gGBsUFgaFEtXqJr4OVc+iz0qpCUjQX0YK
2WP7slyf6OmHa/azHT+/v72U55TzYD34OEPy32rCLxNwnfCK2yJUITAOUUGJqu4F
mH667nY2iHvHhqheurQNUr/fopSqgUbC8TKwtAQOXslkphlc3p692q+7T+FuGBWj
f43s46112lhyEPA2KfJJ6P+azaeKbOnhPwyI9dkx046pY96u0vgslJ6e5i0EKO86
ms+X4/bxGRcySKJT8emVrNWTg89MK+0+jSZmh2oTNnBe7Y9QTN7hiSgVDApSCE1G
Ob5xurSPkWNqolI5BdXISYwUnqi4Me3X6P10vR8DlZw4BYmjoxZesRkIUY+i2x7X
nWzlolJQcR0Vlslnz5B/JBWVl/SUo1TZ2D9OhWkJ642tntxBGkFpMpiTxvPXGnyS
J1ovAFPjP4BqPW7z632VsXEuh9aPafGJNJWQNj/f+tj9c6y5DBE1Bpq128tZqgey
MdgjpQRjRSYWV39RDnsJp+kx2Lhp4SmwKfXRLN9nWtRw2aAY1KMBTkZJhKtF68d3
y09aOTRGy0EmxwqpMc57myYkY+PciOFccnOB2E5cZ1gI/uM7eHlJ2wzlx2jDafee
QDi9JWOZThIUuodLk9I3NpqdDV29PE/6oXqZTp9TXvpea9hQtCnM1np+Rfhli6e8
rHMk+F62P+AhesSh5mrN6L3Kf50CxJl05Zqxb8GD1Ea+/WlLX00vd2aPfgWTtXEu
+qHJ5oE0Doe17Z8n00lvxeVJyJZwma7qOTrnALTZ2mgxKa2zuSsc+e640PmBz54+
ToipYC9hLd4S/uk0HCi1/5znNejrvNlu+DCgyyqPFJixTWZAHoXk01309qr8pD1n
1XNpl/xEhs3EZ7WnRvDrXhzJ83ULmFukyIiGBU+zIfINY3WDAbSdPmYp2ceaVcvs
odpDlqB64xiXcuZXQe9Ly9ggSvHTea5h2XdVEavKJmhBtoct9UpK/mBInupRdj2I
K62VYluFEtOM3dlOXC7kOhp1fw/NWsADBEjbXWXSBdmxFuNw9Awey1HwF2f2IAn3
NsgchCfK1mg4I+6DJIxuaUbfuu3a1ROY9i9tIPrDfL8vKtV57fvztAaqi3Kkghyx
GyIpbc5IymQ2R/t5gojVhVq6IwxCxvXJICcgf8FWHC4zTr8nN8zSyc4yMZRVUsG0
qoeHLi1u37r0hOYd40T7pgsa+MjLSNDZx9zrv/eFhmL3U1K7s97j9pDIiEx0cht+
Ew9Q52DUDAxhaYCoNonJTZAdkRYfn73pIuIc2RHbmYmDM0Q7sIDHI1PjUHljM4/t
SR2wK+BjoIcFWi3Mt1gG15gmrP/j349Hb8hPoP9u1xfmyeq5jznnRJ3bTRrBFyAr
MsjiUr94Tqmtcl9wHfy1IEdd6wYkYLBrOXzWUu6YVyeFu5McMnNsNMSnlRu4kMvX
ZAuoBB1ToyFYMltFtE4qjweTUyHbkl44EAGuleMMT/uz1A6bfZxIc6G+Zt/EAKNW
aQhdAXlu5x/acc9NsDQHP/dtUTuFHag1n/PsLX7Bh/jx4M1ZyqYaD5wqYXNjzXvQ
aPMJpkdEAcwQULWncCWXAyp5k9p3d8nLX6PzMJvUAK+KavQ1ei+LhfoE/DcnBFe4
KXHQQi+cWcoxDv0KitTd7uOdLipV7Z7BKW1cqT84hVSwkgwoDG3/s18XG2BiAEv5
e6B84jE/JdzNd7kGMaBS8Z0fP2X17YiziH2KBcJ8BcR4h9pmFXOFM5l6ny3stI93
kE67raPwJYnyvnRGqmyZ4Kf6F5tDy2Zj/FiW1ljy+njB8Y6RRYxWLMWylC33qwDl
I2UEtavwWPMPtXpzHz58XicAlHgPgZ2A7EZNGc1MqtvSbWb5cESlo5EQx45MkfhH
iEVvxgsZaVlE970LOPH4oISz37LZgJ8a6OiF7Nz6Kg2UDN7nsN5tWS54jyMzpYer
EpP9sNKlzxMq8gbHtoptSWgt/JPFHFxDaVKQ/E/d82xH/iiMvl6JvnI0Ayz5V1QY
yGIlzoGmSL/NjYt5ZMCD9c1t62PBw5r2nm1QVcOOpZZkXBLePR5hfEuE67GdgLkn
uc6MNUsWKmmMlC2VMggvuR4aGRxbGXGYr1cy8+yXtLbdZPj8l9IQ9/YsisNgqkAq
8mlxIwCCqTw3v0dKZ/xx3ldiWeuC27R3HFg4C2EIUSPpqOVmFBHPc0elA7I997Mq
6Ra6KJ/YBfN53tOIxH89i/lHC74bS/1sdpGtehhkyzjJhtpZaO09hvHR8FuI6sSK
YsFOHRn9kiXiOBkrV4F7QqF1r4FA5Jji3lBDsLVQe6RQUKiQqzbJsVsG/oshNVne
em7Ff/pryF9LQOg9hJEMHXjSx/pDZMfoYPm6lICpfXI0ekmQfVNoTBGI/XUvOcMQ
r9nSy+XhrGqumdFJMDX+IE6GBeq5ey3KvGTH4vs0pNr0TsQbIG1r7LDXBwLpJJFu
BglNMDa4MAbfclsk88KuZiC+iTqu6sb5DHLa1y2yPYS6f97ztI8ZMXJ9/YRSlnfW
xAmq3i/rVf/vkdDSn0pEk4MT0GBGjCCg30Rtt41dxn3TS/WJU2klkwHmE2ulzWRD
1/bPn+aJzfkzwnFFFIpOD1yfKnaLDYJajKRmQDFSzb/topNm4FVuH/XMTptPbZMo
Ny+O7J/xS65tZQGYJtZjivhEB8BWpM0ofDhdnxbuFB7p5bnOzQZ86gpoUhGJYtYY
DqzQEe2cYVkz4K2lSe751ZYUMCmtBVxdju341uOtcvc6RSy6ZzsIMUKP36K71S/x
egkxzuIUf8RO9ns7hKVt94y1xUel6jZeI6HTIXbkG+PumYcK/PY82o+VtFP7DAyh
ae8vzPB7jzwqk4KsO+edeYbIeaChJs2PxSTLYS/EvNEvrwAGnvsJz8CW+TdSIvLd
Qh311DFR6hftmK1JMiyrOqZsOlTImoWC/6dmJ0OEXKv3Clgqg8okcHeq1gVKSk5L
LWAFtD9rjrL7zP4/M9kQF1uPjKgVfFzmjjUb4zLVrqi9XHncj61bmn5vfdZxqs5r
Rr6RbHfpF+xUFx+l9ME5vEmogxoAtmeVxt9VHsd7gsD+bRwg5H8c8DsRjwMfW/DV
60x1rCJK3c30AQzD1FWf+q2NgVEl/nVJbsrka0/2hBvYQqNxd8+INMUBGmnNYC1l
q27ng6A3W+VFClNQ8AjsWTHNp436VNT6N0cutd3fuJVL+h7QiX5p5JxiEhMt8U2O
hKyPiVvYqLqaDLLdP4iLp9iPcj9RfOYtjPQFmKXJfZAk0867xuE3n7rtiU+Xj5sB
rGIci5MeSNQNiAIntBVk9wv/UTXkMUjxigGyR32sOgqACHTAHyBZUQgHBaZyV5x9
FnZRmc+tF9uFM6MxL8Tnu0Bys1z3RHuI687zP7FY6Zp56nshKLOeAdneaxF6JXcD
NTBQEa62XR2ZZOZwP/VXDQgnODi+TCG72gGc5sSAgeaI/8TLV2zalFEU3SFSUNA0
hkjKzFEgcwH36iAe6eTZJtCtnezWSFhL3FuHZ0qpt7P8zkykl2k4xtuXX/+rXnPQ
Jv6C1xQhsuzr2DZE2VfqxqlgSR55z8okv5CbKbpbMFmqb2UCwVOZfMa902fGUikx
v/VvhhIkjwqc0OO/auJ+RlTzIp2AYDxt9+e7VDKO8HKT7tjdMU50x6Mhhp21slzb
T/3NrTZpRjxx9ZU6HRP7vXtfkFV6bonvZB2tbnGPn6j15d4kAKF8xL/H7RERd2wd
WPNC6I+T3oMC8llL84p8fe0154u/tsT3PxquR3QNzxiF7QK2ZB+SOtsOQyeEE8ig
bpVK9JlV84035tDtU3Y4lbQD038P+CCN+eGQWCzeUGOibSHUUzzIUPi2ebPhX481
2l6jdJIpD1yexdtBcdOlclIZGBSzTWyzEQKAFV+JAM77aOXWIro0ZxpBb6pY7G2F
l5XWkP7GNSBq7Pq4KobIAgOpxBjWPK57oxtwppLKMRKKWQALDwwR/beEHT5rJjbM
ALP5tv93wQBMrzBG4SiNIHb7gQ/tTvHswBOfskU2qNuGy6FhaXr4okvPBJi9fZrh
2QKquO/p79MzPzwddBW5eBp/HZC3YLTb335eD/cDhCoiLveJRt9ijY7gwNph9U+4
8w5DmHaNMopECyd4fRgX+BxzeQbDneo2gaMXJf1b8tGp0UfgjGdM4LmSZkTT4J8r
gMPy0nqcVcYzaX3XNUrBWFbrbaqNfV8AGpJQdHAwPvxc7QUs8MkpMsgeBAHTsxKa
kxy8qpSeK9H9M88Z1v1g4oTc4qNpFfQWNjGt/NJ3oXHt/MnKlHCk2e1k7h2UHIMe
c+nMlMUnkUbMzDZOkONcvS0VMrRjnEutubzB8Y88DHD960pV/rbwQgO9tWvCvPsO
h/mfRUmr/YauM/VOyIam5h+F5oIvAbJnvCwI5mIIbYVyuO8A90x8uyvz7MtNmXvf
37ow8Lu6VopJnth+7c8Q6MuJnpFbd6pJg4H2R0uoQywuND5JsfXbp1fgYhauXeWN
ayzPMTBuFfXtvCVejx65Z116+OmVrxVnW4THmTEmMihwH9+u+JpkT7DSnjzYrZ9I
6pnUyQXKgSGF1a6G3YopJrnPyeO1uCp4hqr53cawq/Q3ft52MNT9ZSd3fWUOGonM
LBPiIFWTA63ETq0PMl74JjFqt5Fx1DJtyylZgYLXb49Ql8PNk05rBKgqxj8HgU6X
Ssin+eJMOJ9lReOfEnVlRu+j3FbgLtdRy6EhtbXElywKbIBsHSLEB4B69UV4DxSd
rQ+eJcoTTma4RC/93/keeASOPxv4WpKL/ach5s2Haw09BatTX2FpjPVMaEV3/XXd
PfGAcXy1JPqofyza/BdTeiR8SFZRXBLD63Be75ZEPKpPspa5AUm/nX/yj3LGdz/1
ySmZBu69+qH7LCrAhuJao0TwLrVEAhKGKpuRs0rkwRw6uxuoJ5Kp82uz66V7ruZq
q+FBWOU8KCNqK62wpx0yb/dEmck5riCrnJqbhmlaCax1724NYhcl8NbgBwnLLTFB
xvVA2rOfuGTCfadpfIV5po2SxnS2T5tWwc6kkfq3XKswKrWcxOSpI57zpY7tSD6J
l9ooEbjyKW9Wa7jfppYv2npQ8mrzk4dn13Du/H0AA8xq+tdAs0e2NlDI+wV899sl
WJUTMa3V+b/yMIQbtXiMj5hxheMFG9Sf14U9o5EmwUFoTX3TuHyJMe0FozimbQoX
1uAUfR0a6Ob4xs6Z+fKaOpBa0HZlyyP8aZFR0GY5uAm8mOu2xOMfI5w+HkKb9EGL
a5eZ54OYkzxyQ1D3Tng61XUdfCeA8J/4i6xb1zQogv1K6B3zd/7zMzVAxn8eNXf3
hGgwha5l4snZ/f/PCAnxuHhbjpKhWOr7ufgNZCAepE19UEsNidHr+X3gqHIv1njC
5qpcdqaQKW2vR0ixHh+A6lKTp7+w+SpP1cl7w3u7Y7/4MQu66NRR8IshJ40qIrEB
AfjKfX2XlgNsjPv0L6J5caA+AbCpIIcxmFOaosXkCGvNh/wBM64zU9QuTP5cxQ9E
tlTq03wgHSVVuLQdn5+rE6jRX/oQcsL/3K2Qkr89jBnjSQOPNawM+NTVOl6/QwvF
h8Pho5cjA19GMsB10L6HkmB6uzwdIuAGChTMDSQH49nYraDifbJsM5RIaEFiwHlp
ZN/DdU0pI5Gzgi4klhzZxjSl+hUeARxra/W4U0ST+vTT4VNGcOmJzXQNboMo+gvO
ofr3R+YipfvWWDN8lr1Z4fX0E5f6qftlfimPhf5FClVnn3wg2zvR207BZdWcO1yT
sn1m4ppv80z+MNcZyUdu+DzbDZAUUdFG2CZlxthlCOsnEVsS3GOj7T0k3o1jvkZV
XB8kUxQyuq5ttqOym05DuuoQRRvwgZljVL+/8RAmRJDiXTp6lFDgDLLD0O+WkJ2O
39bvxPJtBaB2qEU6QkzjEa3YHAOImLLj0dCZE3cjtoI9kXcXUOxL5bT3YgKz4ueP
U+SKeZVX2GHsDPxQmoxUxoRoB2rKw337UDkuwUuroGKa6dMLaiiTU+ZChvztKZ9J
btv9Dw+ctFsS3yqyAczO7XLjIHvQuXND9ex/OFUDVcVaVISQfnMhGF4RgK0UMfiH
Q4cc0sBJDgimtqhrewBfmyh2FhULljs39wyIgHQJFM4dWvEMOajpyqhAkzcAsM5o
FdPxusBDdmL/k9giCre/ByZM2YdhN9PIoaN1drS6d8045Yxnzcym8wsLdfgKnZ5C
F4DP5zpTEzBF4SGnVNjv+LYIcIXmJmYJwqWBZVW+qYZCrexSw+CZQRkctHzMZNz2
IDPI1mSC2AVZ0RrawT2HqckQCHtWCQPTLGtBPZk3DgVqERxOhk510iHDDjvvYwE+
V2vSD0ly3WylDjbcRNaRFo8ZMmMDQ9/NBZ1LGSLK5zDCw9gS4zAyRgNc+k7GzPX1
kfWTgnmmoZn5iJ3yFhNVJ+VXrG1ziZ4cF0612n+nj3BIS/gCKM00ILMkkjDRYvv5
an/m2FSjjzvi4YjaF1/oAjT9cAyI7jr1rTgeHSndUH8pvTUAQfLvHetPlt8/y8lf
XCGXgSAr1XOjovDnr0itgmP1iTuObi878MNOS3OE5f9JM855wCE+ntw6KOB9T9X5
OF2bdBXvbeKkqBd78HjNcMCYAa24nt/86dwZveH5m6WpaktcoJ1NiL7scCDKcf91
HFofII7Ao5srIyG/J04o/puL1LkZdOrOQlKD0Vtnn5WZJFNyiG7cSyeOIhCM6j7G
MOp+YDx3gG1t/UdDheqpo9+vEoUda6JVDHaRz74IZC2Xr5RWXiFSUYbfgLqHuoeU
th+hpVzJu45GHCXFpO8OOLNXEER7CO8W0qugzDrjTiffRhDH1xTzr1LjjBCJHHTF
07cBAG8NruHUi2XaNU2/REJQsfUkBNC53yB9+MwAdw9MtlX57UeLz1aQMQmJWQYx
I1myugTtvHBksDkxv+JGhGtR2RoPRahivi9A8DwXeh4uEGx20M0shzkVyKZOhRvy
pU4ucj8swNPMLfO6P7Ef/uKfdmVQ77PL6ETx4YQI6MQNETuir5SsverQQFiK6zXp
GhnBaw0YKkfqpydhTfnOFgw4GpJFsKFkoqnbiSnSTcA7XbD3gkd13ch3czUH3uaz
47vQ0Uh2ToL68ZSqkKdJ6bJpSUBcvgGH02TZ/5PG7WUEQ/ZZwZisEvPDX7HWR6WR
rhI8tSIlkbQBUnau5JWoxqr3MfduPLTgkkAl9o0QXHOEl2ak8hEUG23SRIfaosll
kRBodelL826iNe1D9OyD+3PIb9QtzB9cnTD4GU7xRbn8VPaeySFhDTuAEZXLjoIX
xMLkln/2S1z8wOV109Ikg2Q7fKuv9kzJBrqgLzCqyBZdVDpR5zFgvO13c7kVpg6U
YxcdwRR3y/mGwWqJzQ7m/i5TjP0VXiknaNMdfHW1M+fQdYIr7Z8us68R0aFLf1Z7
zUMeUDwN1ih/LVZkwTnG6xydWlkflDcFEdLfN7AqVa8N8PL0cPnrc3MMturZdcul
9E56aGwz/eMMxLQ/mDT776ghKPY75NuLmLw0LYTe1FlT3xrN+AOb7LPFFk+LiXcB
L0TWYrE26e5Jin38BnmtSMuZhvVS+vmj7aEO5OiHuVy8sxmA8mOlpZ2Ir5EodRIw
jtmGTM7Ek9nYl7riVnzyKRm2Od9XtjPCE+YvCvZfnOPhyC8Ij7qvcxiRCGsSieXF
3eTqxlUo/HyQYJFx4E9o9r0OsJXhRj3Di1nx4BzcwAZHPtT4BVpi1JSYeqqiQRP0
UzcSIUpbBCyb8sOJSvh83KI7zPtNovoFUnWBBZuvK76SKhRCd0jB/vp+6cN2yBGA
d/VRfqeuK65lW2HBhsNchcyGE3W3fB18rzi8uPyABh/AhzjqIr07tIUcrAXcQVo1
RPBccnfJL1S5NjWAyknSKWvSoiYA2H4aHq0DY09pBj1aRMevTj9Lt4IWaokU64gk
8vjudNFEbOg75xGol7t0NQgHtMJcEgETe9AMeinVGTOcAu6Hw7gRBkMPdt1XuvZo
zk96gAZ7ehUYZL4FAKA9/9RpDJDwkNpfjzkeAimLNs1yKSfcXO4EcOIaYMeZLjYN
lFbFkSlD1EOk7woVIaZupvC8M0QziSQXhZQzQRrekKX0ITWvKX8IsRZVKaLBE+Lf
+6qXQeU6IMJF3pdShf9mr+xRlY38nI3km3VXyoQmdaLlk1CAoeiELtKeeEeoHpBh
IXsZa6+H5Pa9vhMTJoIlgPi0rKa++CME/Ha+MwLHYVrUMJHydc2a3AS+wh73xc40
L0/10gv8Dl5TFj551rkomqNJhP/BrMG7tfdqMyMLpz/VSALNnmsh4bKH/aUlW4Y0
6f3RYyE10UvuNJQ/Q2qPB0QT2CUe0diQqAagIRJ3h946rzYJVEiGMHQ0YukQ6Bpv
yOzEvV7pbnCq9a9sll2CidoECb6wHYHMBY7nAoHj+Uf2rFG0t/TxjnuzxqlBOcov
2viEPMQHZPYpJxL8qpkns/lRUovIg3v1PQV0osBgANPixsEJ6HqZdJP9TczshQsm
YV8QARXniBHO0mzvEBJW/maPp8U+CNjLpc2AkTfqSFoI3QaE5UlbAjE+Hxdip7zh
xg3qbjLlVP0A85h5RSdQVVp+PjKzqRfebgVMTkHSKz06TICkcUyrk19UF9ZbYa46
7JIm+dq9WItcK8E03mwLTIJe0a00pPqO2VoW/uUCd4KccWzI7JB6TU07Y6mdVjOQ
fwtqPME/nOgwwJFrFkW4k5y3i2fAwiPY9tFlMIX3rW1zXxD5FiIh9jToUwmhEmuo
1QbZu0nmTlX2TIk3b6wMESDFnxMlL/t0tpWR73DqlAx9lwYHwz7vvGpS7NGC4ON2
QZf4TmLRQQPbb9nf0pVdwEijPY4T6Bk25fq4o4QFRRnXADVNE5md29RADiNQ8QdL
y8qb3DfjW49yHL6D5lexbVW35SkkMfpNW0v5rr5WfBbV/vTzQiqJILyOBI0g/OGN
dlxGLHum58m8/FcQ4YwSlB9oL6/FBlNL2FvZFmv1cpiO0Ef2OZNJGJ2WnyeEunrZ
tXgk3w/GogJhtJCaymuNYDpEbBU9+YrewYUcMLDOwg32SqBzt08N3y+0e/cWeaog
Z/Yw+pO2dpheOx7/2W0mRFO0tC5AcIBX0GdXCTJ1PBs39Wr4Jd8zxE1mUOeu+Xav
v30yGvHlL5roLF+VnJ4d6N1nYjnfJfwysWCgTl+/DkJZBJlA2y1tYNytHhQvgMe1
6M43CGnQrCDMhL2x2t/tDruYMG6YrtI437OaFe3ZeJHRnv3fhaH/S/8PfOR+KFMQ
YZHnBQDltoJQzRNsH0wXpFw7bsIl88VBI+CkmrpLm5a0yK0SpQ0vA+iMb8wanwfi
6+fA1EuJhJQL8M1a/xlSqz1UnbrTqCuzujnbwbuhWgBLatyHDZcD4vpEj1rqYLc+
aq4Hhv2ZZobd4pJ2r/vC+9pYmiykJXT952RXHoIlYNfDwY2za2Rxdjxmn9o2S3b0
V1ZoB4SK6b2CxEc60WIpJCJqel28gr49u3hNYpHyCgLKz9L/EbstzTZlAXKRvcQq
WWOzvxggXP/czvFETD00b7PlVt4e5iA9jlrjtba6jbwT3iopkQOmmBzKryIga8AT
/WRb5MjnfcQB42uuMiE4hz8UMi3fFpBPbHtSqQL/bHVd5QdWkn1DmAhQOfaTNyZO
+ASMhxowh3d/rqPl+OBHtN8owcEHyTsRoZKoP9I+lpgSNoy/oyEiNi0HX+KQdw/O
ybbbr2Slkcah0tei6T6OilqxMkSw97esymsHrjSibg7+Xs/e1qqoy0OWbH3CHm+M
VxjYF1o575gvaV+J/zC1410CZNXZrH86lKG26MQwfrrYLe1GyLHAUTH39J5dGeMj
9MnWqPzum+2p3XEpUG7fBSQZWyyGVSTAgTJl+v2PJuG255PeRUQ3UqbnwIKDq25X
z+GeiXaxsFb1OwStR3WoeBLSxfEhZ+pO6+Lrfv2qRVDjhhjQd8wpUXi7yPz7Y8pV
MNzBneykaJ+AGKbMCfQlZGUih0C5lV2yDGEO9uTMubvY2d8ulzHmAZiuuAZK7Pja
bbjpsH/nJs4Yzz4OgGKSul94CXSrkL/hGVeQDgcXpotDn12dFi2Fnpw+rq1g3S+v
oJ4vSe5I3iIYpiN3JaAizUhM88wxWvwd/IuoIVnGOlEhJG/TEQJqBqwRCMt2j+eD
dZjPV+e3JDug6PunulMzeB4wIpJkZJ1xZKL9Cr1zLwVywxeLLJcEhGlM0/y2YMrI
1LoOkQebqC8mngoYO9R85sKfdjA6875o0qBWRa7VjAm0l3iyldF2+/iA7EmuQFO8
QvC/KxEGG9caIDrKFXDe3TrHqDhKzFaaQJ4m7xMSrSsrmAUeikfPQPuHeISqvhgx
eZuj3ndbgzuycL4bGW1XCU1ceqEnlMPRUo4/zDtz3z1gOHcTH71YT9LcVrYUchcw
lbkziff6mV8kCmfbpxeWtNOI9bikvn1wcdvytzWmJxOASwSMp0Gn5EvSR3Z9otem
LQIvE0nWM4MmxM7kRgb6kSfDsoKWXYC661NnjVCkqETO8FA2slDU/RfwyOucJl1R
4XMSpvu8znU+lpuBBoeCuwVYyi6bgBEYvJqBrsHQgbMQy/3bUJ3UrYaY2ABCxRQ4
haDMJJus+1HvkUIST1NLT/yo2QQl/Mk/WhOR9GY19A1NO/JFb9UgcAEQv35FQPAR
ZUhPAtbLzgkdnoGm5dmT9MPIKgV83AZMVHhqkGqCkWhp+M3cPLsrUCZ6oeqRwZYI
Bnat3KRZYOr9Lry3nJpSC/tmM9A9U6S2w7SMNFRIkD3bGJLw7TNWFdnPRTKup4fy
k8ksKxR87vJCFqwj+4YyItl6q0YD6fumNp8ORF0MLBnpvTNW1wytF/Fodav7yxd0
HtPn+uzGcuU2Dh4OycN+z0VFZItaXOWmp7QLN3rLDjiGNkU49lTRx67EV7n6m6po
PR7TnJGfOyMqvHnPT+7crcPISSkHAb5ETHF7UI3Wu4Wl8EzjRMFtcSrb4WUy0eG7
6xd3mgEIzHIXJ2ZE+HifK0ci4m6OOftYmpHjv+EDdIPJsG9B+WuCCU2Sk7t9OSD3
ei5enDh45fPBUMiEXjTWt6mB/w8ffOXb4ffC4pry+0Om2S5rFCUVyNxTjMVbjnfK
JgQmTOmEp/53IV8/jN5m65SetiT38ws+CjDHTSq8tnO2Tz4XMJS6XzpexTJ4tb4r
HgkTrDldAVquZtvst+Sn4DDqc3kAw57MJ70ji7niqZ3qzbYf/atmf/YHXaSbDkFF
bXT5V9tfa47yeT/7MMqQq1MM5hLbPCcKPBc/1u728VqO3iqIcUfGFG97Fa47KGJ0
pu5nbWCeLBq/8XO2/qYqzgsCXpHm60jEUDZyaSAmgVtba51BDKm3GzB5V6MImPIC
46UlvgpaSdypwUKoRtZtDBE6FN/tAC6e/Bi8XxidDlHsKVPO/Jn0pDGrSvyqmpgE
xlNHBK9MF62NFNJsAgctvraazMDNJIUha0kvY1/VDmJvGjEZVE9+/cdOGvb43y7o
GOP33rP8oCh4wgaDZxan1AFPWS3fLlPFCLhMDlQAKHReUb+RF969HbKScssY4cKz
9eekK263rtSq3ngEaMIHh2t6sKac31Jfhwjf+2NgCFHPC7FFNAIceUD0xz4mrqj3
FPjYD0HNcaf05URxN6u9J6BtAKil+ZERIjdgZ03gHVvce5emzxLWtheHxraXt2jt
mg084dAUdjbePSuUT5+bFkJ9zMMtGLG340QP71Q77ASR7IZvkDpuIftWfL83NPwH
Tbo8QINQvRrvvTEuJu/ppiSoF623jAbkSJPImD/HmmOfic5ZkdcpsDvPYzySz64s
sW/5DMN83+fRh/DXjUTvYeYnn6I4cbz/FaufU/r+cQFuIoCbFj5gP5fOJgRYYFhB
nxrE6pNYgM9hjTVQpkAFhvca4M+nRP8xNnfii4q2fnuDZk4sMMyfsTQaXD3i3izk
DYoQOXU9/Dk22wgk4YAZO8uRfw24/YEz+iwhCui2il9pqnGBtytrGInRK5ML9DlL
CIjZjOU4zimdgSGYJNirakNRd6kfGxW6OfwFvTENHj0821Kfucb2vjIW53orzx6p
y9cI8H8rR4ctb2S1PjfgeiZ5U+OPjOBSCj92F7Tnvg2jwABr5PVdosb3dn73pGqU
iHO+YLdynTvUhnYzy0M6iwEfakYr5fGyqwMUTKkFeMzkJVR4uIb0DSafxhXjOL6g
IEzvb0oYb+pp54j89g4skR1dNxJVAgdtC5gTD5nxriBPx0EM17kZ2d9Jdt7A7HHH
xzVw0YGjXwBcqYRl0NrkjiYjWWIhAWebcTJCqjzLTtpxef11zS5ygCAcxZDou2FG
FqHdN0Dkl1X54qQh1BYUaVzmqW/ArAkTuC/fG5mG+9J7m4Kz+wChNqyGKfso/Pu5
eS1cnE8XyGW5NuEB9HFOFjMe4Fu8JqtJaVBKnFSgA93x+6Px0crjnYuvBcp2397V
FMkozwprghXZpGZ6o1r1c4Eq82+05i0+6IqHNWBQ47GJf7utir0Vx42qzdOExTTx
EPMyQqjWL0b7xpt9I86QqgVB8xd2dmEVQ1jQme0GHotaM3zEFrgJC9OK1R0nBl9e
v7uIxA2cds9WoXjL2tGDSm48al+hJ95DEpHG0VDOwd+kVqYlduFJHn56EmeYFcZE
rCAtkVvp5gnJUZEKvQfEQS1H2GQkRgDAlr7Gyw5ShrcDB/JXGz+d2UsDb8vWsb6A
CEa5634CgBdjaRWWoONnHeqWEuJ1/GZy1mLt1QC2pb5PhyP4oCwQ/IwftcMnrGu/
RDVVQJwDwmfGf27Ya8eZmTbtcPEyiGKYzAR/O3JbkEo29GMWRszmMNZNqZKHMpZ+
FEgcSlDYIi07K/UAUnC+XeP717vKl5HMxsTTv5iNfrnZVUjlJVLYiSdtc2iU6dAD
Kf8bsrkBFb8Xje757CBvGksjDCuUkaQpWOGO+IXkwqMS/CY7JaScf3K3ijJ7zZ9V
wLbr3efsKHO8D4R3ZsGASpwiTt8N45xz8ZP8dhj6WAqOhQhR4cVRweBOg1cXK/r9
t4pGciaY+mNdDtz+iyZGq5M/zLNnQZKYnP7XvlKACtMcWKImkP0Kh22cnjLEvOyy
+XqK6Yv7jFqcjAPUqKBJrlg5hrDDdk1SrdJ/bRkKdwiRqeD7hTMdX9fqrwJJxhSG
9HhwdFH/KAYnlbRr71CHEy6kQgqOtrMADFvecgQyyqNWGd38vvi6a4F6TmJdc5OP
sJWKBBZCsPDxLGV3LG+FBckbVGMnFuKJquo6IT0HQHBh0EkRHyFC1/c0gKFhCz5s
umnaxgmfiY90+k+Pl0z5omyv0Zfodk3UqQx5tBpz82ZTLPCTyN6AaI8Jq1Fne0GU
qSl5PfdZarlt2oUtch3UsTCSEwrZnUjqlhacHbi2PJekeuwnO26RzA61iQRxVNfh
0YdEtjM4Tba5PwdIP0IJQmx9IICmELlhZezQHb9ycMKchFdMDmBjdHXDCEd4gqEl
pLPHi/9nqMF445WmTeuQQSRlDWxp8Sb2KzqBKnsAzGvbBAtpD2Io3wT6ntTzvDzX
6CDXPxTbXVDykQt9eIPYvJhHssb33R8D5rJfURKeLyP4WiDEhlDXfsY48vmo7gMh
bCLzPi+0dVwc42ljjFywE+lUAhOgMXtUYM12I35bdld0VDeOMSKvr4ld1+1Bta3d
NLiT+gCJdjGCcosqf9iTjQXeMSE5THtQbH6yb6qsaEueeti1++KGx3+bNjs8VGaS
xC33v8vMVzOOjmrBFCUfZF+3P83Pzs6xBddS+W4FfP6/Wogg7xqM6B2hYflZ99v9
Y+J5t3s7UHawzH3uZu4GNcuqRlIObB/AukMiwFTyS00Ugu4nv6Fhi2KS6IFb4ALm
C700gFdRdFRMjEi4c6nLL+mUPpi9RPFxSDarIjY3eyfcytL+rsqeWKEXXELHCPJs
bDpjMHZyLZMc55bmaa8T7zUZNKY869CZXAftFlbk5BPoOzDIW2cELYniYvyy8HQM
ubc9o2F2K0wkd0o9bR7oHMmmBDoRyomc313bihZ7g321OZkYbLcl8Snhh8iV4TgA
CajjwR+Bdqopx/SUpcZ32TwKHBMNPL2Bajva91RfBT5Oj6fIOb4IQmltBNxuanKv
tObjN9Zz8XKqTliJ/5MvYWJTucE03yg/rDq0tvM4k4kgirzBKqZ3wRAsEdwyNtyV
seCS70r0mn7f8AXNNK3ASUsm/zyJ8xp0sJiLh53t4nfCK9XiCl1lvudoSJMgWNWv
HQ7zMa/TaS9gHQkmCohPFO+kkp0x+lFiRboMZxj6m5cRW2/dKh+ouEC12H6d65v1
35KjbA8pqseSGfbirV+q00yDZKJjpdAcxC9VPmh8WxES+5J1BuwtQcZAsk/2SDNn
RoXEYYVqr/rg3sUgu7TGDJhY0xhCKkxNKjod3XDFLBGP7ndux3h0GzqkaWRhenIR
UEZxwSj/ibRKL/bJl+Ol3BErA54rRZUHsqFGfOGpjpx8AHdsOu9sxm1EmfrF66RU
L3xL1LrD6gz1ZWQXoZtgPjAPoYZlwZdsPhtsJkTzMpQf+LLw4ifCj+tYJgeClC57
YK6V48qEMiB3PgJ0nyntOxD0ddA5i1p8g0lyEJYWd9o+hIuj779yKQz5uZRnaBu7
X3pdD2m7AH7jyf9aDEpERXASyD1APbRk8wSBXh5E+fjT0+mgADxgeXFNr9n8xgfN
LYwEGsm5yOYfSCp3GO6buDZRhCl6HUJTg5zXxbZko4+GIIpE6NPC/F26TfP4TgK9
YFaLdejDEgR4a0AePklN/StD9t/TEcXq4ap4XoaUAun1j6xL2No4tEJ/o3KAaS8X
jWuoD7i9/9gp9nPSu8loLYjFb777UgYnT0iFwUWts84BGGd9axVZO9UMYBHpTD84
0Tkk7JkA9Ib2mUauDaT3Ck8YT3rcMLS879LNBc4Jty06658GlZfEeEmn2kx2DxXC
GClrDJ3oB6MlUZ/Gj+iYsm6TzUbZoBVByIiXFr2nwSe7N/9esumK97gni+X9osa8
SfOdlA7SpmuuHfaHfYuPm12l/Fy8/2XLaYUK4lBkO2llAH0l8LVYZmvSlZMbaPO4
eUf3Qddpa67ROX085T4AW2Et2JdexED637Z1oV3Dz81KTal/lN4vtl/1DQDisUcq
JA2H32wXM7zTuuN4dRIdYVq7LEoeEj0ZaGBxoqd0+D1xNlVzttA8TqKQNEOp4V8o
evastDaqBMDJmWdKouOhIs5z+qu89TBo46Cj2R725X0C8OliAXBQyVtMrocngTC8
u0IeETCFn40bU5Jz2M19Q8gvzmPBlxfbFqbrX+wIVr7DrxowAiOK44YiQfZ1YwLT
QafxjWs7dZsXx763NvD3MPHuwS+L1OzI9uY8NtuTRB3qTdrV22d0ofeMEFlEAI+q
JNp80HcORgF+WPNq7yZjlfgdsEc2jVKIVbivZDcb4YRo1cNdqOeTjKGjcA9junSz
G3KI6+sV7Iq/m38Ul/1O2zGtTJWP3OQIYzRazwqLMxSbzTxMvqNSEvehJkHg5C6m
JKWD3ZXBLaG78h0ZlHKGv3Y7suBzR5H6RjC8jLT3cYDo58BaC2IgQkT0WeqI7JiE
IQ5a6iM/w9PxTKYQrya5mlsE2gtKlVUFNiwLFTikTihVJTD/yfN5ovyi1isFUY6Y
FgBZlbjgUgL/738MU5Ze3dVHGOgBA/RcZ8u1yeUILZ6UKifRMk9EUgHy7zeFVncd
DJzIUFew10KphmmIL0QM2JpFlKTAuuphf3C35lzcO/8MCozwVfRRJ+mJtpUzYq6Y
vVtEx5YjooJ+w4o8A4rIYPLwWytzPS8caYxYY0I7vPEqkxvGOD9U2jtHshdyQO3s
XnIgu6oJy6WvMNNo7oGsw6NiK2/WKsVXbi9ORhVNcuZiVXKfraYOSEi/Z+IlnCCX
uPemLKkZ5PYA1/hs2HvB75aPcz7pFsC60G3SDijbCmeLlyeufohBRxfZ/eSEytWn
FgXg540HKF8NWwlytfa3kSJMa/fDEXtQkLWSrJvfg6Ql/noeSyEvRQ+kw9stBHLC
uMgjTKO6lruaT/8MwlfLYcMCZIE4AbI2kyAHKrwQllr/DnzBjsfum5vcsh9Zf4oe
mvqgtvqtGTXyeG7yI/y6ZqAspawCsuAbWtQT6DgmlSe12KCPTIXEb0Uic/cDKV2q
tNRME0TDzRMoE/l5DemyQkXG+F/zhJ/W+YVjZ9qt5hau0fhYpRCh+p0amzu0kHnL
2+JMVxlRn3oL0ByDO8AA1JFijpAJFRm6eAF2AMvir0hyD325Y47rkLOb73VZ1Ogs
qpV3IwpOlOQ+j409zZd3JFes8ZoFN2cdr98h4amu9XC4m40BTPwJAVFI9YGo7WhJ
Kn7fuvuJoOmCegJ/3Wnys6FR5mQmytFk8L5GoDlT0rUb+RUmbrpdLYGyZ6YTKMRe
zh73M06lgwN1OZ3YflZQSzNL/6/hS8cmO0AxgukAn4v8TsJNh+VBmIwg8rwJ7Iiy
exk90+zQBojTLSZJL/U9lOiSijgm34dhQhq/aRVceeiSaZ4dltdtprfT+N7yjk0W
xIkiUT77u9BwFhHe9i7M0zQBYB1qCNK6ayAA99QeybMXH0xhSvUraJk91P+yIkih
wf0rWSeqoVIoIO+A67urUXp6F8WV8+htsgULNTwy0+Czv+IqrLbi+g2B79AN2iXw
Hvlc3QDjU+Nq7jsuPAKgS0jnNiW+Bsa0e6HQSSWVGp/9U+7HFo42VfFWejqgOnHV
a+MoqZ6kqVv2wd5Nl3ixUPvmwW0ffw9smrecYeZ/9xoWox1ce08r8Y9krYzYo48p
UQjglVfju/Uncnz2KqY9MNI4Mj9ctsKc4srwAdaZDa5L3yNE2bWpqgciVh3flGtL
gyDUJ+UqtkBge44qAwUizYtwj7lH7aNUT3aNOytBy1Dh3JWOQPIul2qnkBNLEZZC
RQf6Sud25PjjcWU0fBKbLQeDWfCdI5/StIEyx0HX5G6nI0AtwHL6GBCgyPE/Em8L
VHI3Oim3GyhhqM/ju7q+GGkmV9Kqf+f7P93bYvKK+sUS+qD2Aw9Lp6nZjv2/XzOV
+5bPl3etPeSd5CX6s+F3SXutkBAaTCm9wWVJg86wv/PQCrNDhpF2LowFIU/9RAjA
03QUSXylf8R5PGxoKAaC1rstBv4uftFDpPRZm11nQXlC+K1qu8CEHUfersqS876R
IJ1WH3Zy0JJqLwwmei3Nyiyq9BC169Tx/DSW0mZG1UoMOzqXtT7hq+zRaJWNfhM/
5K2VzXqIwu2doZhVZ6DgGk2KniB14dkV6qmVzTYhSCnEPMqhq9aajYe6Jt22twqZ
T/m6wPSfO19YbO4mHlYxOlY6bhzt1A1mRxSB4Zd1MlVwnUFr/mW57Ksu4rNkp+3r
ceUGKmAuHHdat5IXCKPsWaeyYpr65asH8iXuX+tIALTBXqW2WBkdx08wDazvmEVP
VPtqve+dEPpPFlYycyC+c+sUR22JLp80tZTjlQsuqq7KN34zYgxAhydE8e6NvUST
q4wzoGZXY5qyCO7FCeiAImwpI1GVQSch3YPaPHTEC7Y0A7qAZquKepJApwgHu60w
23fq0HEX/Hh3Slzvvd4Cm1sreY7lmtZ0Vou7R7hYA2NiejPOCeYlys5KkdrPggnl
e47amKymjHUVG7USAS8RQNXJIpOZNwoA8+EPlrsKhmhpnvNFcbx6Xx2jqQUCpfub
vVguwq85dZLmJSqLd2Ea8mEDBehHDknlWXnUTlrCNVtk0iqY/Ij+KYmsM6hw9Z0a
AsIsW5xzDTzTvdiIxxFR5DQV6Vs8N4olcZBlM6m2kRAo4FgRFEk9IB8vYx0dSw7B
5bGmn6G5Ypme97elhEB9F/oXPplK9h7uBi3qTJdKpBA+KqmNPSvjcFNDMgPyxDIo
Mr2En5Bpm9igjGlC/haoJlRf4D9jdhcBjjwzo1lrvtxkbcUug+HV7g4IVr9/UCar
dzVwBohJo3cPUVrFGgxg30R0A+spPZkmOjE/6Z9exx5dBZqAt17qAXEfY3Xjo9jA
SltmLrHJmDnrU5YYfXszSE7Mh3mlYqubSPSMuQ8ljurCIc+nMO3/9wMYXPHQNROr
j6lBCcsDDy2fjiXes0i3noGqiDc51+5Z1O2XAIH8uDYs2mLOdsMFBZ8rxbnoLSaz
XPnDk4CAOaIEhT44BRdeV3pm8x7p3+PfK6TEVa/8cO/aPwfDLaj9ek8nkVGxWDNs
Qv8D1sGg0PiVDLd0ZqabiLi+5Xkmct+1gj+J6nA9cLMd7iW9fV0nm6R4gPNo40/H
M1QKsSEvtQ3PKUVovqOkOX4GrajdQKnQkPkcrpsboP6BPO5YcFBEut9LXxKGUiZC
7vY/RHKN71S9CqgtzK93Cc491ZagbNhMxNJ30qKfN3ejXgp6+XJrprNdqTgN/dsX
MesUaNrRLh6Tvp38adt/M9D7w/wfqy6cc3QaHtdIexBQQr9nFZOC2RofCYYoQNWx
x410NFQaLxpZi51WGLs6Azt/1UQSGPdE2FrKQ4eTbX9VouMVmLRgefcDRTjksw2o
sVCgc/RgvsYDm6RR7G/4ovCTUnWIWtUBJhjzTZ7RFkjcrs2pG5TXsSghDdru7B8/
5K6JFfl840HNdfSNgpapjkOgmNklHp5XjumZrOISj6zTGVyJODeiTmv3v4nGy4kC
ct8jmssyfjYo/5hUDxgumPqYSHse7IAtS6b8Deop7w275XlRYAyA4ZObV9KlPoWo
1+Ow8HYCsF5wOtw4IWebNCuLHGCpotmWQcmCHLSFMY4OSAIR+3NupPygwftxETp7
7pKim+pBADzsDxUk9apmZpEIibUzhg8bY90iqdBQxDOeSEQfDIIJAcUOCGwsRN4b
oVFDnS6pmOa+5/y0lrEojJ/KUiU3dYAGNLzC8A7e50pZZEQ9ZZ2TqWPiSwG184I2
E+JHBFCOKhPtX07mJDT0Q0meL9AFgyIr5pZbpEK/8NYVsKzKzvFK2qgZ++tDsRMd
C5Nw0ZIklDzj8XDSiN//SjMUxn+QeEtVU/MlPr8+wbbRICSeMNO1JU5XUZcmpbMM
uKUJI0jwTYy48cba/cMeEEzOjrtRn/H70H5vMD0YPGtivHWkNE4DWLgCHZ8tlnKK
GBiQxMsJpXziPL8kFqrRPfgvv0bbN4toObl0gbfhY2TJjWH3sSWHN66sJaHQMJ/x
NMJvxVXqn1k8aAxiR1km8pd2hkmIYYVaN6HZ693gk9WJFZ0pfm+boK4McfMrHBRi
J3CBgP4WA1Jk33iofMhliMNpbf6DRdCjuybNH/G9PdYv1wkeHoPtN3M6nr7grlXO
94o9sPMFSs2f58yQMUKeW5J8H8Yau7zAj7VrRw0Q6IC+oF2u1ekKRKSvHchrdc5o
OB84cApVqxGteCb0/mR/D5Q2DGU4s53k7Me08a16w+CObEuDLz5GwGmTIdiyHD7X
fdlZOuVS7l5p1a4PeLgLWd170wlR4gV4lamW+qO2ygWfSaV9axpoQkzN/RemF98h
ucbLACpL1l8WnIdKepCDOZfNwRxvPPUz9s49gLtT5nZBKbd/5/j1Y6CH2rkKeuK/
ErDnIEWV4UyIf2sYxT1aaTFCQs/uvw0eYlxrNkhZc0HQ2+bMOqJp9pAuRa8xHK7h
kDqAUTXN6M+sBNUsvRqM3TYJAEM7zHqWGdnIZdiwLzh8yXj3TWVT3mypIs2jAQT7
IrOEeb/fDC/PeK8zOZsoGB/+I4PtIpGspaWxvoC+0jRsR6qjwGn6oGnKhyKGkyWZ
cLUtKuK2cFE4btUl8TXJD7/8Hsi41u4oQmGqIk5M3HW2SdyyMBDvWW/+xsR5qFZG
nxbJbitHhkCL7wTjLtU33jJOtwL1sSfks/VB62c4hSx+ryspy4SiEyMuhHJ1NSRI
EEkZIuSRP4mSEdR4Z1Mra120HOnCvul7L5A6j+nBjzQ7WPP3T8MMjGCWnEl5cA6V
W+6vkOR0a0LxvCuG8ngJ7JRV5taLyMqBcY+R47nRAi/IFvlF3yG2sWroQ46mFqU0
ExM2bmBQyEXTXjMh7BqE9ayzenxLEnrzn2kdfit4YJD3G/90cD9ZdtX5ZDW2vSFG
EerTtbk7gThDcJz83bmJumd85TWTlZC5lLyHrJGC+cjHCNEmjhzmdkjejQb5du/f
lrHzv2DLhJ68qc/x2iRZArLOHg9I9habkcWrV7+EASFN0nQ5i1+cuZ5yiaM+7F4E
VSlxP1BK5n+6oJPqiGri+ncUxxKJjiv7I51gDB5ZQkQGpsZMsxP5kd9ct8PW8ELg
EPCTbAi1z3d0N74xR624I71V7jxve26GgzBtZ1hSP0Mk2KOk7o3mfFwqrf9Gerxz
iqtB8jmaKSdaxo27MKgmalk5scsuRIaclw5YBpdYiU4Fxm6tbjVT79OKPdwRQLSE
P7TeHKTmkEpp3ZNLp5x5Rg/JDFWP/IIG65GxPgtzic7nUOoitrJpaIxZ1LN8WKlR
XgN9Tc/lUD/MqLvdzpVXnxuE1MjygOb5Q6YiFTHd+dvo6TZ1GUZB3cITmtxXHIr3
Vh3/nK0EH9FCpSs/dg0CmOWKqiTZ7ip1p458UfWE8UPzpX/UaTGyTODNbty44IMM
/IqjyLMhtI6W52k05vxf3kFHvy74wfFwA5kETfRQMUj6vgkZtODJQRT7I0ucphhi
kSzOH9N+0H0rLydHaHUBY1di82wUD/gua2v79hZMjnKLwrSnrnjOhY4tmO3DkhGx
TPdTa0BROck2zrVqN7w5pdjWM5k1KN86Gzpx6AVw02t/QVp0ik7n3pDPis3/RYqV
lkoLAtN3x8I+phNGOyGgon2bmmNJoQFkIS8lBslzijPwyTc7b14VCVAGoMV0ZeGf
exzOZ+AU9I+SNSgZwXcPX4N7M5nj67MQCcQmp0qzKRF84GSsCqHOEt9DZJloc4R3
xcGj3NdOKr+HeHqfdP7f4A02yVMU3O+G4zRri/waBjxAgg6W2gK3GZ0Naq9UiKAh
iXSYKHqHUg6r3Y7GfmDyKUSNtkym1KaKDaR+snK26R2NTu5SjGvy61Sc/1GY1r/A
SdMzhVSEJqaiALKO8UNyWTph6n+y6fMqZmW3fcr2dUrsboKg99+KHpkAiklclPLj
kVEcFH4ve8c3ldnQiTGxXCkFOI4zvwGYObUYua1Znhsl/O5SN0tmhCcMzzV9aUad
b/vBLbdWfhnh6L20YyBJmvdu0lHCCjpmiLolKHrfFHpyCKqM0dUAsP27kYmXrwbN
XZ/EDs4UqetrxsoiprzdbSkwjcPauFuftTujalaImEke5UVWFZBCYaU47Dq1SmIf
Cc3uZ/uQMs+zhjRK6jig0POjP95DG12oo0YQvgjLeBjWE1+GbU762OWSTyhzlxCq
sw0oKCo/TR4ABJZ9S1ua7BT43TN/v0IGGEubeXziQ8PYUZJ7Y5yr5V9LJFtIalwZ
oXawQmYAAt07dRSzSOquXCJ4HSWdGVkLeLEBJbvTjcrqsNLI/mI6mlyqb4eAOctp
km2GTQNDdNyLtaCWbHQi6061+nu50CL2EQFAem7qM6+C/Dj3Pjytvm7/vkOg7Y4W
NRejXklU7INfxHzjNhvFmfQFFisDZTdJFe2t1h3DbARuV0Om7icN9Isn+us3KUzi
I61HsGXMumHWQBYq6NUn1o5PT8VRtnTo2+rK1EXCkgVd6JMvC60vqZw6SbkDWtCH
U0N6V9N2kHBy5YFUG1A2gIcJVHbYzc2KrBmhOhyyJn/SKmvw+A2jd3TCoTOPRL1Z
jqIxiavzJ0Gt7pUNRll8UNYFMw1onaU/NIvD7IEe3LgdfbEIO3rn1eFAX6GDEe90
GeGm2oIKM2ljG8SoqucH6OmbLcSR36rxkFHPq+zWS7TebcoQ1+J+7K45VlfuyFgk
1H4n0KPFhUgobcSyKpnMj3Zmj3VjF+KYkkH+2M62qH7BSUkPMQMpJC4PP8aHjSAZ
LDfI2Ic40SUk2ehULfKB0Jt9/Nh3KVXiVN8S8IcOGyiM35pAD3RtLE2RKTAfXuvi
guLcrkConQ7Mv8xg7NTlc/ODD+a+om+N1R9Az4J8r/+3sDrehcQdSSeXhmIBWFOm
6zFrJqBZQ7xdyrbSeTChZ772XD56OraLY/q8fUBCmOvrDfNeOEg+DB2bWxycV4nL
7oLsTCqLywe1kyNYEKB3YqYNxPannmiF1U3Qx3cTZjxfHrbSQlJG1XszrRR+YRTa
8H/MUmyTfUO16+3Y5hEaZU+0JKXjp7jQcu8S3EvyDZiw2CRvS2JdZcgUd+YvWRtg
QU4iNViPlVn5UUoz/zWECNmZ2hsVszkSQq3aEa4D5NgZhLbjTTLB0QVwAAy4ke6j
KnfMPSQ1XuPxEdSbZ1JPs9UHdju4OHBClwUDIbOlJ9UKElAj6llY8uJjN1oxI2rU
fBx+ZSibPAgdB4wKl/KFo6/NN8VznaZIGKzM/3LVok249G65NWx1YCHC+sYBnBIu
RPr4+8IQHrI4OMuOH1rvxeLCPQwjR64eBDXkf0/YrdcL1IrMYnXh0V14fTKj+POE
HokNC7pStMNhOShEkzmOaYzp1EX98WKSpQDSknrowoIrLX9eRoxwPiemVCzch2oQ
+gOh6h73xf1pVGAfAhHeQgHP9hwvs6JtDlKN+5E5cdvXpnQgaxC5GSAUUHjSXg4P
8Kvbi08wuy0o3yeFT4yFfWSgt2nHjg5NASZvQlRtfnunJqdETadhKoAU1JM1HeEN
1oWxQ2Y/zrF5MvxP7oVieUzMqkKMKYMY57rTEG+PCpmeMyVRhhox410v46LOgYGE
fyLjvuHYo6VKVckJllD/c0xoetq080HW7OktB2esSWuDUq4746Gig5JOK3yyRykk
B+jb6C5vkmvcqIAwauOJW1C3jRY1qxUT1NBmJiLDFsE/K5XUJHeK8l8ruJHHFSGu
DU/KIqCEGjVeA1vYgIxZlO/pL+wtOa0R3tJR8t7ub20sqH2fWk7Fmbz6l9jjWpab
s2TC8lsYMRyalR3kkAaeXpHJ5yKtb9ojSizZJsXsp6sZiiQlmqAtdeET6FvUeYHI
CuBDwaoJtN+a/R6wMfA5dWDZ5wWlTMoOAeVe+Ec0Aopo+lSw9HFeCYFinsEOctnx
4YR0xPrGYPdrmLLHq5l4W4EPT4BuERuFfdMV1NpRrcISXBM7XNbX59meWy/btEjW
PDkjt7+Yt+S6iQfRvcfGkQGaoMnoWbCGVkLHSc8mHHr/wVXp6pmcrCDZoLJnun1k
3YAcAUunGkgO5bs1/asc1X3eL+8J2/gwFuFwP9Y+ohxabVNwDBkyG+Wjy+JMDiTK
Jc8KC8I7AM5bapxwRB0PZ945vL9rsSsnJ8S8geiEDC2sN3HWc6e0C3CATGop+Kqd
HQUxaQRcxgvA/oNZB7I2J2S9DVHQuE6u3lxMOT5YiN9q2FL2l71/NOMY3rZZ4Onx
OlVSeXAho9Fwo/erj8pZ0pRkZ8NQPjvr84HunbxhJvS6Ss274zQPn3EKbY0rhyfq
qedICL6tYnU7um7QVfM+zErn6v8WKliW2wEWJp5S8sqAqFt3T/Rk/U6kzFNijMqL
B++4Gkunmo63QgfpLaOXt5q8gCWhQEnfHikkKnwrq3vvGG+MOdVECzjV1MfsnSx/
4bUCQeT5zAbkxg8eUHRzxMczS6J9opBmTt3WzgcqZprl9dlUrY7mhgRAIF5N77Lh
lL63Vf+EDkkRIEIVazIeoZSWp8hiRj6R3cmJd7MQc1fxgTs4AjNZwJcR2a+aJ98f
raFBtBk8IOHJwsYAFrSVrDtoewEn6d52Svs9I53x4GsxM8wWWlRSAQ2L3vpUtaLa
baEsNRVO17CdnKn/8STtaeT6JYNfQij5YDkmnYUnY0BciKnJTQHrutqs2cm15ovZ
ocrVyfte4EnPRDpe2MBKMs+sakN6tca8VzJ9tRTa0U/tziyt1/q1ZRUiycn+1vJx
qwzZls/sUuW6LJ95VZjnGAawXRmLmIWf8B9UqnwaiHlMmPxA+rLiiB2C83YudVtb
7mn1eLQpEeC1TuA7er6zGHNQejNSSdFcZ8HSbb817l0giVEHSktCvwIgLHiTZ+da
A+Ny2ZIfGfPQvkiJwEEywtuOT7dfEz+1EA5VWDTRXKYGnovDCCFPEVtmXiMe8ehu
X8jsD9SwN1CPZs3xVjqNbgilGUTdHI8+a7mRJ6ND0hJ6KN2xTwDs9BRmmRW+idq/
+gNNo98O1RfzNWCjOAsW9mz3VYrJmkAVNuyMVc1f1TGrhhWJo6XymL36ipZMm7KM
Jp6GStXoA2AnG5IETP5CctRvH4+s1ztPr0jeL7oBl0r45njnLrCYgurHFg2vxlB4
ycbtpntZslGDnFZzbMGX1O5iToSbqgbbU0PbW82rXtCDSMSP/ddD9KqskK89+rEe
43CRLPtBTFNyy6du4qiGrA3qgeY4BkYe9ouCtFlPmDbjlU8/IZ5xCDl3BdSnRmGP
9sN8/f8eMPjxjhbO3dhW/psxcyl663v/cXC7CveOlXNM+3iqtrORBBEzkV63kxsL
A80j0fSoK/iQeZd6kPRC5SU2FlFlmeHPdF/0++wOqs+jQjmv+WwQbz11OfXbEiTm
e/Lm4ztbIGoRM3T0D4fU6LK/wWJzwDf4mWsIXbrCZ033eiv3VKcDBdSqQMRy1utu
WQ/EU3XOCAHBSNu8n77Xg7zjOaOyNoCvC/KbvMMrSXuBpZKF7BSMiCe3L8sgZnM/
yHQKnFy/4I3N2kbqOA03IUNGpinCw+0HBVf5N3wlUSMfE7XpJ3BSGMNy6Kkpu2P/
jr2GpEISni1iqFsSIMPzOLSFFRkqRVdBmJD1fpVWvoMDy4GugmICafxReTDA/PvR
9Bp9dOBpW+GEg/HHdb+kVPjoe1ooeyGEBcUdRxwgSqq1RoqQc5Fcv2Pq0LQHLn71
vcRxRa65cedrxy84TCMqW2dZ2rOfrNtispMFKsHJiY4DrK5QVRrSedBMxwTTXUjG
KJZotW+6FlyywTI8HIWuBWReh70k7gUgmYwDWIjl4LqKyKF/hSIYP73rrYTKBPOu
LBbs8/xf4GrdxC+vsoCi4IcaIssBPPC6BhxWwPVD3TqYn7/L5jQmMPTam1N1hz1a
pKlzCpM0mbOuTWMI96MYLQiq3RMMm+SCpJjt9tembFNNSMl8ZAnPswiPhBpbC693
0vSJbFRSIiNaLjKE44EqGAYGDKxFZDBb2gQQ/ZUxFp9a7W+kXntJeabNqqSOFwad
XqLEKcx/zEzs/q38E+IC2dCmD4Mj9dlrXAaG2IUg8vZMd0zsgjNQaoLz9vKaENXc
RKoVoGQrCjg0b4XRRz/t11uARJ9WU8vug+lNr3lAN2xKfrYBKkww92kQ1KnmuIUK
aNOURSxDtLUSPWaXWv9y4hgOEoK01RygWq5N3ziIJWFLvgmR3aELGSE2NDH744vh
10V0hs07D/tK1yLCNSxC9yGSnRnNli21yjzcU/JJleZhfpSEjWM288KD6fhJRV3B
CYsH53zkpizgYZ/cEdyF89dweCPCuEIV2miw0VWVQ+oTZU9iGCHkQPTf+OhG2MQv
1pu3NgbsvvBA/4vsR2Ay4eBfB58OiGq016oTls6bLDWoZvPMFtQAb/TkajGCmFLk
n2cFzaJWFVUO4CwAcDiDw9OhRNOuFJLEBk2k+BWAnvgzlysKBWeBZAIaTAzx2iEJ
NQ/YsSS8Z7JWiquSrIdAL23biGgAf4Tym7MvQtqWIHNvG+n0st1YiBN6wSyYPKj4
TDEnNswfHippJj2ae8+kID3zy+SKce2KIj1VafsHvLEEmCRzQ+kNFo1eSO+IBEyo
Hs5YuF9KpNYqI+1WJrRlTxLyPCQjdKfivIPjwERgSBQ2lYWlwlZ1CmobcqDII+gS
co+9WGSn9N3VClHgrkvMaAdT2J4RHHvsTEN0xhmkjmC/6Py7MEbJdgQ+juBiroM7
pMg9hgvQdQiiJJX5fPzyg5IP2yoTJhtLo6pyxcZ9p7cjVDqcQGoBwoFSVxL/3iFJ
TGjePXfDMO50QvG5lsG8SUHr+G1va7zhp3FyRDk1IIZ2JRLKuy2t+9teo+yAGbEo
k9qGLst7fPKj5wpIHQjVx926mZqE4p9ol74nmZlT7KCgVALWXaXiAbswXynmOfi5
6GFz+HVdccsbWKu+NhvFn7/zK2TW9EGOhMftSlDAb555c/pyB0JQZ8+n3Nkizzy/
agVu1bwUL8CrCjdVfeBR/WqAS6iV/CO4f5yj1xR08A64leaSpc2vyzqopGOliuR7
w4vQM752hJRFgYV8gC1xn14B0j+SCLH749lY+icOydG901w5TveOrbnNYWduhILL
xzRBEEp8dBhqxUpeFR1vSl74KHhEdmYydp5l12OLIx2+lGEe52LQMfgmh1hN0wbt
TLlLo/b7Ioooq5XeJfIxLT26S5d8eU2hbX3yvx+ufopbhBd8jucGO+qx+5iR/cKO
KHgFVqZVy094AmWepzy7ehz/cBFDtv06zFJ4LP+VVavpvmcqcP3dA4RFF2Gs/fti
HeGUhe7iQ7g7X+6+7xEi27CYsUglU1YwymC9G74esVZ7ethN0v7X3nVRFmruIPvw
5rB8u7bYCrc68uzwO4SFtRn8LcKQjY25e0P1k7PK664MRUL3Ko4t7rYXpOaEoSgQ
WyFAWB+mFv3qh6Uk1hlMuxEQ4RTWhTtYlcf987wbUAjLfViTU3YoVrtmUzoZ7/hG
az/y5y5AvaXT9Nt95YuARtTM9+7PnhUM9x1DQuf9is1ZHqmA+zYA6xEUbbyulOZv
GtqrHgEi/0Espy5E2YA4Y+sv/BM7/ywdu4KNG5F8CLq3UIBVW3UUBYsF1Bv8WA8b
boytyOt9UcOB7/XZw0RLkDjZZU9xy2C04p1QsynuSaGJeXPxAiNE57Y6PVkSmfAt
FKNUOseju7g+CdLTbHDgCNLlZowsw8l6peQEe2aQkxgkOxn/1EvIW3xxvSQDXlmF
W2G65cfbCR7Skaym9OwsidWyCet/BvqPzDOUgZwFcYiICZ5J6hmKlquDL6MGdr/N
ONerEUf3C3iJ8+MpxCjBSidZOOIy1vNgKaQ1D7+lNPLc1nfo8yMxuQ3go2e8NyQw
7LwBv3qzx43ZvjDAKuXc8pU6BMjIaeo+GzcoE5BWxSJYUaRgKz3sRjHP151WpBZ9
N++d1ecigI6ROTQzMm7+Vop6zDqbihFs/oMrTbqbX4UTYnR+UQiEozh0kg5oJRIm
PHj4kVtyqgzQRwrDIM3/nePA+ks0epY0tZ6lOMduajPirmFUdbDOsbYnbV6E4DIu
ZKmjrfNL2r+52WdT/f0BMVLFoqFzunma6cLV95pYj4KqPI+XS9Gly1oaYz++qZOV
yLmSQK0GjlnOTH/PbuuLyiDDw+PXx8gBdKVXobiB3t1uCGSIZvtju10yzlA+5/8h
YtqM2lTXQwRTx1lY7hK8uC7IbUx4Jmao5CVMEYZf40/FvQLBDnDodXsBxL38cMwU
IYdqxDEBtLOKnOU1GbHaVdM3jRVIZEr/c18yFhUU6eGByFhy9jwVPz6pCwrdXvmn
Ksfp+ym+3VF94UiY8YHS4LtjLf4vCsTIJTbFCcIC27vNIM3LImnRGP5EVz+l12kE
RrTruetZOTEVVrTQNaYESHCe7JsdrsJa/Jl1gkoQtDh6D18QNDZqUYqWLSAluKnM
PzeAHIZCOwPC0idC6DeLajjIgpOOsazY9rKIm3rN5T4CpY6JqXWR2dRZKrUFZ43o
m5EJZvgqBYL4QN5oKEOsGWDTlyGKNr5OCwN/lhmnhYCK6Fl2PyKS1E78FI2FN5IH
qdV7Q1JQ6EhmJ7jC+7W2w8xq4SBqUSYqndLN/O02+QPYJ31wz2LulzBL3f7B/UDI
cLJ00h8V6DyPpVlYUenfg12+UfEOEoAOwob+smnarJW1jx5TCslz/S+n5I5yFzQY
rEktCk/g3gxnMtoLjPqLV+uwn/m2ytbMPi4EKfs9HScZO3OpNo/+AMSxDJtOEO5i
xNyY8Cp1UG5qjBm5U7hajFbec2Xmv4Jls9kCM9SXznyK7t+mJQ3Vmi9MsnbBWjNA
t0GrFWCOQos3uCd45/sumPqxX4T2TSJmO6eRlrbd7EF3ptF4eEaHVXp4pxrHurxm
T3ZVJ3RhBsyKJNYG9j6yscJ8ljktBPjnYvrkI8lA2KcH+2MDwMRaApF3vw/FLnS3
jeAJVlfgbdpjCrMhiOIpCR3wWUC7H8tCb/XOOU3bn6Mgz/wySzA3w4Lvde6uQ/kC
BsVIxGvMtwvwB7AXZIMRHhpKEUt0GbPR7Y4/XwQNL9Uzqdsy6Y/dcEFiywCearuH
1STFpJD9gSAFrUXVdYoxaQfD/EcxxZ4wW0RU2Qme1DqvK2tMZAIPk6GJIK5FmvcN
0fuyMcQ/f45fGR1F9YMXdvq3yZDq9gPo0DqqJCpNtNRmxzr7DQ5jaTxOzdZCie+t
r12OND4Qtlt62KN1t7vEJvkcnEcksX6SOy8ESFdo+yudKNo2RW/pbSFNPHQrle6v
NjpFq0lktwF6BNJZMyyVkmIW8Uc+pPPHmpqnRMbcm7a7oVlhKu80E7eUNK76Oviu
ql2aQ4vtX/Bf+9c4gsgW9c9dRVCV/rPqsi7RNSpBPfHN/ygaIQZbvrqo91X4jtTq
ZxrVDZORFYSKKdt4MI7iLj2My0WJAkNBYcSvX/B/93NxGXW9Fnef218NRdD0Q1AU
XcUcqxo9eg1Y9tK+HTPh/IONK8ucP8ZlriEbe4xjS1YHf23Q3rv6TtkPkh8FsV82
XHJ0As+bnhtQvfMUPeieCywpNrb+qTHgFcBqu/59mXCf4JKcQcin3t+GCfTWkzLH
pBl1Bpk+hfTbPyxpUsSFQqjiPU7il5NyPRWmYUWx3Gk7tqO30ZOlOZMyA8sZ4/bm
c4Woh1BC47N69ercHJmoT9+xqnQnL4R9FyMsvbhj9yFFfM8++rpYyS9ojfDK0j5v
M9IFVJyp9U5iLzMefV/XqzY8WT4ROH3HM4DvR18KfHP48ZGcbMP8X1mpf1VLdow1
u+x10801po9TSnHzq2Y6MGLtludv8cwpxHcmWiE5cCxOna3JEMI/N4Zpn5V/QIlO
C4gDXCROy1HzRzTJUddqWSQ/0QGoBZERnA6Vyh/JQAA4NmBtF13kjIdlsG4NTik4
bpwt4AJz7dvkj45wQlUV+xioRQtSujqZhXCR32Sh9cO6hQAEc+TwbG7WQI8iFZ0z
Y+GWBZkIJUHah8hrdTdjo65VBQbz/NQ9A3rjQgbXAhi+r1sQJmfOyaM0C39Pk4XW
gHY6X4t7cP5PDRz0E6MF4pEdkD9DxDJ0DK9fzAmPMDQwhR96Xs2h8OmYN71C2UBd
raVrAd218Rul8FE0Es3zvVgjp9viLn/Ki9HL/3QykT56SYcHJkobjungplYj8DCP
gbRyD45bRsTNiwwG3v8+JjprulEi9uJ999XMI2pVMAOa0769UqyBAOvpx+E/1lgn
N/jW3oRdOAYJSuTVUItN9Ufc8Wyro5udFWcVEGMRTf8NxSGih10Tt2eG1TWlDIGd
5It4CTHr6vFdfsHB3+VCJX0r4jfOzIg6aOaKPt95TxxCWjJL2o03QzQk5EgzQEQQ
5QdezcC9kmldbdwOS0YxoFBSOY8DcbeXR2VlJcQKzMzpgaxH+OVOVXoLa18bNmBK
bZjMhaCJn/bgDBndOEw32a48j+6L2qQxxttK9XhFYlmXHltXpF+1yTvpmRSaORD7
zmOa+B41Vg15TY17N4AqsGJHgOt0od8QID5nT+QrQlQJy4yKK8zfzMGumNHVDUzE
BCWPlU7WedFnLw9HeeMJGIQk8jX2vrVRtj9Vm/V7xQB7TotKmMYpeg85Y93zLFoA
0SeqslG3nS6MGQewFpnqd5SqLFbSz4liWspmJR4bf+HO+HOX+gZUoutdlQIYiE0t
b4vJx7hpsnPBHTIq7GNlaGIhruwKmv4G5BO5kx+PYKD1p5sfq1Yyq7kyGJIk3yra
fsmYukb9aiEaeneUAfnF7bu6nmorPJAMrPTVBB+P0zqTd/FKVSiyFKyBpU3mnGON
a5ekKUle1wtGynMG5ixeWi4y40P9Pquv5QQ9+i1xSvdmwtZy3qLCQYSF08CXJulA
F4Aq9XgkBy9hVwn+G5Q6nUXi13S8+66nlMGhj+atr9STTpPkqlS6qygzJS8lyHcy
0CTqiZQ821Q441aMRSrnB/mvQwWN/JM7VS2XlgZifxPgPm1dQiLQBHfWiJm99vbt
CV99yrNWtYSn7tS+8nT0FC/S6wTZ4ABGj12xOax+XyxcRQ4kpNA0XpB4hJmfaJna
sMQEP7KVWOgb3bR7spHGVMgnxOGVaNzcZ/FuQHwJ9YH6tUXvK0jroA+uQl7i27ZS
AEl0JFytW7Gdcx/NsouWu7X8/kPeg/ybanst0f9m3Jw4cyo4z+ZoGuIIREmzX1xS
MvS43I4bi7RrTizrXNQTmw2pslO3JnXA/0wKOg0UecTprbemhlpb3vF49Qinj5WR
5Nr/3FJVc2Rdn8U5WtnQ5tFx6GRwMMtbjYUHC88EO7Dc4IIiBeTM93iNCekVYCRb
v3pTe4V3WeeLhb8x40UkjrpoWRvy2PDsvxNGPGXdlxBbBMbpud+ejKQnn/iITin5
sOScew98IcR9dOhY8Z0jzaewRnggxPZV5DhB12ZdZPh2teNxWEc0airJufzkJ5AF
uYCJUIiJSvqlzzQ8DojV+kVane7CWFh9jCAjn/+5kgTE8WPzrKwsQ2Y60FzcD30j
eMdw1fkAg7QTgT9g74lDvdbJ58TR2R9BKMul+UMVzHF7QKgMj6Vmq/33MFn0847W
vPqW9mlH2mPb0QN4f2H1SeOHZVekRkcX/B3AfZFj5Bu1x5sxaPQF/ax2CBPlHq1M
GWjpPTAw0A7oFtQ0UJrmu1al7BoxCpT7JRXMFZvPYZoYoGhLLgReH0PN/HF9dg0R
Z0bMEK25XbinLvisRT5STe8zYdVEg53p7XKEILkIQ+iQ09nU0Q5EWfo5w7t7FXsr
82eyjBr1jEuU3RQgygirl+X8mpAekPABCiYB7o6aLapAMPaDkHIJCmFrtZl5vyJ8
AbcJaOr+5Hx4Wvuiivp9qRHbINbaeqVdQk/BB50R8rodRLojem82LVrcg9wlFju+
WFLjb9A5rSw95GVSZfu1qjO0VBrauBSligYVL6Za6XcGJHY0sOBJsbiGfEhLhzb0
h0R0Y2zeBidIl3m0eI6eJO163+nPEXDPTI6yJe95FqVA8YCb8uX7odBvpzx0fd0D
9sFBot8fE2UfRSm/keihLGZqezQerW5mZMvJgaEJaRtfPUcvcGadZnirvfmQsIaO
iQZCQYL9BWb/kMAaucS27oeyqEyHHfRdtUGiXHoUG/OWqfd8yyJREYkA8QVg2uaV
6/aJ+0djE6E3HfZmVYXMUIFD69cCYkodBuMLKvcrWArMXuOHBxUBOK9NA9xoF+7w
6E828K7B4DbJLQSjJyGj273BsZjmVv5hbfb/xEqK4EDiqYVZJsDL27VWgb4FSoJS
9IJx7bP3Qf+OtV8gwDosmOxFyOcyD1os4JRfVC/BkxU5eyjI8bAHXkrzHtEibMRz
N9Q6P/pZUSvMbU4c33j5V+NIb2hKewMeGRENuTbOCoN8tWBVJvGPB1cvVnnsa5E+
aGYq6pEIdzSzSxRpjsAlN1ydFAya7O7Uh7JjvxeVk8V+IGbNaVgZYqTm+xvJ5gBB
E2tNgmnKjuy9jwriday7jM8PmktzpkkWDKIpedrCcI31i4GAWfe9o7FCT4kw5sNT
x8k4tYkzbqqRhYqC7I865RH80Sl/vpSJTyAo8gIAeOJ9OgOalKQKliXJnW5T9ecd
HKQexnHg8gm/OFBmXYVhsyde/gq5n78ntd2OCicR06yozErOE3svx/fjazKJ1DYd
iyoN9J26wtnrVSarXOUkxfpc3kedbCKaX5GzyKh6RvKxTovAizP55qBFgQ6JYOJW
mgffoWF7crgfzPfNObQVw03UuUF6FN5LuON5Xu8oZax7fjdQt3dsWln//U3LhZ5B
0pw0crKDS+5lTRxsp2LtdzIaiTKKPYv320G4ztlUknBMR+yJwzsNk7qfxFymPuvA
Fc9izhSykYDy1ufq6ubhdvzyYLJ+6eWy3MyOeVMSH97dvWgjRM5zWrc1SNxM6S5s
f1PmB0b6ej+wHsx8/8zUsDtAsToZIU4HzGSFp5SS46CGndYneleoIL/yMdrZ+8p4
mTzcKijp/IEYQzdv6UFKKtJktmeL1WnG/oP9rU53gEokdv9XpNTJ0/fkHVWCsHZN
bgi6oZdh9Z6qDGzsj6+TRM3ZwAOfefZ1dU+mae4GsBKxt+Gk3DTLxspKaqw3pVOu
52mCC59FXNwu9oV6B77yVZYLJ2ZpZ8G4Ti47Cxm890TsWirIlRKkQ3TZ6KnwQ5U6
jXPnXJe3nzGy/gfD/mjPOyJFW4U258ei05AzdPmSFXTQgppfaaD6KTjKjNOmHUmP
5vkmD7guqXPe87wr9PZ7ihHt1tieQXVyca/uGz3UTzcSWh6SENYbgTnntQnzw9X5
DGdayEDO3YP2nUQb6eOEh+KKdeUnFQDxaNCsBIqBd3mwPqVCBQgCj4Cmce1sPkQZ
gWloEkEwrNBSo2LZWugFTJ1U83RYuQoliDkozqToIu+YAyIR/VAAuXMWHhoVVwba
orws11B0OkU8ZyOQd14Fb76dTnKIdQVdQUv2Oj2RYmdYa9PX9DntjxKq4x4yyTrW
f3veWi4aX4jOJtNCtfqX0FYjrSr+N4ke0bdqOcamwAV6fvPkFSdjIVIdNpAJy9as
mhtu6zDZ16/3rkKQ/2J6IfZJcE+qT++9/wSSe6uO2w/K9ksP0jfp1ETCDvbe0ZI6
6C1C7iRuDwOBDBFt3Ya/8vsqrdP52q7lnZo8Zfhesw2q6A6BJZBBfuysc93HRQro
s5GaMTTDu6tgmRZAe9I98Ed6gD8OSoO4ocZN/VZq4XMHN0/JVARGwr086hRgKMS/
FrECAuf4lxsYukBl76MUYYcXy31OTRGDgMxqik+WZDL0QGHzywEX2elE6N3XlveP
vkDZijq68TdDptu472T8Ssq0blbrEhcI/TcxXLcq5v/B05keQfhBR02Jd6Z7cXub
0g3NOk/UXbyMwrFcy/f2TOQTjS/1ngwsahE+5QrEwDiFkBo/CuGfxmviYIhC5xbo
JyGNOfcQWMNAu6jexz/9VcwaVH4WaEbLEogkiLluaZQljr2ZWZ2fGI9gnuCIE/qM
LjqQQ8FuH/TqJEGly6zozFBxoG0rQWNwSvqgzsOEhV9IAWHbyFUmBnrTGbu+9cML
ZUrqS9JjvmB31PdRljSOzG97JQpOplUbBCJKtuIQLIpTSlvg+U5qK12mQanVAP6v
kY6aT/3LY4NBTarOYFkHvxfi2P2n9POFn9ZYY4Ao9jt7erTgc2IIdyh8SomybgHn
AxAeqsPsEdgmJhSRpVfVwYkHFch7wTAvbyfXSdfEv9VPRzx87UB6LQGk9a2swHL5
32covrRnluhiNixhLrchL2yHWhUWPlAKwjwF5modhHJ93FfDGsRqpEyLCZzpbKbA
ydwvhcBijGxL2/VVfvgNaHFUoSxkH8/gv9z7fvb1Idd+41QZGYNv43QXatj+Cbb5
ntNui8KrDC8ZjKM0vWaWq9lEIsEJ7SKEn78ZarfnIgNPohGuEvVJJ50oxhyVP3M7
RvAPkdj3o9JwP3sR119FKhfRvhfq40mz6l+WFC2mWB2askL69LirVKOYdUlmwx2r
vfT+y1gyjPBXle4ITIzGoDoBs/SJoIoRg9xr6YJchRcblkqP6UNY97NJBLszqkbv
0J8u/uze6+2Lj2S9jhQXL+zKqTnXlTyTd5nJUozWelU8IjsqUNtXa6iriGvNrQ4M
EBFreTuiCMuqYY6E1XswWf9fG+Ufrt35wmDvMwHOJcCyjwStB6avIIXo0xASlCN6
4TXXyYIlLWkn7rUomuFn5+nV23pZ622hzU3jk0bAUIUt0Pm1i61FgkK7VF/NC2Yx
K11wQjes6UbJ4fQRj3lyAu1ucM0weGXpu2XesOncroFsNbOpbwpvCB8L4hrsT7B4
om/izYjfzAtrfmmiZgXWXqlZnBGZ9cRd9ipkTJ5TjazpX4JkB96Vk+5/kW3YPYtl
d6bMxnC6cqf/sQ0pKm8rXYIysstzLlASvCIseHX9BsAQ53Olqi5W9roXG+bP52Kx
Y/n0f3OlVqK9+qGWN2TP3aqOaZUyNBRTwY/eEfUljHNdRS/TNQWR3AChVTA2Hh0o
aceemv7bvomZNr1a5X72Fp42s0+l3Rs/uKYxmkMqId7HzQQsRt2LlETdTwi8H+zO
Yj8NO9tWcZ4w4CgQX9xEu1peDRoBghYMh7NKQR8YqdT7OsHISMa4qhl1dzn1myhX
rRVn63PxWMO1Lj0eSsRMufAIZ1Sjy8VXOeDbOFjB3EaAm2ZZ/KsEx/pVN71G2Eu5
3k2vhAXvRYuVyzGvD3r5QWxIUHHgK4qXUjO+G8nKvc/Jm/47GmKe9vYwl/BUnMfy
bkIRpswS/+p8jKbM6AhNKRyIPPIfI+/NgaNudAZjIDgNrb8CURi69HfFUh3NORnD
/GNDs17wJO8Qfaja2e6Q/uweTDL8dziNEJy1yuluO0C5hWDajMVAyuY5RBEP6/Jx
6LbIa15d2HRt7QsJNLUWL300IcmRgzqs8H0RGaZBGgF5aEiPQ8rBGsEj0MTyG+ft
1okByxYSXUoyOPj65+CP16Bv8GMgPggREV5oKDnyDU1IdoTDcwQEeJBKvv4N1tHD
O3aby1PTtwbbVPS4dWUT5FcUpA6tiKS+Ge6ThMVuXavR5jyJdH+NvHzcSkCsib1I
tu65iMRqAGKF48YQhbJxxqsR4/TC65wLBVaoDJ+BQfXg2h1iN6pQRFrW8BhloX17
Vxnyti6i8ddjiHXL5l0wDmxV5JAAXDk7Dgi/8qnFUUjNCJMHsRzN1+Rv/CFleMxD
O9ryYDwrBk58QaxKXMEARW6ymcvYZJHTF8BWW2DWOuMVJC5CQLDvivPkfoWLXl9H
eUq7CBBbhBjmuG6/usHXkHiWjpWtMmueaHME1AgsO2dwFlCJPx3x1xC03+7vc7Fi
60ZtZ6oYm0aDKECRiCvzSP9L996vhSJ+5EYM0EoqlcqTd6QNE7YIrLdvAGOHBhk8
1TRZlQsJOoSZx74Ia4oiuj0EKTOfJ4WRegf5ArpLq6tzxy8hYmi+xYbaMfNr+job
LIypho0c0GuEJzaXi7/u0kqZngtJyNnbygpoCr1d+XYfs9pio/7B6zbZMvzZTZ4h
XxzTpncsUAglm3AcufFrNIbabsEQ3CF1KUaWWhMg4bI9fYGnl6wmpmVM72JLs5F3
aAuNRNeRo21+Rb72j4bsvB7vmDInEm7Oo5qpu3/39wIJ3eWpebXqOesXSBMJsdHi
yaHiuG6DLYeYLvM2a8XMR3begX8FNoPXbQl+eo2ewlGXGe4igCmK6ZEAxJBric1l
wQnfFRtLf5luXJWmKHT6lJ5CSHXcP9fP+rGyW9A5NPVn8DSHyorPt1pk8+fBEZq+
DUuu81ny9Tet2kPSiJRxcKbG04gaCOj8bqB7FiLgj2t2G0fn3BsZ809+SAspMV+K
hgTjDaVKGLjTWq8x810gcEqjLP2iwgxBI2783Xh+v7SyWxdQdelRwbpT9otK55Nv
6OVBDR1uWb6Cz05icyLbf4WBsN92WqQqvmkUBMpFQzg2lq7z4VDyld5UQXVXhpuQ
Dfvu1I+1zLOjVKAgISpwiCKfx4lCSMELpQ8reQHfqZhe7ZfIly5FLqYSUmkmU2lD
XHTVH04qBk/zIi1CF+PIUn6r3bqBgTqkeJoUVJSI+KWdYJktJQaSyZpExR8ACL86
L1fHNeDNPWGoeYHV8FTSLAjVn6lSTQATiBuzfPQ8taJ1dPhp4XUB2hR3nnG2dUuS
Jkhd0DdTMl9FFJ/FN5RQkDdvlw8jRC/iACu9PmeukJpEnl1Q4AABEpW9FWhUAiGj
JuevSStWKJTamAGdFs5fTUOaPT1+yiktmHucXbF0c31Vn7B28sHmHGgJDVQUHwwp
g8RGrYcEh3vrPEIBMInhHyd8KXgW1C41Y1o2ZlBTgvAlE2TMp2TNQDsqqKZt52m4
wagbkHbU5GM51jCU93lyMMdGf8y66IkvhrVFTwPWgOOPDn1nI1fs9sAU/AGVVvqC
SGxnmpDvILZdXkfsSi5XWOvDiuDYEi9cTMuvIblVvlVHWgf3zOMv9CFWSzHRtH1z
U57XRe4VVtN7m0KZbTXnBduWtuGQ0EGHLDJ7Qxr4LbzDYB48l+EXOe+96B3fMTcJ
u2h9LfUrfuKHacylFDrMqRHX0tRsCe19eOP3FHpGaedcTOn7gY25glcxAneFTO5f
NKLUideAjxvBo21oMK69V5zsT3YV97HJX7mNKjVQ/0IatM9u6UW2moVDnbIa7wSa
QsAH8+y/xjQ1Oekk9xNVdsda5XXjB/B2jLp/sJUu4yMcpUhIjxhNca2dQCZd4UjT
QklhsA/vmye+yqxJjVbEOpeqY8jH2WgdpMznLs+gB8EX78977AunG/Pas/AY8C6r
0wFb3gcodYJKKNdKsbK3mRT2gE4dcVWOdx8fk2Nadv6AstEj3INhT6s2a9W66+cp
HntCoXg/yChurGMVAJTiRwd1V7c7xLHlA38dFNJ4tbH54orang0ACOjGfxxwI2Ol
Y8G2ip5kTQPm7R/d4VQSLDQ5RHlhRQmC7FNAbzJNXiRaaNiCKg7VhQ0PJicpmNb6
SMFCuc3YWR3LseH9UF0KJnETuZXIVOAcyuvJVLoXJBcNH8wJ5gHc1L3MsU0OtR/3
cdZMnyQmv+oHRAxfPSfBNMV+XLEtHqXQ2Qp07weT9357qMEvWnE+1zkb1Sqblx9W
tzC2Kz8Wl59FxiQ8s4WRU6BC6ETY7s59PaX1hjzsAMmcfa1mA2obbi+UEVGSRt0m
mDahrCWo1udPEDHs6TlnEiffXU4i3HC0WaqC6xIqpkKddhYa+P4+/G2gUlHSqOqj
ttTAAnA86CNs+vl0qiNT0lnN7cjE5QNikfXekhKUU7iOtUzo9PEZa4wQVebHGmSA
/RUWAPJI1Ig7SXJ3RUdOYPkHCF+u605cQJM4OWwtCvQNOqHMwQK8GgvfOta/750o
QDRjD4OwCbGXVrr9s+SQF2eRQ0XRc77XV9tso9Zft61nsVScQfZx9BkK/gg27xir
8L9ExOWq4X6eqPfUBs4c7YWxnc/cfjSyCBgWhjsERw5bS3EdXvTjAfYwdT8cQpQT
8yOpACqKYKi+Vglgb4zFNLcCKX0OCEghNp/wRJW8fHiiZ3QSlXcqJbQTz8jJBbKa
X+X8mADIy0boVsKfxq4uDILehUuhoDuh9lD6o1PK/aWQOzp3umPZt6U1US2Had+K
/hCp5sVFDuptMygBPG4yOjSSUXgPcah3C1/QTBBUlXVaHdv6HwQK4xUtTMoyb0TY
oqu6q/q335NYl/1m6QHpdPhldXMQfHrW/3cNQLU5ZqPz6A8DLbQJ9w9BDTSX6oC0
27feILt2Emsyjybvthc9QIfHaqGMm6FEiMN50JfOf27T3cLibN5Hm6vPFqqVlYcl
SffovlQN9OU3zuFfq3Eu59hmozdfLSkBo6Kwq9+ktrqKpUDTp1OSVRMTYWm/KN0w
H60VCjLFFxfwscLw3v+dYpB37U8eXFcrg0Ld/3iLc+FHmNlxPr82DESDIBjpeH8i
zT1xKx0dD8oGAO96R7xE1amzlJ2r+eXo4v02J5fYWgjTzQ70zTLUg/vGwXuLJ9x5
1M2R0b0/f8S8ClfwZkRJU0EmANYLRSV/tNB7tTPNTBcIAaOpDJsEr7nio6kCa0IR
jOoV1lxp71Lyu60q2PQyYcuKC/7QmjnTPj8hQz+g2s0wXqDDmgxC0c2CTJ30nRSJ
l7RxmCJEbkfMTvO/e3ayxpA5GeuwtKfan/WMvj0b1acbx//axfer6HQKRrshi7Ud
2AyUHA+UuHrnmcv4JJZX0QoHi2mb5PU92Cjg38+LZVZnawlVnp7iG0e1n0Q1Sg8j
bFHlcV+XQXSTEKZoURxrIsBEJcD3hNRwKhoBwsrAXyAabbE+r0DyTE8qNGGagY8T
3LnW2XnW6wN4P00Joch649DDRq0j2MGjgF6ssHXaom+x0/xaJI+l5ZxwSbpIZoJd
A7Pn/JOuCkwIfx5kqfxrlZJCmlZfdizKeMomnNTrOxyuqDiVcCmi3YjzRaVOtO7l
zsIreyzBrANT/xLGGcZ8Kq+kmXbeIU9MCRvCuCdxmQkhnynuTtQXdlJ3mmVAHoV7
bMsJPTAq0y+auje8zp7jq9wjJRUWzasCWuVKJoiFsAqFAW5ReZuHt84HqezxH/Sk
Z7F9Bzfsh1kOPkwBIvCOqSoIXn4MFydrSoHM0ucWxQxRAe76XCoh84fJgRF7a6Gc
c9pfgMqULj99UebmggKdhoEY5n2eAHm7pHjCJrixW/kPEsn0JuFcU2RK2MAO9Fd7
f6IjDqABzTjrspbDb4HU+T9s7QmHj+IZWyCuGRlSnUDR7dzg7LawJp5amKqXRiSU
L4Ir7RgCkQqS9EBc066aOhDRxrIFV9Q64xHaQLjrInBf8sQ021hg/Qx0wduovfna
ZivMrhQ70K6tj1Hy/g3iDYR0xuIazlHNCj8l/Eg9wug7KgIIE6/ueJNXjMiZxGCP
3c/KhnS8VZWaYKDp09ui8fKR9HSbIOHWHy4NXLqcubaZ822WWboUkBwCQpq3LGvN
im9eujUXtOJMlVv/PmHpII8uXbSLShAWqnTjhrt7DEi0z9DYSIwCJhHS2jgwkO3r
XbLn7xtaWDygEmcA221kHvjjcd4+MvGYQf2jzoVLL9oAGecHoUw6HSlz+IAOp9Ql
D7dynCbPBE03J46BKKxcRj2UGXb91Y7GgHUnwUYoHGDLW2gMhwfrvtJwfd4uxqzt
j3Zj8ePmcIeawAb8kYUGdanb+BuO9KBq4KZnUqwFw8vT22UxhZCYqv5EBMrOurGx
kKRm2SRByIQvpk3+vRCZidJdEkkc2mIxQVDzPg0Hw134IiNB7p+1uy+TeNaeM6D6
ZWM52zQYf4lD53A5/VD8CKm9WKOFssfYp7iVqUdxpmQ+w0kdsY2Td4YKF22eJQ7u
+7tAqpGZK6+aMxWTWUlQ+v2JzyXLpbEFYvNUxTHJ0y3xzbiQbQftB2koQGlLG96/
rPRDVjWvtgXiZy9wWcxilVJyZURyFSEovzxtmp38+Eft8Eq2zKHoOP9MYBvr0FoH
QjVWk3m5y7EiBCabBkx1xWPPaTIzJo/ELgnbuycqm+91YlhiBGw3puxXJ0/gpnIJ
DY3/f4CsjXehc49EN1C/Q+IRNA/isjldOwQ6htvI+nxBEFb1AxhvMc9hr7yOZkAr
zJoIw1QgUzVb9++p6i0OsB/XR1nHdX2/qR9cBqWN5gPXzMrkGDfJlGXRXKrPY/Rf
PNvalvQ5MT95+JXd34hJ/qpon4I5dDphWH1uRK9bxqKZ4PNVMk8ZJ9fRcJrXOCG1
cOxr8A4mJe1izW1WOzgzEe8tKSKmEIXdfUPYooZjHmlIMxhxfyLYCPc8br6YBqA0
MB0pX6pFwKNVsySXG1Rtv9XefXVp19RjtoBkdJRydfhv7kTBsw20zCeyjHn3FMlM
1kaLIoCC/C1hAWOO26WfS+ycaE9fyKE3h3UqEZ6k9rgt1duaImV8z+TaZ8hx1uGJ
p+fJm10Zi8Ps6Lw1phBSObB2keHSfgQG/t2WeYnmWSsSAlWSz4OJyla5KCmMS/FW
q2dl2+lJKVnqROIhWV3ZiEeO6fbJfh+FTbtBqxGqi86AOX3SKWRFi/s5q9pPdv/7
TC9abWonM6SbdYgNRPsTYOTJLa0kWvDZMwh7f4QJNUvaXjfD0WDzOOLKn1TLTi2y
AhKYChBX9HDawEnqClyyQOhhR7Z5/tS+0U17hVJeJFPiPjBXpprKAiL1dzEm5hOn
ExMJlURwQwWKRaqllpNt9CDkXSjsMOt/8Cb467gRXL3wXLm4/XVp/xiAXOtI4Mx1
RVUxbbVFsu7li6doqbdUhi/Uacd8P6i4i2YxDJuGOJt+4hF3wNHh/h2oIm2uaj+O
hjYRx2m5iHVuNrhUq5mjQ5jvdUQZ7vZDnplpuFrBxw/7B5JKgXMKv5l4EP1pX4B5
MHFxgX2eeqDy+Rn/Uv/g988fqJ6DWjicoDdDlsb+jECaogxPTCqLo/1sAaJYmR8c
jwESXb9sqixp5liio6oxeHp2VGYzoxWlHlgWchkKIzUEmNz++ZacJZcZfbuHo3nD
QI1V9qbQNbCD7+2yKlOMGUJ6u6gKmIpdgWszPi8jMg5vxnMEKVRqN5kP6O5m4fuv
zT3p8fcFGlKCluhXnuuYDS0/TL88qpbeZi0h9p5TSvH4NV9dSkV3tr3AwvdUPHh4
mU06V30XrPOKylEQJY2fKZC7PMc+8bgxfCnDSFGavVWBRW1z/eVqbQ52TENFrT9U
zoXVCnRCG3ZalYlt5/kkjvR5BlFoQyajOjF3uUdXBfo01morQJhkImL+4cZsBLwR
DljABWBUC6ozGlQtKuOVSPNKEbbItEGfeqb/vmZ0taVcDTZGFTFEBbPJPSsMxXLc
F1mpS3cT0zaVmUqUREE43a0rIO/vvLN1XsrzyDO18ESBe3P4i+KR1a04BO0MaEbj
8q4pwTgjCqU3q85OY8vix4gbY+aWQLN4ofTBkJW9Q8jena16Fv1NDQqr/m3SIG2U
CL3KNFGXX/N6nmOU//ed702PdZgJHH0G+9aIOsiQ/Vls1siWc0xExZbqk78dTl65
ixJC1Y5o6SYgQH70Nq5JfCT10pyi4o7q1wpbo5aTuE9pooPvXib0uH07jBRkPshu
/G86+to8Yi/saq/obehfi7K4AzoPx1frbP2OrZvyezGsDKcm3+U3bgXINLTRk24r
24WWwxrhGkdLt4YwUYkrz8jIau3XZm38psLJfINW6dOe09FCS7XXTkp6jj940bAf
P5xou6DtrRXl7j6eCaTOpiNLUX5YiFFaP/LSLWUqgQdia9DzCbc1yg0GaWkF8r5U
strXIZ65rmmaOuI6hy6haFkUw2qbXg23I3YPHm0Rljntx/iXf6wlvrCAypGe8xEV
Pg9CqfBc6DIeXnwNPGIKwooBnogTfQnIVBeWVJ7+pGn+DhXqio2pRN9cuEdmr0aq
ed3ZY0AMCnpH+RMsZjgs8RnBx3Bj4pIlqxAyV8uR8fgOghm7FMglz5wYCqExRJsM
EQ8TkMNwx6rY3cwBXcFuo7SKUERgPyTNh76nrPAnb+3QH6CWH/+y6KHo8AmAA6Fg
eT8d7ZVAuBQ2hZl4CvqkjKSFOtTxUFEUhwgPOMdAqkoAY4cJtweTzzBXJYZf9xmT
hzxWQmG9uFLvJ4d+30quPfZdUNpUy1RdzhTa/ad28F2lYHkLHElxKktGfhQBXK3m
9JoCA7zzTg53luQQjau7Kz5nQQ8OX16zob17SdmjJupSGzaZGYtoVugbH+MU5Fuv
BE2PqMC+3B8dgqsVXAEDqHXdMFQLkreJmJDaZjRT0iQBYwMvUk/ocBqp9jb4Xd5x
uhvUbmdmg29o8sdg/n6U0cGbIPHxs+aRBodgyp9k+fNiIU7r0aBrxOWQpbH+CYpy
p8OgFPU+DJW+X9GwIa9Eq8z7rf+Jm9aqxt2rKdzNneUArkVaDZVmGcGI4B0dPBQJ
jLUjflTPUr3T1KKfGE2q5kj+y+DjPaVfqSZPUHLz85W0LRpFbjasCSCu1mUX/L1S
J5T0bxRZJaeLyFASdEQ0kR/gBLQUEAUGgmPq2YJm+4cTgPZU4WUSmib4DyueR5tW
vlgajCMqkC33Wcw3iBYptYTk7K7lhz+pEvRDoobCTVJ3JP8XyvdWvM0MLx8EVYCq
ojSHVPOu9L/irtreFaNpNBUTVT1LXY+0l/iX4f8UgjCK7pQMQjbs9xF1oQKnxPul
eHolJXxrg/gxuMGDi1ru3Yu72Rylv1pv/Vt3H4jdcoxXdH6cRhv76xDg8/3ycqnU
I8yezEMidV2GNfqSUN6gE9scYc/HRl4YQNPaknj6fiFOZOr5PjuMnaQ5UfIjmwkj
tkZIekRHfT7zR/09PQkmjku3poVi5vK7XEGkMn9MxyzXWnXXetdR4ma+4fSRkFMp
cjYenQ5P97f/7IV6mqGVKCLpmksZEeE872EfId4KYKmhkYMS07wX7FFPlQppuf7/
8pvEVFQLHGynhGalZCi83rZYVIS4ab+90aC6EsMX1R9tYz3zw/DhZPKetNLiWl2/
uEOaiw1h/AdOgGQ68SgIjNR5axo4l/32AjRjR7JuLDmb8q8Kd2II1q6hITu7ynrQ
mDT2ldIPnZheBpHGCXbvqw/l9blZ/Ezvcb+pWcWTpG1oY9JW+bBMfbjsfi6TBqFs
H1ofear/GeQ1f7sarmxL6gL5wDtRMDa6zqiJKUrfaQ6d5Pzu0JGvTwPfYoaCbZaG
OhOqBvHE1CaQnNBOs0lV8B9Mjiw3N07vFPgr9HKs182ONFCVJHg7FREc1JWs8dzW
FwKRtbal9PMs3CFw3k4SdG0pOe6DXZjy9vioidqsn5Bdq4DosdKIuwEIkz1rjzpT
eESGaileZriBfiRBvmU2swfxuPQ+a+AjFakqNv5QsoHFJ5KRhs5IQJk6298liHay
87+OSAi/yldhTESXzW4vax8jxj4tmNG9msb/FaOG6uftKsRjSjP/W8eaKMzB4vph
BML5UNxSRRtZFGj31xplWP50eNVmVWCPir34LZ5xSr11a2b2nR3aY++8AZh5awM/
18T7bfWGS91lEjCN7Um1Bob6UB60nzzwViiZlx2oyuL+UBfXno+oaLEErdec+XJu
R/Lqw72s3EKI0AAf2S021C7r3VzLKvX4/loNSKc44rlIeZCR0YmHQXE0AcrsrLJD
fAG93RAP7R/rNVysq9MYq4GemXCPmHneeoEUE9PECINICP/MyLx4i6q+PPBSoii5
HxQfpVJys3ESXTKJkfYNGuavHKMtJDb90gsfrrlMYfO+ioYvbaw8+YNHhZHjVrqH
6X6v0j4ilvvI5pOQbBb/82Qxp9QErKlll7RyZJKqXNtM4jmfkcrnZZp6KRjbQc67
uFYQu0Ta/TsNVJSS2/ybQlEW2ttHRemEU2HXZ/1nTrL2wWAJdt7Dn2auUUDMjM/m
AO9hepFHZRpz1Mr6AZFBLj7nEZssFbET9rNQ2RDIFKm8EBCdulpmbk6LfcuHKZVF
z5fgIo8x33U2QZNDyDlPIH/rNIPYCjvMovdutUC1/CEYohDxelahr0L6zjn4VC+x
+S8Ix/eZaGu7pA6nCIQr6nXwzN8zb6hPPR8iOWl3ctpl5F4DuDINjg3Mxavy0/A8
klkoOUga4qQoQkO0dA1agdLMSFawKZPRg81G8CoP4cFqfFbesjd8OHji/JwwYh0l
l3CETJQ9uo40d6Cvydc42TpnN6oZLljkAPtHmwPLoYGSx2Xg0Es/BoSbhv3z6g2G
VB74WxZQz+VjkE0Z+E1JOyFBT11DzLWR/jlbiPZWQVQ7p6OMxqAc1AlNvhuQL4RD
5Gtrz1SVZWMVe8Xyi8/D5lbq4uuiiRfbPzBckouVN9cy90j/r9HUXUg4S50ACQpY
wkMJLkyaCoM9vInsDMEspFmIAKCEjYC6npcNdj7hgalfwqjfiJkw+nyPK8KNFM+Y
DMxpKdzELw5Nw/lRFo8fkJlZjPZ2POmGk2qwGQBQtXVxhibbbUjuViCmRp+BUs2V
zYth0csr9tKKNGpelvQP+2SsZdBEpLrM+9M+3lF7reGmZAhODq/8xWMoFXBne5dq
I1EY4ALDCtSDiCLyCPciWPmC6TDhHviJMY18gLOX+NSr37BXP0dHwEYY6mkw3IIX
bcsxoBXg4eCt8YoKpO/vL9+RTKC6EXqRUthLR9cYaGKtHLAO6Ixcozz+N39Aa+KN
+WV0mpeJ0r0jyQo/yxla7L1ut/fsOBqsZlFPGfFACXl6KKkZQQedbA+YDTuvj1np
rYwOmfXm+iVLA37P1vCi8UlQQYPNgLRCzNjUPg55U0pi4q2YRsZEzUBoDPmMRonD
VkE3LpcVqiPG2hOyk6FQg+6avmB67d43nxyZi0IOPdQTgcxu4WfwIzNCrp4hbfQE
0ld/lMMH0Jz1kK8a/VGxTsN7K8s/69KhLl06bdN3Ob9ZBkErzH1o7OAjCZet9kPf
tY2cFchZ9ukNGJ4hcizhQFReZf52wSTSCHTUeUc7/K30Nm8kD9Q/zGpIUbKob78z
7KCSDVKF3TjsbKjcC3g71pkMEk75f7Is0k5vrt2Ixa71IAD09suBWSWUbqSTrJjk
g7N97aMgLiIno4NqyX3z8KvDzPEGr+seXvtOjRIKKbiYZH/VXFFeh26ASMt1z+rf
6nPn1BxIzJ2O8NtqIQPxfxzEFCTwmAFeKLR0FehEeKxwiFwVRv+IgnXzCeYNMz+d
E1pXFKzmBcMqhXfIrlJAx3citq+9xQQ6DU8OfCCWlffMUr58/xc0Y915DHBwVsmG
X50j3bhFt7i8licW55YMSPmP2hTKasljmTbA/vfOg9tTvZHwUmUj/hc4aHEvrWNK
6dO0f/TWjS4axoF60yC4hrcIpHa1PBxnw2HmOjv8Rn4hY1Mzu9lDw7QYTgLxbJLI
XMBVnLfeRalcRGA3zJzs5EyWX/iYl4WxHwf1d6aXIEaLeyt4Ugv7J7n0uW0Daeqt
zlm/8ufB9iUawU2NXChSo4C7gDC77MX0KV7Jt0z4Ovqk9mZsNNz92D188ZTsVMJ1
xnVWRS7R4btcFW3OEQQIcekn9hV5ZYoN3vaznLUAJjHM1ExkqLP0QL3O0bJwq9Ep
FCMLPzanzGS3rGdoJbycQ+K8bKKwWNFjjOQjJVm2eYII6s4R6+mPsAnGk1H5BcJq
A0rMcqutjsC3hAkppOsVmH6E9+3IgRJGnSHoID1OuRh9vcUxe6rLSl9hVD8nfFSU
btggE0ItP9O5/AysENMfnawS7OKow82SeRWK9JgqBdMB0dojcHtB9UxhdywcVAiv
Pns9AxDMHW0g4Vyi1wihGo/mu7X9BKRUxNc584Zrh0jLYde1jQkz0IRkAJV2UYEF
Z4A/yf9w5pxw9mMqe9oR5/4YbSOQae0txOWwzu5vYl3QfKj8V883ZrXa92lHlVl5
CM4MlC6+Zc8PV5hPPUwKGawVcgXqwV3APpmhzHiwYmNw3sgYm3340RGYsUrgY2wS
jN7WOj39lyjZ4ZvrxCY872fUv6Ah12YBt/UhVhp+1F3pv4Qu5qdh+rQgF1KHSpug
D34M1zBoMlX0IHgIKBSXE100OHnRoyv9ufORvLseCsCbUpj8Eb002W17u9HbhJVd
6+4xNJDmJ6lktgbzM6afLxsi+WQgmSoSlRwTx2u9VaJHtq9ab3NfEa54Slfhkd5t
E9ymjzovD6TpCtiJ/ttDEoxCWutQhwGM/zkzRBpY7dvxsKvFN+CrDc2Rgshw4avV
dcFc4VCwrAbd0jzUC0HuEeywhFoffogLrjR5OahLRtlxtZUDLpQNgNIFdGizaHef
O+se3+XANs+XganHSwHXcZuAftmmj4U+WeyfXt7aBu84PmRD/S2L6GRiDqkQFAf9
oVP+xG1JlREolSVdixB35U4O9VZdyoiPO12PHmhlbgGDrWrJ2NWum9jGjqF8u4n3
7RAmsg6lBE6WtzY/j6DPzb4/GNx3qxNAudx+yopmu7Uta6lWgESpz0xynaG9bBCU
tbH0gPbaRfUPxK2b8Cg6Yf+JP8B0gy2jV7Kji6iP+mNhAVR82aQp4BTJoRwYACXn
n92oTPMBJdKXJQwj6HQyCo/1Z7kbEsEjP7nYMDU7Nvh/dcvwOqTRTJ7IeP9TiKJz
x8cm0JfAnyIMDq2mkADe+uEanXPk/pErsiKK5+aFrPp+iyxZCjj8kE9oRZh4y4bf
iWVWacFPYGTj7QrF32wAAm/EI3yAy8eem77QQR593XjyWs0qFQXZSRO4bzwSIRSc
8EODy/0P4AAwYJNFNo3FW6yxH4e7Z2GbjjpaDYl17oWF7NSYSOKav/amnU+s8y79
d7jkoQ3RoTbABPOWLlDfMGXsvWnGvjXvAK/R1TNxLHNVw5xFOoY4JL07QuGikjGg
GxOerbMpiUA8VbSCbhyfH9rfTQmFVFRoZ7Kp8GrcZEHB+g+wA0S+RNEQc6QLpLej
g5M4W9965uJTCjdvuFTMC3srVMHTqKunIynjzEPFr9LC4SPIo5ep6qlPo/68IHNT
5XHBFSvWB6x0jO/d8eNZu5K3EDWc8w8IPyN8S6YMfFSzS3E024sDyDzPu6SSUoGe
o+Im7UbU2Jm1lGJvUMMzldygl7TC6WgX1Z8qID8uyInPfbe36KxqMkr+UBHA4ptM
a1B9NHbYHmbcj4chF9+GWyNXJWMKWVF8rxAksq/zfa9M38c3t6MaIXZxsWtlQQId
4UjiPmqetZNrckLdL0oE5eotVU6N/WyiZ3fzL/QTXBWQuEybmSPwIqcNajfBaiCr
9pSrgj+jN+g57Ojqq+XFYCseC+U2ih8PUVnyVWMASv/eTskdGAMD4kXC0sbm5ZC7
AuQA7FFK+HxYJxRuKNXGtTJLhbz20he4qtVa8SHmJuCCwDImt4jvNEdb/dpLUfqG
BlQAomO1Vx4ncNo2Ff4IlT06SRxq+F8vK5xl/dqFPSAzMQcsfLpUFoU813GuzUZZ
Vfp05R2EoAq4081B+g28R6Y1OPKIF7nTVl3jr4ySx/3IZX8T27IHJKj+G2x4x2CO
nwmnhTf8HTmoKtVVxMag4hVXaKUNyd3h5XRaI000iZmczlStOy1JScQNSms2FUwT
WTH74m5LJ/+lkv292NUXHNdI4vfPeyalQN2B4werrCkEIolodeqrbRd9X1A5k6/F
tgVynpIC36eGM6CqF9sDafXV0NXf/otA7uNLMfXymI8Gb/Arn7tYWX4KvVfd+lxV
8HCqJN1ZhOoEAnRqT2YwITAcFbmeJM0/BWI91QTiaLm2bu0BlM20iUpVjFGIncVW
ypjdsjdyTWIyPPZlxbyoe/ygg04xdJr9IhZjIYvo/98pMCyS8d2h17QH5AY6KEyS
Js3fgYCEp4iHcgOX9EFPgbS1yLuQWn+fLw4YTSg0TS/4JrMVW+Zj7hoGT7XyxNr1
8nCyHDUmNU2E9aqIY6K8Z5Chd3E+lFqrirApx3rSvZp9y1Q3tTXu3oYH8jg34Lfq
u9CJZxQzzMvbO8Usppsd9Yq6rtB0jcnQkbuVQGpmXNA3dmVKtVpE+ej4QLmwGe2m
BPWwl3ESZoTEaHH1V80PArUGtSZl5KcBBOIODTI88JUqzPcdOeX5OHX+8TMMxXDv
N7cvAtemg2kp77CT2YI0TkGfljiZxj3SBVTdzQSIFY1hjJR3wENXheaCcsi1+fe3
diSwRzLotOAPZn8gLOgujBByvPTcNspgtM2sW1HOR+kBSW1m9J9CUzQ3y+1sZKip
EoHNTkqF3uoANYOLwMT9NrRsN+NalUonBgEWHhNkPBnBkuwEUSO+m5LKGnWI/eCV
rNJNcPue4o8Tct6UkNtaywRd1fZ0sociDvYITqMvneXY6Lw/6kHtJh4ViGZ3HCQR
TKWD6DGAdLNuT5u1fNYel9z4QtUC69GcIxcIweK68CHTb19mItbGvpqBlUT9pUvd
HYp6Rbh+xBDcbEPFM+EOgv+tICD/hxCkR+xrEI5/SvTpdBY6hYcGOASZgLl746Lf
AXRVy8UToR7PKv9pNesSbrmUuzIz540OfeO0xCYGN9Gtfka3CUb3+2BxSaZu7DEq
xOPMbWRYQ/iqvHXOOjuDhXqER5Nqh+V1RsGCdCIp9YSW3ZWuIevVFRKNxvj4dVNb
pN0n80lzv/XRuet1e9+qgcvPhn86caf2pKH7vdxPgtNcdMQ517pN3we+5erM08V5
8eyH17yqHnW0i3j96g+JKS4Kljy4JvFZWFo6Hsa/LEoMp8aXh4Joj2ByK88j70yr
2I1LfKdTaBgkPwzFimjuCJ4m0pGC7VB99bVHUQDkpuNt/Bzyc2UB5sHQ9HXhigfB
TPlOchYste6YDz40Hu6PZ+5xoRyYf8udPVeYqY/unI6Sm4daw1WmYKPIpeSYmi6Y
T6iHm8VEZv82WHao8Qs2Em9FP62X7sC9OIz0kIGnzeAryaKUPBwUrIcVVfVP/DUm
5sy5AdFZF3xi3k3dFf+I7IOsNluJeOALowhYU9kv5GbYF0BzMPL4cbsXdlVbt7p9
4Ix8VTKHeJQIwlvX8uoZFLrPQgm1GCxWf+EnPO8QocvFMhJq7nbE4absuGIsid5i
RTCDKqh8XOemPQO+ksfKrqsrYK9urc9N+SzoVTad9KMKK5zaKNBB8xy+njceq9aZ
ZX3N8YJjDqwlrBZwILfLpBJuBzUafnqpbFzm0Boz60MUXmQthJnW1W9ueWDRr+Ui
CEggvwxsof3H6zudeUSafbJ04xmrZKDoavj2Ryc5nH0vQDFObtPZz9UHGnmfemxx
hgxqQJS7xuO3nOtrWuiBgHkzsA+JXphkjohAUsL0tor0+nwfZQaq3KlawRUUKpFY
dUAZtC/AmYZAvgNov7atnp+yg5Hh/aErz9944vDgdSfY7nfB63wVt82/0rEMSIUs
Gqs0hXlo6WTo1WZLJeDucYw2uOG8xYYGLAl/6SYs49jUiIHg8ez/VY0NTqhYEv6g
DbsvTt3wZaC8wAN877/UbZB+tkxyCCvbq5s8utKQgz32DI2f+ChnNuOu7z/yF5qq
IYBnjC4yokVZ7NZ1IKXf7xXrZpiGuJXOOGzWUD/eeQGXkiCShYy+sXrIwzMOuf/s
Tv5uNeRqZRueO3UxehwUCFzjonPUzlFiT5YDHmXoSMbjXxDzFZr5YZAsg0UAX57l
1mOEqYCzdx6y/uYXDDQSRGNBV7OK2J4e0Bn2PoeUTY7TY4P5g8dJEyr/+MPeTKAp
ebCQ7uY1Of/oi2P7p0BjawFfk7gsq583PjsxykG0uiMq8bnbQj71XGFO2m+ja6Na
6xej3CJh+s31RPslSHA4CerUNVvlpC/Klno0U3fmq9Ci4m9rddVE28mSEVX55TiA
UMYzEqh0vGFy58n1Orl1uLNBgFcbqJR4DrWTwbaEafUwOdhOePJwGDzqUpOcAeRO
4XSB1R/WUJDH4lemiiSfHbZS95W3Jnw4pFOQ8sNmJ+B3T4+8hVYlyaFfKxi5RGGg
Zwao0h68I4VKPzthqhPvKjzBcxIjaE4gRp1q4VjfIlf20oBUt6Df4kubnysPp8iU
sWumnLI9R/eV90iXY4nV+Vqe4r2gywLrzBr7EuVIuiT4OhZLd1NEzbeTTDVZhgpc
8YuN3LQJH8o+UTIQOQO7wkcx3uH8nfZMBGFppD6XBQVCM/iEI42nMiYBpxqNF4wQ
jkyYV28VTfq40UMHeG1akUawVCvw5APTgHBkeEU3N8UvCVmESxjsPkCqyJuNvszF
0AnQhdjn9WYW6Tt1etc9vCdlig5vFsoVmeEnCCr6DMXRRmQH56e/yWrokRVK6IhE
EPABBS8I8/Er7JUAwv9d3f/pZxVmF8mrkQwciSJM8123r9Pk4t1Jroiovgu+DmJr
Yee8U2gaGr9CtExx99Eb7BrYbMVRvsKllkGWiT3wUe5QYI1ft4oa6WukkNWnzqM7
bVaXWfkqaYTo/rRAPDDZs3Avrd8sL55bROSb7dcSwydOnFf1LqmZLQWXV5Wt/lXv
I4ORyMMaP/1Vaybik6vEE9jhFsqyf9kXPL0SnX71kD2vA3KpVmwVNvqA3AAYsplI
tJwFpxuySBKj+CIDyrZO0hW/8TLScKv5gBzNuKiV6RRgPU6DTQ0inTuIoa4UbDhi
MmZ7ziF1tG7R13f+dk9dysC+p9clSroP0luI4y4M9ERlIk7paCLS/NfBU2jzvscn
Q5KEXOeeHtWDBwDsaexG9eadq4YD0hh66PRDcrzMpy3BOzf1/7oGr9Z+4Dgyg0HB
ZAD50VUtXVxXqyQmh013SrOg8TfWNgUdPrpxWkWSEgBbdO7zLCBPRo7G44TGCfsm
lWJ66DWfebkV3PyIWYrXmZK8ChAkVyB6HtpU1uTRwoyirSs544MMh+FbjZjzQqkm
kki/82t3CMLwOK2dlRNqjo2QBo2bidXAval4J/9KQzvFh39GJxAavDIymhXMIFIp
5ZE7jTzEHmYS/OwBHs+QglHEe7s29jW+uM3ZEj0XwYEqECQCAqk+2joues+YB7jk
pDqYEa0smSsgm/QboH5KuS137ytnynTNWMvk44u5Vh5+jxDS6zEENMhfhlLlhEeu
yFAdahjsVoKXvwN+KG9juzLhxv4V2l8c7+DsdFJPgzvbtx+CHA9YRoQ1cQbqRvIa
aLi9UcjsHLfOQB1vWPEN7Gmm7NtPZazJ555O37hfneKxZEspC5+8a4/6DXnclGHh
rBSqkhQmPoWEbYt3W2Bpbx31sVE0JIxGRiNvJ/4X4RanjLtNDh5hhx9uQFwz5GiT
3LQM55vMWDmcYJUNXc99QqwiROgahpZkpOMAFpFqk6JKLn0xbASuEMvO4iF5h7/v
+mkulco3oDcjsc1Y7iNyjFq+eo5kJmvOLNYwhzLVob1r9GcB6i8bSCRjDYHOXqLc
xVMLHIZgo1zQm1uPbbUIzZ9vPSkmRoC0sYbQDGOtiE6+EOduJnzPx5rZ1219n9lq
16BXqsfs6LlPE3Q5ouM2z30brANKgVZF5cfCNlCjMM/jL5gyU9GveQbB+iCVOzAo
2x+/wX1yzxjkkLI5HXamkSuN/uNCjUI2HP+jRRZ/UlRdzbTE4Sv4T89zK/p4eOL7
q696I6LAQVW/d+NHd2rfXWWc2E3IRiYHElza5xAztpg4TLYJIXOCY1CUY3Bhh5U6
gHdeY67K93OrdZtqLrzv/JP0ROkC3W5TGtHICVlXpkvVY0p0iqYkcM4qktyWgR08
33h9OnFfkfLGHmht3EZrpk+xzDF5tBg019Bff+0fPXHM5MhNHh2X2N+Wki90QRzA
tROv/YFCO+rmrbU1vbKCyjOMCDuN50LcE8cB8SZhtswSWWd2fjUB3M/F/BG004MT
gVE5goTAhspI15pO1uDj0T7wadOtzS7ipXGMwXrja6gbE+m2E10M+CIz/Qi7sGpw
4VNIW03jYaIWMpJdSdq5SpI3mE6PB1GCudWt3SMrUOTCVxXM8iuiVORyG3E3zLL1
GRqY3B5s2bmjdGQwbPhxlm2AvVAmP2BYTkDpv2qEWKM5sfJD69fMOkaI22Uk/VIp
8lmlTTS5+f07XnLbVC8ntWZ7FPvSn4c0el2fZ1PRe7SAHK0J0zN8yq/tj0FJz4O6
y/zhExyRXHBBRGIOa6ZU5H3OpVRDQDsO7VAM8kTYxyfoG46VA1dU9JR79oDjGDQE
RRCpqK0lPtLn27VI+fRkyL7mN4wXk5JtMTeN8/+KLOwFIWPgZCidqvgrXkJIYFkB
vEFmCuU2qeCjxMTqlc8vS7HAX6F89rFShf9fdQHlSTVR7HCCfodQ1lhAvIA3+XBb
2dn+F8w9lSbViIh8jcTDDn/m0O8WGk6nhzeRIaxKcTMP2R+4dpCd0l33B87q/7g7
+PMoBC7cfpcV1Fhd+wVegqTla11T+SVAkGg2KuYznWpHVzBLUPuyJHekLLQcL4K1
gxPtQyx8bM7f6ii61ZddnM85NUxUPL/Gk9eMKuQSJ/+gX0ioX8o45UXHCgoBEtO8
aRHB52xejH11/u9Ia9s2BqN9W1xszgNlLy5f8r4Tgsd+mUgdISWRylRHk4ZZWgdd
IumygQRmIXi9GfUZvYP4x9/8JNZLWcGG3GCkm98bykruOaaCtByQLBz5ankv0Khd
RjVXwHyBWBbj+16lRKnp6zV2EwDi/27/yQWpJTf7POj0Qdy/jEBjCP7ZHgRbPSpj
j5ot/8/9jfM0oJKY542XayboadrCxO3+t9DfVlKEAM5xVzMUSC6zCwQbjsXdzO5d
cyBARARRQWLiKZ2JCui0i+ae2AJMRfnIXi6IH2mEU+pRF+sbpffALasr/8XE0oqE
oC0CVeZHYurjj937UTpaLwiFAfSinIYstLM1Y+HvJ+WWRmJ4oCiKtBMtlzI/pBU5
VcmjtJACIIJT1QTHA2Uv+Fs2TBBuIGbaCv3ZSEJ3XzQKg1MNGkyH5dG0uGnUWbP9
UcP4kwZIOw6on8OymlAQwl5N8ybf7k/RPVMQbxGglW3BnkzyvZenMyymKJxseAjH
oj7BRBZaHZZa2zEUvz6LNE44xrz2OQbrm0FD5WpHVmdcw2Gzlae0Ctsfi63nlxt4
Eqdxkl8yTfocriuJ6fK+7gJLhft2ZSepdNnNtKKBJA9mlHddLhxijBxrS5Ldnb3f
pMoV+fV2muVZaoMDX4IyYi3VTZwPBZ/HQuLaY/E5wVdO8cqVUVInzPveoziVKcGx
ZpNAXpfnOWXlCm2QjNTslf9frr9c+XFI+MNZDc0hrNrqhVD/e3EsvtYtI2MyHN6r
uNsCtu7dM0zi5Zue03xhvWEtdCziWgWy02lvbxpQLkD55ol/1J7kT7ycDQaYrbF1
0biT7bJACOMn+v9221xm/10l5g4Mpu1nVKkEPGuuQD1dnZfBhI3Q37GBIEBehhew
DNh8OGR9ykvUgmJhTQpSPXU1y2glrF9Ggx3chGBUTdI3Y6Q49UA/N1P10sEj+XXM
EDaPsFkBq2ql6ZaDRUG5WlGTxH5bV1tEetHX+HhBCPge+124XgWExjH7Z/tOd5u9
KkgcVew/bMoCsI2XZhofSsMDK0XXX6eiNwOo+VTTaV2GyzMvBbz8d+DsDGGOrvz+
sEWKOUiLJd/ZLxfbdW3OOXI82UzeTX4x/W+T6l1eCfdiQWz1vPXDm+pCqKKUl1kX
n5eULDQYu0KGM4ELHxzzeyTSgQqvLwvE7XTlfLjNxOEvlu2meM+qOe29U3osoGHd
eXm/JY9NE8GW3z9N5bWjS26ItcuG2B2AfF5G8F87eDQjkPqfJ4sae0BzFnE2ab7R
YgcYTtzYreYdJIYNOxlZv+mvgVW6nWdn0Ej5Sq4ZckUmGtKbfPOi6B5iKMgfuNBM
iZEDnHH7w9BTrI4lCPMpZuLOYkYtmkRUmGeOx4AllPbGYChXjE0AwlwbuDyfYLlk
/G9QDCC9XiNjibKYr09igdV90MzT7Il0oBK0jXhOmRI1Mv+el3bBYhUi0iRaAM+E
LGirzMBMNo1B8xr0HUOTFazRRga9fReIvI9dMBgUmoVrmvjhQszXyDmvJZziAqac
spuPH3mlAObtrQbUr3Q2bOMFJ8c/zWfvuv0tulnGf4TYQYGS7hFtwoMFJiBOK0iX
SU3rdjWmpjAM9gyC/xIaZndXKE5LGRRV3HcyeTh1IxTXYIcAIntlQ8DUw+juPcyk
8A4+SU4O8b8hs2SaUQ8jhM3eWc3gMLB08WGecDphmR1mztOaphxCcNMx0xypGchR
gAwBeNC5FCQ5MOMesDb4Lh+1oJivvZ3KVjpHF0xYPNv0YHgdC+91rxduKt7Vz3de
7feucnIOxgjyhnbB52v443QtH/guYUys1iPVWKx4aqKQ8K9xUXj1oo+9Lykjs8fM
3gcpUgc+yfPfBQtiMpfZYFeq6doPBYql9mZHE3VsF23xLU2bz8auAftyKXZpLl6d
MHZFBC2IAIsD4d/UE8orseVvdRwKiLYvQinzDjqRoRRj87oQlEDfI69eY7CJgnOh
kgjVlBvc5Ju4s07u3Vii4alxZtGMIMY9RVO8h7USBKEkvH+sE7fkdL2xu3joVl7S
GlkDxMKvOagiXr5wh8c0Tsjkgjq5Pj+aG7nDl4+VSI+QRjB+LZyF0qvRGQyDGP8K
2jNdWyaTZvfpRLedODtKzDX4+EXUJJYKNfAgH8GIwbuaEERGAjdZBro1d9OUNHWK
Uh94AzGy3T7hMKouqkbdSWeh9Ea7vJX/2Xn4b0RACZSp7hVHNmGuPhheg+qVMvQq
oziz49J3WRQPZmTlz34xnbW2h6tHyyG5V4oPrkQgOlHiEKJsFHs0QJMpwPj7K3OI
oDQE2Vg11+aijiqhS6dAQNy3QIzNH1U4owgEI/Ay+tN9iPVhA+yZLW/ewD6oqAjA
r9L1PQZeuyHmH7NhpJXskIG0AnljIyzlCic+0akG6gA+B4NE6ga+LGX0IQp0zroM
q+tWZ7A1gEmjQ7Q+Zla5/LEs10zYYt++Igb3iW/xnNr3yf3Li6fwEeEqJa5wavYt
vBMw5vUKq0vplo4waNLg9HuhkXsAoHrfo9kSl+wxWXV87lAE6K3jDLRfSzZBj09U
kfKVgMWFFVOqhByA+1bLLEEaS9lCY0Ts3F/M2UKB7EtuJ0Y7evlLU447OZJmg5Zs
xLmYMUURO4bWwFxs3Tw6jC5KGzeUNKx+5VyMyoDXltWsEB0bcWNrKlMLxOHpIDQW
YZmMosjGKybJaCtnqASICZB93FTh+os7kpILE+joI18eb9fQgGuDof3Lz3j6niDw
zP/JRnjCFkMbD+vgFEXSQosLsVIevwfK0aXMH+oqW3dPnF5z1f6wjQG2DjlsiLBj
yWDWvL+WmZ/qAeQ3UxWqgbR5WxDSSKRUNqqg6WI9/JYMHkWrjypy+7EVOnjMohk3
xo2vSysc142CDhzoxlv0QjmYUI3LxBaFUaQ5JMzUVHtRLJQaFEIHGUPFwO5Y7vOf
mwUFPsJgHYvgq7IPjly6iVns7+j8C0xnGQ/RDmikjyr/DIyYcfGr5vlBCaZU8r4P
zpdp4APM60q6QI6QNPdTPwh704hGVzRY71akfSnsOIQLxe7c/5Xo3UuOS42v5YF3
TwoMHaS9AYIBWPkByLfITTViDowsL7jFNynEGbUet0Yrd1uqyhPMV4od+O2ybHww
bk96xL/n7j5tAVJSfNQdsBC1GGVpYdqjs8euIZJ/KVH3GYZNj3wImutEgskFf4pu
yd9Y9hZSF33MFWrgGGqLyjY4nzabR4/Asjz47SRFKuh/HwoKY3x/+JwtMrKli6q4
ufVGHG2EzmHnvRiipJlQ8UezRAtmPfrCml/iqyxdiQ03GzrTaYnxvyvkpqkXRqRc
zDu4Fe9N3mEcCA9/ytCQfPyWUyJo+SrE3tHvb6gf2FxMxpRUi+B49ZCCggnEYHZI
sdMV0nR15zXEhgLef7+OIHGMALbIifksVbdRQ8I/Os4L7jQLxMD2X8nGgwnanL0s
jPuJFUCP/0N3IiG/8V/og4oEZ6c0XqkkeXx0gJQCkF2KZvL+eP6UEo98AIoovq5U
5++nlToez7b9mmGLDEWx/mt7cPoB3UKSvBpLv0BKLisv4bvF/Z3t0Tg+u9vk7dZX
XyGwxYxh3JtWJKyCblBPXvQPymRKqOJzRrgdk4t7olmjt65QxTzL7msDMP4p61sE
Mx+mS2Ss9S6iH1umX6ycCs9nmLt9ARkPiHNsEkkGagvGRH7LWSe9ENJhOEOTkQk8
KIcKM+VLsWOEYOu3f7x9qH0MIxcV2r7W112AIeQJal8+sxMxOD+dNDT/6hP7zciM
wRCxn2KDUJvE4JY8HbcatyfxNLjHdqJPTmU+9UMpSgV7676w9p8RZOCTPE9FoUHg
rAoaCkUQFxfTIRI4yIzOCTpQucYbYVArDyREOK7FPbhry2D42Y2Zpyor+NB/goXY
XYP+QKdkcGd5WK2q4bMPq01VLIoPEvsf6IqjcSDq7tJhiXYIipcJ2A7t7ZugDweB
2FVlGHob8uAWDjyjrrv7OYtifcOhypn6k84DW/pdPDQUaoQG7mIamQ8E+d7InYe2
unr4XRFq/F2I5h06ORoyYWodL1WGJ+Vn5HtyOH5Cl/jE8XUi3W+eLmD/T0+dQNTX
BaWlwSUyT6MTfSkrCSoUhaGtcs7yyU9ByduhKeUKydIy60eVGIxpELmpKu6DkNMi
28ZEDJimq8Z6FbFHhcKt/xflf3TpQSuZ0Zm1W/uDA5oHNjlua19H21CdVwL6x0Zw
1KffTZKkjddpnzPS7OXveOiforD8UP/3aUwutxx5uma8b128HJVQMkCH9zhX8hVq
BONxEA1DpLXZ7zXhDX8rSXMb+J6w81/7wC31fCUpcrKsTJty0WMC+AoFIpHSiOki
fN2ZjKVC6o9wsZ8YbrXbMy9XdbwUOM8twk8PDWVOePbxyh9YBaImBggVLTPpXQNA
bBzSHHxcU3RkRqletWKlaRieFgyFi7Af0Jk5nX4W3WWn4VF/jBQtrt4gq0mUPUTZ
InBAErDEjF4nzXErDWxWorO7NOBZMDcKrp//WkMncAEqyc5bD76Y5HqokfX5XqXJ
1lGc7yD+VU99wirkg2jivB86LehJl6iY8TQ6QT7D03+dju5II+O67qOdQDPMSlbl
NPPpoCz24IQ4/dItcvq+HJp/U1yOHuyEn6v8eAqMIQflL6sMPJsSNsyWqesaYBTq
Q2mOr9p/y0VlzZutBGejjDbdYuBvheE+8Bxl+xvqs8bOhlAh4XqlE3kD8hRjFzf4
DoFF5tDL/VlObOBvjo7XNXbQhtaxJwRygROmj0F2SAIPTr0yQMW0gsgdxGhi0r+5
jzQSwvnS7XA28ToXgSqNJrTja+a/0xST0aK1f1Sl4W0AVGkO5ad+ol/5dG7r9QEZ
A/sLbRJnBHh0AyxOudt86qfzBLSqepE/P58L1DkMHUF1+JFVJMmqfOpVrCKZEAxK
vGiiMKhwpDz+9+VdE693ZU4hnVQp9jCxc8HYA1/ioEjXwS3LohX1+KJVKe4yB2at
jUDBhKPl2T41r5lvNZq2bSqVx1i3N/elO3zehKNypY7YWAIuCPTM0sfXP5HA5MmA
DL7DM7U0gPiv4ej5fT+OPJ17KXvjPlBm0yzvG2gEF31ZVtpJ7xLVSxDCjXlAOSBP
CRGg+Krme8Ioto54MBYL7n31bQX0G8DeT8NYvOcPn97Aqj0mQOVpXpyI3WcsNYdM
s6VV0IAdcZ50xCKtIZhtcj1kf6vTBS/0P07zSVMwRBubic38pzsADIpGXsLLgzjN
pIQvHPeYUCp/U69AbKTMEB6BQPHmHMTxt2MFib+/m13LxqKFlGSovjFAOW8ZRLYr
4zWIfw3UdYtyLAMCBW8TF5IgxI7z2i+XjM4dfWmc/rCllLehk0tNlV5JbAB6cwCl
1cWi59xpuv2Mqt33D6/SCi3KB/Pzyltq0Uy7uM2KuGdWIm5N/2s/j48FjFMZPT6x
MP3botba+LcoEfRjYkth/8DiY2pakgDH/NN6RH/CvJs4LNFPUFaYpuBcA+Fv0/xE
dctFD1lmCX+I4Esba348kcP79okjv9ZqYTmm+7EnPyrdye3m57PY4ARN2gOmrCg2
4Un9/ue5fkWPlNciiIpXSYCGU1VeCu3Y/WULFO965+1FwdGmg6yx+/L/uT4ILhPB
BfV3w1HWBlDjrXbWOY34T+9bcLvio+h9NJgpROdmi5dIni9ELiMF14OuRep010Kb
KdXNKdbEwt1BmDRY4VCxJ0CUjMvkNYXi/fMqT+w+6GBUxP12P1dHxAGjNsEw7SC6
19DBMH005Uoz9RTIgjhVxQt41mUQnf8wa2Vee4t3PuumD0p/CIPxCzvv+zmlXokr
wXhlS0uHXSreknMnjeO7KRy9pgM7DyPjBcL3XBaeULXNSYt1o1ISRarTNCk68COM
sExCHU1Yu1O+dcu7aocrqIhhFmteID9+x/feqqCj0C3z5HqB2yT6OIRxdeBAVSwQ
BzHkhossDcZPBHkGXLXOg84750c6zsYy0rJpL3G3uMHOAxDHBbE8Fd+wel7R2eX5
qkKTyIpxdaf+m0BUkzIfzi5nR0qNBjDPj3ycPsdZf3bmzpwSYs/R2rO9jpeobJBM
keXog32Cm6sLUksdyRnHiUCbh/hlkMuqHS3535lt8SHfCHpeEbRmeoWdOQg0Kc6P
B3/2NdV+EubOWe4zXcn4h6zvZHAh0YZTnodu7LDdgfytyuqtKTfOpaijtZQoNLcJ
dUQ17ewWw0gGoHK35iHSQhkjSwkH1BHqHL6w1ulJ0/A19jqxiV7fwtBQ+AcTLpS8
mKVtj2Ri4G+wPIvmXWCH8glaIft3iintnhAGhuZIuEJjhVCVzEouoQA7cvAsHmFt
qYvUqHf50KODUTaNb/vg4M8lJ5y2+A4fbbtkLKSqxQjemEM3VMDcdtUjMkGyaMc3
C+6Hb1btRJpehlq9U7s75KKx7pEGFfkfoZMQOGYMO/vcE/7hIQHOqSJBCIUu7wnt
rky76BhOt8XZ3UgzwP27suki5E/I/sg/4qmLdFDubONjuTBgcwaQr1ZIphwg7bPE
66nlH6T0K6fZ4rvdTgw1FA08wlaN5AG2hBiAdJeE4Bw5vSmKBRemC/yL3uDrsFJX
eBZ/y4aFUiuC4xZrEK3UpwcwhlXdecRhO+RnFb1NKAUwYmnrb4LVCu4Vk2Wf/uZJ
Gvd8Fe5PPfX7DnfUuKNcW2+qirVmYBqlSUS/cWLMiy0VBGvTRxUTrMsHSaFB2c5G
zro/YDYoAiB2gTMVuFTXWCp/xWCFgKoOXngJTpMpqTOze7t3fyg/cL/5VZIPno75
KB3FxPtGGUxtfrVUhEg+65McysIxEVJ+NkraIzH8799pYvW09Fe1R9KUAWrYv8YS
LBChQ6YIwCG4zcQDUWmMciHkU3+b5acFdGHGN4FNJJizdfrIt7iaAykqLbrIETXF
NBiG2DPZ85ISvw20BIcMBO7MdiGz8T5PIP83VkDOaWpKDPjVM55PtES9h0E8BCTN
O9CdXRgZXyXe8PfQLAcLPHxtNpeN1j01PSlruZ09KFLEhWCBsntLT8lDgluHi7f1
S9H1t8R5xEQSgfNZhrDNIvB3XNDaz1rvhyViz2wpOWsrDRkGu9dO4pBxBz6DxaNh
Ov2mTYPxHJJznfNhf8bwUB3/B9TOAARbkY/wikNW3jm7eMUlMTJ9gDvdwzcwaP7U
RxvJkxTmpe8f7mYcBvt2zSvNCEkdA2FZgPUXQqfccvv5Ayhuwa19jNFKQkAHxj/n
POs0xbOvTUynBDas7vOasOppOPmE2Ir1ZqFVixdaGQhTFWPScJIA/kEo4gnoR3gN
ZHeHCSE3Ze4V7WJ/pwTdgoXP+GgbDrBeHOjnPRp4obESPdJEAYQAxaSVz5tvWx3z
qV+xmWT67ECLG5aUt2QrrxrDuTbwTgdLVTDx6Eq1bOd3m0WXGNaYJcxuSchyLEN8
KuzbHNHkj1Pi8ehBRuVewBeGvQDch1gAIJaZzXTjX3xm3TL/WWhhJ6y9kAR8FHRw
2Nk3lvUld2b8nufSMudhuCdgn4ErtwNolIpaCVKxpgyQmUBsnUERXmqF+MxgZdtJ
XVvhTCnu6eMeRmKC9CIj+NaY5aMlSjMuBQyaHEhcIe/4YBczMigDgU36PsYgyUA/
7DdpXmDyoYTlDY7ztYPhCuiK7ubMNcDIsGRJSLrWljGe+iMlf/YdQYc6hUlGUAzA
lrNFeDQNVLMnvHCJpcYL+yNvMsxan+qC+sL0gH3ysiAl3eg+bZyS6V/Z74jTctIP
W9gOGZCqKRx4UdnbyOnAIVt+17faarOiTwuYx5NwbKKU/wr2UGkJqDz5WS2D9xxj
mTTb9XEk1QoILVMmFnqu79WAzIsb7WAjnmdqFGW4XiBvaOfHVq7ZT/NV0iMv1ECM
1RPocmB/BC4AQn7kupNu1IhOsb9wYPmOWjQT4mylaLDUrhQU3IUrEs5kn/pRChwV
jaWiU4tu8hV4EhYTqwIBDXTNtwN85BqzGVPP+eZqY+Quc3LVC1SXlo/TzJBihCKq
u11o21N32t3fETvLmxuKxXkQqUFq89o8ngGS0J14OfA2+wH+B23Ih24xqjEGBtki
BNgXyI53ecQWVNf+pe4mX0yL5V/iT/8jrduONtH7ctZIM/mcWGjUClEIQ+l56mnt
l896ZFe8DUSYTzbFaSZ0gU2sCcuMPlCrnG8VdYOlXhQe+5qniq0b6BLR4q0cTdGH
15DNh780KzioHe1lPnhy76olJM5nhzJlQJrJUX1v5kNn//q4+0Vf/6XYthcq08QQ
pCqkR+2l8aB0VAxvNHb8jAnMLIrBo+UiqJyo2xnRd1S6g6hXDEmGJ4GrbA5VdnjL
d9Ugb+sf9wlyv2XVz+eylPB3EbNWEYcaPVJCl/x44dngCh0lP5KPsk2bOHz2iF98
WkEH2i1cFwWOCamzmzRZj4BA7mlRUMvV5IzuSJom2Jg7UpT5IWCekshjOYBY7tZ/
tknz/nvgV6tbih4aoGroqXyBpV6ygl7CBXf6ssZ1C0j1QZypbwNUxnOjVGGqgXCw
QVgT46KIIs/gY/dMDnjGvLfsTIj/IjouLh+XqJjflY9gB/hIcUzmioS2jUSZ/HBW
mVyqUGfgQOYkgMhzxqy3ZX7yFdMotZGiq437a14M1P93sgv/R7S32SXm/8oCDEQA
MGYaDhp+y4Qp6qmb/w0KDIw44XQODos83s+oOlhc1VEc+Tx5/ra6+QlMm7Dtxv3i
GBCHIsk1Zf4z6/mF9xJq8d6Hf+SB1AKI3U3Lfd0jY4yCxKm86NXX6A6l+enFsNPj
AulIfpy28+tMz4vQcGo+AVVdSpte8eue7Waq4na2Nx8fDBh8Uyl+/Nh+KebNE+qH
Q5wh/aRNXDVHtHNWhBLKHhRDddsBKKhZih3L8ggKLf/LhgFDUTCIynzcMDvVoJpW
KcvRk6/6h27BkzyLKgdcjXzy1TDYujqeeV7OS59UeLdLY4//xso9bQNGp//vO+rA
Ecz9gMPQ45+3pSzalbjT6DOwNuZjCwpiwOY3YIcXcbhAkIpfb/NiJQtxvpSOXlxA
TfSjD/dKYBS+NcYCaUdw+kN+/3DG2an8YAyB6PiIo8ME2meMQVeDSa01U/Ap40M6
UWMKa5HbpK6okxoB1hG7s+IijYV/3nM5ollWvusnnnlmic8QRsWf3Lng2KemqmCH
zhYfG3SyboFcpM2dmrMXMlNxuzgcXYY+Tpn7hruBnvOIfcf9wGlY34xCHesvk7Rw
kmLFnkGPRbL1I9PjCokUpbbUYK3HMoY+rw80KycSYhkeRQzGzRA7zXyV66pXsDyr
4E72LCFF3zvrih6OvEFaiQITHl+EK9IvErb9BptSzDvYWFuHAGZkRtyL56kHYqmW
PUPD4LjaKkwiKI6k0Gr44xiBlZFK8z5lcZhl/k7B0vNSFxW3c/YgJEEv4gA216h+
w0gsrltSiocHYPecOoF6uqTGOCffFmV3GeSxdNXea3krZR9ySQlTxaKxflFAaU2s
6ulu76Gb/bzCSheob/ehgXvkvsLHm4/KSdB5MYbn5jeuRHu17gak157LiwQY4HQ/
/rbT2gOYqZ5wfYMngFEorp4hxDBW0OvYfw9pM1DeEGHR33jxm7em/ypGG5sbkWT0
Uf+TqkmPMBelD26CbTaFiw1YoEIexHFI/B9Isep9X1ZHkVASdXHAYxO3MO4a4v9T
H+ZeWO4auGSRapTeB/lo4/GHEhxI/0txiPnikURkFCnoNz6CIynT+b4YRkD0DRNS
tG7Ehem8P8+xA0hvlUUluxKv6LbVQoCd5R1Rx6UKBrFwGMgNWG6eBer/+vNf37KJ
ANVgzajD9mYaafw3oWdnCu5//CZ4Y6BqVsWwNnA6GR34IidvwAIAMbTcwtlunWrD
Ly4nTE+BgF7L51tema1RrW3U9Ha7vmbLqozCrtEGGj8JDdA+RsfvqL0evSXo2pOA
A8qnmpLPhOQOzEV6P4QtX142sIezmGpjuycYzWBXJVKu821TyjtOw0P46UBIrCmZ
MlB4CKFjUejKi6iftuI5kPh/dMXSxQlJQmdwwqhjUMNTdKUP3u6v4Q1dsppLNvlk
5zu2RcMwEZg622vnvL4mEGPciYve9QiKXmtS22olgPWJwm9nIRVeVnFNXorxtWCI
j8+5Rr9pkXLGTZEMD7U7dEe928uejU5gjpl9KzOiGcJFESF50XOODEdnSciWUQcm
pBjW6U7bYz5QBS7DecsG45SqgPkiO4v6GepfVgX22uTKcBLIwXgS3+On490grgAS
vT1+3BfUpnF3alufCFuYeihuz+QcBfvV3nl5LJ07NgqQdcKGsa6i1aoe3Ojx8nGk
GbYg1UjMaJxKTsy5FHCgXfQ3kNz7R9q0BefJNJoTXgrPyMH6TFiVnAMbNpLq9mYv
PDW3I410630tJwR7SFZHj7ZQI1/zo9e0oynL3K2k736lq2eWFuFF2JCchiNmFwoF
SyHOoj6zJ0OEdSLC4b2mOxfTrOMJd7zrUL3/mFyuMKyldGrRW2QOz+SqugEU5DiL
dKWRVl0rj8B/qsHDcvxa6KdoNix5QkisGTbeJiBBknlEJugZ1iNAzsdMG04bsqaX
0N273e068JHH1w/irFjXeZEG0NduWHvLFcxcO7eNI0K2Yil0FlFP0MnfyJZJcQ6d
7RcxIgshmY6SjP6BJlv1dbY2hf1gpo9oWcQM4jV30ZCjk5AHTArVHm51JBS7/qWz
5+WUq+SCRYL2LJzOurtnHsjZE2/4t0WqAecyLIvJ14mfbwHs+3mj4ereYOVmq7JP
a8JFYs67Pxa79t7mGu8+MqobqqGQj/hrJ1f2Y6QHrMrTNqH/NLJG+VtzVqq4g+1D
pnXKvRJFie/SsiWZ+e61nLvI5qpnsmxugCBqlcXlgMXKuLD93l8NV+Rf5nv2nGyz
YxnLzAFOY/ymMIiVvBrk89A0+RC7cIrhK/YUdBrGLlZtKkQRgM77/P+RkVs5b5/+
dl9wyeI8bwlQl+wJ5sC7bujyfh1aOLDR6q5Jk65NjsCiDIFEYEBBs9T271FVFUvh
jlC5QPcOBz1WgfHMsOs9IdZMRI7fWdcT1fOZImIwXQFujroUU0BhzF/15cDdi+Tp
sIlmyONNeOHuX6nYGh03xssZ9SXnyZLfvjPMq9A8S1bSepWNzw2wuh4BmO4W9MQC
O0i4hl9mgD4JW4AfeEnzRXhYLqqe7ahBLKmlNLn0pHrrrQiaczyw6JH/+7Wfdzia
Hph/BiGj3NFGRgz7v6Y6f6szQspAtPHFomvHGKTJPVhAAIZ9YMvm3q7mMbXaQwSj
FFVwgUSw8ScMfVwEjSbVL7fft09FbC31wnrKSr8jluH6iLUGR9tnQlGEnUzIwSRT
Hgj2O6hd9wilnCeQAAT764ll7OibdYxHJwa19JRDEsOOPkX5UKZHX43gH7j5X1PS
Yrcm1XAictD/7IedZBxALcdju+UDxq5pYyzgEAd6HngAxjcBSEJUg+augFeiyv9P
V75BoEojxGUkofqp8YjkPnZpHZVzq+SwHM/Do5b9LICUyXNdOduFDydP6IlhxFjK
paaaaxBnmQURTFnf/I9V27Pv2XkeZW4WYTRE3rFFjlmESgFhtqPYgt6jbzX59DtP
4UkK4udaPa/+ATsatcRvwe8HAJ6Ohm57xBgXYZeMMGUfxHlV/MQkYkI/d+M58+je
smO8wg3Ssu5SQ2x9bYH0XQTCqacu0J9MrcZhAV7NJf2g2Tva+HWEvXOlNqw2yL0v
AaMFVTb10aUWLEGESrOL+LbYg8r2GfgTQFy6gNKsvt0bArh0TQBSMg6ULqcXSbfz
NlfdEtOD1lhOa3xqvsFEKu6rM4MDYIVRSu9Yu9JGnKNhcFHic4NVf2Bd4veeLJ19
C9fWpWNBtScwEbg4QrNLFxjDTTdUm0fMojjvOlkSezJgHEkWHHWVtKy7rEDCLvkn
lvo84pHfZzIzAOScxYLUxu0EoYW52GDQ5RtgvZTFI23Rv5Z01yrI0vp+LUkmgvum
cKS7K2ujiHqH7AWkGwqiChT44DfCof2P5VazrpLh8hF2oXy6BLvn07Naykx7zmeq
r2tiVoFdml6ZQGDOsjtre07d/0Wyi03J7rB2ZAxPkaq1f10ZifzRY0zYNd2JIumL
z5GCS60fAzVBP0qDBNpuay58VF8XOHVoAfpQF4Rf8CiLfjZGPvm/jztsJt/a2hJy
2O0ylqOmWftpyBzKDI+BpTpHP8g/EQ6+cVAxEpkRIJ+nXhnOa7y5nL44/7Kckcc+
uxm4XMTYUupfnu3LbB2lQNecg1Sxc6LHeYeaMg/nwV7deHX4QpcFePw6tza6H0om
i1GwDPvZTUJQWmjbV4BJp5kUXnlSMhTEEBL4kePt6WNnWd9hgQ9N41t/EEmS2GXc
kLqNsCWQ0Ol+kqGPSqAuyEAYBzZ7ltE0WN/RnM6BQqhDP2ciHtc6NeNJdZ/pJGKM
4gUj9pZKRwV2r73A2N3g2JaSIZR8GocqflFYeOZt+/yqyTnEwMZkOwcWghpDgpag
ZsK4djx7DFBCgVlNpxl/PXTyj+bcqgir7YLUtktcrvWmXLKI9UjWN9QINoHK7MnL
Zz5R/p5scPGboLeqjR/QXIu1XB7bDmWCpX4F1SFuHGQd7WFnKkc6ip4ancqxBnXF
VVSZ+lfyPU3ND8h77Vbi22vxrAh42Tc2Y9xdFAO1/1MghyiMNX5NSYMJrfS43VL4
r1lfI8RV09EbCtlb1xVLJXkfdKitI3pczpeB8+VGHmBQyXqlWqLvqW4gvTP9VGCe
YUpl7DFSETno5mGsLlf2TI1wTqX1AaejB+kVclzbiijuhj3QjD/qKbstDi/NJQdz
Q7nTnuJIeziDNzEAexalUFUWe6UP2Lts2lbUuWSlIGgDU1cRQCxxxClFfxvUTx35
zy+JxaV03OVQG94EN91/Y9B3Ps4nYteBgLNDPWUHq4crYozYukiN0zeo51P5iv+c
p9zXjpcx9uJXyc2uSvzniSzebA/EdY+miKQYW9xwms23IC6NWllHlNzoSOFOzEQw
w3rkavlKNABjYIaF8ModJBc0xBudO5mAUrJYD7aDpGORYgTn7AS56amv4eDVsVsi
AZH2Gka+puIIi9aJcR8o4GLva0rGQK9InBfn5RnHYuCqXF7c/OXtVkNyHx5b7/Oi
J1t7exUXihEIm5tk7UPM23mREQZjzHKaxw9qiOd/HcmnyHXYHHk/1ZAc2LNHOgoh
Ogl1ViI4hoBQ0FWo2cuN5gryHh4+SZAVFA1YlJJSo5s6YsaBS7Fvp5TzQ/g9f+gD
YphGV+4dUV/+zSzavXRvDoVTYDN3Swn4pUM/d06wFISodcDLgqRQ7o0Tzm3oa0wi
3t+FVn6ERbLMELMDj1mYp9CNO8fxMRYW8bd/TAUt5kMNdD8K+gBYUNs/90ksJZIu
+W0eJCPvqySGCo4ZNlsFLseuHbkMSltAf6FyGHl/kcBAOrV2WfNGgLk361VeJhAA
nWhmxMb7nNpV8JkhEJGC0AGNKIM4Ku1GXn9wCWv+UcklPD2g6iG6m9cqqlwR2fOI
nmybZS67pWtnaeYMhnCB8Z2v1AteuzefyUoLtE+O2gx35gphowjHE2PzRyzn3dIL
Fnvf1St88+WygQxg7bgx1qtQY2Dmyu49PVBrkfetlD7bBhSavuHiE48KIcdE87jr
VuJ9niLX+Su7dV+L50KBkwc8T0yFQfY1fV8BmoNSLQAZfdsJzUvTRtVYMmNjiLfS
vrGt5gV1D691UZhZFKpPbInLBWQDS3Adg2f7aKrzhyCZvDlkHtky0o4YAmf5MyX+
5fSp9EZLmOzKvOcTZ7Lv+dT3PZMHs9wqx9guP4QMb/P7gRDvxtrgiuz2Kyob+Qzp
25xZeNNvMz4IDsGvZ4QLeafbIlsBcvrp87Fx+junrwiQaQLkluWagoSQmGK/WTYH
Zi7Nr5eD/g7mVoQe/ON+KgDVVdPImQSEFDSvoDqfG9qFQ1qg9E/XddAH6DN+42Z9
imRX+xzYa1R1sk7ra3cPdgGgDfiIITI7CFSY/HMjDXyyMVGRYbzIz1K5XHVXnDBD
lrzlKCC903am3/f8jivkBikAlmZ7tmOohZmmhvzJAQ37KxE5u1R3Zp47rFYoRB7C
VJJTDFwbpCTGimyuniiLc3q1oWGYNU7lEe/G3bxcdsK0iAykO9g23tgnlthEtJlE
4SqZfGipLiX0hXNk3+Gykd5Hda8rexFAzF1+TZxa4cwC19+m9FciEUndEotnLgyl
eL3FaxAFjgK+nzfpQw3Bd4jxlL9f30a5tsG3VggapSDxDVomTh6xWpGXqYowp60Q
4tKO+X3iYtZg7ItU4nOZTDY8TnNrU4A0ZS4lPGXxZ5S0YHNJdhx4znhPHtJSjc7/
PIHIJFnYDTNvqO+FajOOJxgH3VuhUo/i1zjKsQcCNWupjhjoAWJPMCEmuHL5B+is
QBHcBjSiXFi6QhB/eaV7XocfB6Sd9zMyh7IYJJxflcQIk9T3tLk2cTS/D2/cTPYh
URUU0jsTWjTG7h3U8prXoKIhKasdrYoJgYPBerM2RAXqZ+lQ3BQ4Re9DOghfj0Pu
rwat6bdpFvRi8abFDb+BItAG1ZK2xG/EP/mOu+4lKGssXxfJ80gGLUtemlrowZ/H
D3L4a+yltvPEQnUs4CWLoEDtBWHdpJy0gP6rYIjZM9vc43/g4TsxwwYSJzFxRAn7
frKRqTeB+YuIkw+hcywqbhBeMplorUWuIp5/HBfxFOGZofUeVrtRYSPGKzqK4Jlo
McWMsMQCkevspetDLSmz9IFb3Sb+vSnNPYIXvTSB2KtZ0u+1SyCipDAi3+XTXdvJ
LaANt6IXk0sadNqJCGOVDjt0QCwOeDuWz20utSyQZo7EjAAYoAYBc8uKiqjAioIU
Ewics2yguwSIeJAJY8teFtXMpgj3eUiNcNPDwoDYK0N0kLZ9wzXQSOyzPus/FPWT
dlBA+vLwlvtaUimMmYfMR0Nxb8Iabrt4A9seseU1q/9y5bGNjMdBtlXq4E5xLWyf
3pFzp8Tt2kw1CIDMgpqiijfZo1yVim+fdM/hrTpFgjIT//kxGa34UGq1LAub7GnX
17kH+tc+z1L5RgYD+yIPzjqQP/kdCd7IKhhLDB/uRm4RS19nqWivJy6bB4aCZZtS
0gKSAyg2istKjFugdqXbDAIOpnnxZitVlCljSL3cu03vuZYgzhLKXYXLl7jeBPid
UUTzQuMtmppQ1AkiNJ3s1QYOfb9/NCwIYRZ+OPRI2tUKHQKriwto6QMZ8fQvGct0
YkgBVxKsV9y9YkgpzQRvcB2QYaduATauzcTuZbpNRVk5RJbn0kkhl6ZMKyjxPwZs
LSJu5GHRFsphH+ZkJCKji1HZpQe79Osxs6g7xQ18usvkbG2ubeKOOYDyvl9SJWjG
z9DRy6fkGbqyROO9M6YYyB0Wvhn73gbKTcpAy+2DN1yjqzOVnoPTrcPzqOukByX7
k/ske9QkNSOfGKsMsfHIOpuPUazS4J/IBpncYz4NPuCQ8hMSYKFSfnjtzftdwd0y
XL+CqrNhWrXATRY8aX+niPMjxHDXZbXt91T3fLmr6yREkdiVfwM/Kwd2/aQb3+9H
WjKdR5fpnJVM9xb/VlDJYk3O35OUhaH0wpIIaSlzobqTP5fc65V2fC4O3RRIMuGX
ucVv4TpNBcVZOqeXhJcTh01vCNKHXopqTg9mcqGSFr/Np+EzmZqlEb29bA1cnpKD
0dNr1acW5PAnAPvrwWDO+iWamFhocWFSVEGUObgFQ/bp6ZlPPA7d8CGiHKejcZWy
LFqpzkj1IOq19Rm5cm73RJY17FmJr5vaTSHaBNB85JIRMDgGaxEfZKJirSitesnF
IZQbdQKhYooWngaGLJI6JiJl2e8f7b/L4riULQ6+tJgOlf1t0DLd/VzeSIcEs1Er
p4ICQDFrOe7L3Gd/h097VDuabIq//yR82A8e5EulNfXRGeDxtjmvq44fXcjN2p+e
HGavCm3Bz6fqQiMVX/z6DURV06uA42GIChGxp+w4JK3oHuGCYv7DbOV4rWGMg8KG
3o56NwAN4e+bY1BRgqOBqLMd6H6nN6fGV5MRWXQoGykKCzkJxgYK2ttto4FNR8Bq
lh7BXhzVbkEndjk4/am0OycuJcBLnJqixqrlpUEE9sv6OIEpO4D53emkysrvsvQv
ipydgVQW8iExUNfUj9H5ydPLpHMNhb42YKIZrNpEcLXsd+i6KZB6702BR+0mNwcj
qW3agvAXyLPIlxEbQdVIq9XAY8LINM2fQxXRTAONVPUaLm5Y8dx38i52zKjpQJ3S
xH3NJyCv2QHQdxHNapWKDjCF1LLLHCfKpn1JNoOxBzv5Xvs0lF0zDnGd+UPw11Rl
mcJkEpnVl6VotR5/fauIl7p1SmOw51BXszkIdfN/TkJ/ZHfP6Awq8JpejGxg5WzE
VcsaLKQ5PNgzxW77UvL+E03JHj7gNHvY/E+xa3ufh16F1j4Vj+d6/775ldB7lO1f
88Vopp/8JTIilbMI8OcdWJ/EReC9Eg+n6WYGskPr2jk2E0BoK4mTMv5RlXKalhT2
w9LbdQv6LqtP+MeZ/i6RjS8sAZETOSiYKKwiWFP46bfmuC1abap/3A6alUZnyWq4
LZ8xU6ua98GlZGNLjqU5z+64komqICt38QfZdw9FxfBdUKyFN3HO3ICSEWzhWhjd
ykkEE93u+YzHr3EgZ8CchPPQ9GGqwm2eMxoYRGCPt9IXJU6jItNT2acdsKetemnA
xtye2apdoU24gxwgtDzrQAZpB24GoPhkZpNbh6VXxzFyunKCvh4Ekd7Bg4VuEdr8
PeBRzBubPBVa+c7ovDZVIIcy73M1x5+8WuaokhouXV6wdPyqrkoJqG4zW3qB4iWa
omKisFal+1j1iQOYyR/TlLEwiKFQr9MqCAePB1NZiHgcxJ59IrCHbhpM/7DiT/l7
XZ8GuyP9f/Gs+nQrtnbEDd8/bMNLcdjcNMGYSbakmzPQK5kJukIo7YM6B7RQCJID
mZmomNnS53c2Sfxn5z61h9SW9hkqED/QPLMvUuH1EeaBAYxWCxYwc9sPQopn6nY3
wbCISNLHvjAp2ZndtCPB6SOUjGx1ekWc0DV3OD5n+AfgPS9BnTucSxP9tQCv5Cfa
R5oKR8zcSrpsqwvvPtZBCIuZLeI5OGayKbCbh3nSD/Qgr42zfE5G019of5JeFZwG
v1ZjjB9qO6GhfCBOogQ7U8Sdn/0bBW6WlrtxIFrbt3U5bx+Eb2pnfimeQXYghFwV
YQ3J30aJNidPGa8QbBo/0oqUzKolh7pHyLZgpT4rb+9DgC8esdtLcInr0U4F3ktc
D9wSNA2vMXPshaI8wjAP0Y0i7ed6XEVXqB8dRdyIE327V9mK095VMPQCNO7lQHjb
xxymg7XeTJCspIH7vNvqFyIsr3dDFcU9bRIGn4xeymdDPsy29huGVAD6ESk5wnTW
5cU6zdktxdw7aZEOMfAW3Q1IQCmPDeb5JAkoTui6fpqWTs9MpFDUcEsaBmC7x6zO
W3LkKljSz053Q0MUJZ8Zuc54GH/DgdPxtBJQoalGJ6RmoyjP+9KAB6Mdxo2njtY6
j84s+GW3fKDVfgUaiMPN7Az4LwwTXSLfjuv2wd/lH8Ehq6KqcAqfrqXLmW+YfZSf
94dwIoGjIcVguEWRb+Unja2jSsx1vkX4wBpdnBJsXrArwPQ3Ni57a76g6mRpC353
jnyQcHbeI9bH93sIbPapHKal8nqUPiH81WHFP2M/BddiWLBcBLjgkBgq1OPFBVLq
1sr/AA8RLcj6rhnAnRVrgg+wBv9WANmWMyyntx0zwG8ZOho9LGsZoieGiQhL9wwh
+giMB+gn1LH4R+fdNDairL1Zw/MFkVxINtILl5dg94vK+uYqJVXbyYYF0afBaBRp
wTt8FW1ftQLbpxdSdBfqiEDb7b3Wj7uXh+FtsdtFp5SoJuTKUY9l9pBBAdeqxxmS
Cq9QhVVIfhDRToyEeEoAGgTP3f3qkS74a9KPvsxrGJ4PKewpSx53tA78pstfoiVz
GDxDS/ciWNIbQl6s/N1w5fyogaOsnwCmGo5MsFCHsIERR1nuE6W8rui40AVoke8i
V4z1jpefnu9vAssB1KxtA1mSTeA2emrz9V+fiAOxnizfBKO159a68tjVjJhDgCSt
ozeXRLsVPWncGXmPfenOjDPabD1ukXmF5Ghke62huFAVem554qhKpE/vtpS83j1y
+O5D0NJL+G4S6uHKt2zfxi4wsIAlbSLsO1GFhpV2zJnKyywJsuhh5G6sApNQfgRI
ENHfYUfQ/o180CATqIj6qAUxCt1cSSv8YsoPl4CJhyiPWjcg9OwmpTZFGj2lqRTs
UacABlfq6UzjMllQ9RacCYLkpIsI07GQIxjI9vuh7nkNnLnwAZ6IQedm9jA92cjl
JFa87AaB48N9343vKXwwqI68K4zoxaFNxdQDyGl314AY7KV6SegX/cPhZDGEtoSx
RAtRG0CQTkzVmoc+5WtAQNnIZfK0ePUqdUP+jKbNbtkUzUUrbdWnIDb/dF2w+8Jk
MemjTjKf0Ok6coionhZjPKSnpdN+KO/lfwoMnvljSbKKyI7pv/P8U+k8VLxcfNLw
tt/azrcyAlMNZJUG2qJNxIpq1D7AVzos+Wn24w2iPXd0flFr0z9FDhRd/OK4i/a2
NSNeqIgK/8Z4cDm2jhQ8D3Wp/XUmt8ck29N/D2Z5gnWGSNrBLKLdxM1/lZ3U08oj
IxDWUemJqs5RARXTg0i71NwiB5WBeyPZiV+RjvliRfWrV2SXbExlm8zzin0OZRDo
9NGGqN6tryMvuARgVhlHgXCoxiB/kp5V8PWZfN36H7dGx1r475f4gPeBw7im28FO
HFxANh/cskV0CCM7TQySMxXKq4ZTVNdyPVXw6gJXDtAfVdxay3kWjZPZYCsxT+NR
kG0mdAzIcV36SWcBrF6u8AbddfBp/0aL9MfhfZRdmFbah6sWd60ZIV6pdHZNs7X/
FwigPKS8I5LlunUJt9WLE+y3PENwXSed8ECS4wb2GCxsqJNcMtPnVXq/ZazGWbYo
smx8A4tYwPd2Bk4cekwop+NN1ZVg60pIO2rORkIBdwGTJuebswPcHnogScwwqjuQ
hMs48X228rVoFBb6xnM8KO8mBGONZwBGwXlpyLvC7ynjUbhFwuf/NEMk5ekrC30j
fI+0daml6BdrsMAipB6cEYGVC/hqMNMpFyUzrdICnaav629dkQ/m4+BokLwW5qqd
B6E5k6sau1pHPveXuDtk8/oqinD/m95vz7StHWEP/ZnmzJk9lNOrezQ04/ixdPEV
ouewMIHUiexT8vvexnVWwIPwZ2TDkDKoF0/tbK1QGoIF+OuPJD1pWB1jxiZG94N8
+ojbsKKJkb1DlWq4+n7OaJSFjXOQgn6aKHk2DBPpp614xRE9lN7A7Yj/YCR9SWWd
SUXWquJIlfp/6DGYWj57IcAbtZJZHdI7hUhMbK/ORsUCDZB6Cx4F8M/Pdk6T3IDn
ysmB8BmZXw8Sk/w3KfG/7+0CdmSAYnJj+upR1I+4swSEBtdv8zv9pqZenutIlHPb
YOvq2oDUpe5HAvVVDsSX0x0F2F+2nXUPTI7xfmPC4k4Bro4RK6ybPD8iiwpXxAF7
DvEKT3SFFahjmPnBn3TJb1/sZUUO66J5rQfGf3JnLbB54mpvlcSOKXsM4YUnnn6h
f4Pb5WQTd/VOhs1eETgjuBjTbx4IFA3rvDGuhh8ggvCA/cCrAyJg67HnqRZT63pm
S8d/pMzSs/W+oeay7M8bjnSyemwMxzBjr0/Z1YlGPvXXdtL00vy15+Fg+18R0RWk
hSfZtDa2ajQCjlXjZ0nZw9FZUp06Rnx5DYOsK55KHDpbqFgpknsgYMpSlNC9Wr8n
2z0tDZDCZazzACuEf99vRmUfKFB5//3bhgi6C5IHvP8fG3WvyiYUsTbFAp5UN1cH
sYfPAk3Wv8gEBW/Fu0kgOk3sH3UxjWSbjSh/k3RrTIApVNMEQffxbK85ljq8VfgF
chdlkZBMlAWeEv1hwxC+tNYJFaogkpHSd2l5mdjDTaz5M8KZ1RH5sMK+4g+PZ5Nb
lB7RgWZS9sUQV7C3MUHBSvaOecdsEqR6QrALijOAY1kh4lzaK9mIFQK0E7yTdsFZ
LPBr4n57nGu6H8WYNV815elGjkPE1paAw6CX6LwvXafFC5N/pyIZ2Xeytes64ZIe
jltyDMgbgG0w9jyvMYwzSSSO55Sa2re9O7XvVBC8kqsFuu8kSFdkY9eoCug6FNcM
PIDPd38j1AYO7HZSr9eCd8Q5BESR6VHRcaE+zrnUHMZIwNdpmGVSAj7lzvI/M9/j
CG2ofrhpRgSLBh4XdEZT0DYndi2lnVFvQFln78CDYr8UsZ+vG5q208ootG5dQU5k
vK9Fd/fsu1EuPsiEvfsJOn6oRh632FMdSQRmgAFnNZfws7B8rili5ZA2pK2ipVvb
dMGtaIAF8wWcTCvc2gQx5INmP2ktfRI+ZEYFHDc5Ae+eU4IkgV+9Cr5A0JXmpLtv
QV51sBeIrxo3LJWoAIkB2SRnNGtouuUYrdgXPeaLN+escpD+fa2ahKYv7coW6qvd
SmAH1p0mlls65ALPq7cBZScBH2Ue/LPQbfnqmX9v298Ng5Vnpd+CR/NvKtw5L2MS
RXPw3ZLMun+5BpNitGR2i6i4mHFwu6NL5tFURXk196fpFELhvBkTkPpSAAAM/c1U
YlQe0++rwmh36xcrXTP/Aq3XUSHdcfkuF5P3QWNL/WyJ+P3lXH2n8pF4ew+c2gpA
hWCNyU7JfMwE9BBFBw8x/TD2Fp4sGiwfKvOoVqRmja6K7aSGbw+2xBadumd0KzUk
MKYFplqg55EcZ6ji0ep7qoJSxIudKTEh3KRSoNIjV5W5B3h9+y48TimhKi0p9ZoB
68UlFIfUNfpxw4MYX1x9NejfPVpy0+r5C1yH0nblfH5lluDK3AxjrKFsABb6lGPp
EySPgN4oBA3XYZ+ShAlklrGhvS4797lGIQ6CBCt+84dSXPt2nl4fF/wdZ+z8T/3J
o+I2TJPHYwZVTmC4oCmHlpRdhyc2/DtF8KXQHUCl8y+WG81/gmCpWte8dDS9HXS5
Uuz8zrhJSI1DMTBdnKLyxIg/GTeGh506cfUgXu4Y1yOskm5khwZ4njKynwBj8/zT
CbyXca1zjD35gvxSKXplKl91R3tDjQoSqExbt4BylXaYxkJk6l7qsgVIE6zBcPDa
2v8d+iqEPec/R+Ra+BcHyG3WLItG0odQbetSJJXppFplLwhRKd3nzPPapqUKXyto
MgnFykc+7cK9qTJ3BjlGT+lRvqwXQXKb/6+EBjVAsA3aTv+j6RnlGaD/Ra3yErXU
CTMSj2clvMhuGzioPia0FuvJ7sROJsbqodH0YqgLmanpEFLmr0S3Xa3SdJNgM1MT
TK47lbEkm3d2Cpapmrzf0qoZxNVf9CWjNWguWPTdK14m7uDcRlq0F8k1RP40w0KJ
lA1GB75zSXLmRqhGNtbHUGPcYf3RcK2wvVnyrIyEgrkTNT8KA7dXIsJi7h7aYx9Z
Oldye9e/FbiGwIzzf3ZNPIqIgEY0Tib9NMURR8zI55UHUzjhh+3GTUjXXKR2IoJn
6ITtsh0FxkDGO16UnKK4Te3M0pKk0UJlZ1aR3xie3xMEz/k3CCES0IbklOOcI6RY
uts+VQCepNUkYIbHcGdVE1qr2FjS0UjsSMAD0NmgUGg0NTCcpmydsSxrBUb5HCvB
1QRIlPV4UD8ZlFmA3MvKnZ64yp/Gm2ZkrKM6r6BRJ2+7mzQCopViWi9FM+ErkOSB
Glzk5jruFU0CuRGGAYbIiamLZPbVKsk1oqpF28h9OGo+dUChTgugNIGEZLmUM7lQ
BZI41Qh0nt/XOoP26eOZCWI8S2baxaPHQatDYcDyFWZHfslCWrxDD1KJsaydZXSZ
/vmQK3bvaS314OVytqJiY7p3/D/URa/muGih52bFf6s55poziP8ZNHLG80Htx47o
rZKZ16p+r+YJLH3cn1N/igL9TveGKoQY1XA2SNBzEOmn9ob58/IglFdPyrmw3G3t
lAQkUV3cGA3piucvxkLKE6U+qWb4XnTVLPQTLCCXcQb1xnITqvOqst/Wx3abG+RW
VA1+dR9c9G8J2RsibkmmyFe0ztrzMr58HL9Y6hu8fjT6lPdFkSlY6nFrdkfvkuQj
97arp3arFEAuJO3K3I0Vbmu5hRskQHE/v2jP4vSvGQmHE1WaP+HjOAm0cKrn9NW8
50/KEW9At+LPustOQuW9ZiMSLwnRT4o/Sk/gKfSYifW80CPVr/rf7whH6Ui1PPzk
XjuvHwrI6tNDXr7cTkZ2xFa2m/zef4HPM04YF7PO4fqmNj4MeyhLQx03XKL8fb4P
wKsbE7ZA8A+V4DnPdNM+RquUnOSC/x+GtB1LYk4KHVteZhbXUFYqKFhkXYnB4J1H
/IVwa+z+vY7NN1c5HUPmLjyvSvqD8JXbSSdqBMxWLbvabrqOzXu4/bltx/D023Ck
4gF/j3wmRHd82MJZa6mx0zr3muoMG5x4WQg1TkME5QPcsU7eiEz0EH35qLjmNmP3
TGH8q3woe1C2oys7JkCIijkLMUD2SIUPYcvbcxDRszzFe0RDlH3m9+RpV6NHYpwO
nUahwD95OHbOhnu8sgPBkZ4V4mPZKgFGZquABy2JW25GFYZwxN+KMe5yhCvMgn4S
6C6SvdVJVTJ5uQ/xsUE9It8BZJZL+faZP0XCqxJDyWn2TvQF3kqIJopwNC3R9bk8
SNJfbzsBGzFww6dxsGD4tNkdrnYjrCXv1lg0/PdtuLQTGOGOlgJMl5S7YY/fZj96
cRYFdD5WN39bXIRq+C/AWnyJk9V8OTrEOTjrKZlODjL2IznnMVr4xNkiShGIV0zA
SzrXMK45uMTnFr0lUqi4f2ztOwpvUV092GRbBwqxq5TXyLyLh08p2yJeNdS7leua
JYo02sh889JlwPFCvMOu0cxvEPmNWi8wpVxs89n3TZvDOx/Gqxm1oYboQlwPgfZ+
HFtkRltPEBItvvAjP+X1LW8bBuaof0I9xbq8WLoatFXBUFfZ0or3NXUeS7b6p1yJ
ERq6i/oUarJG/NdXTkHnKNuXXMPoukJigHm8xfCld9Kt9rA7lV0ENfKbNMEeseHl
UJpFF6tk513n4HZSOpuCokChd3I+k/HwBcHrnx95l0Se9QXLvK2cZ5/xN6+S11Fe
vB2Z9ersuFBLioKD1yZohqm+0p6o917AEeJGrgRhwWZOSOKspXnScDF2E5GRq82R
NGZeDdAJjeXMaAJdpv0ewwvq6Z0uQJ8P1jRt5unKyVr2SqcvAiJ3hdt9kpan7jDu
+PU0xMqFiK4fn7MLH8hT2gJeLxt7IsidNGMKAfN8MuFNWKeYW+EvLebpL+jr27eP
TEEI2tdUPnu2qVHMsIgZMmd4YwOEfJXJQesR5WFiXIdNKo7onac18Qw8mP33AOcN
SVeMyJoVqForsj1aNsA5URlfQxesaHRl5/pt5tw/CiezPenH13MbcENOfwT0i+p8
nn2jYZ0I1DPdNqWcsmGN37vluHRG7hjRK40x/7Tsyf1tTPgIG4U+RVDu/vIasgfz
2Zkkb6qUlPx0rz9feLjNWNWMY7lcMPqx3hYIFypTPOtq0+GSUwnrF9Hn8xI1nvS9
Xmc6emhEj9Xsqr6HfcTRm8c27kbsUZHQbLC4cZxQJUU8CTDVAYAMSmmqRlrNXOl+
lVr4S8n3h417yc5CQfH+E3l4ooCZ+e7srX5/tEjR0WLTgWdO1501HrmfgMsNc/HE
21nw2FE8ZiQqUxNtSvmG7Bw01tz6V37OhF0Xe5pGIPTWHuY9GVBBNJ4Ufn8s9SCa
gbIsqpUMuMcZjMwBk6I2fxEeX9qgnwr/WpDCHtszjNERa9LJBV+0rcqnZN7u2mZ8
tyEDBHmpwiYedMwNI7ymbGlrcnD5ZdJAfyJgSbv1cHf3YFK/aG9mwIVmq/WdH5mw
d/68yv16pcdAvc0RpQZDQvDHUIR0ZCqyF5Ui7jtlQuMTn7nO3wAFeM0Kh5N0UitI
EMyHRH/stHYEaY8TaNG5MbrsdvWnTW+odfVExSiYbRh0kSgBJRQX8Fe2Du0cejsk
3Xpgt7P+Ub52AvCZ6pvI3HGGEZOrofLDtFno5bWxp+na+7B08wxMGpMn8OPoKny3
6LjiMceVtSTCa6FRQjUC8uSrNSz60+QTemDJwP2cIDM8DxhbzuRUS8V3syuYHym8
5SEg6L23ml6hhasgh1lfILJb+Ii63/F3Ck1b2ubeqCHhzcQr+1ZfAGYwswIvW5de
g4pBl2uoCDzAIgmrw+KlLwt9cx0AdlrvUpF3Iht8Dust4T2T9aBeUxzmCBqidc0a
ffd5jovy0SuJwRuOKXjarEYR99cOBWPTwtz/J8DTZr72uIE4oZ6QBarPnJRKHUCH
Aoe+EGiT5KKSl2PzyJ+AVkPXBMz5qmqEPnWAIYlCdHdkM/WP7HEFssoKJyujH5nn
bkUmlEmIclno9cPzVN3Y9/TgtNVToL5MLMi06SD6uOlypsfJkhKmM37c4I1h2kGo
PC3Z62sOn50iWJeyc64rsipvOI47GSlpUobEP6qVBUF4gaLrOakC+6/cenKSSAyw
Tpv1A4m+RyNCqDCxNGieTarCmWt+3OXtbdWwRLZqHkIYgS4RuQ+Q47JpaguUOb9y
p6GlLQMya+UyKkZkesEvW5921DN9mlUz3eOf9Zuy7nKPajjs1QfOMIWWnP2aEwtw
GABu3aARh4hwzxwv452SI6/iOhJyTTfPnME80cgf7+K/6XIq17QeIbTR0gs5qlXu
6ZRODK8z60yah2022zk6kOr+8vyrwwIHgvFDeQbHEpjzUIYpMStG8qC6wbZKPybn
cNLOGsfBSlrZAhBxZz8rzG62kMkoxpiee/PWnLH6026SzS28HsW3Njpw4V8erajA
Il9JaOUvnfzA1h2sK/rh8nkrXeEUyRus+7A8Td0a13Y9RllEl7fr6T6dGlFruNyD
/5ElBrg3ulorY0Zyn76DcfYP0NvQ9pIWFVymZ8Gvjq8IgGkFznVGh53s8lmZp0pd
NnL/Wn2Y+bLYT1tmBYyAQghWvC3S+3zk/6Qpw3cxwjYgcWuG3us95IfRw79yJvXe
7NI/0evo7exPGc1Pcc6gnBiN3kytc7NPCeCPOx93SL+97WHB128vmFzei6nY9l14
ddWPcPz0fZcdUM0hMJQ1VOirHxlles8A0AedNuX6NNqd3FOGoA2WckCKwg/uEMxZ
k3bRj0sSVdWl2eMPxcOctC8qyi6ZP1BeZ1nDs6MxUrX2mSGq0zPdSejDno4Yc+e7
Cjgk6pM7SrYtfRg6mmJFD/yLwho+i+K4U+F9CrgFLFh06sWb/kv2z+NxJTvBZiWz
MDc4oGQUl/wzpUbHfX7rfpuzgZezmXPdVC3aqalDCEF47ZnHStvQaoG4sK1xAj+s
RURFs9YeRFwZ1eZ0YAWhasT9sME47/1ylpGmIofFCZPGK46u3Ps7X9nGV6BmQ4bR
R0HSHheH0/0PqKwpCu7GU3PSbzXKHps64FDWg5mjiLZnMhWqgWzYWdjzzWheKyMd
Mp4PppNmRL4gMW/WcfwEV4Ns/rODCqZj9/dlGAWJI+iq/UCbjOlth9z4Kiu/vhDy
K1dEc0Q2ZM/WzVgYf2khIA5Vb2Uv84OgtiMXV7DLm3p7CpTc98lmJPJ505W8aRui
NtyhJfi+abursLR3/33Rk5chIm4Dqk1cxsw85iOyx4Sxr8MrdpFyXL2dYl/p010L
bT6KXZ4d6V/7NehkutO4zt9hClgR3rs0LkS+c6bDd+Inq3C/6q5DIODu9g3JbVCK
Q9lPkEgsNFdO9ithj/P3y8ysb6LK9MqDNWGHsZ1MO+MjZD6fP19sCGFPUATnwrbt
SZ2Lpqbc6eNZP0/DrTa/AjgDEq6+g9VXDWaCvK0sg/hKlWoJsxrVoPC9M7IwJ6x7
cgQQSJXuTHedGabceXbPlGrUeW/iQIMneBxCYfY1dT6Y8Tct9DuxD8k8oEKwDp8w
3MoReBZfB6W5zZBW7pWaq6ljnapO6THrrBdKoSO4ChnxuzOpeDQgkWLaMM/BszTp
iQVg570f0IahD1X+nu0E139bLGgtKNHG6N9tqz3iKlAZ6H+Z9xgeoLqoPUR1XY3f
Gls4e1KmU3piyxludzx+Gd8iZM6KxoCFUrygf4Or5E95o29uhD+vM4RADAFA0QvQ
ACtSIAWKYNz8q7wBy+sj1SWl8GF+i2MdhjqWexf7oWbkbOmXN/LcZSMYZpZaNN8j
JGdNJk80PG4bXywgsoNbq8tNd8+77OeRWFdVLUxu7RLb61M5y+h8pXblKfgn4woc
J+RuMlsgDIWzQlw5h+A99e8Cprf9ZnW7NPj5XYgAze7fk6A/8V9zNQttP0K4eNj9
KIJwFrfa5v6wU1za2qrEEG5svlWkeCponm4rHyFoP+hgmDyQKNy0eIe5snWzl2le
1P27Y57BZrVasFohA4JJ8aZ2GEEiSN9bLVtjrgxsBTlUfEERESxSLrmjRWMklQsU
R4oyZB8LKtUsiz4/b/KR1pwaZurfMegkLZy7b5y4vbnVpYMT0dxrmhQ6NuJMyPur
LKa+YQYGaYQFxN6s8Nf7K2wWQJP+TsHTKmNGiFmsEIdV0wBOypsjymFm2+GHrg3v
hY1IzZxJ8aw0EdMHaWIhtRBJ9PTc9oMIsX8NmbNH8T5E5vfcnjn8eWd4/iTSF3Vx
RX9CgR39AhLJuo63UmpNHfs11zM2NAcRo5lbqeQ3UweAbaZkUEF8SAtL5+jYGubA
1OGl+EqV3Cm74k4rwLmqGni0BCb01t0aPLUv3ABbnGK1U+ybJx3AcXNRv5kLkWBc
/o79f+vFQQKJUk/dC9pZTFXSKH6WZbmtuFCCFNh0MoG4AVM3LaHq4D6dc/mCp7X5
TOoBFRiG7yOWCZQd/0UH8dB1sshMoZQKaIlrsdA6McwPOh7pcp5l6WDCP6N2PYSu
SDQIjRC4B0VhzN9c3IeSABEDamKXiPRvKiCwS9YmfxS11VmaM6E8RRqr/8dQCw2+
h/LGs+NatVLmxsSteDNpcrQ4xg+NChMZbjaLEmJwYlUQjk0yDb7I4suuhyI8VG2l
5SaJt57Jw3Zxg/ntMR0i9Wtndd8WwxSDvvb25ul0GXcqSLg3HCBP5x6MLNqoDXMF
ZI0ZmL8j9RsKiWCsl8ZtrvbbctBEttL8Y53IcHqDVwb7Zqm3tRBrxW0xxuV+BQUg
F7SM+2PJehK6oWwT9OlCkp+thO8xrlXZ8ESBfQU4OJiWi6T1wLCyHkrSKG70vaeX
OcbngB7mYUEeH7eEp1s1AdxbOiAtHyWbRC/jRup4i7UYHCgcVrEJWg3wGQqSxOv9
lJ8aXm7Mu5pEBGV2D3ghW4zb9HOyZVA60m8xC+zuAezfG/346ayKTeV6mspsA3tq
/4xIx/clZD2KGds9Omw9gFyUpgkmCq1B46Sa85E1fQRB+Kb2LRKO8BHM7NrKw5/X
vlv9knnqEkuCQ0X0DObUXOQn2XxBEGPGi0fDkWb8Y2PPfqoTCZXlLowqztL6kV8m
S8YYpX+W4Mag9wfZUeaTUPID0BBqwuZrGEi1cxE0g8jqRwzsQY2JtHTC2S7Q0a9P
RH0PdS7IrLTMu/s8VqiqSeIKe1cdX86GSkkFTHkw0v0NAJ6xnP+DcQRNFW77IQLQ
3iupfrg0X2Gg44dHXPKR0rScfXCDmcIGpD7EMMH2iJyZBpR4GjKssdSf/C3CbO5m
1spi+HEOLLFCVp9E6OXbAAXmuzU/cNFBw6/lSBrolry74oaYALsV1jJIz0vqtN1D
INvD1wsFiAP/QODzyhEXjWO57a220S93fNoPOoUxDsd9PB4HsqrAAiAISdIqAHVU
cK74yqX5la0NU/mGq8opdugw/M+mQlwz5gsgGdrynOhFmOuBPeodnsPQ2EBYMMTW
SagZRDe3ZfeOPWx3tB6Aq5ezOC/BZmwHhK3tykQ2VtgtdwR1Wl2hd7Lus8okQhLI
va0Ghb0pSJCFcqO5oG1xuHb3m8MkrZIo1dbs3vwBG5DsWHal3ktaQ4rPuJwydpa6
Z5oDoAzsOk7UT2/0Id1d2G3EvxD1DybY0jBdbu3ppHLj0zZDGOVWKlCMGSmv7IpD
TxrjueC6oI+bFWrrVormfVDDy92xmys40Abl8tCWA/zZPFv8tLG5wRtaYl8AaRqS
W9ji1UB6hlks/1bg4y82Yq9AELYiX6u4IAMfLJpY1JxYLhIL4Ig58q4xuGx6QtbC
LKGuWb9BmqyjefPOIWfiF9WaYthHOkPOKCAep6hhJi8XES7oXoGS8jpsxWkaNyxJ
8clsUJRLsPNHPqPkGP/HNnqVo12ToNng1fD3ZKNAFHqinpfOEsZ1tI1ttGXq3Z+8
uqsXoVVsCdtYkwr5fQcYSpVm0Hsmwnc7KFMSkz4at1U9F12Gas2Fh0qrxNrmO7ba
iR0ChepI40WO9wy1o0x+DQVQr4KgQvG5IET4brBuYe3R/gAydh35ae0/+masHNCU
fijSCr7Oes5EE98YdLjoDkCQhtMg4F1Y++C2xckeda2xnsJmIuA7dlJlaSCXpcqn
igbD5TBbx1wuJ+D+I/DDSjN8j9xkgpwRVRnCfJqb+Uibs3zDDDZlm6IbmGm5C/hh
WWEHOBUzqNGb1FWweqqJNGmTvJzk1X28K2vHjkW6vTkhIf6VbgTHU1RPxQuG4l25
YqqfeXvdBnUAdp+c/ukDFrLfEx8JaJEGhTaDW47A2nC63MxcxgzaHHULOmZhdfB7
gLMZzWwu66F+mUmNwePaaSN565xYrI3TG13fdmAJ7IRwihmpW+gCz7TqyO+iAz4r
J/5hW4NB3nnzrFSVsJ9sDfWQfVXK0nIL95bI5aS9NX/K0i4BBiy1l4EgKDUsdJOX
fo5R7IlXC6GjIO7ftyUFnKsDX+/gdJ6GuawSJQnS2nffs+nUHNuQBYPprE+A+aSz
wtGSXUZoamPs3iPiMp7RGs+Tfpf1nlnoYJ/bnH4HuW3mdmOnzppyvv51mkGm7Cyo
H30h1QoEb387gPft96dTNDJipb+pZZL28okRVw9Y9sZR2XUifwDjPFseijbBT5Vj
7gvjJ8eh2XxMHLx5Gu0mMq8GDAiOGIhol0Td42AQ9ZvlSWkRpxraCWukqRrqzDE4
fLdgWLN+mjz958FmmERo+rfhIXX0iK5Q2sF2HErykb/FhL/IxvkOmvkNwls2prIC
dpxaUD3evJlS6O6RaBV00L4GbU65FJfKm1lYEL85fOIJFyOHwEM9jZ7zLZcoZPcH
uoKFih2gK8zlgArAdagMOS2l6s/rtK+2UGu9MhsXumkMg+vbROrOJwQNPX7F8emZ
jPV3CXgujE1jGmQtots3Vvmelen87fFYSIHvn1LhrLMfzlQ9sDMw8g0KSM6eaxQf
C/l0WgAYPvTZDaMGGKAqJe7FeXaZb5Itt7m60DWHhOAig7lgnTT6hFdAnI7aLB4S
iKt7PMOgaZCEFSNGY1BEPo7hbt6w3xHbwHZ+RQsZpuUAdVkYyjOhJZAbhXbWDvji
47MAkiLiJaZwJWKywITvHzeysZ+zqRqnOKJxl1cuqpOTvQ6zNG5jeYIeXfAlgu9K
+S3AsNjAD1yAK6zONa2vOy4DW4IZhGcw68CObfra4KmMioDCT6aNIZ108B/rxaDr
aoQW+jgPWCZ/Y4TZ2AoAX5j2wfKDOJTf3ak5x2Gu9WJFoKwrsmsxBBp5s36Es6du
62EhoyW9HCeMfm4YEhw8j/iNOSe1IUMIkxysHx0ip00bukm2jBLhE7TOT0o5AJXv
/reBEKSM3Ckxct5ojEv4+qgrCH6ZI89qsVTj4ThU5+p6sUmKzTHWupVyIFblz/H5
vYmEM71RGcYN6eC+JaiBtbQKHvSgFT48eybqp2kXF4JluQlguFBQJtMNiWdZ0UK/
H20Zflr0N5nOlegnSIGXMxooIWifa0dU+vAh93dt5+Focb+l7VfznkzHuXtxB+jS
N27vgU1JjMMMkcvHxrhAbBMhsnc+MMsuzGMQF3JzJb4WfJTj+iPBPwODKUpWHzqV
hbYeZZDz6wK9yXg9vNnvfki83UMOPkKTQlLr4ujbglWzFWpFdDOjvTBkqaxweUk8
MRZv/3o/yRp/YR9ijxi+dknJqOUD+njx92MYLqrUx3uulTUnWAifqaiXJ7n/r5/B
JA7paw2Sqnwaygpx9eHJi8wIkil/WylMvZAO2Eh/p3SCXlV6i/GcnLwPnA+V/KMC
MCPSqCiFGNAyH1gARU2iweRNzPF99jD4LeBBbYJchFFCTzc+eyOWrZJko0veZiDI
uGaQG81f83K+nXWfP0Bqc9z9lGM1sCK3lNjt2AdU690mWXNCLYt+OUg/OxcMJ0Z+
F+ZW2jSex1g6nV5PubglcxXSFAcfeiKwmguMxqJtEG3i6GM0gdq8kHwW8CLEta6i
L5hgaLXQYhsZKnfEGukn6PpGyH3oYwHXInsRWf0ofux7omnmZBBew1kzWUyKTV6y
EDsG2fYLfp608fBOewpkd2QpBLpkTpz7sqqisP3ZXhZ7uGuXZmPrWDtQdIzOalZl
TyAMt6fQLUU1KdqkbHS771UlSBD6WzzC0jkPk5a5kaYcW6gWFjEkG+2vp5XQcI4r
4sxMc+oGpDhvs3mkn7B7OqlRU075T/lkKvFtw9pX0QrGTEUxqfmrPYbIBvI9uJoK
Kgj+b7GM5xntXP5XoeyRHPjyBmTdxjYXg0h56qnO6v8F4atIXiWBqB6ri8NsHfIQ
bwvh+2kukVgWoqideLgK0RJjK4qIu8PaPf9r9GZdFCXxEhJd3DkIRYocwJHOtzMO
s1N5jwxTRGIyc3Qua9M3uGsMPeDynpqiUWKZSta/EnvELhLtwHQJtbqscMjXhQWW
b7Jz3Fnese0gTmTyL0RCM+YU/Wd8W2eZKt/8SwAZNutvUENQyoMkt7PySA/l9qAz
jv6yvltwDM3FZRoeBZpuQeDTYVXGBOaDWbS1GmA1DgQYrJ1mBYobQA3wOQpAiV/r
Zpha5a2I7o+KWt/XnLRvX2HV/grP8TZv/dxY4pZ2Cbc3IU+x8oTF+ws8SzLpRY4V
ab+w7PrNwxj/zPZqdAA1tYU2voSP4p1VTXpxrbFNdfEzgemcaya/srBG5gD9fnq0
r7IkwHOfhraK/O82xucnKv1AqTxDXZUNNjmnCU3PIxRafh7XuUvCPLzWcqmSouQ7
+8rA53IQDFu6E+1KeD53yCi+lpBbq9RCucSCPAsz8eReHjmATlG/fiYHST+gXbgJ
Lm+28Av+wgeqWjT6gAOI0ZdzCRUa2R28JFZ2dZnaRNy8ARDAAykQ1EegUJu4KaNI
QgMo5Yp2XCH6TZV/TXfAzVkZUMY1DSFBql4ClezkQ1+4BD9ALJM0hdLIKZ2T9h0z
HT8p1UA792RW9r0pPKeHQfNlA1h0BBRXC1MYbpEbOGvJNiSZQOOJFGhbsKnrVKk+
gcMOFv8oYCZ/XaRdxVA/UWiXBsaDwEyKM2DKoKcueGfheUtdQ5bdYajXNgtiTZl6
SSy/5T/5cG4Xof6/S46Rl3OMxcHEP/NVWYzfOI3eNBjccNzLJEPToSteFNzTwjVl
eWFtBk+ZBmkrqTfLT97KLTj6WHEVi4S9ZWjJn39WGX4h1AkakJWO1I9K370ooXMz
LtdJJHw50sHCia6CE597kMa42Gwy8gMFlyWSdMnZozTd9JrVuyiV1/PVt/EbS6Fb
1Lea45OzSXuKNBYtkfjMyXHlU3FV2FwkODf9PUHvOMbI4AuVvLVy0toomFu9H0z9
vf3jGhXONudcWp4dxejWB/kxoUC6UuNws3gmd3Iw5WK6t0OHYPr4NXRtDP4kqld2
MLGl31jaIRRH27B0noQjQCy+f49t9zuRKZhykNdDmV2KHElBXABWMOrAN1INGycg
+ghK+blT8yo8ajkquVrjZG7MtEJfXoKJp1KeAlTBJ9AN9+XQ+cjMhuVQYOjOdeMM
wiu8tvqCVbhvSTBRktjEX4Chh51hjxYFRiMB+4qrTrOjrETYXfCa3RHdhne0w3O9
kV4ne/sXDF2oRl/eh534RgH+RSNVz51gr8O4TEb6legxpY1LFnsSQRBz6WkyRsaZ
xGVETnkc+lxCQzW+7yFF82ztBfNQEUrHhb8Xw+UzdfXI1rSIgXPQgWXolsN2Rej/
/4XnmCCOqitWgDT5eviii+ytgQ6ZyOc4z1Tzrz1HnTjL1jQPPpxRVMbvsaacnVkG
mTC37ACDKygyRRAE9LrIQKAn+QoA10gOne4JQh/lFWY+TqFLhMQmwk0cuAdu0WUY
Am6aidIBAnqPd968yV/tB6Qnutzr64JDhpJ5d3GH6JYfZXRZx357eVN1fKH95N5F
BFn+GyYnMzMEH6QpQWj8o4EBGoT/HUI9FYvrPYv37VBrLLnE7Pkp9bMh3WQxR6kw
7mO/aB4pd1GOzjZoiQDdXoo4wAdS1ftCVNZPXApeHdCaih6HZEzWYWCGgtQCY3kd
HtIZ94ezvhn3Og+0C81JED92rEXv8lqW4GcmHv+CNueE52F5aMcUNXEbmFtNfNpV
F0QLcP1VIRyfFRrGijSCuWGIoll8A3ry+Z7dHzMPQ8ob82PC+ht/LPR6ezWVVOOA
W+tYMgz7fgc7q4TCM31Luxanxit8L5XsZHTcjHtsmzW3Y1vPUkR+Dg8R6a2aFGfs
B3N2h6GJoaD9tmtXyRjO7b267RDNa9oqo73+wHn5VyvpITbKP1f4CHSWdYSzyS4d
t+VWWx9v4wubaO+9UwK+Mnay/ppVoEWKRMDVjZTAoBNw0QEEDyI6fIFeZtCuXtRR
LVD7TWnPZcTyONupyiA/cBE7yY4c4XWLqUkVymPljlK3lNMU1sq8YM9pcf35ullu
JEs9K8FNx9Jk84gHVWuZ9rdLNg6fEWKppGJQUhviQtwv7mkvD0j7w0Zr16t3gjbI
a5IN5cEN/z62SsYVFHXq+tJ73jOytpdxnEjI1qWTgvButrFu70z3fJU3er4QElxN
MHMKveJ8InBousgFWCP4kax919XJRbWOYABqOdOaphzuVpKAfbJ+eNiI+P1sfJHc
GsPjORJAhl/v68cDJv+6LGP3pgydE/yiK2P8Fn78WgHxlIul6g2Z+rvA1B1L46wv
59Tl5nTc/w0XKQUyqID0qDTq4KOG8yjOY+7WpysaHKfO5LVxvczyjz6ZSng33TiS
413FOsXIRCDr/8b8va5E7inPKr7sQ7zTEe43DiNSVUEPVkndo08PD6fc4WMGOHvn
yR4FBYdEDPRVltc8Gy47+3ZSD7z4tOm/otDKvpoA5GgprvEwuxWCvYGx9VjnlXML
WMhofYptNypxNAXSuCiUCQEdjMQpNeC8BVI2t3vtsfn3uC59TVWspKQ4Ja8PcBF0
uitVCLtjpVam5rPp1xds5Ff229H+y7wtVHkpCAFH1dyM94Mp6NMmM+klULOFiSLw
frKtV6ET6qo0kNWc9q1s2MhHk3QSB/K5/ThAobHggFDl/RiimczdVvkrXZQgDlOZ
EMOdwFHC2YONjJYx1xzyN8cRC6Z9OgW8nV59aIuIJjYb2W2n59Q79EziKPQCbOJh
Dh5phwevH7FgXl7DwxgHRrkRmp6en9rPH6IkuIIsGmaIzT+blFy86IuMOb0jB5DP
tky6GAq2k8wHZnaOciLVnB6fu1N/mZdSzLqYhpVab/seepiAWRQ025/ByaM7r/Vp
ev8yUKhkliytn/S6bPoLeYftDVElVvKCyGK6N2S0MSQPHqG3+mr+le43I5maJ5cD
n/chBMkBinuuiTSt56Zqsmgeg6YrqiBvXxYMQrUgPZorwG4gs7zjbDeIEWO7oSwg
oHPfG/X/vJZb4hVSA2MwVb5OOwybro3RBR+v8mipRAbHTmRGUFBX2SxCpA+5ObW7
TS5PzAm4ISjAbfQp6dgiRRJW7Wv1Oc1i4O326uyqTKJDmxNdsr7qZU/qdOQCkgez
ISp7pNh520r7tcxGRzeshprNXgtwhKvA7gwn32LjEewkfSfu7s7SL33b80Jheh2v
rTZ4UVHBay7ZD7ACucEmM1BAu1i1p3qlr7xqBJBX8JWwIoE6/Qbx362J0KihLZ4K
T1wMxB70zj9Adx0A6/quAKPi2aW9T6Ch6Y25+6RbhrmQKCjPAIlGNB+zdxDAUVQL
Iu3OtAgh2wJ0BWclKgxvMsOpXsYNdnskoG9B4NShH/MsZ92+3S9l8kETZjcReUSE
HDhfwvaM8r51ffR4C7Vugh4o4lSyHVEcLAtCxrzlMfl+B0iyMeO8wS/loTXdSKrh
jK8hzCzlNPgpE8FuiMYq9JAB3o5P63Oc5h0n9yG0AxT5VzHCfCAU9dD8XhCtDKSx
H2+c3i+zbOBj4iOaV5KP5Ki4ZX/tzsSFQVeUj3UtHkQzB3h3EV7yX5o9DJqY/RS+
2ChKTBVjEhFhjIIjAXQQAtQTKCY4VDirZyWYqGc+joSjLfdPKSIhHR1KNir8DBum
CKnoWMSRipIBnl89xaiSfap7Fy3h585Jn7h4/uPjDkUyLjTHzqpk9bk46nAgKA6R
3OkQW9gRySLflrqC+4ORW1CWhtVyj4eMeW4wniEpM+nvzq3F5iNYh/NJ9tBmrJoM
l2QZBeUsRip1KHAVNy0Wp0G7ROMmStsO4Ax4CeSq8sZmHA/T+3LKxwRPxhbCV7ju
KE9BgCnKp/Sd5A5vsZkciE53wLkbIfO9HQUWRPtjpujAjR3jqDqu+/qFsEuB1/lH
BFAjwBYSJVXD7cN1fYoUL0kAYXHrI7WcO+4I0lzGxLpWBuk1IIgNdInemQFBMmSp
TTZ04s2URez9TYvEP4+efY1i2UYvwEr3bSwp5nXriJGC57IqKOa5ugC6VLvDl0f0
tmHDV4isFC7SVNd+Suyx8FTy4MzCDNcZzzhAcJj+KXHHN77Vgb5SZvZJFFRq0LiT
8126Np2UNd6MZ3/xDkEVMw5eh6xxhvCkIRvPA3Z3lWiUPhmgaGInoYJyPO3zEJpx
r8SnHejYYxJMA5eQwbesl7Yiip6kXDRo9zQEtX9UEEdV5jDrnmOz+JlZwwbRc+ct
XtUs5AN8G6pse+QlnKAlWBymPi8V182dMMUgRxU32tEgw52Y2kphwKUMgvdl3PRz
1grsCDUuo2ftRgM9Rjs6UNPfRXC3nzS2F9/WQn6d67bEH4WqChQvKJx01bE1rrUi
8C8CMCkmVmRAWWLYFFekLxjYPnzNpKorSBjv79YM66nd4bcG8plkJvag3syiiYZc
6TS9uIP61dLyred/YGowEdZVqdu0ksNIOoZuvmJxfxemqIW2PJ9id8L8J6+wlkwW
3cdiJTPNWhDtOQRLyGsWkexWDQ9hT/IYa06IxgHlVSg68zHOwcgqw8GzAfENB2u9
+5mMQo8ZwegQ34ULxnFLpM8i+s0H7RdSctNjMynjAmzbLxLsVsmRDRObRGlC5azb
v8M2yDBGTi7Vxn7Nk0couC2ijiC6w7sROhs0k5vO0624m9BdvhD/254uyJzMmwhp
mRxtoJuzTnWqN4zRhfeFFHFKiuR4wgIqz7Dfk6wvrNlc0lAWKDOXtV+KOUqsDgWG
lj/WNEo4Q9b0GbTR6xTzAQfMeWwJ4V+IEI8CTtpLalQO5iOyP3PhN26CntxCooMY
TOkg2/NItq/cKDm87LBIsdc8wHTG2xr4sPM1Zc3IXy+i1JMi8ThA1do7HjC7Mg87
7OIz0NY+E8HhW6DO4mSHXzuBQkZr8e49bnAXLwNJhRaU1lkRerk6PSemALAXUBXg
gcx78zjxqdoJ814RUEuZpbXvMcnaR9Hu5S1dSNh65AtSEh4OUgfodAOaj90/ZuIL
RoOqv0xdSauDGL+iIg7gkZV3T1CWY+AfwXA2GkK+NeDwIqD8i6vZgfpuvhIhkmCO
W7M5gADJJVY89b4WO6OBRTjRvn6pigBmUONElVd/qGeYq9GgwhxLZR8Pu8asH3NO
7+kwtM9ua0LgsCgDMCAcmu3VoUkkkDdPss1HzkJJ5duV4cfDXqM08B+yc/9iDFV8
FcPP1AT0tdtsdJnx7iPgqStK+D3tHXnoywM92tPQtuTWgJx/pW7SN35ciQOgDocE
PJnpYpW5wJQMpoyY7hq58wKavjhpHBU8ZrjJRBP1hMTGaNtitarVnIXjgq1u4K63
esp5YBbOUjWm+JsJ1s3jIc9CPNW2i/2hiPxP5Gcybnga8Oew1zCpI7RKc4m5Iq1P
4O7e4sQ2sgz/Z9CQ8vFe4Zvc2WNU0HJ2ts0XpDiB88gRynaA5wZnPH6oeADBlRes
/jEQdvdKOTqxChN+ZsFtRJ5EmNbBI8A8VRdZBgRMsCfi/dOYAwAiXroM6Fpq+CX3
kcu9laFQIDtkN/S5AABgjw1TCHxbPAmHFV2MwyxAURGVRHfMp1soj3hEVorQSdYc
g5EJbrPQOwB86TNcl5TtrH+RSdsgzkvC+nFJvdWNjntF3qKvOO6rXnQdMb6ZavKw
ramCC4NF/6Z0C+fzLVw6kWgf71ZChRaucv6jcy/IKvynoPOemfJxdVdOLWc60O23
g5oYlBTJL4LYoVt+4ofuSUyvCX7k12GTqh4sATiQWsUtTxUWk1FM+TfkhNqjI+3m
6psoUzSETq70+lhGRIKASTm3oN01g0LYSqzwuzy+T402X9Xu0nr1/bXMbNRMGz1q
gCu7sB+d9VoKIeNXuh3yKUCBX4Dnhxj5EPS6BkVVDLJ76vR90xnZIZTv2YCLlZRY
HYDHFTgAuJaAHgrEjCAmWcYRMDvIAg68QqUleIdvLNp2N1cbAfz6mnz+1+BtH66g
JIdqjzV+ZRQj33/DGeeEi3Rbf3csCidD4t7nEnBxgDMVa3wX2zl3zx9zhfRKsQPb
pRvFbeHp4r2EnF/8KzgnCObH2uG1KFB/zne1FCNZSQMunPRH0CGqoAFsRkfQpNOy
W/G2faxec3L0rN5ePRRKjpR4DzdD2MBWBBN5LQwOmbXtYkU29zXeA2xBreRqiHzm
zBL/R2b7/g1ggW7UgEcR0Fwc+yzrtd0f7qjOJZRTbSa/+KYSxEcC7g/nSNox5s4K
Soj0XlxK4ms4RkvsZ0OPioxJefygrBBBKgcblcTKJKnbA4ljURTPXBF91zfkvNhz
v55qQJwAWC1q/PwQ84VRdXYR+sZoOKqOVQmw09SkOFFz5/vdDyFFs+xuiVMrN3Lf
QBb9pvYhc6IfTqEB+q2cdcygWQC1iP7gsJSb76weR+9EqNatdQB2J3do0I62uLPA
jSeYqf+AJIN/iInz6F5dnNn8e07j8E/fdCFOYIov1+qlt1ayILWEciarbm3yXj5L
uTpEVKoLgNXk2ZqrZmJWBFLws1J6ICIyIKDX1HJXA+PwSQxO5jNd4PeuBvB/Odpt
vpoBqg05fCHYheMlYgmdHfINLtNVMQ4ZdzQ+yQ62uhZtxFV5jnHIrZi2qQvKfFae
fSHSTE1VyyBJ90h8R6yJ3IsXoa8IIeWYFWFj72UEtZwD0lK0f0mYpT4ytPgc9AJj
FFsA6Xi4zKbQGiFm4hZj09poz2Q941QE5tOITn+l0dy0cyv+2fCsn5NcXt1GZrLs
Edz3FhbNvzQzSQhj7bxf5iZl3DBUfwGZF76IIo7bD+qimCBFdKR0y3DdLfj6xtvS
/01NHNEYmVgdKO1iACEFcN2y/GjbY7Z9zD50Wr+eIWs/b0OdeDduFHFKtSVZ5ROH
ifQSSKmbe4dXySIF3KPpJ52QV7x5ShYmQdcmiDQIyyDUPaM21hPWAxyOcF0LKxwB
YdT70WjWUlYY9UZStwpgfXxRLVY9VuxZVJYKcd4hOArjZyllwrgSAzA2kqUKchap
KzNeyyi9ZSP0EkrDaikcBScXfZv+X+iBFtqBlgo+HFoMsoRwxqXzwBVLQC6ZOPfb
PD8yglaujImjqlNPMM5ilcWBYXgu1NvZRtTkA1z8Z6b7kTL2tdZ5LSkcfxVjEV7h
rcJEWwjm92lTQ7Zh3OQEzj1A46X+wLXAHXIl3wubH+PAYSSQQyXchpWSlfPmU8Mu
ek23gH6cHAsjmR3pbl/gVmBvi991fBl+ivOSRchD4yu6VwBLZ4YlWDpLxCnO/ZY8
EhmOOdpf69xtl+j1kSuolwMdZQ4YWF1XG4+zgyeAaQMIqOtfNGluCo6Fp5UmbnEm
A6jSNGQ1S9C6uAA6yJdh5pLCmXWmSEO6/BRxeoVOXWVDwjHRaLJkhq5ecWTjVvnw
jzOBBUE80YAu+HqqjNqDwloWUepVyQGelbV/s1GdPf4ifzt6fpgXdXz5may5403P
dtgZJASMCyo8Hjma52kiFdrBIXjK6NvTAzu0dD78W8B29AOIozTb1NoSODzS7N3P
tqveTMowmyRoopHbUSwveGOBNX0yq91JX23dZRChLnnaK+pKAtk7mDegULOM+LeM
oqPhEPhpRAO+tbcjuD+fU8ADl7Vn04yHbE1svM5BOoRSpoActhZDV/lTvU7JFNYJ
OH6dggj06u0gszFzRqGowQl8qeohq/5ACkqj8wEqgOf2L0ChJmXZhd/mEdYVFU6r
Fd6+5URMvIJu1GiMU41vh3xnCJDM+/5P5UCIDCFxmG7CX7yDLhVIDdvQVqybcM4K
VoL9rt5EL1MryeDOxIdSqBoX1AGSYdeh406efb9YBa2XYCiiFgYj6IEvV5L8/NgL
ya7FEYnz41ZVQUJD/mOdbaRQqLP7FORZzokR0K1Br/nwd+ljgNNwuhHRTpgh26v0
EgcDNBR8K1WHAWjxYbENK1LNlqBbcQ/AXCccRPtC+hH7OgZu0LFRcubLFy+kT9ZF
yKXPVERf5lKcWeEHp0pJFbIDx9WKwZQZWhdX2oxTSKfIWLdG8B7p0R1hS6WpWacr
5tUahBJ1Z1tNxP6L8H2BgySGXtqvMBtxI4uZ/IYVQQF6W7j3Yyd3w0RMJAJmNAQj
5RI8dlMH8A9Gj+oRKB6Jb5xOSFdJ7x2SBaBKuwfLPcjjb4t9Sau3vInl2aK9MqEA
Z/JRxgs7yryGVQcbYcv4OAFysrviBCwh2fhwbdXKDnzRcMPumsNavyFD5l8iwDPW
/yJtcJCaG1fyl6TdMmpYiBbEwoic9ssgImXGwZe9wWyQlZNXtviDTsMDXxy64dWa
sEx474rNQrEJmoHstUeWRQYeTAVuqsoIgEf6/IVXGiFRadGGoyPAXSn+XIsXHRq5
aCfabxYv4H1wfUL1JQSagtu19g/FRuBdKzPmoAjyN4t9dtc4hyXhx7V7lPJQEHLl
JLXmBl40H4SlrqeBwQXgaksd3LN/1VvzAyZiWDpI7ni1bUp/fWw2u19yMLC8rb6Y
B0GyQqYNF2PLtZT2Jm35z6n747WnOEu0/TQdGgeh5EmROLFgqWw6DKxT69e0xxt1
PIuoYwqkgGH3jmRJmoZRo0SlbuCsccufqXI3SXuyKypJFngs51Hk51OL4Top0UGl
o6Hy2G4lur8KyQOEiIcXR/2wYtA3pmTMFSP9NcwM3mv8ANcThsKkQRxBsc6SDIhz
pLteZ6Nh6GZrpQ5vdoJzaHndQUnDNnlUBv84a1C6dr6gHN/CNRP+YyRAZ5LBMwiu
b7K/MpJ7iSBhkVZtKWmVUOChBYdqGDecMoua+kgI4lgRdV3EI33WJQTZQjixhHh2
NON5YM24OPUcbiOpJRglxr0a1wu7if7KOdGbzQyrEZTlQ+n7CYqq1U/2zmzu9cFq
H7rpz95UNghfESlJmnSF8f6IxKRX041nlvtJDd7lUxvHDq3V2x+97oN49DYCpJJX
VW1HI9fGqplk4dQszoCU4Q1ZdL+K0eeZTD9FM/ysQUVxX/Nkvso0+9zgsyg/R7y4
wdjYH+iq34GWEyhVhaLeBpmzAOb+FPhYL6KnwwETGcKbCnGeo5DbYKXMv16HDanP
EdAtSChs00QFjJQdHGE6Dbb8mTL5giYB7XxzwB0XCGv9tOSlmFj+vgoFij7nwJL/
tehFrO5QUvBTrY9MY/0o8idvHO4GBr8JH1JcJehmaKR74sC3OBwV17bmaYr2AvGU
P+3q+EhdPr1zRKBAgty/NBiKY1k9fVMjfy/BqQ3V/Zx3cmha+phSgBZy7AczDLDz
Mr1DnFc7kPRGR/CFpM5+LlgsPHNVVWtRjgU08cTDC3TucKEmmdY/kD246LH1xWmj
C7c7hFPily0IdwcVchi5d3WiOHrgCqIRlmmjCyVc02EUTs8P2GoazQ8zSCY3Caqg
7AF3ZezTf6w5hn7SsCKS02p9ZrSeixXjJveQifHj8RqpLpf4dgb2/QTpRdY3NoZ4
kBV8eevbNS/XUUd2Nax3pDBptp6ok9H+9WR7DCzRadjApUX6g4NeGkXAtYjli8TU
hIMKXuTgIJyjMdhK2ltSzs9AnHTLVf+VZGU7x7ky4BLYgfz/PsFvNWXtOtYlmSEM
ZBtfWC3DDKzU965Lk7wr0VhvP6irPsIaZtDxGtkuoPb6FzgonHeMvPMs3e6IWVHn
eYtkRhfQGEQj1BkzLibDbqilnZ9i6/Tfv2WB+wHQOMKJdtvIFVPSSIs5o1xk/skP
nKAsyWFAl6HqskJe/e2IXtvsMa/gT2Cc7LQtEc0cf/reKXjQS1g6DZEe4s9e2oa+
GVXM9tNforJqMUmKp6Ez1++l0GAem5O2VYdtsg5Wgq+Jlfhk/qgJ/Rt4jFkCYgT+
sfmb1cD4SDoOYrnB/VFcO3ksCnFa5283Pvfkj5jXUoNkiLjYRit4iDGEyZbr3fEI
6Szjl2HlUWjt8dT3wiRYOkZqmNHgxWnfQhEPtInhSBUxtxycoowJX+Y4O5prF2yY
Ioa+5ZG5b2NGCgOCPZGxk4VTEF8dLW2hmJDoKNaCLjzkG974usf6IA5i+ZPrnsIR
eIBKquuBFVZNPRJkWSBVpQKw5R5+4WZtk2KiqIJwEtKZSNuu2Zq8TAPnOp9rxN79
MnBjVR2hmr0iYnykbds9ewhuuk4J/fvMoAYROkGpdRHBlVIoXWLyyzaXk6W2zp3K
vSWhke4DD8TwTUOoN9d/VGlwkUjP4HCtOrIY3L4KF9lCRCnmMz8L+DZgGTIKGcmA
0i94BG1l1HxEEthN1syQzNztmLgcmp039GuPtY7DRrsqkTzsfubCG+MeOlrN5CD9
co3t+lT7p7pon3ru0boFgstDTzRWnFdCWlKEbNV/s5s9JKA1gn9gT0zDpU8A+kWf
sUq7yQ75194rk4jskGQ4om1MKeW2M7HDrJOeqOxyL3nKvrcSSMTv931d3cYo/wFa
ZVYJt5Dwj+D+1rCv6tFYlOSsKJBpqmjCFHLhQ9WXCPJZFU3KCm28mU4mARXFM/yt
DJ3MAf4Xr3yRu/CcdDUj+DfZyyOTI6VLqe7nHKYdVPNhwZgPsnP0ElKaleOu94+I
YNYfXVz7VVFw/okPGuKSTS9vIFcLhAcCxOLoVtl7qTEUtnLVcpXbhK/r0DZ5QapW
Tz9NJ9PWw2F6NIFIzqyid8gGDuJfuXJchkgQpoFRpw683pGbNIkvlVywXgiB8iWf
1+wNRZGSDn25pf0BYnyCz2rqtIHFhyc5zJH+ob8IhOM8lnqCD42YJtzm5CVOj+a0
Ja0nM0gFOWP6xcIOzxzLCitJpB68jYAw0hulGdkYwYaXCtyHpuHEC9dM9sTPEC3I
9whnslIoSLPxFUc7ke0HAjzN5fxyOGIZ5Apgg82Jsg+YNkw8deRlzq/dk1SVLUMC
EaDCpdeYEzg6TZcSHPGbKCzH+ZHC4/ke1leun2SD5DrB8vk0enuH92hcSE/uZmpf
dH9m4LzeDHezRlWva8OZ5SA7J3cD5FLMnk2ZHdZ/Gp40U3gshBOpsZPYfuGztJLU
wZQochy+62JkpA4l3l3IEbIvSE52doh6gUBHBlQDmxKlW9SchZNC3uZX7HIJ2XS6
fisZG5HXuTgfq+E1vOlOikfWfaLITchzxahmMKXgYdnzcd/iGzmNlANlBDt5uAR3
z1WyJNnYuoo49Etl+jXL/3/vxKfN6t7Qd5MTa3IzA6xbRJSFARimteMlz4T9Sorw
R4NcTMViMqijgwQCD7SPXkP7bTpWBONzcAyLOBIpDFShAmqRPX9tPKxEhWZgnKT8
rckchxL2zmVmEV5/T4W0FwYiN0xleJmNBtzF6/bENsFWHBytmdDXx0m+mbFGfwwk
Fur80LO8ye7IEZzOseBCywXVeoqBHHQCbdp0WGCoePtiu/cwD2clEelkBe1dbEEW
P7lquQ3H45WO2R2Zv79kvmgdSh/qOe7eTaTvZniyfeH8L/ZkyYbZwDue0Jh2ieMS
TIxbhNAe5sdJlkNJP2lEgJyKzq/4OzFjbvHo6en19b2zFf9BYg0aoOxGfCqhxexD
AG7HORchNhiWEtOawdnGS7bQtBxCrE34VoQZo1akwky2PFNU/SZ2/KoJb4iGwrOe
G6LW9wr7+TJM4fAapypX3GcnZCpMeeG7zdOsuSiG2EbqljeOB92C6dcHekIy9A2I
Hw4pHJuROIn8fOIr0FpfgTErNBwmA6kZ0yza/nlhVtNBVaUcCMnqhClGlw56QOWe
SXWOyldqiBePtE8gevTBtYvX3a4mgG2oJa4PmvoS2vEnqQC0oAMtCQ7cQiBM/YYx
meZxQM2dVSca3qyLcH8tN76tuRYTmMLQsC2bJH9VeKsKGQ8dAVx3nn5DLWBY7bFi
/xuLCIjJJmBVvPiXKQOoD4ef08oTwR2CrtFfpXh4vhTqgmLyaS+WSFaQQwiXS3a5
c3y04rwnHTmk5s/+TOwe9S+cYLRDClb24W4UBxPsh/JoXtcLFLhfqOjma1Ickk91
hQASs8TDCxIhlL7/d1J76ZDsDtuz6BPvJZu8zTge0YjnGzRecezhUksrCUD6S9vs
iEotrklvNEDh/mOrfAvJz1XOCBBuNb0RYd7BzQFgEa+Z1kpwQZvqGOFEhOU9i/N/
4NIupsQbBHxQCv6P01tUqXtONHoQBO0yK9pUPR2QW6KbyuT9HVXtcY5O+lD+BJcs
nXJotpb7Kc9D+Pgk70u9XuCgKWI127IPspqHX07DMPPMTJuD2FKxQ/fm1a9cRy0S
zjGVO28Nh4ZXgi6Dqtdq7JqG1N6OZCoX5w5spPdJ5GHqW3ElsrKVPwGaMRDCjs0l
+I+s6j2xPfvS5MnZiecxfaTLbMVat2TnS3bmkUjyV6dc11EvKdVimT+S1sfP9hvc
9kHH6QLGujLikaf7udYQPPGAGYs+CHsxGbkmqSkZaUY9WsCLry0F1h2Md4jVIS4B
owg2z/zUPyT7yyo/W8haUTzTrZIuXjWMGg2KQQV6HTTkvvRYK0mDTDccDxfm4vx2
h2ohUj8sHFjIwlsCruEs0hS3h/fJHsH74ES5psINUmWSUGwLfi3Ie9kdauxn0Mrf
fimC2VAwwVVTtopcC7makhb23p6CA50MiQnzvWMwfJjD4w0CPqt82xjGjgS1CGDO
lpgYfp03LcR/sEazPzpUDZU6Ce3poMyNwWmj1smqqPefH6CtCcIt4DRp+tf3nXAu
iTcLceMkHwkp2BRs2UhfecFFFt+M/FZEuIvHbi7zBWYxMsoYXv2uXWNyy+b+luoV
pEvywOX5YWJdRJsx+xrTVdX+3TJPUVOjWm2NDs1x/1SKjV8sbUtJeVBWe2ZRiMOQ
djZ0+HHOxrfEVUPm7E+79kEColqQEnx3O2JqmJ3gU/+09z9jj5mqnSDGe26s6+fm
iW+MiN3Jxtg0LNL4+A1OXi69SWjlLJF5I3nXtDFJw4l2L8IKMqSDGCFXDMv4tT+2
WOFEUsZsVAPTfSs4zh54tqimghmVqcQqkE1e6eF480+e3KUwCdS8k3yMECMwYxlI
rr0fPjRA927CRvktgf5qMyM8Te7T9cI8lf0oMiG0a11Dv+WGFtLp2lHtcFg7qEyU
kunoemFZJn7t2R4sNlJzbM9PhfXIjf4wg/TQ8Bi/7RMNLvsN2uTzo3ajSHeGcnb4
IKtHmRB578QkQaa/cCnP6k/85GKo7v+0EXf6VpZ2emDJC9KgsbhKaqG3zja/wXn3
NNBmyoN2TvJIwi0k+qWe701SD2nUfvabXjwoKwdMBT1a22OpKzCmoXb2v2P7OFlM
qn+HlKS+E2U+smTMJpVPLJ0GsqqG1aDDqauiyZevrZlOsoPz99Lv82qrjC0zXgjI
fodlsLKoaXXL5P6v7PDgYsgI6qfTi6mAUkjPObk5GwEUyyQcXNwDqzK8HJWC21tz
hPcNewg/HKceUIWcfH/dZThqaMBzY4dOFDFGM1MKlJdap7FasLGUbHrLdHmz5Cva
Gu5SKv6LdULOlvi2GJmgd2KFEDRuppnOKs1SBUY1SaHuPuDjsfA8WWPZWz62JZjZ
DOHw89u2KkWwaI3er3dIt38UrIE4aT6X/c1P1/OaVEGZ3KVOjk5tgr2WR5CT1r+V
hvnqehv8kIgRwwG32CJHMOOu3EL163LTi4RyMZM2o4iJCkL2NoygtknDQu7GkrSG
jcirpdYxYlGhs6TeepAWajrDmPnLidHbKDocleT3X/oM+BPG+z977zAW4PZwsvaP
Pdl9518YngY+F2hOMk4U6tTYrP1DwIv15hr26NDfoWLlh0voFaKXZfoDnlfAiQct
T0DLo/rJtCI2Uo3DaIUlSqX/RrIRtrEUpR/27Wp+vekYVoQRs15VnbhjhWNTg4hB
ZweAOxaq47vtKQUmvUqTqlLd8SLD88MKLNOzgN68+PUGdRMmXkoM4MYBSGjXOnsB
M4jMwOw9R3y3PoNXRxq/IUMmTAMCB8HmYHLTyJeI5hI6QHgnTHSeRrCWYixg5a6w
5uZ+Ekg43w4gJNVVCLsXt5205/3K9Xj5UZChSGS2q2AkrG2Bxd0Jfd0ZBfdMZS7e
sTWbFCpas/iHpjgfLxoIND+MjlCjnGKPO3LpEzqOl4uJVWxMDubk0/8UJT8UPOxw
q16C91eh5QdF2+sF7pNJrMdRWvDo7i3/wkfSxtmPjS6nQ7E1Dyeink/AvCBjexME
bzlCPgElId6UBQsjk4dNBao6HrdcYwJHiFLKgIQfamEfAeKCQFtpfvB4Innli4Qr
MI1MSKoOch8aYE4NvUcja5MOlGqyP6mC+C3AXgz60uuwXtzXYY0TxoL8g9H1Kvdg
40usmDi/3xHWAq2/O2z6aXs4jgDU95F20lzBtj/xx0Thj5f0gOyJBhjmIXbHTJB+
PJxPWIT9bskCZTU1dWUG8+UXjv1s1/omIetm2U7CsqgF4V1ybpALh/VktD+/ESeb
5nW7AFZS/g8CHPBMTdgAWObS92HY80+/z0e5+KMmdxGx5sDcksDFvPw3c1QlBdcm
qt2527DrBiARmzw1PuksiBcKrpimmIhCPeyy3a0EtYIBHfFRHzOxXHg3jJOng2ws
icturkl8/Am8mahLukprpNSxb/jK4aNlde1ME52D3U6oy6LIv7XP9vQl/8Zej1f+
K/V/jDulXx7erT9z+EVrhcjtncjHojlI9Uk+ZiP/z69dY+YY39Ft5Z7wHoxz6BfK
b1Y4kzoae/rDyCkPYZqhjCQhZ8v6dD/5UdWHnuZi4y+uSiA5/LkOC/UXdS4wz8pX
7ym/Y28HK2MAB9PgDUMgBkKL5mybw5oYGhwbhrJ1HcPdPlYfXFg6Ji8rK8B7jIAa
Dn5eBa5dz9LSnw3fRyPv9yMOKKripgiS0UV2onRJienzTqvC2SSVGvDFSWcZMTg9
0xrkmhbXw6Iw2T/fUTaYw+cJIJO2xwsaxEKz2uxE738x0mdKTU9kYfohWznU+Hol
ubByAlL0ypZItocMZ+UJa5jQOs1iot7EKldMRHbuwB8Lwm1MjQsCB7ckCNCWYToC
CZZ3fEvuNvGuGKbbdUPTGNQhTbU1CSVB/n1YpMaDppZHbgbzw2YF1BNPCRFwnsno
yzwReb8Fs4BKntqi+aiW5HwiwArbqFENiST3Wao3QgBCrreQ1jN1m690l6mMogb6
+eDl/PjJQfhm3icTX5IoRVT11Fde1+fXRsqyJ7Gmj+RAiGw2tgZ5NWL4IAPerHqN
dmxMYojFh5BlT8ZX2z6sdYAUFilWUem8RUeL8u9ePR57SCQ0WwlsOSrofxWFx3gE
SKn7BETqfFpmKCIrisOzgzR8A+ce0ysLiGAPFU6edvJH8SXuRTn0Fwym9/+lI2WL
9gQ+tJTwcqhKTJBodrRhSnk73vFq1ntIFbMYWpiADYHzfbyCc+b/whNVkgQbuTHV
jMIk0gZydBIoDsCHuD0gCwZblMa4juiNtAU73UDqTuNCPzTer+rGIK7idJPyCxQB
7KhhlrVdkvNzmnVrtKEkioFAv6XP3UKqW6EB0vqT7Oib0Zz5I4DeYyPS2sRcXBng
eVwpSbOUy4mB1/5fd3hA4GkbZKNwxlElEIXK2Y9BASygcd6o91Bl2b6Hgt89JuI2
0WgDtAW5niq42Tz3GCskgz1cMcPpZAW18FUr0ORk5HMf1Tx3x3q8HuVlfmQUACby
TD9o3GNwHKfxmPFnTGkk/jSyugE8r6lV2Ion4Jrs3LZhbRBKP+iDtigkBeUf6VIS
33I7A0lLnbDrX1NU21mCwtwXZOqXMZ98r9/7PEFWMCfzOhVbD00p/tFUMERSgywH
Q2J5nzJXLhvKNlnU3DavX5tGmXeA1EZqv8z74ds6MvhOwnMjsBCHNdOjtj692ihC
ux5w9Rzit1imdwiABmedWgOe5bFO1TR+zVNNx2nHO+wKp4WzjxZLFVYuTIf08tU9
Fnv4zNnIxjxyY8ipbyWDEvpbrqaS4meO5rRxKNKrR2maDg2Jx4JnDZTpMy1jZI+C
HCLDn067gZPcV01xhlZOM9dBkGOZCQM39BbHdhCybmUosRixBR/RVqs19On3agGH
53RQFeMTpkjhcXe6tVq9aZhLaBgAPiUUmjcQhQsjc3gAKkBiRVH0PC7ovue0gH9o
zD1px1dli4qY91PugTwdI3PGpVEa0EyGqgX5VYEWc/ZyLg25WC24zcexxspeZVux
CgRU6bzCdB7tBPSHHkz/0ckcB0l0WrkKlPEvtlaIyZxM7RG1B6AVyXewGFPZwLgU
2Tr/oIBgeudFSd8fKhZRCuEraMpn6DZ6EEguMx5wDQqshEHEtBSioGa6PBLfVuTL
gbcYYcDUozuO2Ptk/i7cIaPA/32DTRrj4Uvez69RVp/uAHwYWkueEnpcgxXoqL3a
xsHVVC5llPkxCQKn2JvRptLDAcnJV1lsjv5rkBT51Cn0ZFZVOmJMZtcAiS33tSwm
Y/Kmdw7XXRtTbG7+o1lGJZ3j1Zv42mTQ8blI0y8pNUaoH3RZRUrd3SixZkk2lxz5
7HMyikJ/HDJ5QGyPSLVbAG7UBVcLuyBnTdFbEuHzGF4UqZoxmgr9KO2mydCDyE+j
cHOSUOChqR6Hra7TrJwZ172twrcgMuuh3jnkFDkA3Hfnt3msjo1F429hgevRpr3J
Vo0cFCzVR74jr0CxHtfnjYJJ89QuuN3l+UvpEzA4opArA5ATrQk2LqE5fJM2dyse
5la8xvpfjV/Yaukx/P5iWPrzx/DylOtY5Q/QzicPkkeTFRxpGHpttlEdbpTIBOgh
o+SZwjzJrQlOuzXMqRWYNrq2c/TwU1ZbJxGHsI+MEiy1opVYPJ890cv5PNeRa54/
9s5/+GbMMG3uUp3E1Ar6aUVyrZhMHTjADA+TRK9NtCLgKaHRuR/wX2N1PxVJ+SBz
uSO20ADOo0wnP17oKGaF9utJaPCDOxgHEF8o9LKZUrZQuflpT5muqBdFFoCvveAG
jqBw7KXHigp/+COR8fE/lli4tVtTB1UTOpapFuZgwaJXQzPiqsZltX8DGtmDD/hX
bL7iCNLcujXjb+kv0Gyh0jkvyyiK0lLMN72LNcYFr0yR5WqnG4YApNUcPluoae/h
wAFn1ib7VsY2QIAvWh+vwmbAOS4K5jODp+OpS//CGDGqkGehtcsCvfNFnginwfHc
0cZC+pY6EnfoS6VBepsPMRLvi0uNC+YCiwQBasXjGWc3GmZb4a3lThjGzgOEuO8V
75XDoR5WOI74FhopoGse/QHQQPq554IU3F3Ob+VkbBK98dl5Km4e/eIYzUI99ye+
Irt4qZhbp2wL8RfQ/Ke33/aENw97Pa3rbLy7HPy/qL0w1SbVheBMrXUlWHZ+XnDc
M6+UyY6gqIBu9pbZ1cM4ZAvd0NeMwKRUsnRN4QWi0v2q7SATppSEoe254z5hTuDx
DLrvouT7Mw3yBErlG/gdRFvTq+G6n1FNqbcl2i+VWLp4qhbSiKD8BveUQGil74e1
d+05DfcwIq+vEBlhSo+G56zm9GOJxGVG3ABULrDbWjTN9tjehbCpDoJvp5cmJEis
MQS4hoCqfpZp1gk1BlrmiRGC4gmvqjEVAHldcAz0zzqkPhigXdLQ4GIoRydElPk4
azzD6XOVrJjONfpNWUaNBKh9TP4KuqCMHZdYpUzIP2N9lexNqMUTvePHff3TVQAg
Z4QjZDOlzahuWXH2WugYEnKqqKPt2D8yWqKMy7fc4U5X46w8d3dmwbBrH88R0lAT
4oQ86hxRR4sGb0Q9EGzaNQsqFoSvU1Vq+MRauWclmYxryvwWBIDISBnLTKXv3z6X
QZjeigpx0gfBEPVPmIgNML3HsVnqGS43/7p83z82dfgyTWWen4SczJsNiPZverKe
49O3CjdS/OdWVqsZ9IT/l0DBGh3G0Ij0t4zGIcdxcZLDYbCOBIxXIyiHYzwQ32Fz
CgK3SkqQBXTBg243lEdv5GWbZXVuGv1jd9qrtbaZYgMG/GMXQUYE9k7Nfx2NE8P5
hy3arwV1rcQ1Nl+kTJuwo23fHYo35hUfdwNv5lNBzCXnBZjsX/orrxZ7OrfZ1Bnd
YzjVivUkv0wzRJo7Uf3pwGBe+UH0OdMOB7FFaRrsCWVD9I+WlLQfVixLnvxk+vlp
6M4nvbCAUXwaalLQrxlyQr+y2aEQmh291t5XmoNDwPBhEzV1heLpFeAT3/rlbmPx
WLoiYxOEY7xwoOH5CadOfzLBmQs0QyHa/t46u89ijzXolewuv/l9wqNsmnRBJo0k
6qak1M4AsdTlxl0UDR4xOuQvK9WVz1ew0PkAEw5laTs7svtSkTnMADs52MnoLCj1
/HH+yFXQlFw9ZfpVqwHAMCmzM12J59M8mPhN0YWm1chYQ2YwGGNK5yimIb+Cso5H
DQQ3QUFGi3OIiwKPZOmec52QneO0NoWp9JC5c/5/omN6oFBVm04BO2gUrSkww77K
jK69FJPdPuADnRRvzw8kEJSjyBpnPdFYOj+DpkzNNbFveOnhIdxTmzJlpw3rnoIG
NPjGuiPdSA4wBxG8vyp6NLw4rhgynmEprakLbm06xS5WioySxnBWrbCxxb4YjOus
+o26GLR/OLWGfBqMLneH3kY9tp6OyBibnkohwovPNHBQ63tZGwygZthcULiy14EC
m0zJkZ5RRpnRgwAdAI9behO64fWTqlG3NgpeLELYrpoeSZaZITbBPf8kVwQMMvw+
Kr62M5Alwufan3/u8cWCD/Aa9rqzzZXikCeZdk0ex23DM+Z9Ctd9MU0u8ISWIhks
7hP7bvh4HR5H+9OGh9ydyLnYXW/5ZozcU14sf1UCNT2r/EtqDv2wm7XYfqM0C1lN
uv4/yJGkWmZLlp9YZljWx1bPpg7fPU9ri8ppnYVPziRowWKPWZUcuzsonrR+3RZK
9SgaKBaKqPP3EXGXr/VUrKTuZiYQiihcDFAbIeWSzSuBX1X0JSv/rgAtnVVDZlhJ
pHf4eszvfMEzrC9z95P7QhvO7Wte6f2ucekhZjH2/V8wB/el9mSRhBmFM+aZEbP5
MaVmyiX0gBg63nEPOO49CoBHzud7WCSPyjpuMDWwvIsqbDwbwFF7MeKa57HzGeKd
7cRf2hspGlZGZnYBBx8P1/CLeeEX9CtD6KgbXbjJWqAYlmeEUiKYiL18C8ACYOJm
hqOZkNLuMkX3r/Vd3/ysHXtIbd2jZ50xnjPnPkgk32ATJaa88DrmdSSaQ9chCuL9
m4uJCTmOaNgzOZXgI9KtiiwHntBKu8BsFXuOnupC8F3maBHhWUXIrp+AcwUTD8rI
TGru1THD1KrQHnVIpMY8FFuhiIFNXaLwDkWyuQ6FdtfYpJHPZYyTCfuA+GMNJXc1
3jHtf2bjGEDYj+kdT5gvmurk15QHccHx41ynFaqm3rnWTWXv6JfYrQQ9vv3MTxah
ES+zznFM/JPPQP8uijVA+YF8uq/G2gWC8y7bphEVQZKmkUywHCn9q/9GpVTlIuvD
SmBBk0mNaNSmVPABI6btpK4lSEZhgqFp1aMBbGV4N3D8LgCcBaKyyLMmQ4zM0SUJ
fiWCye2VCX8st0dKLE2HKU0vTXAsZQ18z3oU3cbdu6zefivMpybTIIwXBR+LSQh5
qH+iKrLru8uLeZOAwDSRK9H0N925fOQbD3R51W81FRUqkEbSM9pBpGRADvnEvbbL
YoKMIiUNxOHMGk+E/+WMBNquWz8tRrZHOS162pm7NqLU8iI++hfKGRgIYwkEFOXs
LsO2pvfEg7LMSAGMoDt9sKz3LHJ3XTRxOBsDnYLVkYm+Kt9F20itT5xChy7WcYiq
U58TWMxExlB+nhkerIBth+3Z8ZxWzCticUqbvjyzJ69PkEQd2M0u4r1zI99eJSSS
RnDl+GVeF/ra31toYH1/XaNt9OAQ/RPWpG/eXT0Hm9sjPg5JTB8Aq+Wir3eYDuFx
xAeQw4jRnODpCAhk9Bk6ItnkAFqNtacLYToBYB81MYcHnVtLpmtE0r8N4+91AJYV
QnifWEvZTkxgM2dihVfCctXfpgJLZs1a9Ov06PNjgSxULGdPLpHNGn3Ivq4QgsLb
qBnkt9Cus5nHCXqSfVp9zNzWPnuHMpZvBncOqT6snaChEOzlB8qDWp6AxQ/pocz7
va5zGPEeA8HMEJ3fXnmw+7BpoMMwyxUxp7m2xk0QH9vEd8OQgichXr7NUhnX2ENf
gLoHVIxolzATqbQ0nSupU4wZslHveY0GgOCChA725X3Qsb+hYMjTrl5RBc/nSYzn
XID4lhnQBjGeHfPz4vNVBjBs3M0WjUfaTDYi/UTjMgQw+IcM5TnlY83dbWEzUBwL
OUWCYRyyQ+A385YqogncHsBxRd+dkjIMk5EOo63Tf2egaBA7rnE3IkJZMPruhCPE
GlqP+GJpVGZuVIXLDMykME8eoUZG6g2aXyRzqOanGd9cCcKRuvpKp7gyxistumdV
Msgitww5SmMMupTYm9u8/UEqJK4OEoBdOf2Wl2c1jOlEkwCkQQTRU8us5kMWX8Ah
YI9TjMnDzfzDMVV3Sh+dBK94ub/t9RAD2v/oIqcuPGDFfG4nYEZOl4MJKHfjFy4d
TES1m5jd06PenOWs4WMKWK4016tW2Iry1k7m+c4ormIRrzZlqlXQsaLaBYlzzjb7
mBH6wTPC/W9WkWhvj9RaqTzCUnyV/ZW9tKBiEF+n1gyvODhb59WpRsyW90YgII7I
IyhmAXovn48qUt8yaFvBQtXH0FVLYNrxVPe74GdrQwuGthTf2ljcnjYLPiuzAFuZ
H3XUboF9CHp5K2HBuk6q7TDV1qkrvSk8ZA12C3gVhRCGnn9FdAn1K8/fsGXxKspS
iyphm7ZBDVFJ3bszD9bX53UOe/46aiSfHDtWf1oUzWuxm5qdMkRADTD5pBf22Hej
vZ8LYQsalyPt85ZuId3TXklBZbPiOdWerOphdbofyQNFyZiWVfNEeuBfKwpxs309
RGkbXENmPU9ksOPDQqZx8hLcq4L4czWXFgz0eZ+lLplRqYGSqmmZ50VzzZjJ21pC
D0t/s8FY6HxJST7duc+nb3bow8+fpJHZ3SE5NcwvdCFWxogzwfdbn5ufAuhET11j
dOMnQOJCXhUrOLRwyU0jnbKekWHa9r2cwhVITZYsQMBo79VUQ4Cz7X4QllaRRk4w
GnQyiWUUGSijmuoofkzAdrgMkkIC/1W8jTFGbOSbZReQe2jWhNGAziiCQSRos6jx
kynjQWsLsUWw817CiKbSwV/zCPPOsuN+iepJAXTYiRH921NsFbTHXu7FkilAhBku
XC3OrTHLS9rPeA8en4Ezi1uIN743WxInRV+Ie7NKaXkmeZGi4pt4h34AKvvNjUzN
UC/e1NQXENpSeYrbR2d3QsMtEqeMNj51Slx4ghJbLLzkrK3Xvb2vy52imW4qU2hC
T9dDCkEEt/GBZH7TM+ncs0LXU3hQGsqN/gV1tNvTTrfOMZ6Dkx8wzSu+YMkSOnE0
umL6Fit2Hp2tYMOr28Ul0/fvilqi30sqSu3gdKw00Que9j9MnzvIg3taToCJatGt
XMzByj+RwXQcDkDg/SEGwcimSjIj/T3SJlY1Gr6AJDz46PgDBiTIBVeomy9cw6w/
M9myJF20scNR2CHQVmY5KNBYYbBe9imsVhkfzo8VRYEy13daTpBY9n9pX2a0C4yO
X7oZqSWOLh7M2HwPwr/npU6H1sYrVLymh9pzf0QHUXLiARblPCk2pqOTmZrBt/VJ
FuEjuH9kTkrqx5QSU2xmrQQ00IcYBuWa14vfgt3fHe5nGDDT/MBozT2ZoqTeyQl4
jv5bPLxSXLIPL02rpfavAVlK2zzTvXil4slCRmNvYSklCArhmbmI4QhgwebubMxw
e+VRlSyln/oXXzmAxqlrtu1f4hTkOGJ7FyJ/P9mhKz5P6C4F5N+44eVil9XY3onW
CjxTYfXaCrvzg0rq+w/uWtBRVJspbJHyqgVGeSo7Y0oa+bE9NatIKPDQSqXhhu5O
EuQXj6YwtBmeTA10BsZQY1intm8jdIYUsBS8VH/VMBzJfeC1yH3vSfGzkh2ew3n0
LRNWIA/LKw/LvlmOHHO0y37jQfqOPM0PwnOiIPzjYk6jFEp44gkbLKBxx/PXVYNT
AaQz8eVSm2F/4z5UkbmzFZCmrLxnCDe2p2P9Ng7UWrfxYzJX/FBl9tBEhB7k4kNo
oY29he1CG30W4vnd2FrLj9juZY2uENDL7lGadX5iinSUvSVWn0WVcjkrZR3dlETb
h3SLJp9ifvU5DtTQLU0eBLdnI8FKr5JWJbtACL/fR1SsrGpS1Q71qWSVb6FLKPE3
T/h5tWPKVDCQqlhvGpAJ7uF7ZSzQjse5TSA11etJ0wFtwbQpYZKIFWv6Jw/8c8f4
UY+OHjZM62+nFB47rNnPFNvbZ1WaMpsrBmCziXkxvfATNjMbo+aIBagmUx2bebgE
nQ9Sez+yh0RsupNRNEl6/KW8Z7plOxHahD3I5G2r7nbFj66nNnSeIlEQcnY5aQv4
nYjY/kLcaeQnyqNd6r5Wu9pPzoTyGzJb77kWf7INEMr6BpQzUwHrSRD0kEOBCsow
tNQaylJyaUpA5CIJws75yfjWQaEFVOrOT9WnJblVZSss0GutC81Nbdcm56jpOIgm
5JDtZ12fnbbY2luGqUBed5b2jm32btkFD+sKBAoIOWqqzRBXmyDreJQ54nOOHpY5
Ojs5ljMCzLph0LtYO3ESmgn+EbrCezrw3o8KZzGvzKDU9QSdKYUqhFDokyLEu34E
vNrNSJy3rdpaiZ+/cygwUYo0/jKNO0ylrSILRGEV3RsZ8srPDnVNERulJPFwXizU
0RzWKZxUXahUtitPbSuQGWfqCJj2U0GnJOw33AkE3lKjOzYzRpK4ZOXejhR8Ga7e
tfowdxpug3kh+05TjWWBsv+0UbJtfUCSV3FJ/PiaBZwiFo5aiGQSMBR1kj6Azad9
lHxA0BQd5+uClttHyyqheHEjciISRY2ZwbvxcTQrjtM5LldXF7S52EZ0k3QA58+P
5d0Ykd1rDEp5nGvGxNWxX0TK8xMlzDAp+hOsGtUaGU04hnQpZ//BYIuMyI7G1s5L
KaUdxEDBUCMMHklhwzULANRaY86IQC2zsvFzU+rIM1OG0jgI+IXM7Rg1t6BPBD8U
w9uy0/O/urIkkxVVrVf/2AqjvhOb5SMmP0CZX7BV0hu6k+xwjGFMncy1ku8aOZBt
+ibFmJPPvdMyouO0psDYpiXt7iKjlm/53LQWiWVVan4+L5zJwv9jTpGINtLUqHIY
W+OXfNY7nyVteIJkxmINM989r81e0pYKhLltfwvgtGWJgEEmdQ/ymnme8MFgq81N
qRCvqY/0FfzekhWE43BOzTnxqkSngBYUUF7h69453OFmjvv8SKY0kV3m1p6tQvYK
+x6/odq8GWer38d1ZGp9Fv5IoR2pjJ2RCizJMdVNkHLDKaMp1IqVhJKY7OiVGAvA
4Z3gVKx3BU3LWyZREyobDK2Czi8ePNzBW2iLiSVGJ5zXTA5aGyODttgtY5/Z+ieM
WnUi+5N47iIlpRIlKUOdEZgSCIBL4A9vPFDM45PXyruLIMJAFerhVhB5pIBIfQxm
YhZj79SzMxLYsESTjvD9OgkcgUMN3HODw6Wi+wtyFtNZm+SPd3ecrxepj4TMmpcV
mTTVdLEmun1Zw+Sx+fBW/YfNbvOwJiTGDXGE7pEpDDlG9xi5UGuRgPlI9jbLarGf
XI4bccq05WgD7lke+5cxX5zzG+k5n+jN2InujHX97esycdhm05VTsfqYAOqqOCca
ORxMc1TBBRg4RoXl9jKE9tW+UFZb3dGX4W+wX+J8ZonXNIOCQrZHqC/icAbJPf+x
Ir6ui3lnj3Np7Saf27o6wORRI29iO4W7BG2Ono9rRa9UL6+yZ+EcEJEmPTrpUp9p
4Xv4dgnf2dw18re9LJj10F8KcBsxdY1/YGgkAH/Ymkr7l2prhEgAonLfszr/bSzP
trkpHnOSA1nxaZHvJqzA15buZ43nCAOmvAaai8t2HBFh+kzVl1VwgZmLr1eo4Ai9
EJeEDhDHhlFq4Voii99JjSNfHqb93qklTr/zq+2VpxHkvqdS9x/19oOuEyKQaHw2
22gbIGunQ31xjtM794jxGB4pBYzOvoe1+rPHMy1fqz92JbCpmsUbQi5XbtH0qEta
op/U6VkdGeGKYyl8Cfy0nuKIc9+TEZh9fgAvRF2L0cCh/Yeb0JKefbqu8Cbq0epy
ErCBP5/6Mi2o/6GkCp6cGx8MlmnWWCgCsUvS0RekGLPUUuvp46ZkfI4rS0yHgZP9
FL1+AGy1RJ03RhXNvhXRsYJYnr7ScoIbn4ZgC21vUkDue+wJhI58Y8HnvvsL31/W
5hFTOlvVLpQTZRqo98JGpPH57PdjAWcaPbMchQda1pYBhf+mciSfiSJLdA39/BBq
Jd4N/KV+SHEUk9RJ0CVaM9vUpzJ2Am05WDzOHz/8GQjX9hhyXwCKqKaZwxb9Gwwk
mSiVLl5WeWnbIkaIxG50Xi7+PYWCIBqJ+bR5xo1hHyBClZaCEPzf8MfzL/ZT44ji
MzfnvKKZ6gF65m2E25ot0DaXofh5e3qulO6asY92D6+zujqVvNOTkTixDZ9E41JA
5khGp9RLOm5lzyPHT+09BBdLdVaBz2nU9z9XMXT8+vZM658MtOAL3nZr5xROcMv1
mM8K/mUr7CEMHG2gcggEYT7RdRz8FybapsK7dwL2KWuXO+hU+1kqWKSO93l6ecMm
ZCjMIN/jo47BVVxODJR3JlY4s/s/IqQ+NOg1SiQMoLmAxUbJnI4m9HdLRUBg3MqF
WkP1Lnt48TWO39efUU5SXH5eXnz3x0iyQStratUb3J64On2ycJX056y7i2luTaip
9qqFgm50pF7Vv9Q3Ruv5s+JLlOvKRZGhlsPmQPi25OuvDhBb1+b6eYf6dH4xl/fY
JZhocIm1N/XhVQ3cv+AsIWz+XepoIXI0ZoaTIFix0JMMWnzio7dajsw1t1vJpYJL
9uHpmKQpvi990y86DkTtYOTLlaV8Xq9v+ykz1kXHHBl5Jr/ks9joNfNtOEhPTeSe
yG2cLaFU2k1J+7XEwMLHKoKBod1ReWCHFP1GuSzLWoz/qI8ZvLZZgoALdBDL5M7J
93H7v2uGCy7bIcWg9UQsCkVWtkQrzBtoLJUbDivEqKWIzrKWe3+ip4N0Nst3eptg
X8Ksz7ABrf56way1vq2WzybpCUBiU8iqCq0m84d2s0XL8edvHA+qm9w2zfK2sb9O
5rDo0oQfEpbURXMx9Bln0rGumSkOfknAVQ22O7zAHq930gEZ6M9KW5ETP3sPgQKt
6LbLV3qTqAb0GqxvRJjYjs8ROIQOkdLZOsrjykktto85/QkudSv0TCTe+LhKnVL/
FsYo25Zlb+gdXTbXcnqjvU8T7lJbKNDPFPGGzDBNSfnjPjznniQPRpwBUF1y4HvJ
BO2zrySrfAx+CeXCUvGQ3uIqfNxT2EisB+6hTW66gt2mRx/Duucz7B6klPbv5RMj
NwwavGiFDD5jHwrWKGWtYLdkt74gnQ5CDwNE0CXSyKhkWwEjxKLlDmxyGSkKvpHQ
4dPOdF8YI9D/YHgiJaMBHJob0K2GHQrg/HqElIYKWacgNihCVnCi6pHI0z8u5ldF
5hbmzUyZmUkNFlg/3GVP0mv7+xRVDzjbzLX0ERU3Yg1vAHBvWqi7oyPN9HvjJIQ+
Llhcri2tBBxSayWhL0XMvfw3OQ3/HtvOeEEDLeYuIHdm+JOUKXgMqt65LOOAjhUh
r1LDyplarf64ltrIFGTlSk6OOCEPZxET7GFtC8JlO9EJOD8c+3vVQ17Zr0XtzbIF
YKJY6LhqQU4nDv1WUXNc2bXQ3QUTyiKx0MOf675Pp5dgrQnHdeS+cMj350hWuLl5
Qr3ZlEw7LGeKUxEbxmEsXHVuUy57zW1+08Dw9nSx7f9FLPqy60TQJTJ5sLadOp5w
1JA5XBz5uqkPE+SbIOARp82VKu2GEaR4Nd2CvJ/TbfEPOeVx4qnUNiKyaV00SHxB
T6pAA7mbiHZ+WBaWMLLaF1vS1IIagJYTWGgki/aNlwQUOcPFp6+NL5McjNeJlQUc
nljw2MOOMv9Xd3UJxpo8X4JCvGP+Z6N2b7SSV/wEG6/U/xqLzOgjEMi3oMoMpA7/
Y9G6MD8kax7Fiy3vK3TgVP53qafIOrr1aTkl6w7rzfDHI54jlf1p6utrbo9hdpNq
1CGUHyVD+lE4aMRLvN5iiirZAW1cxhkrpleYUOETM/cShAiPV1PQ5msGgbGHgr0f
DIhs2Z6Xq0kHi944+/AFtJx4SqZxKCZ7xb11T1Moki44yjJPk17Yq/7BaWQ1iHqj
WY+k+kr27Z1optqjmHb0kZEGYhSRfdmh4vT0UV7hI8WOprzGwvmoFdR2wB1R7D7D
V8XQpAqNT7wk9TlzQg1gQx4vxNFLcfKQPDAKRMi63/ZkJi00YFjNqa+wjIXmDqCb
UwIqcHOttVfHJQ+uFkrnS4n7pe7d/ukZPfzgtnf9gEJJw3uhLtORFZaRNi24/2jE
5CYrRo6H6Y0yhUFt5Kai8HZxiKsJP/zZ+8kdiOpwBkSokXPebEVFKhEtDTIajFu6
buRUrZ/jfTSWbcMcdJV0AiQznAsh9CjMLjJGa4r9Raqo7pGDthFatOfC8HMFfzhw
ExogsnYwdbhpoDCU40VWJxXEU41WZZiPlgPF0wutDJHyx7yAk8aRWbiFhPgtyZt6
znJx28PiSmht/ZcIJ+IFBcJF6DNIo5HX+1G6Ec73GYsbnvQ+zxnkJcISq+KHzS89
KUuCL25DfXoDrkoopgTqaEMIx1RCQZvvWco0rr1R5LkPp1CqPje9Toz5gjstNxXr
eaka7s1LUiIJD9nel0CJ1HiXKjkOyDVFcps717KpnlAaBI83CrrpmXUYOoSo2hW+
3qfpHuWS7Q+jlnd1t1re3762+k5SgGhYeMQJbwJYytCNRtkqY24KJ3JrUqaA9LVt
90bL3U7jbUNsBdQC6xjUYNcUc+NJrEEE2eV4s9KlB2an/KW9pcnzaMNecVO3kbra
lMpVfYDbStspgH4U5QNhbx/p8NeJibkKeMm+P4NZ6rqmnYEd0ihCnOYkSi6LaMdq
jMOIODipQb5TF5ck1OTov7Fs8/+onVqoFVPdvCBrJo7vNWMVFA3PJ8m0/j7QEgKq
pi0u7EORm3rJORLYzpX36DPE709Rz+RJnosRMKMHsMt8M/1WjexHVz3fwoP3vu4l
kzksxULPh/syCNMUcIN6uWRHiwfAKUapKghHlTvWWIkgh3apsieY77YunVDcw34v
N56t53KAjG7vDGFRNsiU7hRGk/lz0xkmMFbbP7J/43BsvmBHAZyq0RfqJ76bK9Lm
HfMgUCP1CjvnD61ywzCnOX/eUPwyKoS8ToDNK8R4lr2kR0Qebn3/G7aksafdDes9
RqQnWVGJRw8jAaUWzTNfhL8+Big07BIyMM5rdc/tJsoyi+O7TPASjej49kXjT0j3
UL32klG169yS/dYXzM9PEfgGN0dYUj+wSlD7r0SR9hgN/2iBrB70DCPjLJEglmbM
B42A3EbYP7Eo7agcpt4nhY0oGNbnpt7WmhYaBlXhsOMv97ofx7Mh3CJKImFKAgFs
gs77iLLsOIgF6kzGb7/5QsFuRbWkEc0nt18VwUccVVitR073tMy2v22miZa/GGi/
bAKqj2pQFb1Is7DWG56S1cZS1DHDtVqUQSUfkYkdUVWqYtDsllJ4hDgrxXPI+h8G
fA0/VjQEG3V97OE6zzzLjL9i8V4vtSd8JK8NRQf8C8I0RmcrZ+bTjgregkVfuSNF
f1u/xcT9AAtc8JO6vLBy7WoQnFEfRK0XCZNXtFVFDwODaa8eoGWA3SsrmwNGrtS8
3ZaK6wVP4/ea1G/UEwEk35lGu5QPPzS2Jh/QFN+/2qccFmjXCMQJAfUixuldIceG
apmDhP3O513JiKHI9U1S7Ub85tPBjfqD84eg8hYoAr0RhuC1I9hRWUOb6EC4Rzr8
lUOBYhY7n02FdeIz4IRYfq3TtAsPuTA62DR0Ge4g+uXy74svUUDQ69a6CMvMxPgn
in9hpstmJKY5ceBcsDixoEbwn2u9r9ce8vQ2hM7SiZTC8b+TdIKZ7jyX1+v+vT1q
dSIuw4GLjLDaYWkZOAyUd+p19icospqRZQIaW2ZHgeEEvJJ9OVUPoLNqAAaJ09Z4
dmSQY6nqyb32tRcsjBa/Uah1AkLF+X8O1TFT1Bp/PDx63ODHdMwMmtykTZ3whLYY
m9gxsJm/rS5b10W5s22cSlSVAOFDJdmnGzePUvjNorcqfGjwCefls0mo+1Qld72E
1IQP9NHWr6F/5+UG92/l1Jtm7qoan/xqtBWyq4bz4TtbMfgyBu70gfv268zPzbLZ
DW01O/ZXQdS86HSsnaeZ8NJnbYzj60If2d/kC+ecJ127Tr+T4qDDiiRUgMsfsmp0
2Fcpk+qzJbq6smVP/Ha9AJqVZQie1m784lJCscljD9I6hnM3pP5wZn7+SrxQTPLo
+Y+ESvvvwfCIIA6AA/9z/sLxofHLZfmvabc40fsu8TxuSEaMHWKxTbLDQy7iAe+K
g//0J70mx5QNhj5paARnsjY/0cT1qrHPNqZNk04qJCGBh0svIHzRQjMCVzBKxmIb
Dp/DZanefN/CnGptLznuajS5nXS7IpwVhHpVRTa3kEZbLth2vtHkR33Ql3nig8a9
XWfyxfWbeXr+TSQ4ooS5VXNekHElQ8mqz4Malp/R9/F+8kMyYuVon0Fn9PgX7PnT
Si8QOrbNkxthtIyrAI0y4GVo31CAdNB8TO70LgnYT/im7gWGaTK9ZUKpiEC5hvln
0gWVywS0QECe5+ahK3Zwtjyr6llUN5iHumDjGhlFyPr3PQ7TEu+IPThvCjoeEf9c
39pFDPso/LjoMz4fm0x2sKFhHoSuZ/LBF9S8TSOeFkTW7lRfQiOsszqDKnLscw7/
VlMNXJ/4NnRW9fONO7VKup+pf1gkL/kiISQM+CRQJpNx+WIy2AH9JXYYPflXQ2Bc
BoFGy4qh/cdOWMkk/vjz57owc1Z7bPQIYeVapMo+Vo/pU2PpkVIAW9WTsR8/v8KO
LQo1FzeMZfKjM/tCwzmoMRODbwJGaVGhwhtxdQFgj+pBbF2F1owlwXXPD1bcv51J
mTDThP/RKGTnt7aRJ0uQBvkEKjXcUc02TTHLgSA4pYI4O+uGP7U9Moj0K6Ebb7yT
fLEqS1mDWAbE26mf6sDn7BV61fP02x7ffTCQQfuSO2Dm0EjOKZEWiz3mzlAAOMrq
9YN9Sm1Mga96ChwhGRHVrNLMg2nliTLjOiuqrxY9JEyqz5uF+wMWQ7/KUuY/JlyJ
yY4Fd9tYJ1Hci2hrI/GVPKvCKpCBTURXO3gMJ56GF+evj6d6tGy4VLRHmQ8Ez95Q
lW6MAj756Xlusue230Wzcn3M+9sFfl08vZFDGHtokkRUSHW4SE0vrzyoXzR7mmao
eOp1PtxCRKlHxPt7etBiExEBDt1mgnKEbq52qH87cl71mUfNCash7ycyA1XWjQS1
WgJlaLg9h2lpgKzdCdvolXmzpOoZA8VaB6qUIoBNNB3qh6ndzoZfiwcgzNu0oDCk
9RkvBAT9g0U04qipbIWADFIfFgGUGMNnVwabP5Z3D4EeYlSAz3XzvZr422Zjg++9
hNQD1eTTmMT9f6Y0yH+gP1VKBwCT93rAUkwNQXES/8kQ5ZPuXXnoMwSBowUNvd+L
UtvL9bc3tPlNA6aP76LbwL+/xqB0a6azXliSnOkjZfZVFUG3UqJGiZI8V0vqli0C
Q3zt9nNaSWMxUNxolsNDNcdl3oQ1p3jHeOs39jPVW3ubfMydJoIC2ZGlc2MeGCAy
HG21mzlc6g0ngVWGiUjJJFaun9GvgiAAkTIxgZ2w8ZuxtAFrLrkCUCJanP/5TO09
AtKP4hKATYN6Ruy8VQ/5jjZ3j3sYAlsHqtLz7capjkO+TJg11yc1J2jXmgjFxI8S
7z51ttyJgmA2QLHPHxeJeY+wm1H0cmv+E1cww0CzpSqJ7UIZafnsm0L1D2YO8nN7
xP6OkU/IIBcS1rIjI3r01uUJw6ZoEztjeE9afLzL4OH1xYxhGL53diUnuFNgWN7H
rr3+EYeFp6pvN78XVYGjy5nn8Bx7YWv+aeflFxTVkx6WmIEMHs6PKwCFIPM7gnV6
8akzMrvqWjw3VOoYkRvL3PdxeND84KuRXKLyTrlYfXXtfeKFinPnUv6SlUbYgnz8
7d3ZogGWJ6Oygvdp+uhSh6ovHZ12M/kHrLKe8ZryauBBW9s49dlQKtcGVEqLtbts
XcU8Udu1OIpLgkGwf7lEIAd5hpzok3DqZH9Jm9iPz1wQMEKO4+35ay+kEfWVh/Yl
9Z+bgSAlLLku0zgNR9PhmDKAzYj1SgeSTyW/5nSeXHCSrIEoC45cTsMBUlGlgY4a
mZyqmSHtQERo8lMlp6NW7ZbzBM7rOe8U8m6mzhTb6HhG57IIRibUvzekdxgutDRI
nuF5L5Gpv5l4ld7E82e0PYRbEklVmZi/WH7paUQUyXDhFTIv+JzHibI5h2bItmCw
cdaQ54pbotPSYNAQxoZWPEeZsbJcFHj3Kvv4ooiG5JSneFhquv3NyV12dg2tls8l
8pQk++YO3vPCIRH/0+q5aSVNrKxoRAcG7YgdgLq1brm2+yeWabFTTER6aK++6XcB
W7tJLQRyW7zbkUeY42qNuP1sAn92l95lc6wfB/FE88385n4HRco6yS1o5Y+nPEls
kHNDXC7K6IHHmOJOiiImkxDow1ZcZ5Z1Z8uCZAmQblYc2IhK2vuzrYaAAcH6g70C
uoQLN2hRxwWzdJ/aWccnQh2uLgWGcsc0bDudgWQaDw7VBXWUsdCNqflhJLnMDG5v
vo+IF7mWSfAQcU9A53kp4QFgH/m4Jkdr6z8wo36JYhaI//lMqL/EJzTMtiu/UoTs
0EYkV9ujM09Vbg1Eaack+/FF0pqVpU8SShxiWV97+UvsXLBW7VF3DwU41yW3hnX0
mLLH7tsRiBOOmmcnxqXSjnOSeT9YUmMcLEmpJ1p5dNtT1JgOSY/kWspr6gFZE4JY
JvxNuWxVeP6wFkjY/1EgBkGloQH0Tc/EKqW/MD8q2j6S++aV7pxh5H+A1K+dKkew
kPQ8UWBr12KAUQnew8CcdmiuMGu6ys9PrBOTdyOAoXzxx0MehZLv1/kefR8qT18n
VDhTe5bknbUAoBeGptkm2hGYETYzMUXl/shn5GIdBi5Cz5BPLSU72EdJffZnoPg9
v9APX3iiaAavdVlgbSCewQMQALNWK4iTs5MyjSPDDOnRM/z6PAHpLf3OAz8RDosB
9SDzokbnh296iUSAN7/iqYnRMyCn+icxSYenFrvxYpaqvCGiBdbdlfWy5uVXaaox
Zr4nq44ZcDUIvEZXy6jNjKdAAPfc24wkgnzU0BcLKloc2H8Biw+QTugU75d2fQ3i
aojDJqWZdvYOchHTDOM8+2VOTQuznIXYmiTJbV0yKUT4hNkySMlhR9ywD0xENYww
6B0SfHiSmpDFDKGcElIAuXuVaeZMejeNrMHxoZlsOJ8LLf986zB94KySJU4Vp8Rs
52IUbisV9ZRo734qecgL+g42y5JdhNeE71XBe3Cohe9npy0jZeN3UXaiTNkrWgk3
gVZjUDbm44lSyfMPwa553Xu789rBK7y2CxX20LiAH29CuT6BRSxgB8hw8IyE6/HJ
l3QgF57uXUhiZqu5oC6FNa4HhXq5G8NR65OBkNcap0J7BnE31dS9Fw3KXfkOH8Gn
hw9yNxOf3CeGBHMjC7SNt3/aKFmZD0Ltwlmyxk0I0/dIkU9vi6kBgIYUgApigu75
kUDT/9cDUhmbc9U9xTe5NA4t4CeqlEsC+P/zuKhtsyqoCed+cpnwEemiDWAve8g8
j40+FZma4uIYuDT+fSTJfgoJLk4u5BsXE2EQdDlYfVh9888c1E0a4X6Kr45Csfyk
5/xtHgbNNX1cN969rjtmthanI/I9Fs2JenLo26m8+uPoCEXqSSFXB+xPY8kAsqiE
jBe4rmmlhkgy//xEF5di4fOEiKyY0v6S7gksC7iK83KVwil5en8/u6u0upgvWAA1
aEWRvU0Y/eVX4h08ic3YkEOVMENWupXEIl6wlnUZyzH2B7iLvrWCtXADlZQHwME0
1FwhXBvBr3PW48MIdHpRnXahZw92bOlF3alT2KFgtw02iT7OlIMn5Bh542CGl1nl
w+q6h3xYMLEDDlVUz/vH9R/UHpbI0E4W9ZG0Pz0F0xsLy0AyYBgs5KNIWCyxrM7e
3vHzn9FkPMDQbE54BxCpL5hiP4OP/4+Bx48BZJwKpce/FuyjA54Ww9Pwl2Hdz42w
FsYyHLGljp2MRMDE+cB7Ty557nzvcaERV0we4e06CVsAUwRNOsuv8xe2CLBd75hd
52PVgCrDjw+S86Y7WZR/NBbW6At7HcyqkDDTY89JPDBsWokmFEqt4iUgbkXpGiI4
ce/W/JHwOXZzckKkLT8O0KJYZV/DB43NklFv/2ASas151DR/2vips+rUAbzWCU0z
m7v645AzaAoknDd48GpaDT9Zp+m4dEiQA4N8gmEo6C9G9LWUJFIgvZ3Hn8+kLytu
ISXXc8WocZ/GHx2Q2foELVGOxzZJwL6pTI2dtxzKbVpqfpSSAs6qSEplYc98gSe3
6o7RqC7zmM8JVePPEw/dc0NNJtIsxpwbuKsBmxYIAgsT6Cx5xXoR2JWtc2CcchRz
SP3RiDKzKtV70AcOp2VCYwnBz6bqcla96gM+GpQAZ1AHKwxeIUxuqbrneqq4y77t
7mfYmkG5igB2g1knd9RwOziWzq5VJ5bemEDudYLYLNGBucslDLih+T2jn3ZWpMsv
ya4rbR4ivMOq2q+0VgBF3OuDTIvTCqMfMq9kS77oztZs6orrj/mvszg2cGnRmeQ8
wP5BcOv1ZyjrrcQxh1zt5xG82JwEON1Y/2PqPdAoYCgA7qCxxr9V5xHh+xVSaQ1R
5rf8y94zDwftr9F8P81K1mJhz1JyIAtSJXWrS1XFJV0JrKiISn+cTIkKk3Xo68+8
sqcjKiS/sqspoTsL8PLJfZrfxQmOk+usXSqQSlmndC/vUK1ruBc+P/dSjEqyOI9h
r3c2JLpG1SHVx1Cuz37rCiRbJUYh6366Jg55Xpjmt3gPcmhkMqjVGKDT7vpyBbV4
MiCyNv28vQ8ce3jKfzHq+z+lAuOjaElXNEZZALhhanyVv29H7RMpGkt/aazOlePq
v5Lg+kfqFwHE8MEpyPWJEqoKEiKowuLFN0xnD/X0+R4FyI+3dgDu+oZcnauOMjQ9
KHRv4ymMxjAUC89Td356ukRGSOBlcWD5GOSd1/vn/B0T1f+2FHJGwWmrZs5LTj/m
c690WlBqL1hUMaMD6HvyFvFIoC8yUXMCN4kdJ33HHr0QV1pduhh5TDVIw16NYx/p
cRQ/IeUpEjQBxtioPVgWm51ulDdXCNHp1tRb63TRXOuE4Ef7J8sr2V42lQ5QEyUT
PeOoforbaYm9IwJQqqzxlKbv15Gx59jXM8bKGkidhh/+fe3WMIeKtC4t5b8fO7tR
gsQ40dIJynTWKCnP5zq/pTzV94HJokK3LfVC4MeIFXWuL+9IHidQvh9Izk/wUaSu
jiVdv7Sy0MzAq3zkfk27X8hHAqBLQuDpNWKkKgLl2D39ZeSBq9O9EHgj6UOFXHZ/
z+HRhHouQQ7QH5BzbNXPkpjw08Yo++ovT2z77UrXRAFDe/Dc467cNeSLCQx1j6N3
BtUcrHOcrXV3h+b7fhpXUi2bqtbK2ds+Si76NFprLiEREVKLuiEJrJysSwJfifTM
ImeYLAnfMfeePXVYUNVB7vWxXIhYeTEeZLL8yH/1TPP/EtBjKB/yEo7R3TUVzOOP
PCkkCbkc7q0UXz7LgXPYB4RqJv4RT1qe1A7JcWMWPBs7EbL2Oc9d4W7I3BdTQeoO
fwOJ9KvV07pwmvz5IDlPvhcuzCc6RpC6CoCXpx/uZNfiWknHRLON3dBH6Fus6dT7
90xrq0SQ5dt2Tr0ruTaT8gdHqJK+Oi83mILwyTse4VCEKh3SpKPPW15DB7lbJVat
F6i8UKBl5eQp/qnpp5qEM4OKL8zjh5NAG8zpCW0pTk6t+vklHey/8B9yJcRz67/D
Jc7nxCuCo5UKk3GTEi4Xmw//KzRPJ94tbSBxjS/mblAxgshCa8gwIyk/0EpClt3n
lE47CiDMXQYnNxlnFPhEXze1mqP3Fja9ks6YHt1oY9cptmMH+uBk/itU/a+ifKxG
uI87gKLR9jZdkS/MYrvKLrsolzdj1JIiM8f5X5Hq/ZTtxNLqI9fy4gHaMvjQcq1Q
p7JfFwvIM03JZxGx/r2SN1pjwSkXxO0KiijMvOeKNGBqMIoLhJtpt5p4ncM3LKGt
fEE6JWRErXryhAdlDYZyIWkCHdh8Phy4mgm4XIgCXoOw/K158n2lzYO1dYOGTnhi
2bNN5Db5a753+XJdF3F7rmYQyKvsyx4Cw8phBbjTdQhHIrWi9qOL9Ea0hMi4w+w3
wMj4EG6rVO/amnxamVgy8C8WBMYmeDQquGI33QX7xhFAJQk3Adm5DzSc42OpcTM+
sJfo10s6ftm9gcXC7jaR0Fe6kkIVsH3QCf+QFSdH3roO4xmTLdGxwBCxgqS2idzm
TFwMWorJjubSfqtGOzL+tk73ELcsOzPt5HosaD8+d94OZcrPufEgzxfG13lYE1hr
GwrxvogGbfQnM9RUnYlbDOmMxGrVPNac+AxQIyoMjj/EYQBpb78mqZJEv9WMhjYI
ItX3E+6JsxUS/NRU3ix1ss2ayyT1F3PPHaV9IeT0MIccDrR91f8PL/wnULWysn5b
MGJdMEZL/Q79eTnEpaW6CoChYOdpZnTGZFiIuWGzOreXFU+zcryWqyt8dXTqHX9I
ht6Ji4efp0N4ErR97DFZYshm8Ydwa4JCP1s9Yk3CFDNrbJWZn9TM+RVS54q0KxVR
HsI592EzVJhfr+MtKWOz8InilTNdTss5fn3jB5dtX+9Dxd9A1mLupeUTu3KNGEze
oY23cV8S3Ien1IRZgu6r64eVHa2CL6C/V3Cmn2ySmTf8OCDG50/R7vQc+ng8jCeI
1UTi1c9s1a/PLfYGy97gK9bNx9NWiD+Ysg5zBx8Qmz7ZkX19yP8u6ZulOokrfakf
FC8XW/H9p33FZ7fI/roJblr7YKs6QMSBMo14uyh8VvGLW7glUcbFRVutyeW2ugl8
SzGsOJpZiqNIZ/0ev183ofRQQ0/jaHMN/6wJDnqO27wwgmAVaWoOh3mfMRy4xoYB
HiT52XsCm7eIQVxNaIoK9f2QUGzj8iYD95LaB+BQ3AdPBq42seMj+n3TBjDjblo/
s7S/WYOUtBIKhv8H6qiAgAXwP4gGIlFmQpRh/G+A/8zfMsxf61qF9Jzi7qjsaFlA
Z/87S6hAowSohTi7qXp/AIkGCtffwjfabqc7dso987XTuqUBCB5xC+hP5vlIQzjE
HJ519qDQa/lNtbgtB3rEkw++/rKw8RuBDOjtaehbESn8g7ZPqBhPJNC9T5JTojxp
MXbOQeM85D5Eu79hdL7bP6hwFfgGRHDkUFzONxhyqt+7nUjzCrpbCFChTBNDRp0A
O7q2X9ZFj0lhNQJ006lWyPJUe79DyXHYYEV5aK1XO+kFLedfn3SRPTOYQmZZLRrv
VLEoKpU66uF6q1n0wgeYULb7+0YpNwd1zfL7DWp2L47tlq2rw5TxYGQzrrL0mim9
G2g3qGi8xITMHRi1RtR/OcCpmL7vri6S+Iq77r17B8BbdLJpz37HFVlNp4cjGbj0
q7wwJuCsMJ65o0eIoXBu54oFqExXV6w28haYRnMalQmyYOA1Sx7wCmhgEMGqEeWw
wJdp4uqRKozcyIl3s56tPNr3wJWnT7PC1lf/jNapqWBa7JysaLQSR79o7zQ29DvP
aDqbfJKJoIgZvpa7J6k79GOiyehWOVNWYR+f4dzYmE8NYrSy9rxU9wwfpCgr52PA
0NC8ySK7SF4yJ/JZrGobHtwZRghCA0Dy95roCmxMkc3AI2/LBaRkXkVHP2eb+qTu
wefJVpBDwIKOAFo8ENHKEKPV9W6YO7c2KVOReCmpAPsIncXdo81twzLfHEP9qwxp
1gP3DhtmJFweTQRS5ewwJvyBvj5ZKIT2WGGkLxUhxmjB0WXsqFnRc2qwYffzLyfC
2m+prLR48zieNVJHJBuOP9SCucL/GQ69IqFRKEwqmPo2fXOb/KXa8X7YXDMPWOj4
tuH+026lhMFIyCO7IFPEInKdxRQRm2J/xI9ZxUpU4S/PwQ6ZNbKd19kRytr9n8N3
hbRUOmTjFOcNSmiW1GDsekh4JC2WPXd1LwJNPcObY0iBPd1Wl7eCqd8osXSYySgq
JG17EV2YRYQw+VGw41/ui95utZR32Qzn++9ryQLZAsspzWtGwzihKKSb1XP4YOcO
g1lGuzK1E3UzKIIc9aCVt0ARHuoBf0pgDAfqzowiO2qHnWOr0ed8gUhttPTo85cG
BhKwm10ItibnsMjhdMx2nkchW64YfwslnhU9zPf8RBbtRrcYftcPxQYLApN2TIcL
6L0Yqcp5HJXMBpA4CbEyKRKmQivBNbaPJwpFHweN9gCcmG9EKBZkJBg/dK43T1KU
GpAHfbRc5ay0hcT6FRACB75SIv5lxMeL04u52tM100Y2cIRD33CVfm/hFyGUEobG
rjercTJwaSf6bp/jICWhS+7Uy05ZSoYYbSxqpuN9j2z33+RbFGraCmTrnTvy+EWV
RuBSCgMUEMylWp9ylUR/mGDgA6H8HTS/pliR577IdgMdXQC+QVo8X4nraextpUR3
rz9y8bRsXC9HGuii69EFLmlk3pZyHkePUTp06/fgIzWZVFAOiaNqJzsd2/UY0Iky
B+u5wyKxibxAJf1zD9qfIZl6DkrvcPfUdUWkDVz8qTUZc1XepMCqYEjGoxhc9JAi
q01wH/8dWv6kYkilXOlHi46k2fl6DEwPwmj6KzxAqvNcJZiXPs/uVvpfwg09Sy+5
LkzxZcpAg0g/6GSXI1CX+YYzGyR8KCxPM983l9SM5VUsaV/lJ0FsxD7FnjxhDOMJ
J5nG+SK4DApsyiPhlc9jztvvj9t/YtG/E0tT05yqZwXbu8xsArn5O26EQ9akYi24
klOQFSIOWICecxMfdciJUWu2FTlSf/ArNLxa7FHrIDvMZvD8fgl5t5oFMwdnLpZ4
c9oaYNHRV01njtWZYPTN4GT53RHsWVP7MKnO4RNbleLUMMaGBxgLfD7ZRE++aHym
hd6C8Vv2uhrx33RKHDskADjj1ODgXAy6f/OrlL/YS2dR8KFVaZqh7vYtvoklxOuN
jVSNVoO9j7gu0Yxt60aRDkAdgpj56N61mY6S8V+HD+AWBP/q2ajXtGS9rIMfj0Lr
LEM+f7krqV0tYczcXX4/HEM9UncCoHYJkFKtN8rbek/iaxOY4KSExoAsa5CZSxua
CE4VUPnoksqbYnkThBhXJ5pMBNR/V399ALAfETAH2Ax4asE3XMyPBWfxuZIPh8p8
a7naJ0G0No+3/gbuUOFtuenY8xOdWzbgthc/v2pZ3homSnn9VQlOB8Y2j19M0e6c
jUdegssS2cFOZVLX9L/Chp6qyIMBsDPLfGX6X0Ju1T7F7I035owk0HKG5PVJGyqY
OeeLuPLcNaDSAGfoDYjnV08hdG8DUJ4pV2WruzI/MdHkg/CmbjUZSJQPhQ0p3t3/
eXSa3u3A07SvhpFxjigGgUpHjrKrjAdiXLMrYNLQnp865P0kUvYaXAJwQuTqc/Ni
7oTKahpvaY5aBq9dwj9EQv/4GBgHbqgDWc5gkODq5CWzjT544arneMoef7+m/Vqw
2Ks+mfszk8uocJqhmz3BIK9OMuRO+ldEXAqp26OCCl4TBClrMhbFGcn48SFoPDA3
EdTMYYKX5W+fZwrd5reCeIRCu6mwRbbkKg/5n4Ytwrl6lMf+xsDi+D9SoDy0S73x
Jgq6SIG4jSCOhVB3TcBHbOH34PEHYe6kW6YubgYAO4v0wqn58Z1OTcVqxDwy4HEe
xnv37VswZP9jrY4eW7zLHEmH0rd0LBU4jAg0IKwMRjIaTUG6IuGF6UndQyD6vzeM
IiEloNKSFHjQFpxESChjbjPABmNGrrcKOhCwntDzMurnkIrWILFqRZSXIAimhNS/
kI/EvtjUTpTLqobN/4xXEtLq6jci0Pfy7L7+cf9Y6k+2r+OLzjYWPJQiHUme5MNJ
X0JC+i4puQKi4VXl90Bzt05Lycbq8FkXGAbqsGzKucQn/tu+mIH07uJ8PHeW4p0G
qoGF0frAndSIY+iJloUINFebL7iLKoPwETqaweAn1QESw9WbKQfAWx5fNM/ZXlLB
epup4a723CS4xoZtjTnzKO6NVr2W5LW4YbSpunzE9zjBclc9q9IjMSJ6QI76xRUb
kWmtQzhF5E7ESlfYldJPSV0G8gNSK6lnoCtdWVnzz2Wx7sK9zAhbIKjVcHHHv+wg
9dDnWj7YiCfaz6uxUNiIDd7POPQ9W9cAY5JrHKRuQNah0tJbqd+eCOb+i6FxUE8K
TLl5XXvZNC/M2uwYnupSx/ngZuJ+f9N485XusEpjoQTNjzIO1eT5Xwc0sQvrOHSg
giPb9fl7bxp42bgaY6IyM7UyLAXJw0oVP+NLCSmCc5UVwHw1H4QyupKpy+qgSER+
jBzwBBSf49F9QYQ9YWgGR/UxyT/Lerx/JR+rL/i0hpiurfBB+RFSvbKVW82cQ5XQ
Upa+vwoOB/MMhHLGG5bBzJf950ZtT/s0nFpI4kWETJwFE3Y5JkXD0/DiU5VEICzf
t2KmlpdnAZUc2nDP575O/YrpBx7q4JH8nEpVZPKf8CrGnCBxOqmDJ/CbdWxy1lGe
8b6n/8VzcA+MPIaOW8PInBi5/cAryO3XPCwNhedDKAVhiVEheEvM2yR9/QaRRUfp
A130hKx3CYdXUSRjOuy5j7b8drXQtvFG8zS+C7rATUW4Jwx0Sfyaxt0krwSPK083
t9t3/ftcF8mFP9sQYX6UDtwfxnl3B+DlaIqEH4IJkbyLvqFCAHXzIDcgFsf203Ho
gZ/hEjjiEb2jJkFo5sSNnu4HDJ7jRwoCiNa3b8mLHS+S1B0RDz08xPBx3ZojhUPW
GS1LILHeBgLLCoQLLoygcmN0bbdL0/Czur8eOZRgcPeLeMhtBn677DYbe76uY4EF
NHoTtlsIuZd2wKN1Zw+ZOM57uKCHXDObSAGTOnv48D2gVlp3VOOwMg9N5NF9nwpB
aW8jhyrPvnb0OeYrxn0q9kB5n8v74uwaDwODlj3fC+Wo1RmuijNApAPZDQXiN3uD
L9SN51c/X5ntg/HIZZ8s+4IVE8Q9n8vFRNrwWOqjRRiM7ZCuh2ZY1RtpcuyN+AeN
PfEOP1O9BIA5/AVO8qtk4ECUvz/Ya84rzBGq28eoQhwbF9opLVn6OBSWfpZAMROC
0EWNo7R9YC1WtQd4GyyLXBme2VrlNuDvA51rSIu/Yx13s75ZCECnIIKUAI1T4TCw
UPQNum5n32Is8QQ0vE3d91z/zZVUITz9aLHFD220AX1s/J5fx8rrNabGziK2mGgu
onuoJrby9eEgoAOwrK57AotY5CqYBjKf+ilI+Ipqsrrhywpe8l2pUdgXbLTgELH8
7dA0SZoZ4mO4wmOTg6APSzZnTU0FN02aLt4HadqWgqenqd7fzeZP9XMY0BRoOZww
KNDAvHD6mx2d19mwCXCEnSlJqn6y//7Xkem5LT4EtWMhJUGmvW/TF9QvoxIMeyM5
brYgFRSJKHP3HqnCmWoxNiP+GEbwTEsAQ+uhRHJNL38AFLcvKNSrVabE8gqdS96n
vWIq9q05rnbo7jRSpJUi3W9MlwRdDbFtKzOlKdBnM7rIJZ/d8Gjw6/l15kQkmwlW
mXMlGhri1OPAb2Ouu0I+Nm3dubcXTDzMBjPao7H1/A4s5+qvL6ziXhn1CEkzlpNG
A1MZwywVd/0S/4/GE+UPqjxTwtgdJ3MyPBodoUAVjelOYY7L+MjGVJRccRB/YH46
y1DyCHZutlsLvnCmu+lnLBPXNXdAAXeG8w7PPq3UXYp/GEooH4SSGJEuYuMwngd6
opzA//V8GUViBEcMVIJVQfJb0dP728V2bn2usOtmWhZXILPssqCFL0sqbhGf656n
O5i+mMCwRucD3GDi7NjQ7+/L3WqAvwkwVeJK7h+iAXh/lxo+dR/7ilCoPa89W5Z4
LVNHi1yomWGVLNEUxUQsCcjjGsXEkV3i0GM7GzMH1ro45Ru/dtmTTREiZcGvhcMd
nxbl+Nv5SXU4trQH5rubMjjk6C9h1yevZfkeBul0XhAC+vyiJadJjF0lmuewPUSc
K2qxgAkfUhxWeiKa0lEtmlrQsFxpfwLG+V73MiU6gL8nywIjIobUFtttzwYL1CxZ
2bUtlSFULMOt/rCbO11UhVQuOJDub4oynrgcaHk2k9hxgHcc2dVDhAUfP/XtDZUz
t5qSO2xr1cHsTvTVdBe+0c8oYWz4bkcRSPJw5kzL9SgRkt2Srcm6bBGRMOOvcENH
hMRbBMDRP/U2ixESUSgNv453wdJTgQl6dLyMso5nUDaWXs4qliRvCor7if6EYkn0
J1hDsr+y4MRLPd0ygcJX/nUW7t71FGvWrxcyOlUumMMQ4m0ezSFWWOGyp3/ZKKjw
29wbqSAk3EuBBpqwtCtlaPn+z9OMZbYeZ/woTEoowsgjsAXi8bBJ26ZUa2d+uV0+
wMR7UCcA0OkgO1zQQ2xqGCxkD7u53mo+zO7LQM8Hvmi1K24qYwicvp0SM2IKX1I+
HtbxC+ql09tL8V01bX7AYxFrlxLMfLujVdSbBYibIpNz8Q6oUVKG2H78b1BWxW8S
ggNxpne4dp/0qVnwWOVYGvm1InYnvU/ME8WEJVmZtCcUbVWigPMnRu/tTFgf5i6y
pEq+aSdlalm05gEi245YM3Cs9jOIDCp1CpnFEAox3MtgFlNeuRKVPioWn/tqmPFy
0fX+t9fGDBKXEltFZqYpKjIpbMmNeyS6d1DwT40FZHiC8VvQlm/Q40zBg/l8O/w1
btO+5wfY3A69BbdJYnuErRF9zxCWoBVKBO7jG7tGsi6Wn274yLTjJ2Sq6RobeXzU
xcBFGKoWyOAx2V2Yje5Xwlz2O++2f2cK0hsZJLsswFgqKuO7eUEQL8htF0ikHSdo
yQg0sI8UySoXWDJbrPPYSpRVIbd/xxg4PFOWvhAVYhPR/OgtEAI8Ebko5kx74+lI
Nbs1Xoi9XYOkeRQL63MgvX7beq9ySZzLJWNbr5VAni6Y6EpfVa6Gjp6gSox4BDPJ
KmUy1UhsQv0wc7Oio0dDiKfBJBTKly6UksEyNc4JX2cCDFzv48r5fCn2XTgYdl12
aSaGSSGoMJUPAgSFHA9Iup1agLe1isrQacn2ZPmCvwTgOs9SuIPW+P/UOb0GlP97
WKOzsXaor0WyX2v2ZC2T4L7tDvBF5xeXtp3OXclabY7coXYnnudTWx0zz1DgrE4t
6gXsigq8Un23esq0E5rSu5cRQe6fzsMsnb6gtzhCzQo/7XBahLlqi1D9GfRr5BPI
awnCT+oOFx2xZr42a100MIxJfQQ6s8Pe4Jyooq/dyH4t7n2XfxYZvGnmY+boXgXE
lm/RyN+VH3Zof3K4I96xcf9qygpxwqKiWJaEaP8M5joFC3VRyKeUrOQF8fC4xTkc
xZewK0mX3JXAzP5MsN7U6ctwLtR1q+yrckCPNQZdRDk/7ZHicgfOKkAUl2TS43cc
HFUySojq6xapr1+iYwykVtGXRJId5MxRXeW92nSsopmXJVfg9oZB0kI674rC6qBE
yzRq/0hZy6Hi9HAXz6S0/jp5IG7VMy3FdomcTnombZjmlGHJlCFILtuuMuLGib9P
Nv5MRL27Dc5OjKUq9fEU4BwSMadylCCub2ZXEVlT/q8lMqTPj6i2VrBqKe6tEymx
8vETc7ojh2NsKhvEL7pcKUgv3ospg84LbrtTJduoLi+5F7zkr0lLMpvtrT+monRH
9QpyNvOSdf3yagVffyO4ZW2+elOVTJkFG94TavBHFWQfP/g3yBNZm4T031RNpq1s
qFOjR+O7SpKjjNkB6GWN/SSsF9Hup7DvKXrbuEcJozHqaUzwqmdghAEAveCoHqqs
qwxXTirnJpvJ5tCFrqnSryCjH+mE1vw2t4Q/CxyqiFx8/7dpuoEKdXGIjEoame9O
UMBUFpSGbXNlNYFaw+XAbSnxqfwY9/pBwn7mFX2VPqZFba/E3A+kkLmbOxmX8fNs
6+qCGw5uaLFZMkxEqcFvG2eRPafzVb2UVtplJxC4VdPl6IJn9ziH74MyQASHYRCJ
e5aV8s3tZgdWin6H2v5QilxdVOkehtn6lN5AJb0rRDysWQIJyrdebVB9qlDsoXr1
6JbMwfFUxFKar2H0OzuJyyfhArSJMcB1VBER04Ul6ZKF518tRP5oE4r/fabHiB+d
0scpOxSk1VCAgnmyd6XXsR1I231f+eW2LTF83q4dPgfDv8FVPDsvo0DKWF4/ILUV
e2qtvNoQPpZRpHpNPAwSr5NkVzsmRWdtJbty2Od9JbcSqvloni2Mp187EjbEKvhl
PqEtMMDycyu9zC6O/aAtX1Y+qDUHBGxr3qw/hS8b0h8CQQyUbzR6HDZ+OJRIvSg1
xd64p/FQ3tIL7GvlDHsKFyAN0JkFBartqpHKs8CUUBQ9wFK/9NJ8mqAuEQj9tMPO
KSEZgOfXBEiYzzpzM+h4Hsv2bDfWxKEvagJfMU/UipWlPGPA0/gXgzJFm4RAmi7c
bZX6XQrW0tGhtuVIonLzr5j1cRxVIUYU6Vm6wp/9zxOx0DWgYWO0Wm82uGaif73G
vvrLcy3LgMKy4CLrEs/NAVRR1q9VSu+OOBXY/WcDSDykcWIDCVlTT5YXtI0RraST
UCj9WzLtGRxJHMg84kAiUd37tbbsFfBxn6gxJUM3r4+1atVol1mGXlysI+YAWf9i
WxgKPdLu2Rtr7TpMod8Knaj3QlXbzjyWCd29wz5iOwotld01oaRJkYmeUU0lme/c
3Zfsnq600hRUvKBjL8lD5TD2f8dsdXMNPlNZuH0H2SYc5Sf15UVGHWq7WwWV3zA+
2N4P8bh9Y21O/2dpDsgGUViUEZQIWNDe1Qlgi2rLzQdznihgnctPiv1so3BHa9JA
/zEbqQLEyjZqy/Ya02LzVTZHLPjZQqLSsZdS1OqG6Jvr/PCTnGv6XIDaOzyNKY1s
Bo3dMm7d+MutGb/Q+5/CG45xXBLPCFiY6EPGOfA3PGsHTILxnopKvmf3Ll+REdSl
yqUAchodKY9wwwgCjvoEW3f2cfegQCC7/RAO2AKw7EC41pxy+wdhIIh9KFTYSazE
QEFHIlKm7tWAbXAtJqdiM4liVnKl/rH27L+RBaPThhqYSs5Wsz0VIgbpXaFACevE
O9+qBM9PHebPM83/qhX5x1cqw7UKm6ZquUIvdLaX74P2Cetr5VVOhOBmaC0MUeve
RUjTKqoEFeEadPB0GVc+Hch4AHw9i1KaivfR+qnDG+IiAVarYS5e7Fbd+UCkpYdG
C8hyCOv2bjcDHIVrNhEfSa70ETeKaStt6XLLBtfQv1mjQDQST1WEZywQ6O/uF6ZH
6Wyq/KbxVrfhiwQejmdtjprxBmJRb25DMQzrFcYmncuYgN5BpD8FEWXoqFOZ8xMX
Q/sA/Zl57maTFSH+1KJOa75YTiK1igEqvMbERWtIz8ZKRJLBXOznr9GNfEde65M7
c+EzPkPlKKodk/UrJ51PzTNdBuloX2mEjdPJJnt0ZR2UOmNtkIgzqAG9mh9HNtwL
uVsPgtakkdvsEwL6vbs5hdjwgs0MOgAASitYymc/VSu1P1i+fKx/IL+qSoNVt2bU
mu3u7vvJ4m9joDJczecCE7e9Ft2iNUE378fJ7bG+bkW9UDJx3xf/X3o8+RV0fR3N
197bStzhzxr5pQ97PWIwtECxwrPKtNWRYm3awjDk3sS1zn0kY2NMGiuGhh2MsuVa
IM7Io8ubfA13ilR9ZYsZvOX0PgEC3vwen9jkz+YY4hmlqhnQRXsfPqd5UJqGOt3A
5YIyKVkWXY2FklU+J7WvAxRwX0SMF4B6/v/ctALhkBUod5hphGmuZIfso0svPGYz
NYQCvcUV8rb0uSM0JhNkMuq0mdsadF0ASheRRKk8r8h0HD7BOsESwI6c09NRc6hc
oWNyymr9GVC90t1QrDw0Xs/RkfzPyIqHLRR7sRf5bq1dn1gH6aIYQ5TLouuAvutV
rA0xU4cNQW1whkSKirQ0BWDUeU2OE5w/Bp1E9wYdY+ZyLMXTCUsvFMF3UPofiiTd
sAlaOeSyirjnYXt51slG70yN9mzN031iKbx+tXT4//4Z63bWvhmXcKkVYyhxYQjh
G+D4eQUsfmklr1161Y5X5zL2svXPtgkC2XPUQyYfibCMqgusi962dNzBOHlJtsTe
Lw5/TXjDTs0YiaY1in7bXJMwJh9aYFU1jQ/M9E3UXi2VBImlgc22QTycumRVlHD6
6/jwEQ0DM/HbC5RsRlob6EDO4w5sFToh3SmVCMfl7L/CdESdBs5D1Ht/w6LwtP9U
oLt2Kqsd1b91wGS31mVx2pOBAvJFzYqSdjQWA0iL7gBLHUCNBlldrzhdKqGwpUWN
6Py3G1pbiOi/v55y9lN8a31+quCFWDpazAF/Z3ckIeMHLZUZTDEB7/Df4/jKRT3S
wXPwb+oa/M1JiDo5PlPtI2UE2S7av/zx6vw4RHslpbbT1h8HG+cgom9CEFN+lTrL
xzRA2QY9c6t351/Trth5Yqoo2VBVSWm5hgBlcNovyN1M0v6Xr/wq9JHopS56tuJw
S11/i3pdo9yQRQMMvbfXXn6tARyOF8Y718jwGy9v9nqYi+1Vti8ENyOZZ2zZ9qVN
7KrdYZ0PiyA8blT8AAMy6v5gsUC2KYutVAItKGiFMOCth7xI1uOdb2iGsDsrTiMA
Ryicatpm5PQk4XD35jeAvG4gYL0tH3ar5e6CWkFkJlCYulZMn3ettssQwaQgFxxv
mrHEgaTSXE0elfO6devdz2QdtZe+2YCwGKmke30S+kQNZNUdmPLbISUOvibyiwgJ
AcZ+QFVBHihciF62wXA6mMnxE24zPVYkGnfJQO0kx31XxChhylNkGqRxiHeUb91Y
2veaKrL3vN8mSlUYbfAJ8leYvjTTN5ZU0t5MBdvK5f/G+tldXIvgJho/MS+qVoCN
DpRI5rajS5mDFb2v0nJzBOCNKS2YS1k30mrI80tbtDg7BjtyJttjojkp4Qn/2lFp
a7/P6DbIS+yHIAe/NcTQgaORiK6Q+PTseC2YnuVY0GHNwiGEGBahpHzKK+ojVI7g
+PfDxVhV2Z8ucEdKkY75ths3Q3kYe9L+G3u1rWbu8eIfSUXrvr3ejnw3hfRdv28o
inyeOQCKAOyprDPiT7wUuRNy/xeUSqt4blBhRtsTd/6j3YUoMPhaHqluJMkir5kU
ru5aNxp04I35rR9tOHnGXnodkTn5l7mDyN8Op+9KKLMeRHmCSNdGzjyF5OFfJUMn
tAuP9jsmu2uU6K6EEu179vhWnh4Ton/XDL49tdDZklR5f7HSFhmkkFSCn5TzLrws
yjLWIg/d83Af/Qr+fUhvlpqkiu5JXeXZ7Lx2K1iAGuTHIvVCRwlEs0u3CTC0XOHt
Jlo3Vj/7wD4GHRVGj80geNLpQ2tbdMGTxu69DqBAsjfl7iDwMOp2AQZJX6PSss9d
rbwjmXqTP0ME6wE+n2TaD5os872i8lcQoKSZsu3h20No5YAXZ24JBxUqgBpEts7c
fHzjc50O/JGjdYsYHoaeX/m48RAt/vlTwvqCZbGHeBCDAuwHUS/u2oacdrh1J5KR
kUJNtIXlg695usliEk8Pm2O/7Lm+p2VwF/2nhuP3BaUpLmcR+HgEEXCOvXU3F5mN
yfK8eurT0hBdxAorGDZc+GZ9ig9PHMHYBB0yFyTLrn2hiClJAav08OHuoQ0lnnW/
W1Z0LTLnfHa7E8ZaUz5YDEZ0I2ohqoOOgUOwkoriOIQaIuMlYpsc/ND3VZQXBeNd
HBOOzNXjejlhy7q1NwbbfglLqgaOazowUUy/xYVwokqXQcveDamaGd7OrlNjA4Wc
aV/DgZPwClBWx+4HmSnWXWgdLJkviDc7qadcS72dvYSAa2LothpnehMIwUIT15rt
5rkpef6gDPszFNET/uWtkVR4XJcycDf9IokN0Fx2YElOiSfFriWdKITjF0kw2ALx
n7RZNMNw07yZON/7C4uGvd/M8w1Sq1weivXmFXQEXTVfvyqcsVkL3voVO426cZqL
h3RF4L6Ox4H6yoPpGeaCnWR6IZjz7sEFjXRRbj1BwfZvnNrdnln9V+yWoLRCWXYw
2mAtWbJ/eS7MuX4INJpfY1ks2G9wwBJxrcQrk7OrMaL2gISikwCKtdPX1Ub1ujqu
L1IbB6gY38KUWKJoQoYRxt9528MHacqfhZGq4soW6FlGMdJRavM1O43TiRRuSZb3
5FKpEmIZKXf5xpOAzreRyKq3PaQQqbBxJU3CLCVyHYzWUqLWQJYacK1NmU5acXJJ
I07i5K8FPXPzByFtKj3TGrgfepcHJzl0nlIGA9W6wC28Hb4PNOvKRaiVzqMjo+Jl
1Mm74rmU4w6qw0zvNOA9+Ax17FXGEcfpippqkahcbx0Irrmc0PWJ4GDxaL26TiAb
CvTc/ZHLQ63jWqegVz6gm0yrR3c4oUUu7QCrXDOQg0E8BFXgN5BUvgbhN8o790s7
DrH5opihgSsljTDNVbcHh2uF+CtXpYPPiavnLwg9l6j4bC0/9mdemLF6y1sRAnxa
vW6m5A2xDqn6aezxG6CpfA0phWoi7UtCvv50NjMwyLSvuklwQ3SVYdPNBVKUBKLF
R7lZ5ou3G4/s7pNboOstKdPzSF6Tf9rcQWxEQkWgx+DK5BON670kkqKFUD7p13Df

//pragma protect end_data_block
//pragma protect digest_block
XF5Kuw4JjchkO8dTEK3RkKjoPrI=
//pragma protect end_digest_block
//pragma protect end_protected
