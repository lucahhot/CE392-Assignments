// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
1Hw6TZBlthgoXmnElEBfQMt1quk9kHWs4Zoi+AkVRPMDBv1ntQCi1rwbb1pllX4z
fJ5bQG8C/djfMJS/xr65dN87cJ+2TWdk548BYwqFEzuC332hWEMUnxyggfkJ7/SV
g3Kj8vr3qjcyJJy4On6s5Kglnp8G1Pl27i34ndk4L8g=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 28928 )
`pragma protect data_block
DiZfpRzhdABo1Q4g2f0FG+CM9anXFNY3of1LZIPxUazsedaKgvtLEwp/wH8DVsdp
0TocngBF3ia886LIMkT9pDNteqn+WmA4eYgVpl3ngy1fXM9ZfXFIScYFAPdJbW/h
75A7dSixQcGT2hUhQcO+s/IOEWFP8RFTNKFeJCv71oe06U8G49IbsgfGoD2crsuP
U36IsGeR5pU0XfoYe9VNzwN91EhDiycQFpXkQJptIa0acBV0wscjoewairVoJ+Qx
dFK0rZ4zsWAKwlUmvr3ibaM9KnbgkMwA8LHretuR28TOdaP3DlbMggRPf2HIfOSZ
1TV4cmZMAmacG9H9TLqoF/nOVLftP2tQu7IjCaIaeKTqHvxovSGPYMTTgFb0Ty4o
fqcUjw+fUzrVx/vErXbsDzqMUGjawx9FdFxc3DvWJH6io0TdB8K4rG9q5zDZNe5a
2lAeCnAnNHsyqhwqQoMCbhh6xbQljzTHhrs8hcoavvJrwo+E7/gFi0A88qjzjj5M
rTpN1syVZ8hltgD8ujXqunC1BH0FxMWj+ayzrL70Q1AvVsJ1UBEwNp30y7qwYIZj
SNQKwYTDv0hylvFjvppjt6l/VQetOwbpXbwT9xS1jLnC0hIJYrsGd2n7dcLyAG6C
6aCx8ySfkrobgC7Dzig9jNWTgiVymtFeiuGaR2ydKwGGY55Mj4cHmmfF7ofUE5+Z
qU+dUDvNaq+Ct32US1Xf0x8Y9aOHh7s41l7Nkj3V+8hMU7bpIUYuDbU5k8N1ysPL
8llNo5OMlfITMmQm8aLs38S6g1bP+ALbOGZ6Ipp70d0WyDnSGpEivAykvpgT2n1v
oFv66aDn1NzK6H2gAUKqbtonYy6tbDiGH8v/jtA5V2oG56xpx8oVAa3A/rkb67kR
U5FZn9DcRhGktEWFsNZfuMqGMm7uyM//wQDzhEhnbgpZiqfzmvdTNYE6gAN5nZT0
tQx3qn4RWsSkVneFZV2jGgwC0KghUv1qrTd9lhYsRDaJeOE5VkXWLlXKc9RdWOYf
pRUT/jZlNtIbowoiO7+Li5hM2UgkXAKlcwqIGL64+gzgXeea1wmnZkXJGMrQhDKr
mnvLXpMJFamY/L5aQ3V5yAWBWH6FT+alYdaqcdCdurv8geiYkHSkKLr0gFfJVdc8
ixFVTg1YhFLFqeBylJljWJKs0jASZdC7D/NLLs80kHNjL4/CsxJ55B+koSzO8JUr
w0HZi55nDCjHxrq7eo5qSgmwGCdZZ9Us3PmpbmFNpJbjHS9XKPQn75VEPkrTMMo+
L42/zpvylvphSO1542ca5KDF3eeFipqtdzRevq2yAdNvKq2t0ztklg6reNULfi24
issa/h5WvfC0l6vQN+mbSWA5pLIZ0OO07+WIy93UOS/4gnpOz6LjXmAFPNPsHQmD
T9K5UuZGoViuUcwoUGILxOczQPodC1owRhDdgAX/yWciey5F2OL1O7mDV2Jas0aP
tqOkS6+VTutTNY6v6jxzhY3k9rxQsXyyRwFi9z6FLbIIUOT2/zQHSMtFG/sqMRkP
adXQdRxRXhqht0zyemAPUiaNALrBQNJppbFvhwRcGnvO9ex/acNzwcXMKg7WQasj
uXFtQnc8NasK57YPq9FupxmYmA/CTKITMJgIYRh4lf83sBWQfdyHvveo1jlF6GxL
f/11DnxlVsLzrS0yAv3WaTluRpO6BfiPkzZY2B65xPNG61fonDkdcRfiDiS9fPAq
JmfC4xmow1tRYGLaVeLNpRVYpi2rl217AfJzpiA8xvmNqIpkcj3z4EV+UA4sEjrK
uG70np0NLCfSG0TkCxAd4T18JnFoopTuIoKG1KMlpuiU2gd00129P0dCtnK02LT5
uX5lXfTQteDSIdq4+L6ceBrmMGemKd/u9ZiKO38LxR1iS2jB5kUY8AI13HJL8n6D
Yn2M0Z+dzaxvYclWF3POAYYD+inEAncAx0bTOZ4S5yI+THwbHp40NULVrnxkx3sU
HjPj7rf1zUzwGvBso8TIGStdvROWczjOhPM7akDvjemDv6aKB1kfVQANLaSDAvQ6
8zURSpXbWGqVR06phhv6rDT+i5oSoR+PA45CzLL+R12HB32Euq1PR6wCXY74gngw
k7nnIcVZi1+SoHHqWqrXCeg5lDPQP3yHr3+ENJ6djpAu90jJWxeSN+OgFfQfzy0v
I/PiIpmGaJ9w6hKK/y2LfwkKCCTwhM52i7k6PGKWg7tpLgC3EuiIHx+24iMP2nwy
Q9b9h+u/J2LsYojOa2pzVfMn7eCF3XoZyWxcphEZtq8zTgmx9Nz7vn0o3MjFlzs0
XFcO4LtQS/mSPTAaNB2lvmLvolGRiueq8Inzxi89Ru4jyYX3h8tES5s5q1Ks3wnV
+ul+TAFrkSLJOFUxu+VOpB8ELtlRxvclwugTbmkmUvSuNfIAAcakJJRvX5uQ+e8p
wFSp3mAoyyeveIhUbiOi2Je8Vrk8GKeRcGW7lEd1VHD1xIAlV134wDXDpOBvP7Ri
8r+of5vYiUHi5/dlGej8zubxgh/NM3iYQNCoj0/Ggdoc4pvogJdxHiyuPkh3ivRq
LzD9rMkvAEZhLOk/zA4CLIWesQq6cXZFoAPtoNQZvnXcKRRSc2nzwaOlb7CvNcDL
bh5wkpebrCcONFighf8gN20PS3RsWRsmRVuU/LLgdy0t6tbD14+6kySZ62pMa0zd
3kYNT/5twUcNIfIjVcVowZp2BMUsBSnebTDAwpK9VjLbhK9w9BDMPOu0BovNSYs6
DfFAyo2bpC3hWXCfixKOnbMXhT0e1n8BI5/IWldpzhDVnYjfWhOGRs0rILXYcsWh
/qBQbIUBsSoJSI7jK46VYkj1iHIRg5WzCJA47e6wdrtRkPXild1Bmx/QAXXoS19V
FQCPdej7QeqY4+Fj2xgRpe2qsdHUEgFFNYv19Jy21dD9YPjceBiPvfnwAgDPaIJC
BRXzw3vzo7qT3uGW+hUT39K9wO98vnf1QHuOtr2phGviwtoS4oe/y2LhzDtOO958
5bXPkN26YY+2SgBo7gANPDy3N6hJj9JgVzFNzrN7Ev8c8/Cawv+SQcG9rqC2tveC
cRCd2OfdgIkC+n645ds51Htj2sRxj5dBCUuqKQXTiyYgtdzEYsuX+dtJT8KaIGTf
bYbzNeOB8JHiSK2XjA1JYOPcrK2blhujkQ3q5iBSueskINaPBBQqaMrWKiwawrKY
FzO/NjGgdhy1Fv3FxKakSusTanJI4vRgExVWJStio9RERqhiMahWawQkX3u8VOp4
T5NqUWsAXXwbyIwvVnAxn6EfcsrG5Piw02depyX7boYXhQActbLiwy1vVPVC+UI5
Bvjn2l9IXV2X8PXIG31EWYjeMD5KICediv2kr+0u4nBVRe1ROgXRPnz8nkhku6Rn
ESW8eSprvivkDgth0x5v+z8KSQ13/nA0moc0/TjEMu7SInuiB2epqtppsTvFs8+X
JX8juKNJH8xlqDyusYTp0gG1q/eTF2ItJiXs2290xB2/0HVbHTmj/TZwRig6Y9yR
jIRv0h2xEw2lk9pkyQUQp1RZzWg9v77lCQCjdZQ8TNpQsMxo6/YEB8oThu+6HM41
5NId68xXIEx1GpvXAS7IvUH2ux6fIQYfQwUaZFl2/KJzE78uWXL21J+CA7RA3iDw
CpROPmWzcIRmKfmwLKDIAL4nb/lDkoUL8SNy+0MRVOgi9rPSNq/iKpRaOXU4k+4A
8wO4WQG9olkBmYjeHq5JOiBgSOGCFFalpEF0pxT0fx0sRYzx4q2hhMToPTXylLzp
O1hBEM79HuzkJL8bXVLpkZT6HrlSCxuHdN5dco7H2Q/M7mzY3bc0KjSwYesS1Ekw
dKMcbRd/+CeC/NPgLZixLxTUTob2YAsPHycnNS1fvr+15rPISI8BbuACVd+f4ugK
X2grzLkK0nxUuuo7oCW/Xd2+cLcFfHyjGvM+zFjpknmGajaQND0C2JDkrCdg8gwC
RlALhIpczgP9HNyaBBc/a9SQvxzx/w90G45KjLS4/SsccNJTXkdphhQbLpe8GG3f
IaUU+LpjaIO8Wz+rosE6bVL5HNbHz41tl7eab9QxhRG96IQlQg1TmLb/dDvwwy9n
Zkt0IndQhgXZjCZRkL/sjVByVj7MEfgaskYzW4C8qonwDqeH4wr0dNaz/QYh8Pdt
i8jje/41uXcKIknIlglwT8T4c+DSn5wnQSBqM4oZuIlVOVEFMe3FuAR0NzuzFBd1
0ptBI6wbDBVrCWF40o/jN6PSk7Ya3EnmDdwl7A4fZXRLar9ZWjwVm+TNIN8MzpbR
CBfeUgI5pr27EbvdHHnLBSoQfHHUETPKqFhEoNfLHCoRsR9lzp/gaXM+3mRxHjfS
SycOlI1D7HS9cS+L1oIwZ7nhMemTLqOpeNClE7UUMIZP8hZVHWYMZi98fZ5/y5n3
QO7U3UzO1cef5wKTpExwh5rxA0cZX0HkWrN6QopHLiutX9ugePyXWRuTJEwZTXQk
PaCQXcXQPNg7O1lv5LeniPJVtEEXdXECuPsywRrMkz6L1HF4e6Ljs8ggpxSIwROM
kJftNPqpffNEK35rEOU2wOXjpfV8tCrHlDPPsZOz4KuHtOa8f/c+mAVcRGkv5E2r
efyVlHdQQcZXGAkFTl6sDM/8Yo6aseunJ2MffoCd0uEOJfyo2qjR0+xOgZ0dYbRu
kXn9BlZzk2pSCtjYJISgUko9wYVIM/ZV81+XXolCb6X+uAYIO+S6lkEaROjpRzpc
Z7kZ6YF7SrF+DhW5Hzy30+pZX61hUboPGDlvXOlbUeCPUiU6Ig09FlH8Qusu8/bv
9ek42PhsuTCxU21GdfThy8T+eK6YhGdZ0+0SZ9O7X7Fhw76o9aAsYCec8vxfQP+V
usO5vRgGhOkB01HHp1XgOvXJ/IQviUoDQ01jTYw9ya7YaJsHFvPUezM5fpy12dVk
0mvVk4jKSXFhLGQPWwTy6/lZNLn7ZvikB5bkhHtCnjBecCd+jiDSKJpmbH4oTBDd
6IM2VQwkemCPmmg6RSCeEUB+7kfcdgNqzUYFDQ13a8oN0+xrp6qDVIvJVcU1hxp9
U0xf6Cwb6mTTmP9yxFSdoSOUqHCGDKKxrcSoqIXgail9K/berYLPHrSX1N1HYwPM
oIhNDCQAHtao4FJkz8bWoOAAVQ3DtiwqtCSQDXcoh9svQJ7pMZTes2MF+tUJSpC8
1TNxC9Q073b5/uhtgdvZbwNFRxVvPCO93QTBys4zTSrxV3AawrBioBPcKu5T78z0
KGXp9vyT08yVOnWjARp08IZf4uM3rMgWXYYKz0rgJzcH3djZPevCfWg8WR0/YZ6K
w/uN8AKL0Tt6TSCbtaDsAGsYFK2hpgh8e219+6iaS1xTb7mZ8aMRtxn7+qMEtOEO
VbiJMVAbWNxPgl3A1Hdj/90pdm+QaZ8GGs4ljosacOu+XRdTsfOaI+y/D+vyEzSq
b1+jE4dlpsc2zlSwDXXuXCT5FQMsXuzul5j3ngdFllUyyhijSe+zFr1bHBixU4UO
AFQMayENZ4L708Ulp09jpqd1MlRJAkHE5+fHAm/53++MJrmBNLH5IBxfy1lXXd+t
IuqD4JbREZpn2ALBJI3wbveW7c2v30sParlBGDM/1PQwlrWDOGJKuhf16FND3Y8B
PX+OjL/cf/T3oZ5wZ1S6ZarTNLH4dZtufrWmI/nrBwbXa1vGLirsGr0Rymw06BHG
wv+JEj2LTTiF0ntLoVZNiKdX1dHLKEZT3/H8NM802gR3vu2p8/MPlKz6ptDw+2+Z
XNG/oslk7NLP53iy8DT/mXkP/RsCV4wbxFYwzluLQzwTbtn5YZRmBPvAEYkcdnvw
6NMHAbVgoA3FXWHYRrkJgF67JI71fEiFXQv5FtpVqo26Vnri1APdP7kY1TUrRHoE
NoIYl78WTM3NW7cCgTl/3XMHB/mkNqga/gJp6cMzaAWsxjnlonqxDYAWwYhQURvq
r4+skYzKa+ggXHMv8oKnv+IrI//pEEVis9/fb7YRUPhLR3EUE3Cdo9BkA0PPfHNO
JEBhM+HwcUCFDjEinXnIXlCm8PgQrQHp7EC9XUWox8gkDhQyCu/WKCHc+FAtAW1I
NlPdRW9FmrtydjBnEktcN7u8OeHdh4WYNKR764OlUtlG4ATKfkpfTBeyiz54uH99
XAoXACBRKsGfV4tmaG4gK+9ufgIRr5lZnEXkRnyT/G84A7MFBr9jKjKacXpHNP4m
zDKXFvFh++tqJNaya/yoN+I3P8iYeAWK3yxlp3sWuvcJJZVzaYFfxvYsmXsrtWQa
AOwohCQPrADR7Qq3TRyAGnxC6beDkCRwFZgKZop3idWPizBaCAfVKsLJ38RJlx4I
HZ8zPiJx4dlNtt4FZ7Grn6LL+byBi9lFn5wlKcJHaM7WLIfykMSGwRkimY2kp4w6
sAV9mHJqpdYL/7Z1JXW51MNeZ18WPA0OH7X7J2/el12yAtPycvF8EFLxecU6XNKo
9h3tQ5A820Bmpr8Qx10plQlYyg53inS888vFVyE4Iwr7cxTF7389hmUr2RD3Zdq7
gGg8RApY7uRVtO6NIhnFImRmNdNkhHXeBQ/fPg1WfvrmvreNK4AZfYRIQve2+kIG
X9scJMH1NuSFDKfMmc3QUwv6NTYToqUSHEjOsc/QjocIItJrGFXu5YoaaPzgc5kd
Rv5kAm3wNr3c8jWZoTC/8bUTUUE4B/fOPdbKYrZW62xRcB45PKKlLM/oQdBsMDnU
UK49BLkLx4c5fLUfNZcZY8zXGlNRMhtrqWtuO+WCYF3OOsvoUowJtvZhvaJR0eyn
kWrHQgXGqTRrDR1oxEoEhY4iO98ThfaZ+qg9Snrv52tYlLqzikPomKHYlgc10dqF
FPT0wSLHZ24ciGZJ1RAXC3cDoo/5Z+OY0wS7c/AjxeRxFmcj06SPtlgYMxAdQPgQ
oG8cbR34VgwXVooNoew4uIxWBKSP/PK9tT7NKuHLYGzW6QxUSNkZw6kIsX1DzHco
ifDEcWkzH2OZ3wp2I1tKtp7Q94ABAaEYgN0hJIkazwGvzPFu8w/vlV3qzXAoxmn1
wxPA6W7gaqNZs2leVcCkUri5gj1YRdTlBMS5Ck4lcGsf2mgYeHHlX7jFIN3BLyPJ
ST1eBvm+C+f/ZYjh3N8io3vSbJaDzl42l0y3np9KdmGdZO3Q8I5vLJvRkUWqSz+o
SC6PhUZ6rcktYYHFrHRgQ1npphTZZyWPf00tT16NuHLSQcDXNqQVhijGygs7DB4Y
kJvYOpfdZkHsZ8qtZXmL2Fi2GPGKUuZZjWBipAsVDMTUm+iN3lijPGAZEYYzSXom
d/jvz8YTvlqUG/4m+mTV7PgkYI3LIAJPzd2G4OMyVKlTfrcz+eDjBpLKA4OL/TO7
/+USJ5d22S/ZsT3cFypCQWDH7If1kdhV9TOrkxriSjU4YVUl6+rQ+Bs/4LkZLZxu
EMxBzp9q98Xv1Ip0Xc3ueR737pGZ9vIrhFsfktycXlv3BGU87HGN1FhEevN+jzZY
vgrqneAsDyyT5Jb0obafleXxT4H5BMnd8G7cGUNS6A2yGPFT/l/vzMRlNx2lYWCR
NC3oFUdBaauIastyusV53NkuQnZUj0sgWXvdR2Fl3MU0opHndBigrONFbBdad7Wo
FDETWkFyixbpmIoasF1LqVxLxlscX8UELY0fkY7aPQouLQEPFG06RquBzhrQst/L
NRyTaQRhoW2i4tkmg5+FAel73Do2rbAmC+QMx7BJmrYQw24n3LQJpPLxerIwb69y
lNCBlhmU59d+Sh2PntcYPQiJ2fWY8jsSh9K/8GLgLtX/l/4J61VDljEe4NYaq/wy
Fn6i0RiiUKw2VtACtZBPQnDD4E5Xc0GmFnTu7mQQSfW4VlolUszcWcKtv6UzK5N5
Th6Hijk+DF5ufTj3Ldp2kUcqDXx3R35WokpTMuatl9Kj+NU0zS2PekCE3Y+MBJ/M
lAjNFaKdNaIrey+ZFnea6TjtHGEUICe11y8/f2/jyHpXbL+XLKhyOD0Zpn1X3281
jGMx9ZFv3BTCqJtG/B6/LsoUtA3/N6FkfjSgb/fLrSSAa3BV2E9PZBRhSEpQ9f5y
UZ+BSrSQcnVJdliHj8EGldjdniTULHcbMyQGMshBxvzlyO32jefREr6Qq6DYxsEX
c61lDyvboZWoIcTg2Nr/GbFLYv6ZISZgxHOKJEG3FP5qO/Izdlp1Tv6txx3yFbNm
JZhrb81Ep7d2VOjwe4/LOQ0AgYruc/9teK7iYQAOMSsYopeoVaKiTtu1TADrLWKG
8bNtLa6npjulReoc6vssodhHMoPerP/aNfbvOlP4cKltDCdwB82FyCDbQtRj/xup
/1hxoB+RkPXwJQO7iK0jhAkZekVUxkr/gV+M6rFRSOOZ3KoaTL7qJ0F1E5CPHN4v
peEsz3PwPk91yA/spoCPF5YpAmMFUMxfzSnlsyFqKWTNCx6P4s3Kg3Jr6hzQ54OF
2CRSB7DR9ihm9rjRMOSZlY0QjBLSLzXS13XMxoTd/Ompytl0UE4ltn+8UZmZE1Lc
ao7/sr4zGLcMIMukp8OnP41PLG6FECCjYEVGWdJoq+gqm4wwE9RKhb+juHalB/KH
Koo8+n5rVHJHundkg39zthTPe+SR+nhHYN14OkPQMm4GQWPcsGZDJ5qyhdpc5jcP
ru5i1cg8XsMg+FGHiVCDRSaD/EKSbx0Ke+kumv7qHAQCry4wdVQ2D0EfuDfflbkR
WTqpjMQ+5XBO0/rmjqFCxzpY59C1i26m8dmHgb5Yq1BBc9rVv6UjflY0vGfU7Hka
HF+J7XomzDDxFsAjOyyQTK6gotMv9Yw+ozpkM4a/Af6cWvZ/p9DD03MZIohiHgLY
2nBNIjUf8eGXnSZ2ZLi8SO6Ym3zwKcNJTOUJ1oMe8oDWtwHsQuJbqE4xQNErkA1Z
y+UJkwO2DTeTcW9k3Nzet7Y+ZZl3mU9U4JwYjCeTLdT+Nh8Rxr/FqofwSbGD3iaj
wZ2yZc+8AzU7oY6Z7jFDilUnuOp4TU3Dw3xfti1GUUEBtPTAs1HJ9pRXAbjGwiTy
gbtRff6EGIikl+W3By8NnB/hQwuPEte1w3i5aknm1e+h9niZ5We7CteqdbaGjpH7
FwWEtB+qSYLYOuHxX1kKfOpuij8y8Lm8VMR7xfi+hFp2AHFHEZzR+4RfvwmYg4Ds
MK9dAUOJ6c6HSDYtPk6uRhuSNNXdPbnrBOYkPLFg9p4LGys8t0S9NdsENi/OpW5k
DVz9cmHpOCqVcPSJAdC/VcZalged1nkJNxRMR9eT/wO+RR5VulXYvXq4RC4jI2Vh
CNf3ukszk0WFoarkuj7HJcbGUy8uB3R7gJwo7x9yM9VmlxSD+8Bv93DZxjLZtopM
UwUF9PmDclcXRfRlPQc6dlMnc15gMdq/AhWUkBc+lrzHwrpxULYxMA+dCvij2URa
yJyW16CCFi9NW4/lASF5d8o0Gy7c3RRUEWCZOtXYJil/vBTCdVZ2WafEIJ51Lm4h
iDyDN+whkiWwWNqC5+6+yE4IAJfdRyHBn7NUtEQH4APtOySjA+MCuf4FhSkWa2B8
lvmkHyETUMyL7bCjl4eVTd4oNScqQyr/HlE2eu5nENoj2tGbigPXpUazB+G+e1rt
RuueyAAg38wYLVL6odJz+Kpbsju84CcC5J4UMx/xKwtWB4q8OIkASL3lNwhllFxH
Hdr0HMXW1xHjquOQzTacYoL2PtYiUUD0pWzlEg5VvZFyVryTbO6OqVWKtvH+jcgT
tJ085yi3Wyncj/MIuDNSDgRlWym+bIR9bTUjMZ+JISWcGOprMXnBrbyfy7x4R84N
YNwUrF9hVZTjW0s1/j88NfJ4GH5BFSFUFok+LFm1ZWpjaAd48ErmhTcXOw+Httpb
MiDzUxXX8Yr6hTffEsI1ywxVSqoYCB+dz/pGVKALNPp54W3BdUdy7hwjFel65i9a
Y2C3qV5DF+K7EZYOqhT2TZ2uZ0MyzRPz4T1diGMY0l8b2osu6PzDELENVqR2qHiD
qIxhEeAM4DTWMy+60+L4WeCELuG9h0g6Oz/kLucqB/Q90sfTcXz0C/tM/QEQazj6
5sJeDvOzA88vxb5c19/UlWGONrfzONTzWMRpEf+lSc38r0WlkF2PEg+Wc72XIeD4
GwNDShAvgpKrilul/1SvwpexaPnBPX2ih4GpHniMljZ9uOYxOt+tT/vSFuDfE+1e
9lerl1Skqz6i8EGsUWJCHSFiGr1NiqaFcZ+tGNbepWrxQYiu58rUoPQB7qK85XWW
VpT8uRC4jLqrd+U7ZB8V4wbWfA6w1229ZkNgetDhDRVdQnVawkHeKpcR0BwBYJA1
eNyQSj6FYOo4kWPxas8JOP5PntHieaZlkn3QGkfJnCAQS9d6mpvgF+HfWx9uTYna
XCJ8mwadoOJljWKjah530l0bhaRwYTFcwmG5sYxzOJOQWk64rRhMMN8f4cm5Ewz5
HBcDfMlV9MuapUCLvvcTIJs1GamT5HpzKtLmsG/pq8Zudt2t4obhgn3CeBwem8iG
ERuipHvIRYKyW9nnlup33yuqQJnC96toTUMG4/PZgF2ZWMSrCnEdQQGOaqgA/V9h
Mpvus+Ks+Mmb55g9OYPA5xU3pRqzdYJ2GradGkMx+4AxWCMtbQcxPh7Gq43zYnwj
Nhc2YjTyhQsM5m4NujF0lvlPcg7Zg1ls/6rmSiU7zzHPn4OOR89NXOAfIEQvgiB/
hqd1MkNhAsXe7kmeOHl8BmsmDJkXozcAbP70qbez6ytAlKXm6ni2G9/M1VAD4msK
pKirxIf/EtWN4V1IzhoqKHPVogmBZYqe0hR4Vk2XLppuI6jyeVhfy2LVaORQSDmb
y3ZCtLDO6NLhKuuhCwmkduBza/Y19NVS2ZRKOYPZu3bIjD+rYh9VBMcpQSHISN39
3ZW/lskeL5DqNOQS63uCW96itaPYCcIfLUGNZAUhhsrobAentYwuTBIQMI0+dnjF
2S1htOxWDrN0pE1Z8Qz3aEb5e7eI7RFHHWBoV/1UGPRRAYjEMEuuYWN793C2ovKJ
u14TQJ3qlMlWniIujWSAH/kTjbaT+lRgQmz9PpyQIdXIfn1MVwSb5OUjWHWCoxgr
wWzPnLJQc03mi9Mv80+dDiMHFjD606l1nPpMF/qE86wxYC7lPR++2DIlDWaykaQ8
PAPUlmxUTkVAn/FXjMhOwGlm6pSqKCds7TN/DJxdLnXGq326/MLm83viP7BgTPRT
bjMgr5GKnlipu8PhqntRk2w0YRZVSRiig5mB0WGiDr/pa5rSrwvtkn01jC2cfV2k
56CKLORmJC3Blp1xh+fPonT7RJoW+iIhibdI6sK91aO4tRrTzNKprT9Bw9uobPFY
AWer8ZiqzJrofB3Qpk31R08ytdZ6nULSEdOZEt/xRh8YTzC2U5xBe/nz5ZScTcgq
nPssnDWTLE5geLKkNxVHAF08a/JE98iTJHruUS4BQqXE0imeJ7y4jIHskgp4wKC/
b8aahZJetG2dQn5cK6LxvpLA9hAQErBoUOdPaE0jUmit4GP/fB6y47T1D9NRcuxX
G9ClwTRlig8VR6adeoOr/+ddXRM7g2O0my/Xm5KGTe4ucQ1C4otUqOnz4e9POAJA
/QldSnKq1wCPx09qdRgfqhsijEsdC63KKokOQgvI1RVUx9OQhU7lncCeCTuaqslz
m/5OZB/LuWiHQjTy+SfFJvs/6C1YoC7dUO0nTWGOiydyb8M53ICO+wFihu2zEHKo
d84W36ItFnVC0ByApWuD/beLZgKF4cOwdMdHJ/TWwmuT3TTdHgEgTeB2YHNJkSFZ
RFc2trNZ6Vp09rfWLcrMSuL2HZqI9OaSvfxoH8VZi/So2/VcqdHyOxYE1jjl94gW
zZpR73k2W2hcnRnsRfZnZ8RJXRdFW2IfRq1LE4U4YWtph0Fx/BWVkr2fKXi1+NGU
lEpdeZ5ffHC/N7aI6Y+RicwXWfcPOKdCt02a/zgEbOpRsu5M+Rh3xGs84gwHoL29
06mxP9RiIPOInpUBO9aSrOBMOWJlEgxXfOoFpGPWsD2aziVrPhXW2qSqOZRChwiX
PNYZEh7zTi3gEnA6FhAHncGCxr7QFJ00wisFmXBbusLlYzbTtPrMaLs4lScc6sbT
bEZk1fLQNATx9TxLdLIFLfAOsmL8eoL0mTbhOV88AHluI6yovfI3k8AbC4luiauI
BCXTRQ+bZnsmxsfh3chy3BZfNupDPOsdvvcICPmI7zIZ/hZ2HWNYBOAcOmRxWjwH
POGdDyIav4nNyK0sz1ATnSq1hJz2BaI4p6JUTovorhAJf/5xAxJCSY/rZ2RZ1Xk9
90FCPxF+WW6tH/jtgyqiKDEv4GKtdW2njoIz4Fwp4UwIr3wBXe0s6tDH7/hSu3Gk
jhcITK4ULRf2OJv4g2DSDqRbBZem/NrfvQQroOzuUW1A8WMNxPyhzGUTCi77xWMO
ggJwzFrPs6wD1rJaCtgCJ2OQUed3vIQ7i4PWcYaTVKzP3YYKdbsy3fh9lTNf7hb2
im5ZrG9a1ap2CgC0WrEFbCdDbWbgtvkIQE9oyyFDk1sDiI7T0B6lGYtTKGSN89UC
XYjaUjYjGd4qn9HgxdB8nrafkMYW13v2x5Q1/9LblJRrlZkZpYpFttvlY1uzJ1od
rQ6Hv8yUb9FilUpH6HnFzVCTHbEDsH5mznKe/T8lkyKhRmLl7icEidqtUZP1H2jw
1XvETMyLNQBnxlzGvbGKwIETbOLP5JPPyldXmDYCsICB8MDK7B5Cy2+75Tc4E0W7
VlDUtYXb7UVG2fndnBGFgbpiQ5vWrpYcTbgBYs0ZsUd9jBHHNP8/FnsUrihnoD+i
XDxzbYnuSMjO1AJoGWi8gn+67MI20u8FZhrDvoS//bcIES3Zf7NFgp5QDmZlyFdU
5b0NKc5Kaw0O27yHGCPnPP3L9J9pJoO9ZGFoS8KKHVm1IxceyRQ76KpkgTWHyP2G
xhfJFr/qbthxJlZ3uWlhd9xxIRv3hyOMq0ETmXk+57DOJAjBMXg+NX+04wFQVNKV
1bgEsvpCZ3cjnkZtrjQtmfOSn9lSFoYepmjM6bDntz27HBqHDknofyXIuGtGyNhy
8Bxn+un8ZRLnbjaCGoghbJ4xBN4gRB94Ebc/3IAhnGO88SM9WY1NDJOtheMBs8Rf
IsVyYEozuUwuB9gBUxFRIXv06t7HhEYCLvqUYx5b693qfL1yZYfM3PtTVl7W8q2z
+DhdFBjAFEosJv/AmWVAiJvQmUElPOWR9/kyDyxBxuzr+u+P0VTNYtprVvKud0d2
vb+8Tm8zgomO9HltgNAq10mqHc1iYcb6Xm4ebeSZCkx6StV1VitZyEleYdJzrD46
FOB1Shc3vPHhHexHuqry3PKVj81JPDOl8P8kNYaKah0d7nanR2G+qy3N5LIlbzoW
ZITVSGfNq6oc5rkjr7QwewZBc/53UIYN/tA7sPapeR0swlPRbfmXKxvZO/Cu4p5p
X32MA+y+fIFAYhz39QeSGF3S97bxUKimqdSj0j1HQwtmt2B0f+3JQkw5GDVOS50o
jdD6stcx8eHlj2hGYb3zQ6d1wvS6kt+C8jzC9lF45u3lTRWVSXnxjfUCdsosNemI
hvWMq3NvmHZq33CJ+g5Lup49dxHbJGioTRtJ4ctUCd0hPZZ6ASrekK6KKI8ZzxLw
ueEVXDMMKHKuk5nPqWPnJ7Om7jB2Kvy/QfqdN/xJnNfC/LBfk1Ix2LzsPLd1qAnp
wmIQ3ueqJVOkItiNFePudfSpAjcLnsPkvRd9ROPFQoUUbZHaWPmtk2Kr1+W0ymit
l58ySo6E/Y054Gtd6Bxc6aDEFKnPSEDtEZmWyth9ENlIVcdb9sS/pX1J8b83R0rX
flmP3uVpkd3HIkhPEoYMuMR6quUPCsu5x+KwXjYnSHUFQiMncQPE3RCrZS28Ou4S
HEmdln2iGkBii71XT52276mMSaz32s7R/d8yNXDZTJjt6p0updRfZSjV5swZggCv
ta6rW33i+9FyeSzODv7Iu3qzxygTV1cunbl+/vpHolGOh0wxVfT7QjzOlhqPchdY
JDDOxRiZXq/AdO+4gzStyrGL+/uO4tMylY0ytNuDqYSwMGAijgakEmI8hye7U6WT
jhErUyTVaDrQjR1XxygxoGTU4CJV51FdKvD24a5BTxIHzSoSSm29FTg88KIlFzCt
Y/lJIVCn96fIMfAzNu///l6MHNG8s84Lp7AKOe2HdOg0lMnUYJNR+6Lhb/ctblFc
mC+2uI8DLblygYjdzfV8qxj4f7aDKtu+7e1OKSVwB7VP5r8cpAyVi3sjy4uOZZiX
JSoyfXfgbdEoc9SyyF0MsVgeaNc3yI6i46jv1E/BrEiG49RauXRaIQIzJPjs4ToY
n7X7+3cPAzSbti6CdCYEj2t9SYLnQbektOCkdBIZOVuUVyZPVvLWjif0UYQ73Mzl
fNKQjehTM5KYyyy2/CLyU72VjXv/KpWuMP7daI2ypH77ufQXV9tq7Gi1uuKwSwHx
KD44TOwdeoBvbcAWaV+Wgi9MHw+peh6jNSgaFVDKrVuJa6ApkNDphi2Gl0EtXXG4
ANxxmCw055KpzIBRMbxXQkeQ6QH3yL/No0UGxqcOTJCswcMas6/O1v/f3i+xspvd
kNX9AlFgsGZ5W+d6YkXWPOhmyh+EzTOULSf0gWX8TEAhfnxX73EEY6OXYnQXXmQO
xIplwmuoIk7zkfo8t5TjZtUFMVSIpfuLkiv6bl+oZ+0oT5STK+psDWMRDPETdr8U
KsBWW3ZpYZXR19cXkdmYmzJlC1LllRdSgacYtrO1V395Ou38NJ3//jXKEIcpv6/Y
zSBoSTqcFQMSl/O7GzfLjAfX4BQLb+29HNUY9x9fsx4IkDeJ19uQBoRNXA7i53AI
1uUQ9ue4FJFtXTE0wyDRmOusDtV2zuo04VcMvpbNg5hvJbWAnWbN0YPIa/Ap7InM
YXTPChk0Vdq2ew5HzLRFiwhhyQYN8/gHUrZHNIm2CM6ipnzW5c4EKC7EyJECeWHX
CAJqbruujKEL/jvPXILNwBanghaxbSy6GtIbeJfPSAVKrSfti17a3Ic9RXIaHO9L
TzfTZVM/JSpabkkquhx67tILoD4JUao4VNoPYHI8OIwudWjmPkVfXAue4MB4iK+E
hJ8B6rurrd8vehadXctwAtsxCGbrchtbUMj7TwnJTnWLP4L3bEXWq8bzCGreyufc
3vEcBlGYVamBxz7/UmIcLg1QQDfjFEDUJvCIEi+wbkuMQwFsKPxLi/nsLgpFo2Y5
IBMWVk1f3RfTM531UnjTvMNjnNFVqPOiUUFkBztLz68bAT8Df/YC2XPcod+gS1Ys
q6R8Uvvs4xmpWUVKi2hBlKVLbvgRutQ2vgZgD2P7qVdc/XQVq6quSd2ZM3pLIe7/
SyRPEJUyLxwjYJBpyYKchPB9/vq5ZwXTuQCBn6eXAGBpMsEW6+aFENqLqztefjCP
J6fUYAEL2sThaSQs2YJzEpVNllpdrarXBW2pSib5Li6/pI8RwdY1y98AomqBw9ED
z3g6hrf4hQJVyoqxD1COqaL1l/pxCaTs36fKRLjVDhiHOR2O5yEFGzQk4k62kJfn
X8CFqz5mYCpn61z4J0eNMtNWNNptT9SR7ylB5x5fOVbnTVUgApMG4b05tKNkIOUR
LO9EDQCa33rIhyHFzXCTJkrzyS1WXFWy926pC+CZt3i1b1jSIZvjbXIiTOERjhwy
hDGSOc8KMrb27zej8KAYhdySbjxlt+TZXmv2dazRDScf07+i7kiV+Ds+Zs8j8hMF
IruKGDf3mWxFOEaFhqYxaPbhdxrWms30RfD2XGKwhENMGxOlQFV8pbvn5kWYmuwc
/I+I036jojAY/MDTFFz6bVzZ9rVhfXk9RmTkSnOEqIelWZ6CrbDJHuSAuBFCQYIU
yxVbwBtHFwmS5UK/oOxLzS+JkBo5RNmYhIH5Hz24W063DVU4zm7MxEfLcb3221eX
YReCOTDynrQeWCx8OV5FLUdVmqmVLtJnJ4bBrBELNcjsb70YvyGO8tAituD5iFc7
Mc65ftYZGpu2WCfPgNOJnNazb7ZE7KpOHxuBv3ixJv/JUcMQPHdh8buIvBHqZZ95
kd+NFrtLM1G8dpIHNkivp0IjtQ/xRkwBzt7a8NygilwtjrYPXg3nwJKq6zQ58WAm
8+IjRnYDt3gZminxd67jLAoI8hlcy9s1SoJooMP9kNcS0Umof6xY607KidpliWuv
KF916K7FwYpWvofZ2gX/OtaMKQo6RMj+f15LcUCl0jcVyJZULWUIkSchP3by1a0b
rvXsrnNkr/D79HhOuXMabGTz01dq0qP8rTwEb/693ZJg8xV+jm50899Ze6MC60OP
a8DVlYSQm2iXOK6zCxKRCp+dq8QcZtDID1gxr2Ng4DMnQSdrm+ipNOQS5z4VW3rP
ckkdAKV6tEY17YXd2AKGgp+1TV3YWETp12dI94a5JUlNA9ZUDapIe73rwZ+ZDghE
5mPjlYlIEqmeTOy8C8cYYXmfIhja4PHe4+E1ib0RKLnyBQxYsstkVpUzOno4Ji4k
OOFyil7NTojX0nSOmuQ15zEffF2ouUVzf6ZzkH1XonJwa8+ESGFHZjLnUayroWCf
ojC0GF9K8qZ5KjTKCanU5RQ/vaDrOAaY8i3pWyobbtrUuDh6Ynj9XDvuSuch2L1t
9ioGbL7JrYp5tKC3sv59b29EQB6f0tu7S+tTPN4dFFEhB6vekoCn7GfL3EnOi6Su
GTHJ6+ywzGOYTPGpqqQWXCmtt9FNYP0g6NqmjKfQTSnPl6Bf/muiKJowHVnTgIhP
hhzDrq8xZT/GTaAyh2/+8xHP3QKCYurSrmWVbR8tnYQQEFssJzTTpqVWF/l5uvrs
j3byjqzqAm1V6+CiTSer2U/mQfvhZ6fL9UZz4Oqhp82r1eTjafFoioflJYhG6HW/
RDdKj3yrnaLTBV+QgiFbGQd/gTScAaZHxDQ/Wakxa0andtPIdlOhRfH79NrbSUQP
t8dFD5oSxb1YtPXT/t0Ly97j65+MjOzBzeM2Bs050Now5z4yaCdCd4n+CayGpKA+
VJZdFExb5lPp5aU4IUCPCxPUdCkskejWtXRfW1lF6LjxMaz6+WKMHuo7sjR3LPTA
V/DKrBhPg1gv9dIK6GnlhJqdJCXnrRIZwlfiNFNySX7Xz1T+1VIDwLp8yOq03kys
ow6u3wr4TI+AUXvAPntREEWNVzGO2Lfa6EMJFcEA4gbgDC3f+MjqXA5y666keH92
vd9uCmieEDtqhqfCUzzTfmeFa+nS2iV6opESR51HFrIGv2vp6dX1uawYtYISzW0E
hN3uQDxi9Zz4NyEGyCQtlFkAztzO/M/BLHji8gXdXtyt19nbAbFCC7B4xiLT46DN
0HMI1CLdVF1CDNPF0OWSVdXeZNjVWuWOXX7qKrDFUe1Qxt+xj/7niWYt43I3d6Xl
XW2/j+tNsqtZVxA+KTjlwaf1kjNoT/BDhtf9/d3CrRH98pOvK90v2T04VpyXUikH
ixnMXap9UCq8n24KBdgejIKtfKZJMJsDzztuOlX1Ip3/n7NBTn+GJPF0UzL9/c5I
c0RknjPiUJJjW5s0GwNgnsT31HfxEFGmX8URVFk37oM0BpNWcnDDfr8uv+BFfKr0
KU8smJBMAqZeaa5NtPubMgCrYRfhjusH+dyX62zBVwreiBN7H3vyTBPGZUba91gm
O2LtNspy1LeBGy25TbVQp/pmBNt0YGgf+wDmV27Rwr4+LBPJjdUg6bfSkSzyn2E5
8EE4aAud31pOgr0Kclba9Udp0aYB4sVBVIz0kozE2poOK7zAKj9WPpncD0D4LsSC
FJPfh20xnw6qhTvDAGl8OjskZDrieXt9NwxJhZowmtn331TBWrV0zkDk/MW/Ekg2
BnJ1o+EMdry6N2L3emi6cYdLd9/U2ROVnNuRSOQKjlQnjFjPTTiGo53/7zrBeJUQ
6sXXHI57kaMdKh+WWmmTlcxRwhBaTT6A4xBUZ08LmOSEYiTuRJaG+NSxaEOTf/IW
A+Y3xqzkk6zKwGo7CsefDs/B3doT8aacTZmrvDpGYX0v//4t5M9JlZ06aW1yMtQJ
Wq0o0du5F/TmUcmbXQgcdecx7suuQWABDAoGdOkPWtNgUqQp2SDyQV8OUxss7Elz
dDFPvlS36rWVh+LWXJuRjN31ivV0H7nYbWkx8+gHlyOhsN2raNB+dC02dhHB5zRP
POwB6zTuAwCLTQOM6mdo0uiV4V0wDgyBjounbGQkelMhR8GARa+8BDQNST10+blm
xtCso2jOt6KuKTbxtafWXIvbd3uptEQkMGN4o9WI/sK26r2ti7gE/ornlwyEUmcI
s5p8tWkGgI5OrjfwxPG3r23jzNbgFeaJceMmbQxPzkMdQp7uJKbp9KxDtxPW1weD
YwWKxno4fRNTNSXb49luGOwWz50czNICLWQoe1WUIJqnI+kIuZV6YFwA5Re19/SH
/vnxFJ3415CrhllWXBOARkVF4TV6OPo2pwAqeXeAr3/41R3yGq1hEj3sXFEh6ueV
vdLFYIlBylQ2GehO0I7Zc6/t9vuayMU2Im85dock9OXNM/U1j8zmNq8+t2bVZ9Pl
eUZtRZQ6K0exnY866rPVD6q4B+d406R/G6CFS0PfdyBLPgP/EnqICmRUn67xWKOI
jmjekJnLe7U4ue25XK8L7yLappiWsm7hLNBtKZhDUjuquar8M3fgS0gyrxrBAHHn
sp+BDzU2hPPH+3JQK2ZT6BmUGWvPrv1wPK8bcmS7rDkR5Toa7ZIjnPkei2xomQsX
Xvn24lEFEYVEcsZYiSnQeK5Jn8Ry1GU8N8YnBzJjAA2kCJdSFTrkje+2k5LIYGrH
18DfraWh8DkEh1i0aumaOr1eiYapKOHoYrFFTnoNMxQ5TM2U95xgIZ3CA+H62GF8
MhlrOKPZ5n8NKvruNWJXVl+exsi5LD4FxMa/nY0MzpXbnCGPVlzXJvzx6W9Df6S5
wRmbunJ9exuz+k774Fjm3wkU8lZGEmUwx09fTaok8wxojuaj8yduTrh/4Bhv5xJv
P97lTzCLqJw3uvNn+FZR6Igi5Gix6WCOGmKtqsH+Zxm+mUqqIfrrnqdXoMRUTB9V
qSl9HgW86eFwkmFzy5PyPyaueLrLSJlBeuwngiewESsOHND9qu3XW7NsOZautGMB
xSlF6T83Vaju9x9Us2mOjohRxIbfMCa+yKBIzxBySX080qURJ9oOzC7YkT1o8ZWt
zcWirilSZrIp6q949od2vv3LdTWNBMb4gTf5s+rIptQNkN5WSLf0Nbl+dfqORljm
CZg6DWOiWd77ZEQbIuj7usR9Y0GpEW+M+763N53lirxyxyAAwoO3xdQ7VfRNQQbF
/cWbcPufaN5vBSDRhq0AmZykzVWDPnXavz3O2bY0aIHsKJFkLj74lEtVQ4wMDLA6
48Yax6hHHZsjra/07zIPNXtA+rSaH3N3ZKLfvcv4Q5HzGATXpYrJgBevPQIGgwZ+
+4z3ZQQKpgfDmIUbvW4sIKLIaprTl+pFjeILB2kg78h+8qerQVNk/j51Ij1RG8uP
TJyR0fxx5NWBtrwmwF7eatPpGePQN4H6ik/9/nRNvO+fOyVsVZLkTXx5QY22RTlX
SS3mRm0oHPlsfNPxfEaQMYORZabUrQWjPHAWUz0++57Eq4S/TP0y7a0XIFeNDwx7
WMrDJVLuJINaT7ZSKQaW7xaAKhZwteklUUC1/n9yt+Z9UZcV96Iyfv4bLKc+wdZc
8bcm77bbScvhEKVeVzBzYrSEJnWzOD0vXEsIiv3aqkPIdOwZdOwiexdZUcrwKdOW
Pl/yAAHiaKVor8Mi/6M5LCjt0Z7EIIIMkjR6t0H3lc6vBM6rjtPyehIbIQEKVazo
SikAmmBX6qzLPpcNlmnmE2fQRJFZY2SHvDKjWv8GJ8c9P1fFyKhbMI3MsQK1X01k
ecDflQqalBD5QzgaIPtqyqifgv5j98ENWkTNTpjDqoDFMLvL/eBCq9wkubBqpu15
Ks5zyMul9n1iz5fbsqprnMMc0AeoF50eARs74//znFNNczpPOS24KwcoDEFtVpnd
GG0pDmx7p8kqoEXT6cPD6BEsK6dsLIHRGmin6eecYrgiI5eDam/AcsRiZWZtfn+8
Moe/v8KtcV0Et6QFjbb2fMPJS6MgoiEnSdlV6isLI4q9Zc0GQ3h3fe+ZlAGUULgL
tKfl4hGf4p/xajK5+6k761QzfteMdaW0HeWfbFcjX//UFSf3gCj7wd3Dp1u6PgV+
/EmGU3FE57xObcInyqOwwTAlndPYrc9o+wOcAbcyJQD3BwNSmKxt2CZdyYqD9LgU
N0diwGemZlCwqBUkOVHGKCiUvqB9zf103YmFD5bYMcmZd+CSeE3E03xmrUzOPQgU
th3D+rL6635tVp36gzEwB0hmaImbU8yH+6JsgUrGOybYqroNXLu2x4Qc15skydqu
xZgVbAy+33AFfuzAshRStm5vfA2KESALnxK+XfrGC4cAvkL+QzQmpaeee+FNBvlJ
J7vlVSzcZFA3AOTLUU8sZ2IqrJq0PR3vr/Z77HJR0t924A7+xsKj0V7A+UypJ9Aq
yFt347JoXO09ZjecpFMNhGpezm9UHv6uW8X1XO2o6rWQU/GRa0U61W0mSrlM1qin
mfmLTdnEKFRrZ6y9qP+ttDcxeQMiJw8iq+y9T/KO90It+ByHGAqMZI+dPlvii3eY
U1RdFcYKduGzghK+OZb6IUGYmrB6GWQZL2vKA2Vwnz4YJA6ArL6Eh7P6fie7D1tD
W2ROQuj7idUFUeuLnoqS+8jbhogTgKqxqst8c2H94vAj6L2PWjAk5DaDR6yLE4x4
9zPDW75n61rfPjMcpODBKGSvNv/8KmaF3D+2zLCOWgGZQjWAAMPfRr/sw5g9nHP/
3qMVWdgpTN4qih/LtxiVdQ2/SvRa6tsqYcKi5LzMNqGNTug44yYLv5VUL2zRXH0X
jzyfYundJgQlJ1rerbu55ObnJHF9xWsb4at2iKVJq/EGEXih36F+00/4sJOKtTKL
uquZWDXoysgRkRK2v0ECS/U8dLQIsWbJPeLhkE2BADB9hDnBaNtMvA5z5klhj/Qd
KTEyOehECJZ7cYFGwANWre09JG6tRb/d9Zza0utVvYTuuZz69Rg92yBy93LSVWyI
TFKIFGvebOA+TjkMrdegZr4B3Wm4egMY20803R30Lu72RIevKaiSXU9WxWMWNVS1
YTTNs/2XCcqZX+StqdZbIKTOvBda8kAZFQZZgLB4pp9jmU7J2tTmk7dFneSrFLS8
O7KRMKQg25+UbUm0dn+lawwzCGVW9M00q3pTJ7z7wABA5hDvtEWANlZpRWF8RdXA
5H+1Jr9ymIJLiselc+7a7mtI/uluxKyP7bcRSinXfsGNbXFey17rJltqefQV5xUR
zRP2g8/NPAxYo7csMsvxTRuzRS6kFfX1TOejxAYeWBwC+Noh+RCRj3ipPCgxotO8
SgDjKA1w92T/sn+sMfp+4KUektjp3+9R2npLQ7LPbe1fVDWmvtsT0ZfQK2/eeMYo
3ZmEISwDcHzU9DsXKFW+78Zh7QYKihxUR3Vb73g+MLbp8lHI6mXjC1slg158139M
cfbARRraeUIX7jAw3oIOUJ0MDip3Nc/sTn7BWyJGI/axNtF0Q/XCqNMxz1I5wgGR
SSGCKuRQFXcIxliqSJlBMwexr7/qNhtxw3HP0QS3UzruOofwnxYIIraOB3AZgnTu
aTuGjiQXz0hFKcQp8xLc9DFO4TZdXJYe2La8ES+uVtPcEY1oKK6+X/+gjzjilJbF
P+DYuFJNimagiifdg0aNYyKU5v37rJXcfCcOkhUdYnQuGJ5fKNNineAtxup9kOCR
bmgINAN8JaGCoWTgHPMzTtV+SEk298rnO6MwmAj/CgFPayUi89APphl+mHFYl8NZ
dvkSUEs1nI14uODeQ3PBLqMb+zSJxQVXZQCb0h5Jwbjths7FRBRaCBZ41/NoWAqn
Rk731bb5m/cbCTSlL7ieUaxdIiuzRYKW4oGRzmGUCft4xEowYMGc8vv7Msn4nKmr
XX4BZMbFKRWEDTNFZ5KvA9UVTTTMGNi7e1Je5imjOcsazQGQ3sQywyukwmw0daHT
GIIljQLrgoPsYMxBKfevVikS2/ak4pKaRydSrXbH4gITK+mPQZFMOHdb2w+fh9pt
1Tz5PH1ix+IymRfcA8u11PbMRre1sLJq/veBKSpMgGtJoXBa8EI+vMV9mRAZwu/F
I0eCzccFI9+BRxmEUeaFUNqpcy4+lfL+rh5iTLEdrDU2bWft2RkmM1ksQK90Se8I
2enJANxCWBiXyRivzdSYgV8TY481aLA5dhexEG4h37VaDFLXMUc5jnbwhQzf6SwE
LDu4xBjyZGpgwiWKa3ceSNYudszePI3BwUerF18d48xH4ZudPTCNezvkXxsVqgWx
pLBQL+ahgSsiDKg+h+I7c6junyovdYXGXJCT7wY8wp824y34MWtqJ3+NM3g++Etv
VOeTqIuBcgA6fxhPceYIkbm+7QP3FujOMTc57IDNFGU7ui1Y5DKi2Dzfh85DapRz
piM0+8bYUVFVChtlhBT1mKltgJM+z+NZEq66f9JOXXZeaj+aVXVxZu+AuHFGpbW6
G606fMsaMnyDhmuCNE3jdZ+XpmviO6XCZmrnzKw7H5gKtmxGpWSQOzJ+jho4LWCO
6MmeH+Lk/SXdahBs9IMUPAVh8/hPrmyzdysL5NS3UxvWy0paskVN320COFOqo5uH
x2HKFGNjqv5hJO+gHpUsPwN4luSatqn9WbEcdPWSyi9HneLTEZNkpzRcsd7Ei2LI
YmdzC0TTcLLyeAE8l5+eLRs32IYtOgqSlSqq6ukP15KnEZu3IdTn9D6q4gvnik9Q
HpD7jTeE4AB/akfogdIk09J5I0rLBrGuyvSuFD12aerAC6G39Lujz6ePasbntS/r
1OZbwXXxI1iZIcNXbqxZc1VEi/8IsuhsSoAxpOitnY5tBTcVAlVhZdWM6ARX153W
p7srQ+8+VDwvh+E8eQL6n5AysV33azExpONWiIoU0HmVwFHoNmXeFb2rPrBOC7oc
UKM99ykVhXWH2nDOxrH0Pju7vYjHBvtTqRN8D+PbhLn53Xw0Aawr8ecioNbNViIm
hK+6JIMNnCFgltzjFLuTYXnPZ5zsFxn7o20UnQv94myII50CQANPZ12n6mbNQB44
ybk82nG2sOYUkuUdwgs+bEMwORNzEeP26J1gs+Aehaoqn+aoPkq5ZhqbCvvN+XiM
qjSNJ/G31Sjqkue0SlQ6qgUXPk3nb4UNkF5vOMcqKzROzXIoin6sp7xQ6i65lM05
aL34KKND6UJJA8dVcgc6Tv9bebvx8xjY8H7zm6z/JyY1fURM7MW3pHePXOur34n5
vVLkuel7GcFMI6IV/ZPB/RZU+RmtxffQwFsz8VIr5IuxHDUrVvkriR854wuBVVHf
qK1LN906uLbbMobTx5rZNf+pt51dict3Nqh9+AGwXTZwPvVTM7r+iKSWSkjxHfJm
0XUK8K0DaMAg4eqUgNaazHtKqHxMN2Uio1T+2k+op6DJOpNOqiSCEmqzJQqJU5mz
Z9G0wNaViMwj0zSih0DtjP+6vMFQwzWWAxQ/kBFqvRTW7/V5hbmfFBiPIJBos7bi
DeKn2z7uRxA9HGGhI+5PCs8Ck7f+c60NgRMc+L6HNuKQvRYJKzhHyT/tQo1dSIrZ
Z9zWBpD1cBxFmqELjjXHvflXT9iJpAxyGcMP60353MQ09x9fto+mLoif/UCU9uS1
pH9iPwLikTaDEKCJ+yb/gk7mzrRJH66ZZVQqwe/p6CtQMgZgH/63yZgOWULu5IYu
XID/Z4t8j3348nAoxjr59aGdQy+nDawGoTM5iejfbnOFtOGCjv1fQyLdSDTWaHQB
lZhdNckJI+XF6V1kXFHpTR+WXL7DpQhfrGCyoYEiPqT9wJ54/CCey+lySaEeCq9Y
QhxAhwBw7tNOL0+ZsuKuLD47rBplHjxIQdrSisoCLPAFEROxab/3UzXvs6XU74Yw
cxS25ev0bCPTm/6FqHDl73NRwpSrWGFzUzFZ1jInaguxnLNNykbWBe4r8KKJcM2r
70Ghi9RbfVHMfmFmor+hJUiR6Bq3dNrplqiFKPErl+2ULhfO68Cn935V5BP4uSic
fct1T48NrMThYpEC0bE45pBmUIfu+XpIlA+jmzp1W4aGc8Cp3nXvC945uzF5uYny
65B8nvs1jzMlS3R/JTYRKHTILBTJx+ZCan1KyyJQoqsIocKbMCtQmf6zYcbLh7dY
flHHuvjkPtNSCo9jOEyIAynuKkCS4iHw/KQH7ljqiGPueHQq40MILTZlR0q4Ah4x
rZ5ovNylgz5RCBdP4JrLzHbCvhRmaz0ojCCmHXkWG7lS0+SHxNcl7Js2Lc31wgN5
n/EsgoTyx5wadUsHm2EpVlSQ1+BJngEs1FGFpGJ2zp2SGCVm1enPWguoLbZ2e5Jj
v1E9Tdw7YVqHPunIGP9J9Fp4v3lq5xuY/Wbnm9oeYrn91rVls0+IugWhtJqMXl34
+DW0UZJVonRWlGqof7giynao2Tl8tYtldlB2xdLlI+UYZOHMFeEXyPJ2cJ/v4lbZ
5DtR0Wf4oiStpjZrY9XEDAut0D9fnUWhjPc5x4D9u1jBHxG23L4LClJ94frStjlx
aui4RL4/fJvYQaaK4hfjTJsOe4Wva4YN3M8CxdiGWLblf54oz7clzBGxFqOL5b/D
Y+hJRiCUUdYlwGPkEdfoUcKz/tqfBl/eYjF1Xx6U7a301Of3O8+SuqyA7JGIS4Iv
mNOcOaIcjW28L7S11KTA+YdvJR77Sdg6xKPvjBda1GnqmqZqciO/oezJVYVfXOMK
qh9mwRcv4pDsmyiEOjaWKPQoqv8HxZpuKVmebahARhonG9+AzhuqwwoELex0dw4M
X1w20LlsO0+BZoBK/StUrnpE9NRXJzYlnFscYLP+Ekc8D/pl/40M3lpnJETPKJkL
6wgc2YL03O3uMtmfvKq4azTdH9dlvSSiH93SiubErI4jC5bhZ0TOFfluEYOMk7gv
PYA4tVVnO3HGgwebp5wOGKOTIE9/m388dNrVP66RjHQm0caIbuE03PXTP/57OIT7
KPzhS258Oo5nmpopOBYvTpRZuV2taRfKgrH205xWrRDnAdccv5yM3V7hsQWOEqy9
xJ+fyzP3ZRvzXa8e0Dg/qXMo/ztQB/t/JTMdTrJgxmbFmx0ktLkigcqnfoQdkKef
u/842C4aJkIkpQJbKar+p2qyL4yKpe0VBpQb7/Vk7oOMEtEPIYjYPTyf/vO4YN7d
VXHbSurJf+MggugY6Jr2JAu3wAXLDLmwEB6LAfgUiSXxEkiHxV2rbT23izHVRfqY
BpVygNpcHbYc/6EesuW0rNRmphge0Mv/8ohz9aMBjRgxx96gagmDWORK9vjf0DNX
UnWhtUMKqpueoaUobZ1D/me+9KsJ4EFHkV+uB5xTCCM1PsRMn6zIw4TKP3JVjAtR
VdcMoFSL4saLK8vh/oX9GHT75T8knNA9+FCVwzPPDb2D1iDwYVzbUcV8hydkVxIs
kJ7LDLWVUoi3w1TNSwtaqc3iAP7yG49UUQAPwKFxe/JHlqsV7zESaMx0kOGTbyjF
ud7TpDmRlGq+717Rys+4/mf/pMBicb5NEPsu5pf4SnFMkMDYDLAg2ZHlvqrS3hSw
//CuAFcHq+PanMrWhxC6IeamhFl/Hm6WYA4lp2wy4ocVORYrLU3D6OoDTQf2mKdt
785mWCDkG6KjQw9tkIwyFW/rBcADvF6gIb7wByzSX0zy0sFV3qRTjL7DOMTPGfEH
KlvV/33zU8bQcIsjJIIbtq3Fxw0+R90h3z5dROTzcITQhdNhLW13+QmYvh0b1rZ0
8oR04wQ6deEKkIkum3G6sd44rBM5hp3fcjCOq6ghU422/xUtatAOCc+N2nY4BD+Z
Nm72CgJC3JbagHafpB00qb9I8qzqIVZjRc2jmytTl1vnv0LgRqb+IB+u8moyT0aL
Ig1ws0OS+BxGJkpzXt0VpgAo5GvgL15Tk8JLRPygb6/8vRHyp06HmOuqtSK5LYHV
EkLltaxhTI0BmG5aPFEQN7qlJKEgnMEuO8ooDk/H7Yq+ma8t19gFz56XXFrKT/tt
qJ9HH7jxxwSS99aaBt7BTcZgw5TccuyOzKX6nnsV3cNDJMNLpj/B5ZBxGSJOopu9
QNoOo/WsW6VU4yBzoO7PWiSlrbHCX0XiYE7cMhaaA6euKMJcDMo4iyF2qUsTJfeu
hNjBLRzmSLw2HBAmVaknh0uTF8aMCpdrw/tE5d/3moqyRVw4yrcrvhInQRsi1TSj
90gCW8/rSu2fer/SlaPdvmkXdnaxJtE8vHGEhtEDIi8WU+UVM+mk2SCuXldOz7L7
p7DQfSsEiawaxdtbqNaM1ZWOEH8cw3mJxeLbCeLYH07NQJ0bMhSIIuID9eRPX0/0
z1F5/1XKNvV4i494B6B5uw+qnLDHqPwDxZkJZCJvqe+7TRdFPHxEcAhMtCy8fX20
evlfuwZMYGP4yXVXt9j8x/3Vlnt/ZPuHklXqJr6yEGGXd48fgupptHe+jfl6WkGD
lhY3SbOwh6GoTkTCn2b75ffBMSdTL2CFvJArrycMEobWIEuGldQEF/KdQhzJ3KwU
VcDh5+/uLz7VDluAZaezwrIxyNcWUHVdL3soixpfA8NUQiOodALg0Hm3rVjfsrbr
4x1j19d4m3hSrCImfTqq7hCjD5bGiTz+c2tGsyVQ+oSc8ss3KUIf45Vb1L5yROvn
E6Si3/9iQQV1rggK4BIdH9Ts6ZFfkd7o5nH52ehqpy8E3kFSfVCPumTCckyvKrh7
zbYyL+mzXki7/yJznR2xqG5Nks172ow3622YPeSb3oaz+C2eobhnWpfboZ9NKppf
CWG4/8gpra6xmCi4CKzxtYSqUBYh2qb4xp2WHmDGq0yrwi9OTwU7UoIyZALKPfjt
e2V9pXZvJ8ccWA4HmHYJ4mHD0PCK8a9c+N/jWHo4SkbjEq8EmtW02tVCSaoNZyxT
Bai+s2Bow4fOd79FcgMPjs6jHyh60Eq9c4MHgPVUoTNuseFY9iCRxwYXjyc6Ix72
UrEb9FBIl3uPdZAJTevVTERFL61R2RJmpF/kQEL01WOOQDCy+mHW9TbKpeM1Z41U
QRZy4m37TKlKHaBD543A+GUg3WMK2qKJ5SM8+xxf5M2faWHETh/tei8oLx4OQ1qV
oBCfYZ6eg26x0D+F80zr/O+8RXGel4pj9LKkquNYJJmIslxAjFdO9mpEatJB6szz
eOJeGRxA4BBDA3Q2nrZFyDziC3nvneQYYLnfzaZXPf90e7xDAdp/Vn8VaZ7rPjAz
Ex54dcJfWKHh+5Y44kM8fZLL97doztax/Z8BgKnJ8Wj9lDI5HkmZzFGrkRArIofo
1HkmpcA7CQvB03iHlNTTp5K6eoC5j9N5+r04lSeyF3U4htwLTK1OqzgFTrrwztLP
a3DPXfpW2zzPlG5Qjhi2bO+Wn5QxySOLK8lbUQv747vA/yHRzH/L0nm7XBLOn8RN
TchsZSnyfgibU4J8uISsUthb5oKL5usnqo23+6Nep8lCtJc3VMFvuHormxEw1Tjh
TiTQmJ6j8jgAxJyp+v529gi4KJzBByASQqC3NYv5BvodMWymK57rDfdmA9pnzG3v
yQ1lxMccoIBZk9rR87L5OPvPwAt4MvFyFm8tD12uujLD4w5AbdhijryTejRwFm9G
iWMO2ydw52RT3su5rX33cpsqX5uBhytWaa4Oite4Bufg2RnKdTcP8jY/Xwv5kUVM
RXIXVaR9+88pRpowx3BmBmbsfOg7k2dfVQBPTW5Ju40LkLcvWUyTshb8qoLlq8B1
DXUfE6v+LcyEHEQ6UBu8qAdOah9/xodX64WxG1hsZxDNR7A8yyN4SnZGANzeRPja
5tGNyqdCh4Edp6o5J/3JhHO+D5Cb3qVD4KPp6fFM1vs1X1Xl9kIbmfRD8FPlRfQx
dhMd/fvn9VNBk9ON2NvkfuEXqTCRRD/DnW0vkoumqirVPSQiO6QyurkPIjkWfLPq
Jm/YrnT1w1y8+dKUPFGNH54MNZMe2koWbgNKVIv1SJzal+/I9EJJyiMMzkIC4i/e
YWrr5P1iw5WozGNU9I/I37b7gJr2EjSh0o5FHbJYjRPfUSiwYpT38uNFPrcOHNOO
XDHeGW360k5d+YNi36qnEfVcVCxkMj9S2KNgSylsQnzcdskUWttHZA1kLtWUfGgo
4uGRFewgDTetuCi+K8N7nSUpwpw1x4FaBQSeTgelU0M4BrH0T/hzHO1nrV0F/DoD
fgs/gY0Mo4ZurE/sF+wWALQYUJQYZubJW+oQLeW6zlLNyKfYlyXnE9lFRwO/elmU
joRvuktKaF1n8KOMl6lz5mynYyzQRkC/ANuhg3dOfgf4d52JTRXotZcbWXs91yVk
ErYPnnmOLV4zn23vA4vFHkrWTBzOLYVN86FVlJIVD3pUKTATeNp3BgdrRgmh925P
n7dikNK2EVK8IIHg74OY5LfKyPykvC7VMXY58FuDYtr/FAcE7mtAjhnJtwubxN+l
rGvRCcZmZ+NNWa0fTBbLObl9qkkWvsViIHahOU2zRSUbPkGG/8q9NmWGbOBPoa2E
oRzWpsRkA1Cj5k0CRbMbQ5/Xyzxq+p7gqtJj4wG2zrhCbqsuGGQVmOMvKl3sySEA
yOTuCg9nbYld7GRrvDokDRG+xfJwbytMptDetuX39Uk9VRlWRPC2uzXO2OEzG8VW
cyHQxiR6s7nUywExe0tELiJKJYrBy4TXzij5lcLeRTlz2vH0iixR0BcdPQGNhSJc
A/MjCwZ9iVPKkQvtfRI2i4EKMs5EuB+6nbQkgERJUnnN7fAIH83Jqwp5815jWcRo
BLP7qbnggWeLS2/UUob5NcHc1SYohNGu7mwK94TwWGYfN47KLZIqrQDAydAc1RQC
PAUIqHeDetGd3Wdc2FygzuFQH2SfoEQrCgcIf1A5plDrg2AwOIQk2qy0EybAUjme
kVE/Y34U7UXr3AiPr6msxJB9hJGOs6HoD9vXZzXITUFGppySETOHRl7u+9XsuQxu
T3ax4AUXoJLES6bi/qVHM3tOluUp3IDIqgNAn4xuTe3hRDafhUGiJ/kgieYTmeMk
1MD3HLU0pROBvc4/oGwuGre6lyuGctgKAGMfWX4bthT9JEcXw//RMS08u6+9YLXO
gRtd1pLQiP7vJ8097iKbznt7OsrUF6WDP9F1n7vla5uOjQytkEt5qBSFrMYJPG4v
1DQ7sB2X5/5+iX+sVIDa+Umz++NLF64GcixkZ8FSfBRxzgrg9GdZuX6YP6HcSJFH
a33xkSso9iaJwx/EZHF94qhLb8RLod/EzDqfLdG7boWq/rOA/ajDC1U8yto0pVpE
YfhgKFQhvahwLD2UtkcnTOMMO/C9twhn7DmrEPDDGVsF4UVC/9Z4IZq034PLDddK
WJtalFHqFr+dDzgRGifXwpSVFem/8/Yo/FqkU0cRj4FCP27HUL0dwAr1dHQ58ckx
D/sGTYILRRimLLcLlImXS9kMioAWhPDZi783vxDUuYYpwS9PaaMHCBeRg1m/y1AW
/JZ/bVQaEpPqmGrv9ADxRx7cuT0ARjKvZ3bZRJBYLYDFhXAXnf03E02CrLoXurrp
sOz+5CTWIndM15w7ceAVO1SoytY6QARIdp6nrFnhTgIvap33oHkzPVbQ7Ch99+Nu
Xv/7fZg7tkAOATzVjypDAPkYMDCbFXBhPL6YTzgxbL07aH6Ec5YJq16yMIVd28Uk
XLMQkdg2auqSU/uDqANYTCst0TsSn8basF9hpcnrUTYWI0M6f6dkRKfdwXS/LEcQ
ovItoubeCQL57eUeBTdByp7IeyJrEuZGDfHGmrw0VapEBXTLg5sVDjt7Ebq7cmnk
xPuXFX+9wL8T+nSkIKVJcHfDNn/zLpkwGpUGj2l3z3qeiUPqbCSIfihd2UQQujFD
WvDx7FBQ+KTUBI7YwltBwX2/ZjC1EDhlTV3jCOye8tPTB7NLXdOEK30ePhUFzWcl
xGRglEwrDURMPTqxV5FOImblcSY4TR5nP4OWEouHJXch+d51MNthZqLXaT/wGdEj
IVmxCsMNMuNm13ixGr6nHMVJ+5dUB3GNYowTcyrd7CVzF7hGp8os32Ttu93C/xYo
+5367G6l8W2P98vjRx/47GHKWRDr/CxxeG9l94W8+pVsX5D3ySQIKmbX4v4Xy4m9
SYtM8LgnRDqM0ImTmqNiAzD7uFhXYwmrBZYEzVJfXo+63AmzoLkck0XE51irXmEB
+C6B/vHqkQR5bQE1dIwyLpoxhUwdtbNQ3gYnYljWcnlimeviCRskt7Bb+xKmh2LQ
kiTbcy/T5nYYK7ztIR6GyRqpEiL+ZWxJQo5ALlXCt8sQE2ztxYTbsyQqds/zHbJR
LBqxI9bc7mDKeeOCPIm2kMNpOy+ek7PfeUrYXwz9apt36X+eIuPtjbeIqiwNW+bt
WVbKk94GOvDESnWPmkmh4t223iMpwrQz2RlexdZPtPTwStB51VA/BqmO60KMVdy1
ld7NkcOQx0wov/olQmDI3++Esd1dh0CPn64r9xoRgI4f12KFE/arPx9UMt+fQI5o
vxVVcbYuHE19r26JraGwkDuz4QNXGErb73iryDWkPVG6/E9Ma4a5Vy2gOssLaGg9
xX+1HB2q/FTX3twFm3fyKXotkZFnRRbsaw7Y3ViLQ1jbWcGYsoudQz5npnF2EqjC
VGIm4R0WsgmP66Sg+q6KEczekGDAprnYxulzESQAlJEk7Xfq6TQr09vfDzC4HvR1
3hvRiwQOB6xc61Wo7Mr9RXp8ZDok/R9LjpD9rCCVfVjJOmzHof9UmtZaZv+8dWYs
nEV4YSPRGB6DMxW8ooSN4W59PlALZFD7rOG059fzZdRlB2J61CCL0YE0FC3qXDur
bNt0MB9H8zO/L1xwKxX3Sp4DB+ovhkrlvsvXTB7F4rI1VjmBWsdxKruCHUMlai75
lDnj7xBUqD8qD9EHEKOVj+PBvWWsKDbdSg73lURIlUqp9fA6i0Hz17o4aRVvEwZJ
2HRGHpTNSQO3YyoWiCqUhUOJ1un2O4DHLdQrD7ErL5GhfRsGsD7BabSAPR3t35VQ
fMUh8nhchBzoWlz+xk+00oPD4F5X0gC3B9h6g8yw7yshDoEWf+tvp4QBQWZcYlt4
qyxeA3dt+heVO9DMay2wSMfWc4SibltmZP/a7LFLjWPKnlUPQuerzj4IueZr0vWw
rrU+2sKg4g+tZVLewHWIF8hJFj08j4fbJIq9qy9MLvY7ZcT0pURzJSogBv1bpfnQ
qe7rnjk2RYA8zp7yIX/GGtMJvITezmSSqXXN8YHfl0fq0d/7qzAmp7/idgfHwcxU
ZGgQkr4D0SmgNLC5FVbzH8i+eoUiullufpn8WJNoZxbEBvy48uAUwnSMZ1mq8KhC
MFARD1aKtAvHF9FzIHuickU4oE/VuEtxygdHXUgPhRZjVdMZru0lDT+CQK2PKGyD
hHZjNVlxGjqG2goNTxm0w5RX0NreW1l91Pipu4RPbOA6XtFv7eoxX66QvNvHQUU1
CsbhVIVLXrnm4GVSHpXOVNMhal0bG7ml2l5nDNJTmsQalBwkW+vRjk96+Cv+bJIB
0sGJ99JYg9gi0oUzcOe3FaJ5OdQBQtTQrF30Hjw0kl3uANEIXc0kPmyJNssWqrIw
LcK9ti/scr7BmSMlWWdQOUQCvitSuxmpu9VTsDyscg6DEX7c1aWPZRGtGz/gJk7g
gGX5MMEidPQu1D6K9H4nt94RLpU4z4FPBl91C7fI2j2QKQxrEMW7uOaIB9YFEAHm
ecpQP+63TlJlpJUJbfAuflbFbEDtcYjIL+FvVs0k46vaSQ6E2Ny79Mj+eKRC07/5
DgCq4gg/yLxOoaMrIdrRp4iJ1MZkGRxqe8qRlfmXSb2j7EtOZvhOuJHEG3RFJh+c
VYgdxEE3aPO5jFR/t1kyfMN0IUiOO8Ou0UkTp/WcqthlcT9OtpcDhuk32slKqk+x
3Kdn2J2Z4um+wSqPwMdxVkDSPgI+ufZslx6ScG03g0iZo9yIhFsqkMg8ob0XDOx4
azJWmNS+xdk3KZhFTyKAA7xfewsr5MTLeKJeoquYm8TLkksdOaMlCLkEzixxrlhq
27EdWtm+TNwfyJRETAh16xsiMZ8TGulElY7695XfRqZAmeLGdywLbN3ZMg2kVqvd
hfReAg6X6LAhZHsd9oAxiG6CBMIXx3yfZlo9V0gIXJIDT8ltok6d6NWrhXAoGfIE
pTU38QcmSNkg4VTmLoKboqlN+I0mxjQ2Fm8DKrmyxmrn+yOTLd9i6zRqrFiAU0dn
vXDoHQgd5MomZ7bcthNA7KoOhECg8P2wRIUH2kgijFdfeP9zuuAQLfBBqPIXcbny
dPh+JGCLsjwGwBoPLbYVeWgMQ+aBTSCGBta7LhRZMqwCZ8LkYD8hE8qbzgHMr6vd
m5onoqkbQwWX91SefoPYI2J+lb/7PCx6DEqUHZ1XloBfD6aI3ZzRUMYJaHV03Fw4
Vj8tXmpU6U6FOy+Li7Rtg0S9oyuSzHaQ/b3SL9Tsn4i8DV424Ijiep4UOZsQizRX
Z4M7kz1iW+LwzDVK2yIUvcjR9gatVxfJ7zSdVsBJoU8afs6ULlRUwH59X88WRLkM
aMl3+DXM9k9P5N1nDsf5hNEA48gMYovYz7NFY+RidjrawjgD1J5/teJezddYTNd9
nHou0KYgs/NAkSuXT2NeCUfdi7eU7NMmivH4enR+g2fu7oZG37V8wTZ6EEFWpXgv
55SS+2nkl1Gg4y1PTlt579MxZE2/+437vwJhT8ecO6oN/onc2LisofHUizWCAEny
U3j/3EiYHlvibh07uuQ35Dia2VaZ+Jm/OE0qDwHZl4hO+c7Y+I62t1N7b9ND9iEF
wh1IjR16kV3I7WfdwhPs22dfLXSRX3uUSb5+VDmPmUmQeGan6j7jUU49v5w/zfZS
oTaDWAUJ+dr8boGRfJP7bTLVek0yG5DRTGwD1V7MfdqdSSLrR3odwf7fLtsHD/N7
NsB2xC0EtqVxaaDxvnofE+Xvla7hMAXry7itMm3Ip1LdcRlJ81VMGB5OMPBP8eV7
YMKPCWohmnhrV1794dbqXnCOEm+YfzPovk92qO0tIEJP3uTALFJSHYiK7ykQFacq
DTU6sK92WphEmdy5kVwC/bhFKcLwDeEMiNya8RfGxYcVF0jUXIyM3X6fI1r40ZMG
N/mJ1DcBdRvA7mfSKe8gYae4ZZd3L0lRo82ngcPKQas6M/0KD8feqwiwsNZdEbiZ
VMuhzv8xCLjPkkgFcLOC4mip0HJw6eJKhg3uTNcfXIChhLEWLF4Rgw8UUfddhvtu
SHpuBCryU+wZtIMynsjxD8Auh+7ZWK+ZD417DgfLwnDUc4kvZjr0HzBtzs+4dnfo
zC8HDgjmA4Or175ICADvwr+5DhRwO6wwTzWfpBjGZQ8rn40TTnDJ/5fLVdtWVSGy
sdpzXkW7Et6EbsjMyH07RFJECInMAjS7ybuZwcA6DLKJ74SulFVyNz6Zm/MaXDn/
tbLItqvKaxaG/hPrjGtzhS/60rELm/6V3XnmrfYDmgnT7j2/EELzsY3MydFXXjgh
xr7QqzE4YURcN1d7+pHSPSIMJ2joW8g4z1MAS4k661Bu8eq0xy8+LWxcWjoDOxcF
XD0eHoG5EkeYcETP9l8E3se4Uuw6KvbC1XLlKmWGb7T2dVkRecuQvjmrP/EusEfe
BNa1Skl6KoWOq78Bi7OGenLZR6Sv48g+FEYNOEFN0elkDRk6U+bbp1X/A6+uAR8R
CnJr12VnyfZKB9JMiBw1OFpnQzidK0clzY9YVpBFdD7Im6EGugEw8s3eKLM0xaWw
jEvg3cFCLdeLi+PLnBOf2ABnEfd08gYyDNHFUSMlLHJBnr/wDfjop9J95giNhOlo
+WqEqJ96YGLkO9Kd3nQ+Rddlo0vd/9dIUh4SRb+9CFueerXVGSiEApG9nzQ+6QUZ
Kc6W+Zpm3DMqEYSb8mP/OS7LOaRw7fHd/Z1HmdhI7+y0gg8UNMt+s5FJRFGXI8Ja
5scAY5/7r8jmjaenlzo0eIO7bS8bPjuLfq3REKqzF1sOdp/osVO2j965cRHF4k3E
G7jN4NLZNUsQmGp4ydk1ep0smN4nNu4fpI3t2Cogv7JtaaM0K5xKmsZ4xYU5oETN
n9ziPr9RlSIRdAOVnQa82t9vDz4XsUS335TZvlkIJ1jVsBxmDFzB8GWj5yK+Yus0
sx6UjBWNmKRM2xTJvUlRHE+WyA/Zc8uUwsbxaaCc5YGlXDlsz9zf9f+t2OTtpNn4
mv11qaWJRrUMgH/5g9mVwqm7JluZI+5gPSnLSrlVtYWXkXLV3qJXDfsx0wUlDQks
KYRauNbM10GeHtPZC7eSLFuJ9sd2wMtDWC2zf4CYZSEKXF93jcmLWu0P1N8mJSej
6xhLrzinjUsuXiQQkGDIHK36fnTjoHnNTFAk00Cfu/MAmOfMQrW129Myc/gGTxWl
zxJfiB3RInoagMNoYxjXMTWRo8TVvuqu426sODaEiM5iTIDfmHnC8//KPYti6CA3
XdkgRGtzFttUDiZNOt4w5QqDhHh0USrPR3vjv1b3HnwalO3M6m6gG3hA4qe2uVW/
+nyrUxDc7G7q9/0/pYhpwsyY0e1M1E5BNZALlXM+8PPOG/MVuXNe8ZeCpSaa0qcy
hyrvLGGGZAZzLYeLt9ItSydnvQT/D60O34bhktUR1dPI6+BgK26P9+mzGzZsivoH
lKvwnznsDRvr7Gqia9kxZQG6p59zgNQLSEgVk/9J/t5A2F0eLlUKAlbNkj8gvjLJ
uP0bUJKr+WIi52CGRheAygZhpV6yz4loeuXFHvYKWuijskLOtVqk/Xjg2KhR1PgY
AFsknsNUQnAGOUvYnDx38ig/fg8vGXXTjf2V04NIpDeIaC+qTGyIp4i1yHr1MP3S
dY8V/oXQKcVa4Hc7sLFw1Wh5AimGXYcVHp5/HxXeVaBBw8jh9fL+GistRabkjZ7E
imp9WOkHiPrPoLohczgQUQyExRwN7c0lvjdJoCRgKVJV8Bjy64je09TywtVeQaLB
f/iJPSZ1H5FvXwE5Xeum12Urc16Hj1J/nIwrxsdbv2KgljU4xj1lExZbmzOrID3N
NlAYci/WnnlGbptcQjmWgzQgRWldPzFYWv9Frl1W5BYGuQN1R6qAva3Hgu7jTMIn
4RpUfBM22mCxWsKoH+krUcM0yqQWqasGNjOpSHlVuB7fF3FQel7fqm6lrJCbsqrO
GYRI2V3LfkjuHcI/Reivnth2HsMA+EMFR+r4rrcbzbMJg7y1suRpGiJiNI1+WUzB
rMXVxWn6Ui9joF1B31gnRjU2iijyQJU0rErP9bbh/njd+p4eVw6YvTQh5wB+AScY
XpWcvEAWv4Yfy50w32ERShzCGnUrhkid8c4TzBjIrdNaEQyCsHfbfhYRD5CrfjRG
p9aLNygnLM2kP07fdEbLXduNLm8pqEAenqmDGXp/JNFQ1GgijqggYLX/Ptdto53l
b2bZ9q4o5TNaaavbg19NOUpX/6GVJDhea6vF67AaeDNUGK7wheRdAI+aGSG0dy8U
hAyrm30E5k8FGZmnUPj255EKzEwU68Od5ID61qCCry3+GkD1X3w716OC0D2dIiPV
RtUHyeRm/Vq9OxIrptQpn6/3LTT1lm2rKI6f2dprZXzIBmjW/RnuA7XhkgUReSQB
eI1uBGVp19pkQCZA4/agRpirSbgPpRoPudFfrw2PkDygIRj36bIBGaBRvUwkiaPR
nljrOYa9Hzy/khHvnC/IUFCp/OXq9TOH8Z/FxAYgd6BIfpfcO1UnJTEBR3USlSTE
e+OgKYsHcYXWtcVTFr3vONQt+a1YM1SHXk7GZyoZw6tzFvMiWDsWkxdHVwSLA+Ll
Iu7fHn5n5hhAAq80NKI9a5sQxqvQa14NvyILwZ//x9q7EOUwwJu6zlSE+CKKfs3s
VMjntXAp4+oE+whX8uTLvu+X0W7mqsDrXXKnozAQd6j38qlXvKs6yIg6eUhd+85J
G2foabJg43LNduxV+hwxzAjzYxoO8ebxLoqAMl0pQMKDDlHiagOmRaM0PrTjp05Z
vd1jTn/zeLOPQwR5QDXVOM1NAonVzeKlpgKf9KhVrUlLAIzOd6SIWcg2SvtKMnt+
/iFC76iCJVaqpKrA3ofoGuzK9I1uRtU0IOFyimTcK4r3PfGe0v5rFePG0ydkqP69
33HcVfZt8WIrQ5kgbQRnj9SpcwRBWWiwjhBilVUE5fTYjbjgvHWd/NjWGk+hlMrT
c/nb3HrHXMAbGgXm02Gv3VYeXcb3N4rQ+B8L70O+LQxnhrjhcxFE9qcJxddgRQoC
iBaLtFyMbQRbBNGvStZjTPzIomRjCOoXPbH+ICUpOCqPV8QcMZvzpwWmPMHJ932L
ojUlmMygTZRSl7SzCFHweLTsgd9aYzN8A/g86BgPef1cTJy6dwJE5ni3C+QSxx2J
fJSMbqAtHJ+zyHwVcuiPHToKGwVDp8+D5qd/oqVHjaIrkjwsxZ0E/nR/7Ue/rYt0
TG0YjGCMY0jQtN+Tk40P4E6LKY7qJ8Rf8XSdoq9XcDdqwM580a4tlaT6TyXcaSCK
7kdrRvMP0PteSfu0fi6uaN7gwB0SWTS3x0TlCaCBe+DFHlpJXhUROrLlK8QutCWD
KdlMQbZe0vde1Syj9fnOK3XD0izuNqsNEq4APdgwruPYuFmZSGpuVYsPMaD/d4LL
tdPWg8wV9l5Rqt9ltrh98IF9suLTDHlcHsszdz+Y5p9OeEm1Dbn9kpJGo9oN2kNL
D5hdmQQUXvbPJRKPpfScPJIHvdCaZOqdNVkszaHT3ihpw8E0B0uzcgj5z1NxG/Yb
SQkiBHE6bADluJLUFlV2KyiFyXtFp7dbmBeect9/KvmNCIcSx1FwUpNZ7XG+iBox
jmEZiu49Oduu89kDLG4CT+frOXne5fIm0MpD9mWFLNtb+dWsf223u9DHODBTWRJF
EKabp0+ZZvmqHDfs34HgLURdwiAFT7ZbnsKB66+mydelUDeexWbglulbIwCwmPR6
WXCNAynPhhRLktdyl2LU5PO1X/fVlNQhkpUd48tU6Y2PXEilOekBmwaGYLl19Z/F
33GSzMlSTZJw33Ep/RIm7kZkyV0QQTviU1KkCNr/LPRBLMlzWYaWDfwwRnPZaM6+
mz3VaRppzXMHHqloI4EJ4xHKq0d5/tANExjJj9kq+GT9EhEZqw7Swh2Ixo3gpNRL
sbC0vngmiR/oirUjQvkox+EgeimAr5ggHoiUYFsnos264T7lA9C8WoDiRYD2KsKs
fJujVq/akXMQmVO3mvP7gonZ0Rret+oXsnkutuWx80GePg/DJeSfeyo4exrIP3s0
pL4FF6Ct67nc7k93V2ifBAjmEq8Xv53t87KtlBJ5U3W8e5wHngwm2c3CmW6ewDgs
TYyO7IijOFPPLTuGyyHkmW+vrWsOPnvm86tjwPxnzFzWs73skcSuBKh9ffFbiP9g
3J7bdZtKdK7P3CmkSTfh1ewdhmfbjz7jUG0+CboxPtqTL+uBA28/9iIhCKQNdqlO
oXwP9IbAi921Se/Fs074B2tpRNlgdxm+riCcQI+5FPsp9P9xYXRb99gI4ghVVmqs
mK0KYBA9YkMPptxRKF38HNWA2//Y3IZ5jqjqUkZvWXJ0wy8gQh+O1nHcCWfs8a6T
V63eic/AYZb0XpzJY9RCrufmxQWikkc7yBCQA+6gIkGgg9ue0NknfAumBwvglGfF
xzwKyd9QP51icjHApOWVi5e9lpdvajyTeh8LAGpXl6Dl4X1QIxsuO/0k7yScqQM3
uLEpXYRC4MaFmBnm6OBQegOc27aO/DAFeRmvqyH51CVD3lTH7UpaHH6DnriV0AmB
mDJI8xLFT6c8ltbSKOtO1bBCgpeMztepeJp+sI+QAPDpWwYYzoiU7AIUYqQ51s3H
erOGtf2Yw6iok6d9u8MEstMS6uRFZFCs162vqYETfmzJLsI3/4nyLsCNxt9xBvQY
gnOYm/nnUL8mJy7U7r2abzKPGb8S+axCTWWug0/jPNLqL3AwHrSWM6rXQIHiFTDp
10H5Ni8ZO1xDpR2VpqqMFctR3tortXw5ranEo1KjMG+VIYj9xb04ykd1ukAIA0d3
vl3cbFxz4uBDmMt45Qp7roohB/vVjKzQ7I8Ihq8K4AEleewnqtIFhRV5dd4e+/80
s1F6pc4VI/4EKsfZKmAUzKT/bhuTizTrMem6Q8AHo+tOAXHUBrScenSv4ZkztLPm
OQ6LeU9oIwEWoNlA/HNvM/qg7ncRBoxbkLut1bWU0vlyHMdDF+3PzF6kzXBMm5o9
m0gGNpxxWT2skGHxmoaPuqkGDZV7YPAbzKXC2rXdPbqWU37ohBCoDLOX9B2fSIX1
KNXCY7zJ/l1JnGLLQM4nnvJFstz+XxTModKTRKB952h6fpxlXOiJudaCdBp+jEqI
s102KfLmrXaRtip2fwp8McZF5YKZajB8wfamfJPG8iBNHWQxSbXL3QQ7D3DmyvEp
N1RxeWJT9ZdlFluDRyAVCs2FNCaz9xCwvSURw0/kb7w=

`pragma protect end_protected
