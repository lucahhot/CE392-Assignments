// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
xZZz1xaHQxkm0cVQFWE5sQNU2F4qWuUNu7H/bhqLEECTYv1MAarc9VpsiFs/w5xmcXc7LCyjmWaQ
U292hKRh8YYmG0AAp7xd8pm52nVaenBpjEiDtusCIT8TM2VqwwMxk1q717tXY/49AqTrb6v+pKlx
ihJj3B1ZHsZdGRmjFOHn8fiUlNepSGJRyGMjEp4o8//wdPkjt1wfoQXC+tkriYtu64Lsfikcslef
eO30pwUlz3ulb7od7SSIAnU25fv7BS6LX3y9YfTCu+yNUi4/Yrb32dgXXyO5PK5ZQjljfi3TGeki
/1HX1Pq1649mJdqMaZYQEi7k/12FWS9xOLIzWw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2048)
n52DNd9oajVrsymcvfcuTOgN4K0q7ctcl4kO9fRpqAfQVcS3MV7MLf3FmI9P8zIT31H92UBUJ9sD
QkD+9zgre/tq5YMLFB0TBRtbA1g3mWwXrJ2/dIPR1Mf+bQzGYjjMco6Q8wDRa1WTEBHkwwz4DgTi
UoRpah1EnicUM38nvNMPLsTeW32jzdJzqkUxecWvLWxNzRae7teag3zJg35GwEuPSNSMqCT/iKQw
3ofFBQIhDhrWBAlFnhYcx5W55ruEavkBW8E0+PjzYIARXN+3wEhWzzuntHirtHSFGVbv43m9uy5K
+Kr5InKNUgH2FLc6TL5TVJZBwhRWBPB2G2HSSm1vF039jqXfPLIAKcX27xg/TnV3LyDc4IXC7DkU
EbO4f5tQoA3woC7Pa16NBGvCwZXeF93LA2TdNp26Eon7R0Bg1e3ENuI3EM3IsNFaCCeX+kzfEmcN
//nEwMB406oODKNpoxbt5hdjblyZX4DVzPdQd0BD7EfVUnXvI+/BOVYHS8h9SI86Gcj1uhdaJr10
1n4UvQU8mH3jFfGKO5Pkz5MN9R1PYmGFvH6EKHkAUjfG3Za/Ev3EUD17S84H8xfRY8fp57g+CSnh
3aEkHWBCPdeGHizHn8E1nUa8+DhQ6VgjA0Q1ChrpfxYflUxMNsmiOnI4jtepI5i0cXu8lYIDIWbi
nh8qvhupbV2pDKvcvKn9MO5bQ4e+D6gMflSMiQbRrF3QsdCVvg+NZAV9Rj+ql5DBeoYQECCXenW6
rSpvoEHbYXYcGZx0wX285W9fJ4TCVbghBdjbwfVZHl8aR7DGTi+M6NuN0XPjTCzttTMnuYczhunw
KGxJevfoRzjpP1fZ7bKDHdMy6iXyCnJKk0UTCpcVavwfUDN09xjngZnWY7nbaHxxmx3/+tWKl3lX
CV3hIofJIldFY4CpX6g5NkFK4h4mSXLCy7F2HGyNiDC7VqBgt6uk7jURI2F1UWSs6b4EEJYry1Pe
Hu2StQTooISgg9GCMG1VYIdRVZ4H5YcMKPp8zMo6itW0HaqcGgGsbR7U+X1ForT6FtJkicuEy7c/
jkYmJg5ZOLZGOwvG2bmHFJvGQYme+IK3aMj1tFu71YPU6WbK37HSsEPI44COPM5rLNh8eNl/z5Ls
vSB9ivpgJVVBnX164XZqaofIJhxZrzHSzH/iXXtKPVuSCZzPIwI8Rr1roIWt7N/it3vpeWasOXE3
2bmHPmlYaulO3xbypGiC2ds2xMXg29qo7GJj27CeI8Lh+nr2HZGfNpDL038qY3bG2avPDzu5RoUD
x8PlDzGoz4QGrostS4kvrS7VKK0bGzjVDKjxQSaQIDkFEP+3IdKiyUvgtTqcSbDNJhGlrxIWl64d
ENjYe67kXyd1Mg6pZQtIwGZb6nkKpo3KCj23rJO5rgTkdshxj62uO2XmZxS98Hzo/VwYX40s56SY
2HZmWn2VcmldB249mlkKW+egRrm/mPThKLP2N5GeDmqQDFBUce98zraLWJ+hQn6jXE9vvNj6LMF8
tIhUkt3y7RVT1dUFALMS/JFwAVuyd2kGcHVmMjD88rWGqlPTpWC5i5tjmLIdYDkzRJoNHvVseu0W
Z8yYgJURyZYhoE3M2pVXzMr9UxgQNDl0XwSdhFXcLZJjZ1SWVxA6bnTrwzdID97K1E0Wh+MTgQbY
zM/KtroB6VWzVPADs2+/8crMOnSGeK6Eg/oobV5ZCtr+f+OMZYMODid7ypOh2+zub4XiHm/pshWF
CCsiqyqT9I2n9YfISq02xkVJVFSo+fl5+otUmHxcaSptFJ5KqzBeWv9GI1m5BaC9BTa518K65WFO
JSUAG3QKtWMbmGJQQ44hzI+mRbR9Ic/f8AE6w+CLQmckXFjcn+dWwyxFeTdvhQ6B8gJUWdZFwtH6
AfXmI1zEuSVq8Td3gGoC9iXQspxcLyhs5MGwnVaiR8jiLClCVz0KBi6ntX1udK5TgxM/Dbd6FhCR
b0bDz0wZVR+ndz6RpyjjY8tG9mvyFGuBBx4oSJUMjWKdIvlib6S+UIzky7Xz1YEVbcElOci0gjOA
20+xmAuDe9meywRio12pT2RFmQvs4f2mZJTbp+2tgnPCMP1haep07JhGDwWFUvlX7CxltT5YQOSP
8TyZYdZ8lD7C8jqN4+fosOqzjqQ3TDq3wQfzRND/boGAeTUDQxCVxT6xsKpe63ERzyqzl6h4Z3J0
pMqG42b0P/ICUq/ZPy2raS+Zo17HXVv0ehLVvGFEDVBaE5yYJZ+7nw3PYmX4ppO1I4euPxHfhAat
X3Bv4LXx2bpYHBdP7VafQZDQJvX0Kov6OF4gE+AV8Qn0cnkmE92DWyJO8xD+LhJiTXZhzFOBJ4Bp
8RnEjHBQikDFXJVR8cjlIs8NzqbqTsU1Jc/HDBOx/D4bzy8zfFFsx65tEcfFql73MS0kvESe5GAx
dvHCzPsFPf1JafUtCVaNiVpwqI9WsLimcEt4MKrmJ4TBQrfSFK/bPtsl2QVJTlR5/v7E4PLFcTQp
M3NryEC3GteNKfH7F+vc5m5YSSAmYfY3QS6sh2l6XrTGZSV4HBuMmjY/o5OjjTNbyx4nPMPx2oRd
bxXLAYRM7xYUogv8xE9AC3w+we0wnDrl03ttxbqBPvbsNJ7uLxumvc1EvLgQPZpx66ruHhT8SvTb
g2BzBsdwEoFJLh9Tnq56O+CL8jUe8aPD9FBHd2I4UVELhIhE/E0LbFryrlN7rNdyGHmgfvc=
`pragma protect end_protected
