// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+eBYSsKOJt+o0lBHPkSTVrqrw9sUU7VKzzeN1CV2gn4LoxGOC+12LjofOrK9TVt4
0JZoq3L4wh0FbZeRCKwB5oSdJ0+P1qoOgq+Sdat55vdzDeaMGXX/rIwQus1Xjs+e
s6GZ84Nhasj/gacRTWSNCx2PmQlwDFpJqvnlzlOV7781SeJZUrimPQ==
//pragma protect end_key_block
//pragma protect digest_block
BUAHZYZvYMxdHMhTv5jtUJ3Dess=
//pragma protect end_digest_block
//pragma protect data_block
Td7SuXjVo/hQUmYeg9hiR6VJssMoG+0mYKeaaxzVSymCDGQtGWgN894TH1qYDF4h
A0eSPEDPMeF21xZNTvxDRithkq/CmV5L4JMHAYWrBLcm7GObSE2d/lBnApSPNNop
zUeBJNs/upThvel5u7+dipyjPyodO7yvwV5mcRYVYcKDU7QGfgVAKVFTHD+/h5i3
eB5dx9Z1dhqrIcmzed4MptSzguK09LKwDnHmdeJR+HHzNYqlQWKwU31zyPBiAVJ4
wyI/UeslJnlIAVig4gX2c1Bd1WjrkG3tyw7YF+bF/Ni0IPw2OI46IkgZVzgE+pAm
NrUK5RdQmU5lf/Rq1KiNlfZKaNGLTv0Or2dcwP31beGYIiHyD67KGtDlm5KPeXCi
cRX3nsgCmlhedq2J/1TaLzGOvN8UMEWKmMv0NO3EwAkZFtR3DuJ5uWRwQ7UkUVyG
zoSohfx6fI5Bjb94AQfcvjDO7kVTqVViNGEhvYWrLrPyFbcZcQ500u3to/khWS69
pTQYD6jVTeqA82Xotj6/8CJxa4LWqIA2rehIEfzNh6Yl6V3P+v3UiZQLqLiIc1qs
Xu3/PMnt70UGch5izOAx4tRObiTfgy1ucaQ6uJxGIvTRUD4slCaiOWkH+5MZaWWL
foCbQDpRLiWFhzLLgRIH2NJn1yHSDkZUUTLEMRqLavTSYshT0I83FlYXXZ6U7Ixm
FqK6HMMD12ByN5zMXWRFX09uWt9r7XaJnR+P8o1tDThAS2yHBObe21VFZtJ6LaYr
vwJ68OkurodRtfVFPaI2llfI72HZiNksO6i28wqm5Yn4VJXhKKWYLas7NZ7jkTat
a+PVz69o4+LSMCzVp8xS7L0GZHWh5Z/jZYzUsfhoCiJnZDGIWnzPgk9qM79+c3rQ
x0LDXDH/Uu7Jt1VB/eyKL9R1zoSBIes7Tu0ME3urlwa20Gv1uHGmiFHyCENfJbvo
FRyuVscrVeA0DM255/9LvRqOB6FF4r4Vj/HaeOFqJ5DoWoT/Yg2lybIBgPTNJTQH
OxeTUlx0xM+e+DNFlEguo402jKdsAK9JPZXvjmxA7oDeIVmfgjwpn2nYyCwxcMpH
zX6seNaGCQjejEv686dHBsILrjZsuY4YoTpoNPNe6Kzwvexsz3lsrZKkoiVXOw9w
FVkvvba5u30emuCYYgSYqChP45OxwqlnijWxuL5sAMerwUCCV71phTXC22cGqhlb
Xx6OW6oLDJg4oKGE91Ojw58WCMcYdGgXIV7HOxyIwlqBI6yCVBRH3bTD9SA0HY3k
r7FLASD0ASqujPijgoymuBmBql4XvKSjhW6EMqcBBsw4qV/GQSEGNh43jiNOoho/
8pKhxO/uY1jXBp/s1TdKigGn5YiVMP4eC5wEQa48e1q9MYM13uY3DCj+sMIiKc7U
n1FeE+Dw/hMEUXmzW6NSAeKEEIr/XdGgE4DG7oQo0L5WxQG7adIIzuKwpcPihnJz
mmHA2LrxBbSjxUcW5jIIq6okqRSqTstTuQxqA++eV+gjStiI1deybfY52JyfdOj9
ezHj19B6eZWndVpObHjS9DNUk0iHP/ZpHUenU7mgY5en0TJmHJYassXTlk+Tk9N/
jAd2gW+FGGqDvcLSHUFK5MCLYFLDAtRNxQ3de1D6nCa6ncMYE0L5mENOTAYkC6Bu
oG37/xV02vemY1bfNkqKpFmqiG53EykIHHi3M6W/pkjRkEMcV/k3pjnTy5w8DgIH
7ewdEB8+ja3vkHNxrUdRvKEnlqxs9JhILC2/LH+4QffnNX81+XEUUabesx3IugcC
ho4JVcqbCBAqq5dsT9j8tECDA/uE0j5QiBreSCDVleCV/IcFU83jqpae9ZCC4LAW
eQjaOkwoR8zxlc+1aLTuXkh7AY4Gu8hIk6El+fgznY6eViLM9AOkR/y81xcEAk4a
Sr+aRMN/ta1aVYARZ8HGRhjNInpLb5Sza8NFdTK7r683aS/6zDd2v6KBMcEAmG/V
3dmI1rt0QcEbmgGdSSWs2q5UAiriOP5swfFDw8VXUvNjrKDYHZMktkBE/i1y0c4z
74h6dnXhOeqcLa6gVKXbX/+eVn7k/CJZxtw6xI0WqJ/k7UkdsSLvX4fD6S1fCH9T
MAcmR+rz5gtWoYD9x02a2B/WU6L9P6Qn7XifIgfUkZfFGFuO6q7UgGYNP+YhLKE5
vvFsHkUil4nncVbAVMb2s8vNj/+uKcXkXULmOrwkiSm+FnmHSsXbePE/+W3bJ2+p
w/zwxL/TwKA7uGgoFdCx8WdUVm4u6bYLzHaew+JEIPPxPtmPqGNhhT0kLz6sOUvu
DOFQzCNQl3TWhDLurCN/jkB5TXaCU9OxQGiBn6TosDDegtp56MgNSJKkZewVxho0
U2qwhVmd573FnVqbIuEhL+EX+Aw+laW40DgBLlePul18KI0O0IiahL1FygnE6HsZ
/xxgQViPVtVbBVVg8UqN6wcZL5XZhPNS/DkD6l2894GqBDPSIWk741XlCG1+RT0R
X4PleEj4wdAVqHY6pCkgUtKoikovP2pYHXgBkyWqTDVh9HmZl06QG9m/9ZNIOzQH
Uow2tJGKJKBWhqrVeiJlZBmSiKJns7fqhbHuTdksCqQ4Qu8Y2BtEeMP5KIMEN+gS
LzIhz8GCFJwNnPucQ09thTkeU5Ss4qzj9DVBxeBvxMRxzIUADBsV0bu0gPcYaEh5
jz8tTIMP3J8dly/6mQ63TlGXk8I6TqBrYkktODmaSctRsCkYPmqcFhz9fPboydIw
a6eCRjRG0GCMwbHJPfWoQ6LAy6ObWbRcC/Jd492nC6gjmvQ4UvzK3iAtr+52sD3i
9A7EvGc2OP8TbksuvtXC8SaYzicZgrYJ6M0gMQZhoiWDfm6k0kX6iCaoKYzJa/ta
fqTxxHKtmxWvJ6DH6+gtEWEHF0knyDKCDLhQB08dfwQNOT5gqllg7aHkAPZ2XiTA
KdJz/LDbXPgFuKQ0apnf8E+F4ugu384BrSFeCTtF4SQ8Nob6ZscELkGRgGQzBcET
PGzA+preb4s/oqhzBEANUVepboyYeZec2m/Pr/4Q1+TuVRu+GosMS0RMq4bE4GBE
g8pq5EN3w64uiHGKGryNXzYUhVL0JbU90GpcXg/FRAejzKc2EkML6s7z01EhR1Wc
XvBz4rYblfsTghreh9+3qhzkMBrmdbBdTPdfW0UT4SbKrdd4ti9L+QEEPU3lz7Ao
s56X5Xf1mrZCFclC7qYjGEeqtOtx7e4qgf2EldJnYsH9+CkrGY5ZV3nDF71AzAnX
xf3it1iyW0UjDqgEP2z3FWJy90Pc9DRuPknAYCvKlQYacEixaXIdGU/aq+VeLp4K
ZvMGuZsNJT9tdkjBvHFhDqd/ApmUlj4YGz0vq3PQ6FZTML/MQqtlS4uBTuImvhu1
1K7pKhvtom6JuTt8wp/6cDOip5CtFkzfWKyPLj59CS0YhUwigvjfZtEg7cucdGnQ
gWUsjeFfAyH3v2GPuyCtvcNPdlJ0kRkkt9evTTJOOHeCzZoKxartV5qg0B2QVe3h
ThgBzfC8lZF5FJC4idCWP5yhCABn9dnW4Pt9tbAjhfn4Sej7qB20QI99SDoZyKYA
u+f5mbuWCwmi2nZhNoZzbCTX4L1oUBPAbonm32rRRNIadI83f22i0AG6w88tbtna
5BMKSNoceLy0AqS1mLY0b15KPfertUXQoeXoHD8B+Q/j7OWlcBMwaPChzauVcfP4
VQreywkUvEGC/O9YlRm8omSno3SHRvky5XjPNtQgyAr5xxyeONyazE0DflVck0nw
UyG7qWtSL6+qVzMvsEArQyxxW+UjCevHBIoPjloPjeXAKWjq9VUv8w4FGuX33xlC
YjndPzYZ7RNjHG+45qDJa0P9UYCeY5yGNr/Fy6F7ofnVIQmjm5XcACt+E2PAhXbK
EhXoSI3WREz3Z7XV+l4LGedL4kp+y+YHfbzJR1ystpUMNpAKJZxZWeSrJbiG3DaV
W4uVKW7ACZJZDWVD8Bu2xNF+glVwIrWjnLX2CiEB9X1M4976rnNJUeLn7h3L1dAx
w7CQyUvrR3EiRwj65iQk+t4S7FFi7MCQSVAJU8F3jBAePM4+nEbGNr2JcLbgR0zx
O7H91pfaS5fVWtc7H0++CH0hk3Onyfvj8h3c7sA/jo1K6I/5QwS9+pIO/eWNXz89
5ge14nDYlTWvLYjUfUL1hYV+Wa6Ipvpm5kGJJmpuaziq3mEQNyTYkFSBQqEOYfqn
PVB4pRS/00hoMrajbDEuyPPiV+qsIft8FuXJpMjV9fWBBOjUMMR2sIwVkB15TIxs
Hu8fcjWZsnFyS0sL9RB9zEr/6w0O+z+nIFAjMy5g4vKkSKg0rV3M+r7QIofmdHyc
P/kxO/6b/4ezDBniJ7VyZJ5aiwWB2injOS6l+Nfi1fvZMC+P+SPOzNLqKpB4kbkl
hRpxT9ZOGexlMRKwQ6WnUO284uJPR10A89joQPobSqVD7UbCHN68Gla42CI3GZ0q
3yiu1HLTJ2pxG94Prs5Cmf6Ka9uVwBdh2/pEZRbDHCwOYC+AnlIVQgKDazovoXuH
uIMhoduGNk1ZR2UWmZDJNqokKi0Kt75+ebtXTew22RrJJhoRNnqVvYHsvhqKk85y
0q3mMQ7JVzER/yOQfsaup6+DZ+/Rqdu/DR6HRthdRRYxr+P/ZsQ73WtbdIX51Wgz
jfYmkeGAIi3znyOaDAvB2807eNKw9s7X4UecPkmVmk5N/sjr95pXzwXLt+p4x403
VYdeMCSpEdjHS5AXShmh/iXg4QohOyMuJveaDGG1EnUl+LbXhIALV3Pi95RRkQ1e
6MuQIs2fsNyrQg4uJkwKpvcykcTyd6cdYbipnUaVvO3Bjer2FpaeIfMAobOiVGm8
ZV3tpCU12VJJRL4adSQTqNZv9FJAo9Gp9oyAsnt9Ebz7CDh2Xr5lI0qDCKWGCF5M
BpYV77QGD5WyyOtySh2l+ilqGalPXRla6Pybla5kfly+H7XS3z3H/2mqMnFuZR8/
t8lZnNMqLFk1MH6BhopjY2LC0CPOtWqNkn1DbHQhPBnpzGewkm4geHGE7UuPDDrL
+jU7/RinvEMrs1cCB52NiyiHXEEeHm99u1Nf2N0FyFrpmVuFkFA75X7t2WxIAkSm
6GxBpblQWiY/btKAOFav1NVC8c/83jDethuO3bnKbiXQ/zr5ye1J8hNoU0hUAcdR
0QY+Dg0YPQqphWgdqKYtfCHV92Wt3pUu6lqPjrkHMWuAPjDuUYIqhydkKHlbq3QN
dcgXYcMdCzHZxcrDG7dvwlO3/qh2xhhBZASBOzGFq7/LT0g8iwxQJJLEmQnM2a7E
AFZaLTNtuRcsswxRCHwHHxoOHCiBUbUCNyD+lzM2AxMD4WtYoCyNJzHI5LlOVqjy
h7hS6ii/aXbZYe/iDDQ0POkxkGabrGKGkb/hVogDOmlJU1wU9BLweLKKB/7pjI34
iCjMPPNoPjBAmVZGt3NJTXcd/Tb09HjGcStq7XOG0QaLNXAH1giRp0vPNiTll/Nl
bMIKGmlKanyRmYAhYHqXVdfAOI6znf33ygaUIZrt7qzxvj6zZRE/ofOGIiZizrBw
TSPAxknOs2dYM/zmQWpUGUoMY4imaMWlxEquUlA9x9atY2sJywV4kElFKfPcEBsU
3lkUmhPZPQs5v9Qibn14S3kEejRRhJs97wPuJKfjT3fEQJD3X+Yy9FlsLNkIyzxV
Ew1pjQMck/hVOie5QpJTonMlFXxTwRkwkzCuyDslBajKqwm2qfZ3G3HB2KSvlwT3
GtY4wRDItUGg66nHvoFsv1fN/vPtvMIdYEltel+KR52SIBbS9BV3I8CSqbIbypFD
0pJOKyq6Meo8VHYvrTdHgGA8ru4VaAoNnWwjzUp88wb/MlI5A1mZa46GtcOpS+d/
XsIx42lK3H3CbNyxAo+irxlDAIjiXy9n+nvSLvTYV87urNVTX/Q2JUTBVsHSuzn1
CT3xk+MdSCVn+UrctJ36ELtqGoi53boCIdmBtpTibYoeO3KHz4qcL/qEKqWeKhC7
pQJrhBpWk5ouOSbpfW6pTAPIn/j5Q2YiN6KTUCZLnJg6bcAfLcR/V1izJB8t0Bye
+v9G5hXdRogYX78T9hFHakvOHXJXW7ULhVp8sjESCTR3Va4BfHkqQIuJHDZYeled
ObDfhlvg1XbRuVVyCkYEmBopyUVXcbEu9Mc12k25aGX+2IscRzV4tW36Cum/OEwB
fu9ABPCRW7DdWu2h9/job01JpP0IpX+c0Ktyb/6oT1RdrHZouWUq8NJfdPoTYXwW
t5gYf1UHFyCd10/87G3wieW6mFk+7gFeJBfMuISmYOYwxcnoPfQ2HVhFWIX5m5pl
c+s/NvynULZS+pdczZW/3QTkn2cmT7NZVJkC3QX9rxbUXbmx86VFdharIbtvN7/p
s4EmaJP1o2OuqnpX+UtTjKbYqrn8P6GB2swhFv0/i5JEnWaa9UYMQ4wYWcvERukN
papLKRX6ON/F3THSVtbOlO8nHDIK1KPR1oqFs9Vv9vNhTlQpbqXXgg2eHA0PqIhf
W13fVdOJbz/R/HfflrzJKuyrSM8GfnldoxjqREFqMM8k+NEJACRHESUmfZCWKovM
xJzLTIl3hJx+fUIqtyTTU51tVCB8xZ3dD+kSmrGra7no2Jht+F6CewF6D39nnO6L
XoPu5uEZxTAY89BAl+csG1y+vgQ1UTMCf0lw3onGJNywVsh8tT6W2TUou8ijCLGD
Pmez9x1y1deDGf2l4X8+HUQkF1F+ZUL/hn+kCRphlCzIwEENFDeEARJmh/RL11YR
nbWuhtCH/NywLSs2d+QJ86rjiWvK+Vru7SAXEDjNi5SabXEKUpksFWWpVURAUUXk
bywm6sdkSIBjD0Bx+RDVESROcOWKmQzIOyd82TFWasE+ZaOUnAa+s9k8tAmlE4L8
huHu/SLj2Q6CrC3l1cWWhiwfNh3GKAyzNPHBGdRVkACtaKCa5cnZiH5fMap95GgN
Qom8ESqOmmShYAHi/j6I9eJQM4Y6yugyrOIn2MCiGxhEtPlj7p5iQ6JuWwyLnPf7
mN5aRPnHo6SonnbUk4EBwHv0TzQSKiE09XuoIg/M8lJ++pTNSeJ0/Y5FcRQHhW+u
7gQBwFeEJ8aCA3aWsowNYesjBNuQUEIpAKAKg8mMzVv110X8PNVoajCsPtMtqa7x
AEugFvdJgyWnfOhLFfa2tVRQMc/5uWNwgq3WlGzuW6gwf84ld6Nf6OdIgfV0Ftfk
Xs5NrumglYFb2tp6PnJKrI588BJJQ7Nnzxxj8rFYF16nATLo5lMjDFWl1dfPfrU2
YmkIEv2VaJrJJpsN9uG2dedvVOnDd/RH5FYWKpHdFlxT2hBSVr2i7mF1+3++4exH
UIIWRRwP6aI/ZAvFQPUWAFtupYBGe3kOuo6r0IulkzgD6Uj+iZJof/BpikOIkqRi
0vctX+0aHoF3mKkegVzjrNZsC6E8805kSSEiOg5smd0LWG6xNLSBwUBApZe0yP+Y
FipFek+5bMXowdZkEZn18lQj0V84jNA1xapK5cV25wQNjU+jjS4enelDnzJKGUUv
11ElohpwHyrbqZBXch9P0MdG7WZPV3+FRo5jtcj0lqkr6r/iJfshTiaGfYoRX1UG
FvVr3LgT64IfkYn9Q9DOcxAJR+QehTPzXDah7wCeWmOhsP1Z88TVakCcbcPW4gl+
/qysF6WhPXd8yIJswfGre5xT/hbwD1hO4ht1Seu989gBI4iA6UBGi3vig2klxpX/
cgKD4/aNsJX128hbT6X2ULdWPQ6OvpIDr0VBWa+GuNqhG+WfGCiKID9fgmtMe2qX
zUz4mo6qmp1LluxxbjVPtTyCi8Rk9uZLtE+ltalz1+daw3eB/F6o4RG9aZO+05dl
xWYctfGJvxCfNmOb3FmDZ0wpX+1/DisllvKYOexpqUhZ2ZsPUfVPZ/UL1crk/LwI
U63yfvUK807DW8anHhFwTu2IOSiPjpMFE8/n+Zzt3uM0FvShoOwjVW1EG9m8mfm7
gfJ6QLW4mRRsa+OTKV9NvbuQwk6zCBFG++VuMwaRGCz+oCuc6NpM7+v3nLmJ6FP7
vsVAMHqitYtTTCf+KA++k+IjTiGP5hspwvp46Nf2aC2jpHm9rvfJJsMC7gH/UDU/
4nZn99cRoAEVRZvsyPbzerEqsDstkrvlRcCP2KEWuYRMmOZt4KiXoKTTEL4kNjBD
JLh+B0nErkOvYDox9tlX3HJCVXQYD9ihIZs7PEG+MBp9cTGbVhrDNFDMZhkc7bz4
5fyX8dh8wVLLLB1NYN5QWK/SOE0UPvWkgyyjsM8iNPC4S/t8CAbgv1hA6rDiS/Ul
pzKM8JkAfLGLDuUVLhMaQo88YLBjOy8m3JkrIcZCavbR3UjRdgbxUhRmtuuVnalB
52nfsfUlOMbv3vB5+PmyTPSUy86SWpU14ouLtyS6jCf2Tk9qnXWevzp6TyE0yspW
7STsgb2Tf8aHKW5llzUEx6drgGcAAl6APy/DHW2aPgylngyLjYCslU/SJlikLwI0
tm0c3cWDYohtUgvgq4GH3Fx9+SPG8bFiSs40SiCcUQFweNat+4P4NH0ogOJdVgjm
e3NRAnZ8X1n1bgvpKVl0y4vj8rIEMSI4aLOmHssYO6WeCR62QIW80yacdlPEJ73Y
BNv3mvbtUFid1fDMHwStqn5nF3N34Z+zFeyR4kw6KFWkLcClonrodh/6+UQR4YN2
iibmxrYrRWr8Uo7F/gav+a9xz5VqDcCOn1SrjNs6tIqeFUc7x50Sd8tnEjY9M0Re
3mcRdTvq6CMhRYpokqSRSxbvY90wj7TuhOv6Aa7v1fKQXawQA5zZfFrMpSrTdOHE
9jblXx1+LIQ+ohWo4FQ38puhZQwn+pPAB9foOT9z5hCPC/J+uLxuoAJbz9bEmWeo
s0u0wD3kLCQcQKqp4H0zSrvO0OQvyshlJqsTsXYsUuZ1uWcxWpViKyfgpyrnlSpT
Fw8Cv5Ts6D5v/qHnr7nfmO8xFwiQ/sj/WDzSAtzTj44yF1eoY8a3a64LvOBoATCP
lLpQEuVKQq4By61uTtNSSsfPRKuhpgJpXMkgIdBvXYE78LrU5RMNSFn8nysvaY5Q
G4etfAdNSFfUKXDdUANwP6wcYLVAR7pC2UepfzZsUn4gwUtiplro4qaYJbVkrC87
T4vyIPrJ4EZ71kljBDjWHTy1j2TN270jC0QI9LNztyP77SGiebKfkjYTziRF+CiG
a7TeBwqisc2xf4hb3H9M6wgPUcz4Eba83DjnCytIIOsAByT4aREU21VjTlaFkSZt
pC0Gqb7+lg9Ua/3oOcJXFuovr5kdcUGzrGJOFNroJS+G9jRq72Gm4Tx5rBJY5fJF
3+7rxODOK9Finh1iMVTSKTCgf3ddf/2DrtHieMTYvI23lcRw+6jeTxu1xBroBYsC
PyuIIVYtrss58YXIzALdtyCJ5H86KTsTplRr8y6eS3ZE4sWll0lCCvV3Tum++PaK
JjXZrKka4B06EEntKntSqtygfNps3itlRYjaGxkzUQEDbs51sXpWp/z3Zi80v5LP
QAAt/AY3yAFyhqiIirzMsQA6/PjVtdvKBbNLtJJ4M4PHkEW0KOWF1eUgDuwd3eH6
lT4CZGypHbHJ3RD64NodBKWrC9XjfUpekNwQg/b0Oyx/Ckjw03TGOP8vUcxqEg6x
bQ3R0X1z+8XNCy3rOP1Wsil6ZczJpzRVCykikgN2JWJPjBbRF1IUWL4VhK8vRUGH
wELWmxvx19dpgJj/vgA3QbyEkkn7Nj02JFWAZDvTBn0HQTRFGpOflMcW6FwYd/2i
4DEdWFZRgBaZhAXyKO4Ic1tZDjb0prgHMDeVlwWow3CuySW3cBYPMF8FCqPWK+GD
2J0U4gtyOx+PApQKK8u3D2WLy9DnBP6LlURE+z3YkEj0dQ+80vl9NrA3ESJ1moeV
Pzfs8jLPeVZpCD5icez2TVs/wadxIsYRz9e0tKsv7W3O+ohFf63YWu2tMSvC7Zmd
32ZbNT1Eu4fOp+tBJUsR105oo5JTtvE/Fu03I8a+5buyyQBTo0iYpmV5+BqT5TD/
j+KWfE2sVUYY+BSUCwZaNSgojI7BRypgpEL6e340jfamr+xQUBIFPF+i9LBkNc3F
PyBMvWDQFhmCqN6SMhfcCOxlfF+ovJdw+GK8mDKGL8cV8nkqw/swpsZeZJ4OxLeu
1t+E0e4e3s31LoL41ZoeXAraV8fEVrmLAc/8N2eJcRb3u9wbybcFzCvR2roeDQAw
Bl5E9c/JbIWp3ZbXO3mC59V8GFe8OW5bToiWdvTWEd7ThtnDHRzwn3x3ElKtlEM4
Tt364JHOSi9qUVJu5Jy4uNvpSLp7oxsaQvRb87EV6uuLCYFEPWdMyXWXIaAi25Fu
c2tCsmfzuNGYD6OsWNRHmJzDhWUhgHicxwX7N+cQNs/PzbOfWZBCjKs5NlvjSTZp
IdsWq6DbAlvdAxrs3cnnwfoNvMYQLgLnceKAKaFT4D9Et9BcMctODrKHZHO9iDlN
KoNrG3SdIyBT1as7iz8L2kuHPYUe3m8kfe6235f7KVb1FCqLP+OVjWY5Jzdprq8R
AUEs6AshslPQhuBv9v6oGns939VK6IQkFMg3gVKQouqf/ld3Re1bWJNI9Ii/ry/d
PjQEFbChAQW2Gh661xF/CL9/D+98aEKyGlT0Q+g7qj8bawzu68VUootKUsPDflLk
lLRPTdRc4eXHtKKqodnpZP10E09H+Rq5US2u1qOFngoEwaUkbjxP6qi2YJ9nNLGb
M2DNk7iztNTls6J9q7O2sz8oayLlwGrXmcJ15ZVRnjWchBL1VH89i20AX8dJM6uf
CLZ6tNK27MR6oCs94zLlpykARVcmCQf0dkavCz/bWxmK4HQn2rOiTI7Xkp5ipkCA
UU0trbB736WWBle+ihyHdUhc2RCHbi5Na/I83LMITbbFWIxzeXlhDNbE4BiPAAMC
Lm7z9TQc71w50GCjT2kTN+yudBf66PAHrk77pNfGE63jGSffpZpRLDxmgC0SITS5
ACsTK/KkTM8x4GIILbQdcOdserwR9Is3Et2cOsyM+0H1NEjdvPzvEQl+UTJlpb9k
Tj0TK1F/n8qcA8SHsVoyv5dBNyK5DmElK4nbo4sYixY+IpgXzc8ScFfiaeaOWl7T
Wrd076CZccFFkQ2qPwfoz2CGtKDJvHyBio17xRkq5hyks3Fbr/VkO1vpVlnIvvEr
yoGAaEQtcFTbtxB5gOHN6fltHIoNPD1MnnxlKCpCySnZ1GcayB/oM6kKKQZCTN3O
bQo2NOIhjvDFQ+qn30xmK/FLBQ5I82XKOg+qKXaO9pyToiqVwBBxwK7EaS43PEKi
V1PZEqmWSLu05FoaZjqK2vyMkyKnAg4yvOui7m3BBV/iYGSPXCq1YzGiuxpSJPSz
3rQNwFNb3nZAV8c8JOgaPV1LfeCv9emn4b6XDooxm5KvGlgIgHAQcZ+Zl4Sw7du8
UlfY3cHPKiZ5+WDkL3zOQjRZkEmETRuXmDcRTueusE70MesCmQhcXs80gM6G0fuz
5tFYXknSDCFwQ4YlxP7UhrK+htqZd8zMJWoW/9NnMKIcRvvWErlMXe/mhFGcYcBJ
2lxtrQvwDHt0Zom7Eu3jxEAYVDXr2RAxAQIMqWl1SVVrgSyFtt88YC33yblvTr/p
AX9EJx+3M0r/xZNE4NlncZUiqJeo4JI7U+02bg1JJDppxwR2TLvjMZHC5Iau875B
FxDcjLy40Wfl7fJB5KTAi+yf9hkejhZjX3FEn/+ghsXnlRiJHwvEKXjl1NZB+roN
EaCRLbS/g2AiO+u97vTXfNBuOaafqg9XT5WxO6xKv6sAECQjcVhr0a8XNTWDpx/Q
Tcv61moSgIbXm0VUnubcpif0uIyiJidx/8Z8c4ntOmzX20o/OSkvEaGUNXxyLfi2
CaKgTKg0X1PjEx40s1elWgmRp40d3ZuIPPbONqUf5L9UUcRnhgb8gdFUVhtPFK1y
7Jq9l2N2rLx6Qfy6RU8EZfrKykSgWSK4LXv49s/t7q4r4WL3B5QsfPu95VCVJNIZ
jujOnmajgdWOdWdqx+dj7LxRng+vbo+w7sibBOkg7ZPyVKUVtM2n56XdlbUpLQXC
OXE577JkGbGQ12Th4lBzLrGourSnW0gpoq7do2AtVTlR0hMqzHscYqxHkW8Yddkd
A25aXBJon72wBEirUA4OR/YqopdjM4V52UDbLSsIx6MQsq9bYzXRKJVKt9SjNYnx
rQishC353ThLGSmS/OLgRySgtDQd0DkmD5vdS1A9QYSofHUL3QgJbt5f15PBucoR
0nNusruWVM3UCRAYS73I6faMpvqd16pnwMEAg14pSrkmYxltThMX1XEeXN/NKkQ9
w10yHzhQXL9/tawscInVXQH3dZahT6XXDsra0lZeEsoR3f7vhEVzJ4HqZz6wSE6+
sCcn6OnzWxywesvlZn1iM9yrEq7UJz0AK4G+KiPi8sQGMDE7smoT9tFLiJq1EYvr
UnKw3iaYzWI6SW/MV+siwa7sNKhpwDhqpJHGOxmG2ftkR/MRGrpfQ3iwmjFibG48
Eqk7M6EO05hNzN1XCr8pOHOjYPaj8GQeL57RlWYAvPEtG4XxjIzRN0WCyV3zz+FZ
Vsk+v3finlNO/nNBGhPbMeEOtEfZSuX6qB0Rw8Bf6U/XnKyObEtMuQ4m02KuxEIA
i2SAmjd5kNU3D04XVQtILQLLIRO5C4W4K2z+FNBfRAuFVbF9os2QmkHIu2WoJm7x
Vi3rMsbX9+Nu914RanBL1KPSbI47QO6hdhQYeH1hpqNAwERnYU6X5trWDXqAGwGb
HdlJJEHHBRQovuR+ucZk+NJdoleVTSf8h+eNJBZf0p2qY3Hx9lT1p0VDT5WlDtxq
cXHqGn8eYZyFuLCFlnWzLPRL3RFJO4rAPMl/4EzRq4KYPmV58Pw02qxxJk+t39fI
o2KBXtxHvB2fdEwTGxITXd4AoB95IE6zXiLz2RssWid5HQSmH7A4AYHBOm9t73+X
u++TRng4jxZT+88IqfGFAjjXheRq+0QCNuYJotDeeInkELK7cyargYQnn/AkeD78
N1n/Cgo2X4EK97qbO0r1D1pxrUGOjWDEdiC/yeWCVDjZWUwU75/IU6DOof1PhQYf
75Wotry1ZW6BzpWZ0XRUG30DLrEfuNMhKGGPQkT9ipMQSrg6QbCaXkkLeeCgGjLc
/Le1a3PkApvhHSjmwSqqW53lqvzfHjI/MCNaTNgWKnNl2k57QLZJoAyOyhyqnJC7
XzoPyO4olWmHCaYhs/LcehHOnqcE/xywMxKkvKDve7bmSPILyVHJT1WdORBI5L4t
TpP29tHPgaG2hrCp6r/Ov+cfLresNUZRFm65hLM51Tm8fS4YykHJwaE7c4wou0Gz
LsWFaSdUv+YkoYUi9bDif21jiGeQVK9KEjdVV2ShAhwtzur3hEBltNprxNxS4YB5
4zm/CZlgw4fX9A9MDjKPCo6xaueYjgRiGYV/pTEGEc5/L999EjQBpAmqCNlFQ5Ak
iirw9B21KkwrbfXxo4CdnYwm0NYt6xoyz1LPGWMLyV2pmeC0yo6Hted9mNzGn97i
JNh2DLqkXVJVcxTsuF4tvRK6UChAPSgEHpIbq31JA410U45ephmErejWpXHyLXg0
ib7a/PMT+tGWNxmq9pBgv0SAMBS7wrnt7e9UwZjZbz+MGjCSBF8s3HrJYFMTlKy5
77AWV03ekh4A3OVlwOge5wkqHO6sVhF79zSAahw6BzeXtHBNlwd0mCVTcDnMTygV
z1yOrJ2OwrQChSynjCIXLpU55SKimc1djxrWItpjTrx/RyqdqYoWqpi4XwDRbW6n
x7JIu9j7tT8PO28gSDWKr2kVE6Aexp/W8SjSBpGmm+5zhmnYpfHckQ2G4cYuBh9W
5B8gbXuRpsDdMPFibfKdswhwmpqfv9CBwroWUKVeMNBXUCey+IHOYaKTa8z3nlYV
LIHqEtajkh4m0yttk8VExHNAzsDZD0KOMeVQU53GHogSA2PkQw8t0eihrLs/BG8Q
4lybXY15OXtsGh1OLTRVfHFRTtDoaqtdgTQINH+Zohof6AV/4aQExSlyyP9FFwtN
QnD/rA4zsU0dr3dw1tCeccXkQIpMYFmtPyJxSSxJKhG8SGnLgRh45FcczXsgG5zM
GetS4aS8xHSrmliAlMNGSd5NKsoi8rV1IzkR9KsVH2iCYf45dWUvGEtJwJpcLoHR
yqOnqLst3FA9YDQ+2sbrsDEc2AV/zSPLG3BiaMkU2YIzM+FxQg+f7WOLNSStAxML
vIfe/WEG3GfYBBoa1bWedP3JMD2YYrhunoyGunUlhsMnkL5i1zsaNpWZ2LEkDSe3
fGulB7XnZ/eb1jZPA5+Y7NVHdvvunKnT6d9PVKLxHrd320ngcNJ3OnTXlljy/eky
K2ucBOaImqk0HsGH78WtbvM5OJpZYmKVQUippDaVykJduyAJv6RYQVHELVfn/8qy
wbms7LPVcZYqs+sDt2R9sO3B/ULUk6kTzqscAk0dB+4JtXUY94i6vnXDX7BYD4sS
KglOGjOofinBl8DqNnhaPzAVsVmcUVJR6jaHqwNcHdbBCTlchLfrLNv6QKJC+Tcn
A390OkNIyIudMf4lRso0C3Yuuv1wPHJDGFEO2PvoQMItfIGGQwwWWZe6GxPFwFSx
krWale77lkebyCZ9bIlgr14VRiviVvYp7jAwMUIrw+4S4iE8L2E1dtCRgmHODvaD
R07HfdFll4x0Sg3cwEwS79LwfGvNlst6+TCI4wp35QFQ+pj6/viuUY4Uu/bhZCh1
GTUQdB944hHt8FdxIuY7+ixMR5qI6IWofDtzhMl7XCW0Fe3kp0dEmt4hTEVTYiVN
V2LgV9KY91r54D910iCWPAPDIuhiyf4BPYWMkq7I9BnSmnMfaGthYGSC6l/iXwNu
Zydj6kWFR8B2smARtLaOeDzyyttMXVzUmzJpJwC1Cipa9xy+ngbfK+XVHCTUIKKr
KFdrXDERtjnwnr+Z0PMVBrx1xZw/lQMVF/IDu1ppqq867rRcedJ3R/h4c7MqLIx2
6rSFNeiL2LMmWx62vo0vKWfdDtXN9hN2eWumXPxNVIBXMTV79ij35AA2caO9oOOQ
5EcfFOzPt9SBkwCDtHHms2x3cC/VtPGLiijp9zeOhkroSKOmjfE3H4GIIrS/7uLS
678Rd91qj0OUZj7SSfBADlYAeAETs5ge4YnD5aLVlDaSGvhApc9U1BUEO8GUjlRu
pk5BffBMFDrpwpJz2beNJzT4gmlrj4ycaivaVWTjwjsGymDnIWvqCXWve+HQyqvB
FYDEfxSyCzqZ5xccTFIpZlAp0jT6UmZ48tBs5/ok7qK8KAtkdTGDfgLsaU4X6WtY
NUjk//sK2wPHtxpk9pNJPNehvgdYJJvirMomTz3TTbqjjXtmG1JPPMtt4joB8dda
WjpjJtd3bqilpKvuphK0dWMdWrkrGUStuxll4dqm3/AT2B3hddmQ4zs88QLvPiQ3
6cuLxyxDQQZ6RTwuSWCaRbgQSe9kbH46np76FCfbmac0IxXld1NgQDOVFlhKa4sc
aNpISqPNJuVy0+R9h9tW7QqZ5rukm9G8pWnqRnfSkGm+gKC2Ndez/9aPMYyQUefz
N1OHnBewqlM9o6d7L7Mdodb1ZcbE9H/bcoEfF/BfKiOurFHXllQaK/djXSAvMB4o
KzFGcObv728nrI+uPMUhqqUC6DO9BYbx4qY/oGONTZUpL5eDS5+YKXtcZsAPz/Ag
+3JnWwlXnRGWm5qGx9u1yGFipcEMhMyWrQNg2CNz6Klsf5nRXUCIhQ7sYCq+d01M
DmLCpRO4jMC8mVQ+nTzV99+MA0N6zY7tuujiUKiqX7OsRTLHwgrwLHFaIKK6L0TH
ARzO3krQ8rkcbxmh1g3mBtAybGWhXB3DbUq08NpvDCJBAtmyNH9BqZrXuoelOHn5
tCi07RkDwVRmoFxrJEpkJyLuWSPLNDiOHYmUO9eXu4DMIc9QtG2glPBH1T9xDC/r
injH0mmib97ZvmzAIUKxft/aHbmbaD3TQLks4XALcx73BkWP0TmwCYDvGdBKbvHt
BYb5tH8BeDiMu4Yum873nVrwRS2mpxG4xoVCR3gOWv1C5M+HRNhpauK+7ZJzSWAC
WnkYNii0Qhceu1fP+CrdwYJU0gqLE5puj4OTd3AIiy9usVtBuHsgHd0BtYzEtSMz
8d2/AtHmeaA+9vD7uAqRiVWCatWQ1XF+A0gWgr48akNlXzgFbrjZvD41f2867FFT
t/W9W8bCaS2LGzk1TsD3ZuOTVT85PPH9L99ol+vLFPEF2jfzKILKHqKvkCJyBLFQ
cncNtjUlrIbenlgAfMlAgiPvy9KG6g3/b8k3P2Y2fyLaX1HoD9EoqMMqMBlUf1yy
c5jK85b0lw1FO9anL+stGY01agzs8GWrYykhuW3Z77uMiIibgtQhA1LjYrRcE74m
v9eIdpfDz/7sf1QNzRNTOIME3IFyJ35IjJAKnTGts+eVQhpWkJmErbKyHfqNMVLj
2JUltNAXNh8PWPAtdJ1x+goeO9mpjeVXh/t3JMnhHtkTFAHRiXyD9rbkDWfzJbJJ
sEanhtIvRcD9Pxyf//s25SZ+zYZxhVXU0Njg9AhW++N0pPKqXBsGKVWq47n+FqTU
70uIF82CngsRgRTDZ86BOUs7gvGMrE4ZDtBU2C9rxcBp8bHOI10YvbrSy8SBvYcV
P7V1boyqu9WV5DsXW8/famMXttONX3/xre4xn0JiWiQEzJa9LphgN+PCNFUXnAvs
fCk4+f8q4zv0Z21L/TiBUoFtb3R/RbqGcgEiQ0fU6jqZBTdWlK73rN+CvLaiyHEr
K0yiZFDf4zxImoYa3lhjWI1kXYZoiS1WVFVVi6ODC76AKGxz5GIM1k+qXyW+pKGs
12dBh+HpKFBpzD/xZwTSKmldPrCx2bYcFu84+p2m6NSRdRXnRKF1AgpxAOW6E06G
3eULByWPBtbM/F8ODUFz+L/Z2zMk9u3T6jthgDOPT8cUaz6L4goFBJTOsrLjtJPS
oH3xHg32pWBCj/AMYDjf24/bnnH5OFhaKuL6WtLjOkRTn6gVilSjXKMQa98FF9rP
jo4ftzGMdkJe8mpjouOfUVnZitX4mlRs2qUtwbsc2S+Q43Nk5efHP3r+9MZLvPhs
S+BrPCURVu2qPbzFr8z060o53JSqWF2bNs43VxLi0KyjzEiEb7HW9rPP8tCDBbpa
vZoCp9oeEhWnhB43t/ecwAyPzfW8ocrwXEd3ayYIm22KxDzHxyuv6xQ2uiQAIEYk
JsFObhAKW3ud1yHOPh0AK288+DSBfsnLNUV/3Jsc69cE6yo++2vF8ArTuydLvc73
CiK/9MHAfustohnlrPIe+IXa430LKUS5Ye+8mEwt0HuKql45maspq4HQZeXGz5El
IOBv56ru76BCbUI/06Gm7iXmu3ILT393GPtG1kRxagy3AxAUEL1lxomlCuszwjuq
a3RP1fIoxTwcnmPl2/QRbWdOIHf7VlGPWnuaSjCMNt/CLVjpkH5EIQZZa4nnlN6u
kPy+zgutm0tGDU5++iDUhdAxhE4vbwXZRpebV/kqL9dZJGL3i2VGgxwZigtIkfIJ
A+EWqqHpwLaMDxPYegLJmTde29JJaMarhgS/Z5S4d6O+l1Uu9EsU3dldqbQSOYEe
uhlysSm5s/cvWgK+6rkHrs442uZw3YGx6GfRlia+YTk7l7WDLjV4QMaEJwSQ0nxQ
G2c+OasNV2L7OaEOS/im4EnXHQVV8tZsj4cQDXNITAB1QG/o3r+F3B0UPMNp++0s
mcwLmwGx1aJgnGjoLtVNANjepkXZUmiqCD+Gxm750FU73n3/TILcUnJo3vX2X8vM
pST7J9BwUS/muRlNqCBVVf+1USPiEYiyAUHfcWqSzsWVMKpcLrjh5QsvTa2usGQV
dJYtIQplNrLoSYfA6vsslzB7mHRL03V6Hp4pZbZGddlFhVI5mj9HqNsywpmqKwOG
Y7zHYy3wdqPRVETA3iOg/Str5qQB3qWFN0mBNueNn0LS7LLkgNiwfXinv+Odv3CP
ZqbnI8qyzn1Qf1zJLhKZbyNYAT+Q+Xgk8fbxt8vibpombpHohYAP9x9N9XbgkvvU
DAXYpsUDuJJ/3q4TXnodJSIS+yOeeeNqjW/IIk+dhb3Av8iz/psVfiCXkim+J+oL
X774PflBwIUS4hJ4LupPdNbJnagJNyBpCn/LNGwgq7GGnx157DDB7YXaLmtvHO5J
GbxbbikrBOwpgO2cX+Eeb/mP7Cm7xX9mI8zE4pSV8tWRUn0jNd3jyywXvKKTYuO/
zIjvjfmncCnw8D3ffL+jKecbT4Ec25mdFqsK9iMzh4kyLZHTgtvufeorvO+tOR3Z
4jlTsdE+ZEfyICOWYTPhjuYxg3WCH/d5J+RB6Bp57eWxvch7tKeO61U8uYvpdRGc
kAkRPRkT4HjLj60OpGZcDVZFSDV4+e+CO8/3Pq3dKNJArt6VCDwai5E9Mib8ltdc
GzEieTJAHt+42w4l2Z25DGD0dieClj9DbgTAum+CTKhKJem5oxWn0VMHkiHXdDfB
m0jCyvrh1mSYSyKveCgCpEFUtc7s+AdjfW4lMeD5R4zGImYkmYxB2SvrMoP+HPQe
IDV3D+a6CjOIhGOC6/BQ0zVDA2eRQgube4LFADbkpha5QWgfarP6YYukOzVwZ1Y3
1MY3bYU8gGEWi6av0ORsgUEJsi8MJ14z73rRD4jAhKfEkKYDHea+cMbPDu+icH/+
w8m6p8eL4yj1jFQ8R79NGhf4ekcAQIAwmH8EQE9Fe6DtxM1CHt2Wfq672rHE4+E5
a+dparZfWq8w1gtbWVyFZNpD1Afk2AVLeWnvy1EPL/KWRLh061GR8cLt2eO5k6Yk
qOiiv3L6yZlq2iwKjMPA3kC9Lv+67/PJYk2tXYF5ur5+KBSdoX8uKQWo9Jp64FDY
R3TB+nVcMYloYj3uQ4g6Xd0Ga1uJjETINvaeJ8LNL4nJ5c/yODDNZE/TMyDjZb2A
iG1d9HVErhbzlJoll//LZPe7GXxl5/GGb4nQ2xpGhC4mfvzk6IGLPpG2PC7qXMFx
JZd4cr1ZtQ9GWdraQkTYs2+NjRW5EGiaKhsUCuWv9fvXT1XH8xJMI63cYCmNqdAb
vk+bMM6xFcEGjgFbZi8nmhrfr97pATdiCNvnmjeRrKuKHd47cV3Tqn1IMX+a1K5A
sm/ulF2pYqIpJbfrJ2cluyxDT8Z4O3OY3i3v8h+GI5wnan3mT5d9A9j89HWF8LN6
0mBqRr57Q+NApd3NRPce+7GAFbWlpk97Px2RsAn8vMHODE4uwXD57qWWB4aWHX3X
DqlTStP4uL+CN8ah+zz93WMt34mSmFkXM1aRSgr6bvWcwp8PzYw4WpKXjdpBNNAN
KEjhrrbkC/yqt4j9STQ6lj2fKCKaghrf3jqBa3p4+5Ie8K6Rs4eDWLbgNln4IumM
rc9DZfRtKuJneItG5ws0Mm6KbwACgH15IVX6yau5aaqooMh4HiT4mrGdxsRV12rY
tnhD7382KGWFTdZ/WHyjbnvNKej7X8Ny7DsUsTpi1ViR6MOseFvAklJTNmu3Km1P
k4aIXh7ApTeNQFvB7IHqXsVz5WG5HFKR4Yd8xfHTOKP9YzzaCjTvrBqhzOoMA9D3
EF+Y99yDXIOrh2utZktHfOVLcOVB+umCLJXpLvFXu4lhnkaPyco4Znkkg62yrUTh
YmBRA98kPm1J4eWmwgW9LXAPoFaRonEfAfCUdfv7EeoooYEoyzCQ71L0Qh4GzBPw
sXElK6i/DgQ1rPJfCTjAvb7btxF3t+nJzC2MMxfM2gU+UcLxhy9nVikYSVcJSIUL
fCQkX6KPh4yomVz6tAAW2M5vuMOXWXDEJM/UfyRt5HiOMcEfMmTBJISG2e9D5+1A
QfomYUlHSUAMRpZ2ujJvxuk/YNL8mImvdlfegsDov01NqFjCYZitFK7wXCU6Wu1p
ULbik8eUfoWEO1Bl38kzUGLd9o1IC9ZK3wsSwH6NnzfEmCPJSOyC1Sh6Oha2TVKo
oHhGIftbQh94AFLxsvGghNGonHP/V9au0ZHoLDrg+PMym5JHQp/wpHnfICv3QWzU
1kVzTkEhpWBHbamQnfNoZ5FTdBxijVaCVcT4FfKiIqhP7Uavln50rceyVPPiMS7M
hkftV11zu2nzyAJR0trCAanwZgJ+u3arrx1F0SNHv5MGx2mXEYEvt97gK5/XFOrY
nOGlxbDaxwpedq/pInFmPPIUyFY4z3CXPfIoYFyMaSKIh0bRZK83c9kpKcRwi5V2
2yr0UyLjodcCHWD5ficf4SDdl7UC1X1iuCFsG1zl82bvo4JJD3fO5ajLfXEyY0Mm
7RTgoHmdhFRbDmRj+cidoRgU+ra05R4mkzEoOLemtRy1a0v2o12t7TJ1ZcvMZnAv
DmTOUaQyy9A1/Ls4wma06VLnAXA28IDok/b65w4TveBYCSN9SqTh1HGzfsaUfJFh
SqmyAwl8BjBXyIuiJ2ZMomP7i4fr+ABxJpfOg86GYCUlf2XPD97b+gXyoI/GBXUx
4cKaml0dzycJtf1k6JzyjLXodx/SR4fYLTdi3MvTqwJDuV0BXJfXBL9BFxiQMebO
THtu3uWFCVxPid1GOtB4u0jUEPRrB1tJpn36/8SMK0NvsVqY0TBgqyRNT18L681u
Oglkny2MFEW/V0ZSIxuOlJduTP3FDpKOZuz4yAn9NAB4KRi/4N4AbsZcH8FOusfh
RnZ4pDHZ1oXmXcWew4iiXpzm8ByWRwyhxH7yanN6XuzpDXq5LISFsNYbPwSlMbCo
6crFGB01bnB0lbBTLbFF7zOVyH55PNduDdjjl1QTbPpUgZtwyUIDbWJSYoyG5w4e
5FGiQnTFpkq4YCk47r4FNLmqTS0br19v5jFSJtOEUQhRvhE/rekncXgORatCLZcc
1VdzFQeBr5pTuI+0RApjjKi/9ZONEJ6etcFhAQkAWZyBVKYnfBU/Np5IxX554oWK
inEnA0PQUQMGpPa5p76ycFbCGcoFIwb+HRlCilOnAL9MAVZZbQfLW6SaGg8BFlIE
hpOe9+5J4p7R6dwwpKglEqgTDLVB1zLGatC4G2su4fTp2YVw8oWOu/WlR3xi+4Yu
gYk6aHoCL04bJQF76edv6NqWhqmCnIRU8/iDN8S5fjplYfENA5RAZ34iBIA20V3d
gWulkz+0lexCGwv0CEviuegLk55p+MIJAKx2jjR5LcJecr0jWB2O4xzbRmaZ5Ldx
KapGXJeyljcswYi93LStpYXEBzMnHKmxkvqRAkCWE7mHE8JY2PK+CtPMTUt8rgd0
0zuOSaq1kbfJ+Djy8PupugBDMuJfSmjBTltSwA0gl1fM8FqxV9K7GOW5gUwZlV26
XFTAkn4e71Ie5BP96159PaAhhljwzJvvqqSDcEgwWe0HEItwEC/Svhc74Hlb01F7
aSKBC1daOlXYiZ9ZvjGMqkWb7CQfEcRheprNGNj//8J3lIv5Oq4C/aDncM8avI7a
0DO0DZF9rDPUAD2pGc6siCYiO0AowZXsiRBjGptsXD9E8tfsmkhM4ChKoREUdjnU
PGliLEl0OQI/SOG/ap+hqFKEcuEkLjYB2qIyy5Ty1+U5ggxm7Zxeldb8ApGStxho
n0bSqY0x061NapOn+2gcfAuillUtm8sDASOvA0oxRYUmBxLisdgyJe3y1/CpqZJX
mxFvgIsSH84pq7M2Nk0s30P1mLQx8hrBRb603Yd/Gpn3Gp12pa5oOxq3eP5qOtVA
MwA7/4bfB5vHQdHx4E75E052+F23LMSxUVkQmWmJtRs+ycd8MMmwNPUuZhJJBqPK
7dEmwIM5ru0ARJRtGfy5rUoXOtILBjflA1ZvmxL6FWqsiurPcnKu3OP+qG2VfXTT
L1DRo0MITTBBUBXjhm7WtpzOT6PMkpBC9N1811FhXUX3DD3i1oZy7hVBPdtx5K5C
rE4z/rd5LXW4KQcPNX1ucYE89/tf10vrBx1yNNR9rpMtnfqI2j1FC+RWJqnSg3nj
3WSORE8muXvAiQUAgiUVfkA+le7SDDi3ZaZRvKG3qjtsK9M9QBjuC3Me8eT1JoCd
ovVUWmbYMATm60RqvD+Fu8Cwd1VS6rCF/LoyP602GDyIfP6gq7t6carczQmoOdgJ
zaH9Q1TUjOp1A96Z0dzaxNn94RpnIU/xKQEqvIoJNjoBO7P8gAR2KXoEwsWIGoZU
+e/nkeS9NcBzoQIFefW8rfRB9bLzGwZ2P/DlHzhp3jAglAp4Sfvbys/sVHbNMH7T
K+w17Xy8xymyq3h+m+5QdSU/frIUVoEb68a78h4estO3tU2XbToTvBE4B0Igj51g
cYPKQJeWprC5vicvLImb8Biji/52cFgfvwPTAXz2NrmqKCh5YYFrP8pkp1t8mCNO
rEji59ifgw7El+S9dXu8r0aVs5D8aTKWBNjyiWHNhW9aLPl0pmGJr4BLgg5mtrBx
Hs0q4gkzsPlQKNUCnIlX+HZ36BEaA5kKQkeL3ht0rhJvYSTTpgAbu7eBcYc9laDu
N1mgjPu0vTXJCtWKKflGSD4WHusOSRrSbYaLx+9cAT2zAERnuUmrp1Wth4PH4sAr
5O/6Cq9gm+I7UljHO7iD04Javikyto4jnwbhxlhnHu9W4F6NxBEh2WnoPEm+URz8
Hw2JDsGO5iNZmT7BvY9SD2mxk4QRgS58b/TtQ5Gve9zz3ZsYiqezoCXvXOVs4ZZF
vc8LrkqoNIHA1CsiJOjbipUXJVh+HfcNyTPsHhqMjytkeIrJfvVnC7iFaR863mCO
HHkNxWKzkWY7cwOa2hl3y+1mCpIz79eG52fFbeTCiasdE9gyhgzJ8G4S0yQdHk7L
BUG0v4zDqHi2HV2NqN0g5WnvS/Q6V++LwAoAXNU4KGky+0Xb/6revsgtqoYYGukE
HJJNumdRF8DDToycJFoICzcNnQH3Q+PzRU07qGwZYTaa4O7YBMeWkwKaelvnZ2pT
uuSGp4UZ5QOdBCmvVpB+OuAer8qXygCv3/pogk1ESiwS1wfMAiJ5xQIB4aW01x87
kECqqneT8XQbjUEEdYWkqvDeqQwgWaG4PJvs9zy/08Q3TFn8UdSxyfBhEzsU6tcU
zCwIO68nT2qVXFMVZ/b8s5SH03srmMajXP7dL0EH7Ztn376Nh9wtzPAcOW/gxujA
nZ/VjX+/NHQBbsImbd4e8qIui5ZGFQkmPxQ8Gdc1wIWDpNZzAO6KelFAfYBPfUwQ
ctlXeakg3P13fawC9qIcAG5uXTTFc3guMwh6fQbQ9a7tiZ/NC0zF2uW+3DdGMyQo
zHQq9+Q2rc8oYdfJLXQtm7o3aqs8FXrafAoI1worWurhbd1bOGXhSyoXah98Cb+G
XJ0h6FDv07bEF8pSmlo89zobBhH7zCKOfZ78AFMwsx41ryDrMapJNVVPnB631JmM
DJVwPzo1dQLx9yEQgMQI0G4rBc8iYHwUmNrGwcO0hg1MWC6/5kHQNLuUf2H/t4/c
3THQotksObZN+C7KycJVp+BDgBksuEkYFkx/u3kpwwYj+bNi1Ewsor2CbrKOm49R
k0lyw37DzGsPfURAw0OZzGTIxLwrvBooCcvcPibj7IPkl2eDRSxMUWHcEJnEtkcB
fcXRbfLy8wkuf/hx4xaHOftyPPK8L+3tZ6W5/Uj6UsoEb6Bx9hjAUghm8yhfKvLj
TjsVGToURCWQg7/+dT83/2qwq3TW10keJuEszJg6ySoaOCVvE39HLCeX8T3a4smT
IQY0N155KKICBxpGd8yVAoEwOFwuTHeqa41QdE/XM8areWqFJmOMU3N+ir3g270z
AaWUhnCc99pcBlb6eG3hNTnP0XiouHgfF6zqZ8tZnu4x5YFwfI/y0os68RrXQweD
vac/Xza2P+JrcVDaci2hOpXeWopyUSJ2qLjpSOdkMXbkHoy9oBy78zYmO4NCWx19
dnSUMPInO9VNvb4OXyXVuCOFuT+2LbXNDbsUAPvwM1nbDhKJH2SGAJXPLhp2IT+s
oTbHofx0QUD+iLh7kKdlZQ0mF5sNdTdr+w+6cLPxDPhd2/L36MKnW94BxXyGc+e+
RxMxOfDxZmHU7bJ74AOdvKZM3f77trswRz7A8Lth7SmjQ3uLyCy/2cYQTBT7zNl9
uzzsRsWKi77nfZEg0/eaer91ibsXNwFQN4lpLD/SzQodLIjk6yLANYdP8mX418YE
kXympiUALOSLEjdUcIqQa3S49W9XxEWRVmY79/8qMiy6gwcmk2Y6XycFfboWFy8R
7RdS1YsIbdqYw/2At+DQfmEj1mjURo+nwv3uXMHTJobyu3LcSgiHz7doAvOsA/or
CH1a+Kl9h2LX3wlm3H6H+cI/K7etZp87VAICj8pJNNDDdCmtW2D2oJtAUgvXRULs
YjlDq8F1fjyIUs1HVqa5Hh7Tm2vic7RoIDUjvnihojGRcTxt0ZL1sZpdt9z77Qfc
2P57apVBBXws0YPowS63t7lpykZD6OdeyEIDdqdPQkJ8QePr92BewOMjSkOcdGLH
9RLG3RAeUwlvvEL5q81+aZF2cGdZcBcSzrAmkpVmhB5/ALnw+KA4kwHVx8BS0qx6
n/qMRleIZB5rYyZuSnfXcvfOaV0kFPfnhrsbvyzmJVz/BO4SeIfUHhe97J0EJUDk
CKbWRbwEo3MTZ6YkV6i/i5FCuDgIAG6865TBpT46cgxojoCEecYPgbdSuhQEaFok
2NMt/fvmgmUtyIRVLF9mwCE9tRdQ0Q+9Rafz6IGMNJ+puoeleMtf/YrmTxs0bQ1Y
0ns5cOEGzuRCJIsAwILp2IVipHV664w/ZT02eGOZursGyuM/JV9ceafmWWB5IIJB
Yv0pjndcj9OmPuTBiIjzkYVwpORezNQ+eHgYTi4N9owlYCw/UhSgep94UZwI1UUS
XT6xoB2gZv18kj7r/5eXTxZxxXuO50JqzhPVpNARu7SbSzrqE9+PkGRDS1Ex/K8p
zChfGHBI7AJ5d026xHF/ZY5udFfxngZuBvRQy1dr3VpXtuPqP6+lob7qf6POEJEc
h2cFjvFTaEZ2RmPM2ZWyY74VfqPG9aZzukFtwu7pCrCw7gwQy4mDudLYcTaAR2Pv
LyxxzdM8vYdgcoktsrylTD4ajQGUjV2xfSrcoXsMgVwBKMX7eVPF+Wns0vYnafEZ
rzMMSwsnA+rpohpS9Lcht3/PWrVA1Y4nuzOJ3WLmmNtJDq3Q7TjMmEgXttK+r+3w
sW/cp18lcqShkqe49lTFZTHk5aeWBtXuBzV6EkZTOSv4W9zi1fUFwlgtlQpEhPhw
zkINwsdto1L9cgR7Fy+Lm0Hp6vjaA7ZMi1ylMPOs10TIK8iguaQrk+m07ALw+y64
yFYkJ/2oBA+/6jC34bvPG2YCqwH7awYQK+h2tDdNFcKzanIYBJ98ZyWPXmzCrc/A
mlN3itK61apV8ZzJBddfTBTTivikQLX56kBtEITU1vlfchMl7SLBC3LGQFKmHSIK
BZSz5jGamSyV8za83TtRtn9wNyuoDapJNbgQ97PJNXWHVq9uyjuO5apL3G+VZvpV
CqBltn6aUr/kEUl1coXi0wv46ZaXc0obkW6a1HaqlzpfSmkldlwvFgjq/Utd5KpX
5JkdWDDz9WWJKtNW1C/pfIGAVXxfdzjqYU7qrQ7f8Glv1SdzO8jR/H+wBLTyDqTq
AiIU5z23svm5NT4W6D4triwXEoSxIxLbq17CAA6FRK6FF045QkHIDhRVjd9EQD3e
a7n3EQcsXYsAo3EUrV82lp18GxFqSzwBfGCQus3fYf1W+onqCItwdg8j3XRheBIz
B9bQH8xwU0nlDG2nkvLrz5UPf+25xPh/5JxzBwLu9dziseohIrSQw9f8vM+6adtq
l+Ai+W8smUwuIs3n3Nm8vLXu+6Fx4buDOkh4+oQysKuVGhnKdksQvqMFvub5CNm9
+v/vBrfC9MptbPEYu4DzVSjABfF1Jz6u8rO8MPxH+XImrSrIcRpnsfybAcwamLPl
YBBPBON8ntROCSE9ko2vTHAe14za3cpAGd4xaCHGAnz19l3Mr6SgrKFOfCo5qaAG
hkoB1qkMVmYmT5wuMFFO4PjFLRzSfbo88IU1sy0g1WeVGSJ1OvcYo1uAs2dUMdDV
XqAaIuSKmr3cgK0XXv+mykqoXpE5fN+tpP87CKLK+Uc97G3SbW2mptnX96zSkVdX
EOfe/Ry4eJjUdwOzZy6NBEcS+l5lF5H0EpYh8qBjGbN29yo0PmOduIVdYm1euH7F
lZxznZSbVXxIobIAakUh1002owJGtHKBk4sHR16zR+dzs7bMu6zCWYJK81B1Ti92
ztd7HpgxNBfx0iVF85ZADzS86FzuQcvmWuMFzdArUTpBZhCyrpm06qijOYyc+LGe
0E09PFHlBx2AUXFud1wMSgnGjshNyhjHr49dbgpaJNahzkqOQQxYjKliEE0ancov
DAgBrKHSR9rvSRPOCv2Aka7ntyOZqYisMIWdAykDkN4+Jh+TZ1vHIiPwg/I0y5vW
DgO8DCC1wIenR70cgTI3mfXIEkicf+iCSFXrh2RmPEHt2JfUw0GsN3BGS4ACzVyv
KKw3m3DGTbZ9AtS/KgkNT6lv/NrY9EaWuh9APxfIjPSRI3G/22S2RDhPNZn5EkZG
Rd60JnYnidbG0TsNdXJ/SpJ1bYsepmFvve0ysf9K2WuCM0ZNJHwHpqbyAWYofYWu
evSfxOmPYQkkDShiO6zwz7Yscokiu4pQuf/o4x4ckDcbXSp96a691vEYbNcHTNT0
Wc4IAxsQEk4uJyylzLES+PBwCLUgDu/z36SJrA7rYkdfM9lKnwPR/M8xNP1UM0cQ
CTKay1BIjysyVh7wUB0l61QeqjdMQ0piRg6tv6SabEW1DViBA4Cb+QfyNmLGiXJY
EfaSsXwK9ZSBRJu9gn2YQMizTwM7Gau+bq+y9SfDQSFxJ2+feJfrOwk4zSZ9TM+S
ys9bPoXLtbMMn2Iz7KrZSyDClqjumML6aVifuF5WAiPBYGaAQMOsb+rTGcbZ+txi
uOrwq5SjqvngbAk1HL5E2JaqnKmAi59H1iAb2E+1gLKh1FLdK9lNmbF/uIB2Fnj6
qSHTcG8Iuavvi1FL6oPYnlh41pXgjZ6PwRX4LzNW+61zmQ2fqq52o//kANbQ8pCG
s3Jqj6t0aW0IdkaCJFlaDiZhTa3WeD/Kd2XlkLNkyuLEW+SakUCkTfpWCsuTG+bb
sMyQMgG1r4CFB0ZZ/vbWHmdj3V/GSoX73PDPH9loj98/mS/mcm0dxlS4DJHTdEIH
Tn7Vy+wCYx9uxWNf50H62ygna6O5ry9/27cJQ0BkjWijqS2ZdyWrV0G/egwG73p6
FmptQW8yr3t7nm4p/WdXQn5dOTm+uktKKwK1867Xc8vISB3IY95bMionhKijTvcx
Avld7KI/91kS0981scazf+3R0flyUlLNITgBDsCVjj5qHYzFcd0pZQxnPLuekoo1
MdMyEpEDvLDux1g6nzXbx+cqyLCadtr4iOwmynsyzpF0YAEhvmLfE0Ia5q/utN1Y
jaqZVA3gneJTL5yneMA9+wxcKcHLerKqvOmnjEfQ7jz06khsQtAo864WDhh5QKld
8JRqinqnaq+MFy5JBuHkjPHKN/X708MS3vP3jiNaDpJAqOO2okbM0MUDdPsHUc73
dd2N++t4iyo/3V7fozQ2QIs7lqAJimwZjSXEqU0yaxYBtJRmvNEZzV/PyZ55IOyI
Z8xenI1/1bnNlrfg8huuYsLgzvuF3X8PgFsYwK5MTqw/7EW6gp09HCo2XnQYCmmv
hBXmBEdUpU95FPrNbPeNpMRDMY9lchnxYXg09PkJsgtC7EyDJvY1cWwPKoWWJITN
pJ0BVcpmNDwoiqu9JTY8c+iSP8ClXAnr4ws/GlNfucwLrmizHMIte52KcaLHjYhe
WFoktUMsytaAbIfzdRcPotNdR0RqLE73jBno0s0mt5q0FaJiyJLqtgfkXLkEfv2N
4tE1DGoqGgCZwzMKLuDIpHNcTV3O1ruBQtYiysb57zvBkHEIB/TzDMurD3vkGLJB
WBSfITYOu5IbHdPN6OBD+bmyjOC59iT2mpU3h7CKSVROjvf14uVveu9CQnfhrFia
let+tbB1ehTlHH3i7cGymgG3+i19DIIrXYqIymIcWX0KlTPf0xyutHSyVQcjL4ze
zdpwNXEMHSFFZBGv3Gq7wL03uKwwzKvm5iKquAXk8u6Vzj9JZCNzNowkKnMN/InS
RyrUAVe4imPb+VgTfeVrJcKHyf5fQSJr79aa9nLh5o2uJqKu8IypS1NblHlWKSOR
V5gd28jzSGbhDO4WdLuQEetAFfRl84Q2tnIUAFWC/OAczZAFFDLv5YmMoVQm/9P3
49y6V/y7XlwJeCK1GfzWGUTd16dv7TzScYmFMFZvtom1wm6uAeiQCYbzqiFIvcRF
thip0pAZH1Y2a92Dk9cP3PbVehp/9iRpVdSopOMMv68D8IS/xdfP0h8USnHfUAk8
cinHNWY00/15Z4AE8zPRAmwVeR9NDp7bYL98Kt9pcIInmsUYJNrV3lm6nsnKSeND
pbB8JeTD2gjakSXk754fIZv/uH+WiSDSNUa4bbwqc8FDRoL6GhR3ePXocpnZy4HT
SxNxeTEWptlIOMfDnrxqYys2ASN6AAZrqhD6TsQPxS4sVHvbyWiTaaXkQJjG7P4w
ByKGgqOnni4f1EPJQYPgYenfmjOu2fS/mc5ENwei53uKo/kNbyHf/EAUvDomv073
26up18rpZmsN/7sZSGn9K6bkeu81G3+Ugz8BwwiHKHsbd2lv4xhjbxTzM6Gs7PVi
l8gdb5ZlTmqPdZs09Ae1cNe0vDy6+7DgdRk2hMrbq70J0QvzO7U4EgRymqJONoFM
9ZvDjRNipBkbHrUAlnZiprHxnVx1N1t7V2aoHxYV7hDIvOfnIn9bzukEF+AcPKLW
z9lpuvuViroeai2fdEnnqq0CITMNfYYnQnQ0xzSbB7POOgXsEDXeZ+8UVpWIETRy
SuXtgD3aWhivU87y0JdHNK/ZdzxVIJBbVoHLsODOhgQX2keaKCoAen9BeAG+cchZ
NR7VBVDs+01j+dZvf1byN4cWsdVmBna0WnVp1IK6fPmCO3XBnbxxBFjRmgWmO4U3
UdUBO65BwCsUjVVx5SxyFrz6rgC3nwQ+3KbZAFwrXNMG7rscSSrVNljs5YzhVU++
jFnMe6GICkEYGF6KBhAwLiapXPwOg6bKrGxPW0A818DwV1lh04mJal3d8ywqirLF
4FXRc51+VdAfokuWI7K33ZsyBNVOs7NIrnZdg9d6fcPqlfFM5/iImuK4H2Jwnzhw
XD7AjT3k8XICWsEbiFBP5ERkz+SGsavbpQ5h7qK7l7ifuItsXYL3nn8ia/T98hDs
scIaAlpc3BvPn0Qi5aiWKsH82dUn0mOV//+H0UP+ZvmQex14zfgXEdFLLtC6RWwN
zXTCORgrxBCRFnQ4yyr60RmjPl0s/eyv44xCQteMDc00rOMDvQPjH2eC+Eua/q4M
fyDho+b1QWbDFzxAvaz6hnyCbhRHQ6vVCxTw8Kj6CHn0kb7xndBJL6JN7kGx1+uX
gf2m1En8HUj4DuzNoGTCifEl8FCy1NUImEdWsa2euLHqjm3tiMRvvT9MvFpuKwRu
U6ok6LS5fT8N37hCROiH+Zy/RqHEH9+kRI+16KTvZw0QxKGjlNthlnSKJH651X7X
GCEnkCbl0wUheROneNUGb/LUJH0LGuQvNNr8qoXtVvdByt+BFUZB5rZ5ve8lI6q0
tV8usRGwm2R0hyU6t5GuBr4znXbYti6LZQohxImso8c1+lq2LaPJwajXAmFR+NXN
+c1006sS+oJZwPvq9hB8b4F0xyAKjakynfPpuw/LBEFh/3gFTYMbilKIY05girL8
ytD83oLayWQpbzXLHReozRvjdOoo4FZnrilU9q7vQC7ln9+Ds5Nn4x/UWVYIAjn7
zWH62t1dNL/rd7IrtFm+J+f6ZJz5Mxj/uIDk3wt3W9H80l7JBO/GuIxyV3f9+aI9
yOe0D05++la6+ddwykJxEPvfbK2UzomXwlTYIw72eZthAktZCn3ikINYibnRqefB
arYhH1D6KGLUq6VfdG+lTCqA/v63PqPM/+hBfNs/c9ld5Va9yaG3u63JykUBt+om
02pE3BrLBIcyFZwZScvhc69g6YwO0kxtMdC0rtPhOCbbQ+xsPwW/fl1cEAP+Cm3O
vqScIp0omL61DMNIk4PunfRVwVsSLW3BG7quBnLSDzvrg9Ugju5ZmkUMG+VFyNt2
wUa0eadlZQcMGKKB5sK6ma/tCFr9HQ6D7mf5abRWXqNPwsV5r/1xo7ecV5J7Bwmu
FpYLeXnd6A92unfvxkQ4byy7I4qR5wa7xFumA9z1Ovq0LtKXe1xcjEWhykGo5/RG
tWMpogMsQcwtWYR/QwQ2Iv1efLXYYY1mcdVXY1ChFU0A42FglRtM9rzqr5rsJYm+
8JZqI4EQqIv0xnU4ZiGeBtK1t46SSh5sHS7bjx7BeUw7dxnI6cWSoWOPd/t4sv+x
njrlV9mxnvYbP7ELPvqAX+mT8uQjD7+xnz0F/RiLv8BbO51aAGUf5RFE1pWKmxx7
NIEq6/SMJ49Dpaiv5hXkUUcB6cy8BmOSC63ClliHduXdR9z7Ap07Sx6OEfJna3vp
cdFFjadPGzFCB7KysappkjmYj1RNPvqI3QzjeVeNeS54ZUR1WnU5iqMXtxQ/rQ4n
mX6A9uxgLDPbyx28jQqHibH2Wbe+uqw5VBPjtsJiEhOMkpqKCvVHXsbC89qObCWA
KBdc/OTQ+tvu1aG6L5InmLLDTuUVPM2RO3mBzRkgKVinurRMrVVItNiDclje2GZt
heeQGnxXqq3B5/3Tyz+OIr3ArL+b4EjCttUDR5dUmJnZzwCmBT2bKEvm15yDfLuN
7sDKGYY9zDnevZs7zTdEoZyg22ibj/xfLjL4fQ0zs3Z+OiNmL/ULOo93NampDCXI
7vbJxhcuTC1jwkOHLIJJs0vKFckV/a39f/IWQyryuRW9hIfNqmHHDbTCdT9/vdZX
qaGE4U6nS/Ty/Hs8bcPsElSUdDEvRfNnTKIj6FRJc9kW13aHZyV2BrnpuhZppK4D
WBjk/CObQqaE53fOXtJpAt5mtklH7lsmesfVIgaEQOCIQ1hu4cuSiy6IU2ofUdYv
BESZdyD/z3XB3Zq8T4U3tUxS5gj61Z1jM4O8C/C8iNPHsXw3Evp0i/2oiT3bAPyi
d3XbDBxKXLD93eGStm2jvdMiCLhAJf9YpAGikECeQmZKg8r3/iroeBDuRjpcH0+H
mblKkrxohcx4wgUH/W67dHPoT/3uFGe62XOzw8EQhZGrAGoaXXFQDK0obD89/uIk
CEt9u1Dnfu2S7M3Fnib89Qj2Y0OEoYEFz5oG2RqxUOyCsjG/TTWXWufl0UouHPbj
i1cD8POYX4e/NbeGill8ffq3MAv6Wx1aAaz/IQHYDrEG0gghuNO54vpb65Gi4Zv7
5LoW03UHUO67JfuJ/thALjfCK0SmPTR0yxAIUd7E6yIv5++coo7XBW19gTkSlvJM
ZSnVPTnFN7dEGCYvE/ejrMSS9JjkjSyH1ekabve/Otbb9IyloQQ9Z8kXwme0dUps
qKMJZSKSNdgK/A5f2fhYsQEkgI7hgC3ItKPplIeLlLdaUGEtRgQyrGfbV2Ep9LPN
dbssKFxhR82Cf1xEk1xCMG8oo/E63RLPVRPpfwuVuea0TRTK2xqJCSXC4Xqphw9I
kdgJCjDsRMXoq5pWCMhMPVd7aFv8OTV5IofjJ8KcaEiMW+/nq6zZ2GIQ3GIH4j3f
1/R2aQjrwomzLFGRbLrjhYq+bjMQZ+uoZmFzfruZuM4MhShgFPcvYIN5HSUzx9Wz
IOOuZY7q5ariTOT2seirc0EXR+ykWm5sznBN+itbaZh1DRbeqj+hz+b9E+OiMa1D
T1UI5lwCkBtn20fzsB/FGLvHywNBsmYIkZoveOpLqHBo8x7mZQINJKR6iq2Ssefr
AsbLU+MBWdtcpysk45Z9zjHoi67op960guBkltjzmHUp6Whc6zDOjTVy6X6crX2Z
go7sntZbHvlg5rxdPrSxe1EZBvY8Vp4FDPx2KXjs+/uJtRA1+iSgtPx9gMb4F7lT
pyaBuY06j5TBndepoI4QDI8rDJFSweNdRXvOal7AgD9Ytp/XhCy0QFqnGPZm6UkV
WU239s0UQO0QTTczHl2Zb7GZNq4v9TteL8beK5cHkl1WwC0S/BsC1naj0W3wdGzc
8qE1+qqqbsvioa/hxfEEKuHpFhXJJ2X/YjWpEhKjFzUhObtNL0lmOvrsnpA0F04u
NiTf8vsWb6FirRFoUNn0m7IxSF1zjRddVqAne3nNGWKSRYDsht2+fWRajCA54EfV
xuBja+rWxz1sKYihvqdkXi//3FBjEr7+pMh60UqReZc49az5uFSiJL0Pbdx3IEPV
zxXZG4nssHb7Wp9dh/RuHEqw+S37vipsl1cEefrOwn6LCdQNmVHkEYMb5YBI02II
hq9O/AFrUzX2wc4o9dMXrsZzruUwKrgCnYhqsagqqep6zbGepQ6SYL5j2ylzTiaZ
oWSAiswa+DQyzATFPgHGjgUz3Qd2sUup/b89Upg5uHnq9ZkmcFuJssB4IS5izVN1
mtruzrbpBimiUJJgdLKAIvVUj3JO0M6KmiWa5Oob+lmwkbDUvplvZs1dreRdUXEs
mmBLdmD9QEosZww3AM5gLBwoS+elE2Zeo8SlbeN8xTuCbE/qg0PZ1e59nUOBllly
wdC2N4kYKwxwSF9kF2hi9uPhtfw6T1icUgh1BZugB/PWbC95rTI/KSD4VK0nosFJ
5Eiacywe0sSbY+7PMSLSfrPWg+pM8zCwg1zWjPNtcq9jWhsmwbeQv+5Qe+ui+4NE
MjH7IEOxaj6+YlQAGDlLjB87Pznvbp5cjBQbdLNq/YPJd7+kmLD2DFMW/BuiEY8A
rsmBZ+QraLXpg+/E8q6TfpPFvI7QRwKIYNOmnHac3/xagMX5zbVgX2h30RVCVXkR
mJGJOaM6dC5RE9nqza4dH6oLapOmheojBGUSNK9Pj79nkgMQ47G2RyJDcBKMW98n
kaCsJEht3PCpg+ghRNnYYj8ZfhwOBcbkEY1sZeKpyf0kAvRXKoUUOfnGvkx6W8mK
1+ltC3o76NTGf9YZpySxzwtc9M/u/KOmfayHbUzuS6Z+if6ZcvFQnHvJkW3OXpYk
SXLkt5LJN0Fo/+SnJH4by1K8FGSdsw9hnwQCGhuzYVC9+8hc4M72R+nF+knugwGi
AtDXuLFHx06PfYcJOpuZ0eOddOgOIAOXvqCBVaLWux6GODLymQE8xOqiS/LLBg/k
QNCwL+2w9dbi7cIjzoVXACnao/QZ81WXfnycO8J8V8sGDqwDejePrVbvVSyKYyK8
0oiHjdfJGuXLZnbb8kntq7q7uSbmjkWrmHSnYhGLHQL9J3XU0YD7mD7rpgOnDS91
znTUkhfCF0DLLgFALG700ikHGluzwan09DQLMkpMk35U/5dNF1ZV1V4Yfs/NUH4b
61e7pgDOczRy/TEIF9ZKPdNYKeiNfdgF97ul4TleFIfsa8780TaGFP4u/cG45U3c
i6h7I/YM0A8AnF26RfpPsSvTJnSEzAe3n5d1ZzhwyZyRy7y8dDN+7+xEGsxTHoq9
Bxshoyl6UcbJaJx2ZMOvAVAML7T0cOiZcDq2SP7YMZN9i8EGhP0VHKIlzTd0qD0u
wx39Jv3l/FtZuNwGILXcged4Kkw3U8fVjLV94+M1SdL0nhn+NqX/ogueuOdLkNCZ
ekvEyGQdyq2WqI0oCy33ll7LFLar/kwvwzeEZX7euxzi01krx/5evNWfpb0Q4mZA
lyge/6CqFqGOfj4fFpE8jgf0IuR4WhHtT/VK4CIVvoNjxJF5H0yX48jLeeU0ZfYo
xZ8S0c1ousmNPTWkx/48BOYDmK0KIo6LdZUh+A5FQzLfAkCIXnfFzFhU3cQA24ft
B0UtFpambk7RsF3CbPnXY8tELSiGGIbSARq2Gy1ELnw4UDPlVHtif3UPPX9SE/+L
7yfDcFgkCyyRRSpI6rmDCWjWubM1TbWiHU81flUSxXOtO+vK//OMFmCruByno6X4
FhMSiSFw4x8luHz/WJQ4mHOcl9r0sztRO877y9KcfiDD26QuCIqnRfIBg/VfaAEe
uAcX3wf1qq7zuVVIK0s54lUxnJufYTUFHXCmgq1yrZpWZjpbgPuv7qZ3IAUobEXP
cFE2JA9jU0jnqysv3zH6sp5hoeXqE/abJtPJ3Puza5rNVPz8dCgCZEgqMARMk/F0
dScUcJYbJuSHUI590Q+k/IkRYpPq+68Pf569zF41EpcHSJtAqx6ffM/g4VpQNzw4
3PRCrJOJxNFnRgcwHFzOJ7dIjnmhbekWwBYV/AEpT0RCpTn68dpcomPMkEsSfQnu
2zY91fpihbX+sKCpHAIe7m8bsqxMS0pDI4ZT1tfif542elskhekStneO60Sholv+
40QYTBC4oieGc0oZriOJil9VMdyZTYrVHz5+fDSooRKfG/SDDNOwzllkmN8A4PI2
OJWzg1wGQlz4Dc1VLiQCyj8C5XkVvd1PGgI9JGP5ZV6oKnJU3U/V1RSB3KYsdL7E
gv1Dsb2LhpB7L45beU2WFvfkDuoWLWqbGrIbS+G5yJHTD6ndGNGOOuwdYlMD2x1k
HvAJjHW6KSk4POhgKu8t6hEAVJVxEl0l6My+Cz1ebkq4jWuPrASKLxR+u8r/5hoP
p9JFUUYMd3DIUSOKlPB8HH4gk2JXaDFVakg+WbAp1RQeC9G91tvI0qNbsyHyOqni
9wu3M0C3kxT4DxjcetpL5AlI9jmYHhJjvyM6Z7KyunfMa5FUoBnQXyK2H9lHb41l
GgjxUVSlrHXE5Wias+c6To7/kH0qJRlI59jPxXiwSRqaQohEKkQpkVMRJLs9Ad50
eBKEO8uPcZFTRXHnQyQVnMlKZZM7KaDDICvD4DJXODF/9tIhAbqTAd7DqzRX06Ki
fQj4MGH03BxJOtFlJPMBbcdg23a1STgjCTimMjW+6XLNqFB1vczB5fxTNXWh1N6i
MEkLVNDDzl/Pq4F7hZ+60sb21n5TISny5/DCURbSYH6WlUY8In1W+4V2rdi+tQ4w
ElVOMDNFNcOvzB/pmD58Csjn+Wum44QQ8uWQQI6COKpR5NyLTNM7OasIkz2AMYrJ
NbTTeUeEVTsgMiI+lkTvRQqzCAhSfX6K1gqZWu3Rxee1YcC1FCxlq83n4e+TfO4c
00fFlGvo5wldtEavVZSrMznHSW8W/G6BwL4++l3Xp9JP7ag8iID8i3KejbhW3gi0
tdXiwuqIQRu51C4yPcun/13OjPh7BwIaaCFc4HojYxxP1tAr482iXJ9DMb50jS8H
nIhDFbKysirWnqnMgVrDiSgk5YG2zKJcFxzwsCfJQufUCprFssdU2u2FretfzGQD
eNrh2nIFoVEPEiUkZ1dPnIh8+muAesemfT0vbEGu/iUlGoJk3rpuB6tp7zkLsifQ
AcV1YsAJaW9+MCoHZ5N+SBDj7o25zkLLrYTHlJuEE4qMf7vzokQHkT9R77DCnHWp
LcuneQ1n6L5KU3UEpu2DS1HV6xXFCxMgUwrjfYKDhJ0h5PQj3vqsslO9XHYGfQQo
1LHJwOGcmCZTH5o9meFiHkGaj+etOM29TW5f7CSfBAHAeFQ/zoBxlHTnalCbl5Xk
QW0wGc2hu3Kmcqw9ay89Wlze8bvYgGPN7MUv5UhKSNQpsp0TWrjTzNSnJ4AEbQS+
0zh+3cb5k0jy0B04KyPoK86MVtpOXvxQ7UE8VOYeru2HWngmiCBPsjacLw1S17rd
I93elX7hUmhbAvPbJQia92caxkHegQXGmC/4smh/2+jc7WoccGUhiXvlBqA1HdKI
9iUmyp/pHyHHJDNLQ+f1P/AUrbQbnEeF5mlkfAOK7f2E4WHYLmN9HBu797ZPgKvP
7+wAdvTSY/rs+vRTXzQnneM/EJB5yvF6UzLcM9jrbKnlEr5/TZOexZlVcwVVxZV1
goe4nMPuE1qzGSYayd3d2VC7RkHx+wWMlUfh7nxah9En8yvrR39nHbCNUu6VPxBS
xsOABFWbR0cg7txpG1/pxaKSR2IESKQ0qDfipKWw1YAhWzzgqFGuTcBZO6V4jx57
Ydnr5wIxN2+BNylRr3ilxuyDNymOAByq6e5yDzU3TC1fQbfRE2xDaaWkHg2SEBrB
kfrGwV0mhgOxS7+L/vOEUHCoJ11lqpI+mhbt+rvaUn0YTAVUppsobNaN2Bz/fS9u
Z4eIr7Gs4ktu5S2pJ6d8fIeF+iTGNgvIfp633DD+ZGCB23akbJRZubEz24oYxiuo
/O2UfH765mdHoBgZ40kqW2OUZB7gHumd5oQt0iG8Rhu42o3ZbXwBhZnh9wg8I0nY
eN/Lg7hfL+tN0FED6WIisUUO3P8mFRx8hM0qBvbbWoUlWhm+biPyQcxRpW0vIbUD
YYviowkp2rVT7PlqzqNCWTCA16YZyX4OmvuZOdRikeTnqrc9ZmwW6yKZ47kSOv8j
WMzFwYCscvD84+8kPXWDzAGr7rAG2zIj4uyGljJhw3hhd8kxbJOAIaIXCREucM3D
MFx059BDvYqYWtUWIFk/DtL4f2xh7MggfBO/0EYQ5DzN5HZi8Sc1+F+uwXiul6Y7
7RVoS3+3b5MemXiLN/CHn7Itq7Qg0atOr07NtjldPFArxR9KP/Qa6xf//BDBHGrS
U/ZtRA8RO7PJojC14W+UqGiLPsYq9mMBkB14SxuBa/pFIRIQnL5a8uhH5v06S4gU
5fSl/p6A/x3BKJdM/MFYiD6/8fd/FvbQqDNC/rnIQ9N5FQXSVORauQzL3FPZpXMl
eS4CJoLjgLSOGh0GoKE4SirXmVmAyZsLJWiIj/UEbW/g/k92Rv//GE18QvJFtTIU
YFw88LSgMAgjVCaiaL31XjbRumcBrck9qhIwcPAUPlF4mlelryTcR1W1AeMt/Wol
gEF4Lvtd9LvrL0iujHQJUlWLyPVu1stOKCYJdbNdUQD4UeBh21pohlOCrdyDhDAz
rlMWceZPJsJRhQF/RGRtpWty4J2vQ/dFU7xdO0fHKwx0FnMoAZCXJbPeuSUIVz2d
jMITWIpoxNjcrWvZf6OSaW8okqZKZzcPdgunr9s9oo8xeqPOZpWuRet7WXqSBZac
0w+YWqpL+dFAlpqdn27ozA1vEbuAIbHUOOGS2yqNRHqOv/aRFD+JXDYWl1Csh0oo
o/vrC0okjbPerMMO8lEWIXOW0SnuD5yCEPqjXWs33kiOlEWHUfx8Q4wzK+W6ficG
kcWO7rEx7+s6OzBZ2YvZY6E8u70OOzBpf8Cd9vOFOXZYXTyRFOE3pRh4RngqiM34
lwSYrygnUDPcMwsC6Qfv5Z2dp9qZEpUmtXkAUS1vcoqrO/ZMnNTBvlViKedAJtNt
uqkZOMJkDGmT1ouvO5ccvyeZwXyPIr438AmSSjKSIlGEbi05QlVCe0MfujNa4yzx
LiR1o8nOPrXSj+WOrqnomW+U5gEHloaOIOMp7F1Yd7Piz2DyC3C9j40NcrY2ojvm
thd1k2aGk/ay4od4RdVSHet9OBRJ8nig1tzdErVggysUDirU20i0I5c9xBiLFnV1
/s9zjUSclAScixaW3wXRvFhFJUanJkyZpFKcmsxa7Bk1dun3MX/aIV1Ba55sP3h3
disC60T4tZnBCBv4PekELvE/hgEc4Ly2GVLdHGcnLUu6QZmnzkhK9O925WVLA5gS
QCLeLE8Wq08+qIq2kY4kbREOSFLnuNIOvMnpxX3bD59cL2C7Q9SCnPsYZz48eo3D
YsS+IBkR5vUNgEh3WbdzteMOqPEVGLhg167a4Vz7XWpMNpLhiIbYU4bSTn9pFvy8
ZRg1Wmh4x0Z0sItDk5n9khW+zutvxLoqVWc5Fi8yOHBrDM19R1qkLwAQlhJuJh0/
oRF/hL/w2BfnzQpAJBRXmn/7AkIIN22srcD/62fozFl7CniejFBNMn0tpd/G521Q
sMJiolBa0HkKZtMIkYoRFluheZrXtOQFobGyuMfnC12Oy4GNMH9cKMQPbTm2WIbO
TzK1R7AC7FaDmT0w8ibAkGlueVSjEEaf6SrcZV+BN9S83LXi7LH/nKYCCk1wyJ7w
qv1e99VbLwc6fzAM+l8UZEgnRGJ+k+VY8sBuGeWmoG8MURX+05uYqnCW7ZWYE7wZ
LGS8tw576Bge+Uf9ejFF0dzqCCYW3sJWPNYOrYagMw+4HRbIC0lI99lev97mCK89
dHxwPqagSJ7oDAyrvMMtlTLvoZy0WLWgunb+8/6qY+MKk0QERMWiJUFNG0Z105W4
+p+OgwgsLWJJSbVvCbEE9g1eH1vBNKwrqKlg//TghAcZ0IKJ7QlObfbeVjGWI2ZW
ChLYDMm9CaVS+1uwcrdPv7YZaGvGMEuLM2JSMScO3xYn1sLreozmTZ4KSzXBcD0c
iKZIN26CY+RGqbIXbWn9kTLhUVOGirr2Heo1fh6bbQ69o+ysjtZqKt/1oS5DNDoh
vshkDTGR2/9hylpSuicIFamypAuJAkt5Dk0H0Y5H30eqfdWMeEviMhvE8ctLBncW
kifiDlnyWWBWljaddp4dV/icg0DEbdQSPZZPhjJ2Fe+FJcd4ul1zHeqhJZtacwP9
9XV06JVMtdSxL9vhgKStHmpSlexX3dXpFI7K0zsZr16sVvUJKXZyE6ZKE9FvAfVR
eW21mIAT0cOKpOknVQPKs6nBVrbIA+SedH+Kj7NPMbpvNXAwyjHLd4K2DmJGDnKr
aYWoEDLOM9WurPRtY9GS9s0AYS2sk+c5grGSuvb32oBK+MYEOt/wVEHywCU8JlqL
UNam7jD0/vZt+NCIbpbhQATB7bJTc7jHMOHbItqPy1K144/Gt3YzapoJ/z7cOmwR
mN+LXWrE1lXvzlQr7njZo8+Ym+oQocBBh7HFaSR8D14Oi1wYFInphwmITrusAysX
MFRNWvX79HzzrDDmdwgMYBogQmATyY0AKa/c1lnzWOFIpekUsJefkZmaR0BZWqyr
8V1WcKA6ByY+YblTWRn8Fgqn6CjjlhdZEBJDwMMw5PTkiaHgBkjdsTwIcdRGXYf+
D009TFRu13kZ21EVBN90dvFJvtZsl1u8dKUub40yNjXwgckfSvxrI+k7i9wD9Fbt
GjT9U/cGVHnyxzYvg5z5bqUFakIFZhKIbTAfyFBMwjZ29S8aPhG1Re1HWgj1DHX1
u/GzMrEYsjUiwrQyHasQDa+yPPuornLnQEc6WdQk5Q++BX9KtQJHIxXYHmV6SzJR
8U1kthiwkh7oaW+oq9zRtQ5WiL72oq4uVS0xhFV71UrEXzfvy2YXoEcBJpv/SDKh
Kdm6rlG6T5GDhrKYQDVDKrbsA8xVbXHJW0kyPLcTKW03J5Q0J/TkIxJMkENhqXA0
wOZCEyrrAqNkwvCF8Iu9CuiZnQdxXHYSd17CrD1lrKMGZpCQ2/yWvUNS5/397JDo
k2mFgU3xXyxbcjaBvSXzpYtnSu1dThj7Sh55idnS3PaKaAU9E+6zqtbVewyft1lR
mrE7CgA8XiInlI/71d1Bx8uhiUWER2g7fuxAhG2e35x0xH6zo5a2sTPN9IeJpG6b
Iu8SjbC2wYZkJnoIGMhTq09atwp7Xdfro9wGCgWoIgXZ+7KzylgjkqnqpcacLkAh
jtJeJl2qlo6wF2LOyq5PIF/7J1rULpJdUQ0Z7yVFNsKc9sT9sihfS5M2QVXkp15U
8UhRdLKp0mFSzw7bMxRM+w4O6O3R08vGtA5nQhK18xsr6Kcosfe4Bzk+I52zPteQ
AeYmqr/IADErw3da7INQy50v7gBt7rkr/GiG3fOMhe9s0Lko1zifglwMRuH6FUSU
TSBZgCo6HwX48aQJTf49RhYr6MS/0mAdvhJaW23YCs/+OWX+jpEuKFVOyxTg3EMx
JTOdYFTzTxZtrjG16s2AJKPyxLQDoXy0Mf+14/+pclaVwjG7XpQBSz5ZwScs1g1O
rCXklWxliFR9uFgN9VzWDdEqMVY5iiQq60NPKaRIxnPg+N4hj0yWbNZVIy851Vrz
lIOD00Tz1Ri6ur8TEplXh0uFQFSzg8+C6Z3GOjwfMgPPqRFGZKTG1fDiZE9GLaJw
sRlleHxbnuxO/ExTA4Wxa9Hodz7RSREZBejM/uIb4PeoX6kWvuRmtRegF5AXFWty
A0v8h864aWX07SeKHilU7X8zwm410sXjfsjTSaPTjY0xMjDK51zivhH8nolwiw3C
V9hjW8ONpkGmgDd3cuMYePGcidgFmLAB5ogtVySOY0salnK+hOJa7dAsqgT3fwty
OlsgKvYi1Uq3ted1RUkDCCR068S39EigRA1tmwjKGgvlD0uyHS68NPQ+D3saRT7v
RySKLExgUrxUGgR6xL44tDrWpxqr9B7HKM6peJboL+oZ2xYqkQmEnY7oLifw8LKh
C7gnXaGs0BQcin9cx+8bITEYoqsZTPjUzvUYIDRfy6E5EnQov+bnw7sow77j2RN/
eDsdAeP69i0v9qlYftBH/LxNhAhbc0MebWfO+8uD+qHdBvtD3rGzhIbmMFhFAcUO
vW1yPIXKpQSHFQ2hZSosde6mwFFRjenXV/nyTf0z/EX44myzMRxAfDLkJbp9EZSQ
ydYhpA1i492Q+hVMkhMuZGTEhR8URawk+unf1+FLxGaQm8NQCVlD53QgFOQPLzDZ
qvP4/a6UCm9r3iRVYfHEfVvkb2jV5F/9zX6/P4L+XivBbkJfevRKLS3jm7TwF+YE
rYvEhu/dV98ea1nmlmxe/UUdBARuan4BrPOV9N3C1NND1N86D02NZ9gE58ZbDO/S
Nx099l4+WJBAsdfZNXaJpLFk+qV9Tw9SntC7Mu+ZyLEw6jsXCO0qRfpC0P2GcHQL
4Pfay+/S+1M7m/z48Dk3JhmpkLQ/Auno1aUuFS5UVCzCFRg6Bp+/Zo6jfy0JZFZh
ywPEp6ZLLp+SHloqMWsau37roUik3WCBtVLjBuLcKfMjrTKG3h382R/MQWs983Pu
/UF8RwHVuPLdCwt+2oDfypkYkVCH2mcvPYdWi1irweF6Ou8x8V8/dq3ogzts3jJU
vIR0uC4j/TBnL7NiDI3E2I+yDWvjVY4zm2NyLToY5hgJuKAMlKwoCZ1gTtzgv0QR
EDfMVCD3JiWfebT8WGvjHudZsNDfjK1o/0RcudY7YLawZZzCWWOiIWH/M0tm6VRh
GlkPgC1k/HRBKDLhV0kd/tsJ/rYVKAzEEnhUiUCQ3D0j83GUpY/lufMdDUhvWxT0
TkLJ7+hGiWDvVJ/TZ5e6TQHoNe+aciPVV+s9mqIZaL97rG69jQRa5vnIZacbiNtw
aRI6ZEG9RBq9mj07cUIC24jgECq7EACyUEDxhkJhTU9IUhU6RtUUji991pdKbmTa
eBiVld6AiCVEmQD/4ev/N1Z8svmNNgChfMN91ZPc5r2QBwyFjyZjtA6b5WOEIq7j
k79k0lF++cincKmrD7n9vEfFXkHA9F29Rrvp+Bdy45GikyHM20MTtNGsZdlNIkcz
2u+dP43pddkYY9u0+EY/VddVh+PJHno7y5Qcqul9eC6jAM5adDe6E+XGkfL/qrUV
spllarbS2loenWhatiTDXLosQuFap1yYFlKbUKN0n8jMJ/xd6j0GK15A9JL0AgUL
D9+aVFafS5xKzxOXb1t9ZhsXry5e+wc/Iy9no2jh6TYFNpSmHGqfCEtKaIS8DCNI
WTkJowBtxKO1Bi9BfR6xQmKtO0EJlWWkmCLDnMRxnGgx5+Wl1Zyx6+s+DoPoGGq9
ndiAe4/PZWwV9Vn9P/gLDCrhlyOcULi6Y8v3qR01YpjTA+PB+Q35NezblJX8+ryZ
LcAcwWDAuj1nZOQ0C2fgoysm7xkEj9SfYES4OVNtUdlQGv6xpmwZz5+yGvMoGvHa
pkcNlLBX+gnaWxnIq/ydiVeu0z4ZRtKY6sFz7npOVZWpwi/pcrmegsTnUr7MuCxp
5H7J7H2D1aLdKFo41FinTPz/HRsmGmKfUon6pR16iXFdB8kPYrbQeisAQBbKR5EL
XfuU1qTFasVh1j3j1c/tyKF8V8OCmisvG8ZY/0Vid2z6o12Oj6FReVNZm69mwn99
R6+3WZHUI2D9xlQ3M9xPfqhPzWe0V1BuJmt9z6bB92EEzu5meoAJLnF0Co+6sJOs
ziDCtrsr0qgvwgBIAGcAy5UJJhS6XCIBTbj2c0wLwIEq+hQDb264SjllVfCWKdcV
WiXjNRpEEz26gf1rLuLPVejE9yvuHSC67TqGffKhhKsBzm1PSMYElfkVcZJbM3yD
rkWltEPZYSEgPlWfPocW/iaRosmyfAWBTHNoj0HSk2tk4uRDjYKl9jYbHKe6gVUf
aXqwpf3wQK61PSspGiUy0kzGz15UwkiwPlPXYRL4Ov/w1IxREURcy7NBVGyGKZjc
m2hNI63TjAS1VghAFIcN900pFXstCO+WDXJjbJVBDHkPuDFxYHYonwTh+CJG7K4b
x3/rMEbtxWY59qqNMFF/C+oLwNIThV/7uMHtI8+ImDXZEgP1o5F+lalaB7xO/bBP
CZvlO4Xv36OTkvkDXlC0KJX4+LvWhO0bMNi4l9euCe2XGE29tI0CztIFslG7nJjT
7pGQdaa6OXyG8GO6osnraJoABHVK/dy20V9j5fpHWt9XP0/uXXBp1gnys5j20biA
WkoF5e3xi9MW1RGmtXFPnfcMrTArzAikZuq4C8yqvx1kPVGdKW5LE0B0Ggmm2z6O
9eMo356eHh9P1p7JvC0LnLqBM31ADO0BD3rh6prWxGrhrD6VstvA05FqHux0DOqB
Wt/NbjaOvw9SblcNAPYEiQLv0BbQ1rGOqQR62eblgMdMGjHLIEWrnvpvYDbmLvL4
efRbhjdJUfpsUj9E5hX2SdNHm1BZC3CYq4FuuQSsy3MBOQkJBMkvkZPo6caD3Bsg
biKYahZuW0RKswH4z6J88+nB/+DnQfZzYqVBBjDC0rLXLw6NFlCn7VEuU9jS9/8g
or/kFYV0Nz6Pdv45iwYJxO+vMfamKSmVX+29PPLnDARhHgKh4Sgsn0iQPYBH0nn2
zJYURay19MI3EliYUqfpeuP308TMWOYHdjYAw7E/WC/l8tbRSS/qoIwDEZL4Kgsw
hRvPENioY7tgVwEgRO3VXtTemtCiXfgTgyQ2/g8iVUmgYmcZRBFi7ImbMyPokzS9
B9CQFMDb3WiepSXTGKanXiO+wWRKyAxmEzovZg/wCRS1u1oKBv+iAwsQXKVOCIIq
wvYnXeyHfHUpp040teffnMQKH1HJza8NcRLlY5vkCXQIYpoF/LvocBm7fex1VDW/
/5Mq1is1WLDHW2o4wSeiy8e89cV05jsqmGGDpWM2kU3PRO8hUrRL5zYIOJFirym5
ruFKubI5uVu1rP5AkHARO+mTZXKri/381s62OjOkFBa0QpQrI+4Ve2AuG+0R7bDd
LixSABDCnnu9czTIE0a7IhVoXIbw0/jiILz3lyf3IxvpvyjCK0bztGlnVVPNBoCq
hRKzb/NMLkkqt6H8c/9+oon1qsBaYvRegVuPA6PllUawSqylLzX6lPcwcUCUQu3I
xA5olnQOd3gnwOzRHqjS6gJ7FyWpzIUv6CkkxlMt3/eA4PMxJSecxWAvgIBx0fBj
6skxTcWDXFXn/ugoc0JLYYfBoSQUTVe+WVLMDbAq5AMLbIPOHhewq48uXKqMQwyo
BipTx/Y+1xsOjb4TtqYB31Nz9mckKgHARFD0EFcD9yJABrQwudd91O+0RCqt1Nfe
6odrKy9uGEMsI2qcTS4o9pWrlYXCyucGIkjLcRGaDYRTLe6sIiRkqy6Uq1Hz8xed
osk2XNXUcU1urSEQfR1/wYRu3oFQLpv4K+KB+PC90zaO7I9nwaOtetkpfYGXbRl5
tZsAShuX3JZnIjGaOMX+TSMPo5McMd3jxFO3VJ7Vzb3iZF/L6c8YW6LToE009neU
Z0BNzVdcZj76rNN+c+Adv+wOKzB2Bdsjr5ixvc/ZCSbMfRog7NbEOeYr2yy8xsp2
VL/Ne4LIgTs6pLkQ+q4gw0RWqMHHvtSDLFIYXdj1EvF60+PLynevgyTnZiAUgi05
pB0dwe4x5lZL2CdPSuVClVGMd0NXY6PHTkT4Tzrcq9OU8HI30bAk+CtDhkfngM9U
5XiUUQJJsLu+zItMPUqlYl9fiRYzmUFLRnLis1bz40+gmAGGtctICuDs1PVy9dRu
W0DL+SyJWacsU77uEDYVsu6RNLlWVcxMy0Cp5NzUgrd0SKnWlJz1VgTc+L/OiBYU
dSz8ex6MkmBeDGomXyEW2rtwlJ7EQ5wmfsdeaz4kw+JIqr5GFRJvykxQAYsciuM3
AM+uBiEVdDeAX9JKMcYJ8OsVlmmwpLPX9vJdPzPAyR10b6h4vRR6Arqgcxp7waWY
bdPZRMl2E/exeeN7Kjyq+nBP+NfwzjarmsbZeCvLMJjDmDoQYN1u6xrJmoCXmxs3
1JHMswsQKXe+fn2KWUklIrOvrzIU2Bb0TurruUnxj6JAGHXdEP5uqjZz73zThXDb
PJitcGhiq9KfnAAklLHCbr3OkFtDCT/o79f4ZZ3G7Ocj3PjGXRwVjSlWUoyfSkUv
X8O/7DVg/6psJ0l62UVpvczQoGjZnMTHWEX+cJQjk0OlbCt/0dpGSkkjEBmqVXu9
WoOHw11NGze6XiZwp0OVT2QJsQ2gBBnPCvnAyNdKANN33Mx2e0/pqtyR5Y8U9rNu
us8OFZrRPqF9czeIW80Sc5/MWZEWvBG8UlsGA0WWTtsOrKOhTGSo4BNfLgePcoE5
+iI0fI7C3c689DzdmrsTPL1amHn1QNie1KM7cCIaYK+4XGMLqSBNnkugzHB30A8K
WVBQ07J7NLLlPSHFAPNGEZRpBkTRjezz+/2Nw2dZQiCjAuYxZ2xPubKF4CvPOChf
rOK8kJNa4zR92Xn5E6FGPMLLwvHB4Hlv2i1T36k6LP9s+ONcTvBarYo4THzOColQ
+3QbIs9jl7ycn/6IO12kBY7xVzHKMdVqS41EwV0LlYRU510yD2Zb8RSRQ0ynLZHO
LG+hsiLlLazfL51O27EykTQT9fmT8cRhhWfcP398CO/ct36zabZ1QmE7oWS1cXhC
/KfAfO1I9N8r3I+kMIinMNJg/+Yhr3v4xjIteZv6kpmbLXOJilpjWysqMb0DmBkv
LCJGa5lIU/9bsmeyjzNvQlokWoIf2CzPDDbcsZztLiMWlVlCGWaTWId4Vj6bLH2w
ci/DWyPKsbg7aiUZWBokKpwdStdSacUjE5dUmXf86kg8/v4gS0sDupgH739/44YR
GKU7BMj7HE0Pilqj7sLW8EpJepg6MYJQF/tS+NcoHzEobE8+tp8YbvNO6hNlOTzf
53oQeSWbeKZ8y5DEpK21HY+2LxxHAeh5pEq4CJ68hzzAF0GR+T6jqklpLDOaLCSq
ioHgYG5jf4Ok0XdEeisQqDOcqceOgEyb5DCc5qweEv/VKUcCmXNeCgTXluZSByOe
97O35kQYWBGAjjsVACtZdnBaqdDlR6+kow2Hm8o95Y9tT1A37PWjjG98NbCGIdmO
EWbQvMzgZna4PdZ52Mo1hnbYxrFJP7kVdIRnhwxPd9IvwFqbZdWWy0g5Kuw0RouD
DeW3sjdgRzV6S6A5nqrtWwgHeiiszXPo/0ESKs4jFkNhM0/PHXvhQKGVnLRlyLg/
IUIdpjpVKQQysBYEwhmYhkNiqunCrYoIrbNuGSHAiqh1tKo5Frc1R/ATtP56gqlJ
fjIikolfAEvML/fxm91h/336/g7glb+vxSkZ0c/rbYHNlvRtb54o/yWoSRISMLni
WpOmwGLdi/tfDX0ibhA6c0Urw1dPk2VJ9eRIO3xoglwfDi1g+4lXGobmUH/btJqY
BS0o30tFlgcdclifUh7WVbpKFixue1hyZnIdBoJf3CE3ED7NMNOqZM1+eGHB/4wc
ALp7ShVJKSzuN06K8jlVoEiIk/gLd2F+aY25+c9mSkhc4rNeGCMmDBK0NhsXtsGt
lnO/ud7wdNksinHFI2TZL7IwSI3R4b4c6FuF+HMDRDnMJUXj4NbK6d385IAIHNkp
j/d+cwfFO612u2P0frrP6QiHJBB6cwMIOtI9LxiM5tExmYcOkWY4RWS/W7sJBi0x
Iugo2dkpd3qW80ljLzEJLOJcAhZF+mSl9ALM9GglAycfiErr4qxIdVrtTad6jmoX
A+6KNk6032x+u3qyWOooHMU6v9LHKnNhSSNNoBX4c9iYjbn/NgnXGTsNwxZxbqIY
Q2hn+1jhtCtFdo2C1SmdaNMra2QPBs0io7gXh9/ipNMcYKXpAHPPHBlt5eYF6A78
OpeQ6sIOeRNqB7n2HF6eNLInRQMJrjrGGeuCKNO10mxiG432N5bJ71+/sIa5aVRw
gsuXAGGxbjqVP+8BDHN37dVGk/jaSlFZjeloEyWF12D1/WbcdY6NC5Uwzs8cXpK9
g4O6uKalpNt/Wm9VTtmLi+dmL9E8yCah2D/B3L4shLT0FIt/LzbJF+H6GnFUSb9o
Fsvx509RyQkiyMTLhznNECU2E2NmnC72kqDflQAxxQV+p2/wJ+giOhWpjBVofZ++
I39q/OvoGr6pqkBss8n6iO+dmtvc3h0yUqbtH0x18QMzoct9zpiZvYybX6SLWKUp
eWkSdYBAMsm6sp6A712Zv1Xghoe4AbZw9NrkpHwm3iTtUhSNOBlQzSk34w3aOVDf
4MA2D7MhhzzzUx4itfV4XsOKgzn6i647mt4TKh9g/Fz1N4tdOMpoyZ83HqGxFxt3
AInMZiNQmgzzrZkMrkAO4CHCHXBhmofQeyBNYTQ7YSBnVcbaNjC0qPkTjr98InFx
f37C2BookBl9wZ+Q/rPZrpKJlHs33Y1D3gD9b+n/8D0IWh351JDvILvEZ8AzRh+s
tcw0WBW1PI4RupzLzBZbJH7FmL/P9RuRuoJ03oMesDBdlIF0GIjDXSdPQusViwgY
Z3ptWlQyXicHpWUuLo+FrjIydor+PLZZcZ1lRLjHslqIpT7XOCqcnKXL8gTsPpuY
i59Rdvd/x0hXF1zWYY1IWrDxLcZNPc8IheVEBEmANMnltXWkAw7Wk/DoyNssbuXy
ZmIxsYy4Gv0JKHTFjLe7S10Sb5JiBMpd7+AEPzsgZ1BfkTWS03UFgyRhpJ9BDRZ8
XKWXkI30+ixS7Mi9Juqk8eA95BsNHvaDJ87o1KliGDgwD8iQzygr4W6Ml7gySKFd
A9pUTZnmEpXhnfGCNAUQL86N8myC3d5yzMcm+/wPW6Fvqh3tNM4lpuR+5u8ljF/8
S/LG8SwPjWTULhIw8JiqX0lgLlkzvg4Fv+27egCOGkZfPEcJVf8M1LQUTrJnK8MH
cpFQ2h1o/WmDAdAh5LNMq0bP4bbUpinyHKWSau0Y7T5NtSjiX2LcxfJUal413xyv
HXssVYVLfbLt/asGiGZRcb3/ph7FEbmMiR84qrt1i0vRy096U/Tg5M3C3gKgcHRu
z6CYAekZJNrn7LOlRkxYDUX9xiw4kH+OpkjS+rLWoD0LeUzNv4fvEUdEJcsXFQNk
yyUVRQdplAmS/itpENGDq6EP5qxHzlyksDFatJIPc+wwsSTBnQPYrh2xhqhoYgmn
ZeKHnvalweqqRAPZF2jyzlwMgz+dyHWksmPbVRrpVcljEqh+KVQgfLIwJGLxdz/W
kL3SHc9r0y7Onbx+gQ/d1o0NaB1yVp+GOg4FqKX5GLQN3vbJWamaTO8najH7g3tB
m7qssrgpSZtHq3Vh4VN1LarQUseGeuZt8gzqc3W5is2jvqAHMRNafJ862SHYRFRN
ICWO4QKnlj5HOKqSDsO9bbJlokEzzNG320Kk6VqvgRiB4VsHGFZgT9DQxWQFIAgs
HpblT2Adt5NaJv8zFrE6CnT259SELB9WEqGm75pEwrkyTgidWiM07E5ujXGNZBfn
kbRxfzk/ZCky3avAa3PdAYDxvUH+ndukBGBqejNgeGnWQ1S4DwXwvVtLxJi1wyCx
qgk5sS7EQieKjRyT8c6LkJrm1wwE0lsEYgNqSl6FE6+83s9zE49zCPyRpU9fvNXa
y4c70/WvRUjzTXMliZhHMYgPCL7VFdWCcFcuwrdcT8R22j1DBEDkxLu7FhgzUAWV
5F0SoPIYt7l8BFQDnAw1GqHnAxyH0VwIvqOXuMQae+kkQeC8SccDoiOJvfzH7XU9
I9wOMBuVCdfLP3uD8+EzN1kOMYb9Lou/fxJ0cHWYrIcAKg8LtAfgwUlfFXXZkhs1
/6MmjKIqgVtUR/GCXUivdjJKywdZv9T7IrE/QiTpPm08GTIPKzq9606Ii7OfVqHP
/nG90Lu3hP2hKql/VQzWRj84jI6AuSQNfR+F6Ot3iEmYS4ittNvfFmRAPbzOYjDW
thwStpbQsFBiYWXrkSQGyhpuhbZphpSCUctwfjG3SRbOf16ENYDl0ghoDtOQ6MWE
CMNAWQbOWmna0jP7mj81ZE4wFoybf5wbVZC1jjFUnlwz6/LIRXokieUoL92At2+8
6J60tvvmXAkkNNdw1BLT/3MIfVTI2AqbujDy1kOkUA1bDZ+C2AwVDeUW7mkVjhbE
o7Pz+C7fN2mqtsrXQQXvXheuezzQ3oTksevnfI3R1ZMRQqyzwMT565BuRjiEx5eW
ZMFUY+T1xOuP056DDBGQFmxo5qFPv79eh0bwjj/ZvqquY17+jMefkli+NrVOnMUW
4M6yGBxrSxAnX0+9Lxkxg3X4un5rCHNUSwo3KST+x8cycP3irSg//C9cCQU+fsyN
+4qhEBccML5WoCindHzME0ZZFFrG33K0/QHuJ1Z0jdDSUfSfEnLGgSd9k72lI5Hs
FIQtFNaVz0pkf9Xeujzgh826LP5OfcQBvclYMvynad4I0j3Ek0zJj5sVXNWLul0A
FF7cPcs5YZpkFyzCJedQ2XOkndukjTxJMfxhksB/v2k04W4qty7GwjbQnxBiFGNQ
Fbp7qq8J5Uqbe9Wq4B5JMxXZZDEfmr+wjIZXISX3LuXRAPG0oBCi/Iyh2lvOfDPc
c1qlHI1mWcrvnzRl4jNbJbZVL3x2pI+IMcwJ6hO+1ymXz7cnFtjwa9oNMOGxUZ4d
inbX21NjnOYc7PGmb/GXwLobnXZP2uUommlyTI9+y3+Qpx7UPTEAcYC6wPEy0G0h
RhLRv53ig2BUwoSUuhjueqfeZlcfwmWofWPiGhdqOiFK2gRXJIhr+CAiEtTasqkL
J2DIOB/2J0B9n+Z9GjeBgH+34VgtUQfMTh3u6MvvKiJUV6isKs1qyUEy3zgrjvBz
vwGib7quFFxbyNyYNdI2WRyQLK2xMmHZarUTP0RKCMGjWrRC6SiFpZpK+SyFAZP5
YhMURSm+88nkwbRbVNGoN5G2Ah7v3ii7XchViWO1doI5T5ohNjcWhSwlt2TC7/Lw
qnpE46u6ecJ+UUKSvVh5OWz3fV0WvvLcXuSpbyXMCixvnsxnBlo6SNMU3CJGROtW
eVAl1PuYuPOQqCvwjjshrANv0rn7pw170shdzposopPhSEk8fR8FHglYDEfrPHP8
ISwAJdvYjWy5Yh5KXHAOEOeJK0JDvI5D0X4Zo7qCommfIcn1wjwpUX/0SPhJeZlj
O2w6E+TAeauaogqL1B0ghZmubdcrfszmhVdyki9qAj/YRrJNkg6y93LWj+EdrrU5
8XEzvkMtTrfmX05Q6GHN3DAxPy0QSbYPe0XlUndUOt6JyXr2Wv3MNJSAP0iwvx3a
mmuqG8ar9O4Fyuo6jR6c4CzDLGdLs86wy+6T4A6v2cHfLKGab3+kGggA90CjJPHn
nKHq7Wmi2LU9THJ9p5TBQKOVx3M0crQsiaqYoDfXTYLebefAcL0TFUXYmlyFBFGt
E1ijXj7nbnNVxsbEJ7fXKqKFUIJEN4dx7Tlq4qS3iBjjYB8lz0GNsUdXO+6wKaUa
muPqJ0JGGXp9I2Bbi8IVfBNiJkkd1MTytAJpLv/Kb/c+1QE9NjnuOpjsuwfPSZ2z
lw8M+4EB6kCPWGjFFS6f34NCmoytNjrp0lHIPGBnHhuzpZDrR/IGyE3aC8KLwECI
toq1OS0W5ZUg0SdaTFL5vRfc9WUcrSwAqzLBRvkTQTPFfvJVAic22Grm0cFyTFeX
nsn3GfWf/+e5PlUC0m7Ozn4LHxB1d2Rx/LPszYvTPV3SnpC1MkvWmWDe9ESDZ3Mg
xbMjP4tSRVPRMr/jz+uUZUeYbzQbE478+q4JxyKssLL/Shakbi4KE70/YZYb5K+v
5lRLFnYdGipEkPOzfYQ6bH/xdPaasLaguoAFQmKQBP7fcpHjTBTTctCwy0Q4hUG0
qAe2T5UDI1JE2dNozt2GASfaHMOMlRAsLV79DtLFEte9dT0TPm4Fj4YQNaYA25L8
yRgonb4d0bowSV1dagI9a/EOZNWt08S4Gw7ituV9BGaDi0QQF12dfMC8L3deUw18
W3IF8HRzZVbwVzjpukn+gI+patmQLQJ7Q2r/eHdkAlvCkoaaGomlPUc1/t3J4xtY
YRNk+ql2lJGiXyxiI+qVzYn2iMYlEEg+Yqo8E9aUSIX5kANYr7biMAgAJqXwEroq
iKnQWiKu3PeGJ5ZPMnjyvhpeMPynvivmBuBrFfCOwSrJX1/lWjGWARUNOmIcApf/
kyXZGzuXYx2A3bX731bTr7bbRVbRWjPAr/K8K5D+Ru5AeyBfq2gsaGJFxKCcb/rN
H6zLr4xSgYU0alaDB8I51wZPBfIiFBzrleGHcyCkPAqcuh7nVhlgePMDRm5VRNbq
sQq7FjQbw36zGlFbd2VCOi/LuXPZTlKkmlvHreG2nANfCp+ecbEh3QC955UO0XXz
YsR6s1nncJ+viG7qvUz7ymTwZE59J9s9T5YSPeFPRfsxfjNTdoNYrNcY4xyMSi2E
cwIp4Vr5XPak53JzuvrDk0cTNGYa7gfjeS8sZqRFKZAB3wnWaNJfBmE6imB1KESD
UE7fw/S1dDIxKcfGCPnbQyUr/ug8zLiag/EZXAnB/mKVBm5h0kgd9iQc5YGHJb9T
slWiiQvd3FjCzBUs++2E9+YuRjJcmE0sHd9S4bazXrRgJNeRRtIQUdDWk9Tv68tE
bmGUmUVLBFrdBNYhNrN6tNaqW5oNn48Kf1Gvic1E8bWq0qyVRiGkGmaslUXsTwON
W//moWOMzS40x986nyHT5xgbcTNGOEkCOnVGs9jhyAJMI/GFp/MqfHvPTVKxPgFO
NV8TnMYhu3m1FdZI1tGqb/SYEFX5FdDZGURH7AVxpI+t/82PEpzbdRYbsNZSabCe
DfOhSgaOAZDS5Z2bfNS2gGot+Xy/bqbgG9gAx29GSam0PZHkgKsuNrO5VyWyCzUo
Uf3/hzlYheddP9cSxj2GXM2DhLsazlpzOk8bo00bck3E5BApdfr60ujOvHWrGiJa
q2CiKebHIycyA61t7Jp3bvE0a9dIDeOZuSwOedSmFLbk7hRJYLRqvxc0VE3tZqeX
ZsjZVmDFEUaDF2jJL+CvmpHJ8UJyXSY1DLnMhJMFkZvSrjuhKVaL46ibQK/An5Do
TQvhIlU5LDziDSakf4rIA9oVCXlfQBj6BvP1xbJ0VP6zYMxcaqrEk9v357XjIszI
JfkzDjY4pzjZvbWRwK0iQEutIRODDGBkm5Sl8uznS54xsgxjjiEbmsu3u7KiaMaF
2OqJNTlZEiGwN+nk+39obhmd/G+pn0r36sTtNM7mmyHMmQYOROxytMycky2Hd86D
t+SZ7Hx5PRhVpNIN0An7SjpAlz74KiiUv7bIw51EjimjohP9dinUfoL+dtRDjaQ4
rFp6ZXkgLlNhyvvdM/sgU5WyUMOv4tbTJsaLWx7APxShc5LLgHmJKXg37Quq+euG
GPE3Vw5R8HQe7qAHZnjZx6nwdoavBivTTH+NgpRK78Ybdj4luRsZWF3ga/aql3Ag
qCuhksm+gqAwow2tym8QznmIoMtclQEI8pClcjE1gaeeLVJcO1lCJgDucEcuhyzt
WpUxXtwdRFYGP7j4t/XZDCFY9N7EmbtJ2jgkrOxtB0Tj2LhkfkH68nrA07WuTPZi
dJNltD4gLYlc1YSA0WCtJJvpegH1Ue5PIQ1TLw185SZun+uEBeWs6sWl5PL+4y2P
zOR1Cl86GpYYu9QaRkjr4vrLoiDLAfYAxj3MX8D6VvFbA69zOuRCa/vNBgjPjCLF
3ovj0Ts/UotgYQ/w4rhdvRGVujMIDu4N1x46I5QZ54Kz1udD5FWnS+OGVrI6pAMI
L0Acpzq39HjSjddt+XMqBIQI0NS3YfKMtudZ0SLHI9EOECPzvWnBYYAeFxTTQj/S
hSAKjagUgY4l1pAbq4DH58xlkUruuSoekcj98kN4K0HX5Hu/VjwcxrVkT916882P
0ohf0+yvVOTzBCe9aT3pJyrnRe+SpFlJJFuuOukIzU9jlOtek9z1Ewho1PoOn8tA
DV9XUB65hVxNQn+t7P03Q2cRAXlMyF5FYT2S+CKcjy9DsfDAAyarmvvFL86RppQL
XZcrh6+fj/qPyGCYDvtvRgdsyX32zTqbyCjM7bH0NUU65C7IQxUURbSPWNSJRuFE
MBY6IGmwSCMotx/nO+USgfNrpMEOOzmb3Lna4sVXRubi2l2Fd37CDIuOhjOcLmYu
Wkij00GaQ514xbKtBYCad4P1bmkaKDpoO2hNG0UyUI9oKZ/HX0+tehgRXOq1Rrp5
c5d1Uwqpb0jmDWoAf8WkRDT4MbiQFsqdf2y3UgUWrvFfn0YSTFoSI6puboz/Y1Hd
P++/7maV+ZEA8cMIu8GyI33lPQUzm2t0m1J3K5JGQbpm3qmaFTj9g11DBRznIR6A
9hoc0NhOyc9b6tUaBphAJxgAFJnic1hRI/tuuO+pvZnlqLp0jFFAWVgLKIzXAorm
0qxCbLuotQxSxzJ25t11GuoXyNWSpcav9wn5HiTembDl7PkfPPoXpBHpUJEdD+vF
yrCMOElgAyCtvGDQBNNjgSLPqHviNjYkrFKjOgKsGimAzaTEzGzQ0cvU2wrNkVfV
s/2UMnFuASU5FQQ2EBNkXmQQvou1MFtVhuyiONCOzWDcMVq7UBo0cRuK4N+U56UA
+/TMegwiJY/iASpfey937XnAKeD6rPDYXxypEBolffLnc+4BMROhJkSvM6NrZvPn
9ZSwfoJ4LNvf2UmGwWJcsx669teuP6cJ65dPVuFBjxGRiwg2BQcUs0IEIpf6TRg4
bFIepZyI8pWe5A1foRxDo0BmifEbJweLTtWWgst+fsqcp3tcIGPC5G0Gs3v1EWtK
ji3tARp/q9C1v/2vXA3A/RU/DF17v26bw5Dvhd395x0QbadFfqDx2L+rEOyS1OKG
qTXPjBjHq8iaogVDufbb/0/ooAgOZCJ9sCVsfpoyoRs/ffYo1lA20LlRecy7XNzW
DR++T5B2+Rdthz/hze84+1pvNevn9G1LY4qB4dOTQuSI+g1F9QE333HuQx+OTwz9
87ahQO3l4j8MCAw0EUG3zBP2zPH8LrvD0E/cjdo9JcAAYvhnMqCcVJ2RdRsBfds9
u5EHPayvNCEIswEDEycbj0PSMCvoxx3r53wXV0LoQijL40FBLA1HUuUMZRpNqujB
4CDFe4lM+7E4P1o/Kvf8qv+3saV49X7CpgN6k7Xq1JcbFsvX7l+99+bv+X1bHFJU
cT5sn34wAbamHHdKU2WLYLkGppgfrdIqy10Ey9a2sKG1duvlGfU5FAdfKg3XlxRc
3rgPr/kLBJg6Ii2ut64SgaLrKdG89HsJhX67W7a+OMwLju4+do2tz+c7XLO66Xgm
TqcWwB9kzS87NYb9JOejY8feIUdCPkNElq+fdNZItVW7yhYG2WxhqJcBzrDEqykk
uBLBpM6VQCQx4JxCjEh+8lvTDia23kXISHuUMDDPG1+tnZ3fIfMaNnbP76OAsrc7
hET5FWmYQOjeVVIFp+l3LTS61E+r1vKsP16X8NgM2eIXEG4bHIWlzCxfx47PpSif
A6HSWnSyctcvkTM9vkv1Vrnrdo+DwNupgvL2Ln2eHFhI5nJ04Qn8GtiJMIe+sYfk
iCxXnzHXII1gxUHDS1ixhCBHh2NXD6MA4KJNZaWjZxO3yqyiE3kvbcgWAXbiVpGb
jCJvd0rb9T4bsj/LC5bugLPRgHfzveRiJ9ubZbAbKkFJHDT5Nf/DtuD6AhfyZy1D
OL0jEbvLou6PzKLfLUYPBiOG7xQHwVD3w96ZMXJiDjVaOFBp346UvMZxZ6I9RR5m
ROuEvNRv2YsjNj77lsffes/5M81wxutG/glLIAtMB0OnAhafjUP5ZHBnc/oKV1Et
IyX7Z757Lrb7eeGHeGVOtwDuI1IH6xuL9Q/cqbMhvGhbYV6SNpLEm4vJ7BNMlXtu
KTgnkFKvIqM36vH1MnazW5nNT83yJ0Bt34IXh/J9NkpIxOKo9meDjVLS5AizlCXc
EUkECZaC8UHWjuJXJmU4eHtMdiGGw8gg4SwwkA6bh2ehbi/CnCNaCTTjy9gTgrYX
qFzLXV/p3bZ9ESzGqH2OKMGcUIw4QWQfRFhp11xXQJDlqfhfDTtD+PGGrycEPGsk
kbSzeBJWaTJLWa2jwRQgf1Lki/HmYA58NvFyWEA3GBc7G34eTJ8QaW+oRzBUACbX
p1VvdvmKC6OoiG1CJ+qxUedG2jvhMccnzSNLzrI3xZGZTTNn9Pe5AOP+QxZ7B1zs
Ao6SQr0FZbWkgNUsAkH0f7vnEBslWr6W6fjgCYf1VfTK3eYQyfW0Va37shrJKzI3
ab/D+a+qWCN5n5Z40bUpD6N3KGmAy6YJfV9Mnl+s5CAIyfxKLHo2gi00NXin5Q7S
e/8YVD+qezAbRqC4SXfRhCDPGwwm4zP4aVm3X5HW7A4qDIQuR6jFA7fDh1bFYWE8
1j+WsQFQmz6x4CzRB7R7kxVI0mooXerTecR6bIYHVkVb7eq5LOqfWhYbuBgrkA23
vjIrwMxoXxuj+7zBcJWyCSj7Rg1+R4/C0PFysxYBZyhrWh7T7MgSC5MEYbPuHVAN
oIImu8olRc0I37SyTW92YkbQXNiBKrtK51XzjSZ6aTq6p8I4zOLSfrTgnFFBonQ2
Thgpt27PoPmXYSzo4416R7M4AHf53f1mVTp3H9nDkwtk7FQ2YaK8zoOKAeXsK31T
jWhGcTT1Mvnh1M5Q2ao0HMFcMj4S4kFdYHoxxGJeSfCxwy30vhTcHBnXLwJ0LKo8
7dgo1KqohuILD7fK3jx6fZc0WLpcNmzD3BJx5bgnomLMpU6RcPyKHLR+JGYjiwba
VerJasN90ka0SuTAC4KF0k98NM6ZWcLtOT7/zMulVBAROte/LM6WwYAm5igfr12J
NtSM3fkixpeSbAHGI38iDTzIOVtB3WHxZJ9ueWVADKDXOKIb7tM76QL6yzdUCgGD
RSgo8DQIOc2V6AYFSAyloHyBIdjr02QbkS9DqpOUdWnai4ap/oV14c6SdbG0Sa2d
ZDCsnE0dClbTkU7XvFI1izWqWLZoEcTz1UCbnJrq5o+lrsPbxs8OHVDDeK6ZU/Gy
J0f8pb38NVicDyNxjdsHcUsM0+1SpYurnDFwTJhHfOqQBF4EBsguPlEjmhOBQeyl
X7sutWvJdIO3NK444q5kicbBEwqQb8bAwqVbrKu3fD6TDzp/+XDE7lyEp/NoIG9u
RrvxpXwUZ+RKRDEXaKdiaeJZkiZQnnhT5LeJ4vFJ6+suMJQJDNND25/Nux0EjsOa
E47OJunq9ZaTX/ngGgRi2wc2BtHnuVaTYywyjiYQAuCgB++4LFiISkQKJCmwYu8v
JHxwGY6K2Wnpl8DV0FuXzYCcSYOXz60zeiJjY9EmAT0wFMW5y3ZORAhiZppquIY1
Pcy4iEtIS0GJRmUHlU9759uWeXxO5BgkMwr5qjn+AwkA3UCoYm7UnV323+wc4QqI
ITlTWGo9TL5mHv0AqIXeXfQCOLtL1vXyR5su8Jp7KSHg/lREA6hc9wVjlrQUiHR5
/zj64QAc9FM4tebcqmh3E6eTXukAh+goxqieUkj7qss1y0guO1cvKZLn1Z6eZUed
z+zJQ7EZFDNSQy9x18rGdLkwsWTI8m8jdGf+uKiCmqBVspnc8pOad9vze2tVkHkh
iBufV4XcAVe/MmD3H4oXackKifONTBcLiLdWDO22P2SUM9+aKhA6U1wY1ynRODYG
DI3lOREegp6qE+2B9qYHQT+jsQo/uOcl1GLm2eetXE5WSZwmofMyLjkV5fcGgZGd
Fback7Ds8kYU8HMnn/kwM036HR6LqIRV2lYboI214Ckhnd4MLFsgnwLksse9vu4g
zMxjXJ1iJaV/JIUc03Bwu1kkAFz7S50Qi8G1T1N+US0uIxYnZosYes7dGQ9hT/7k
I+1QbvsAG8elVsc8ixqvt3ZGcWgjBArbFi5uUAb6FtTBQRE4hG/EGWlz5AeqJDmL
60vTjl6HLeBBE8aLq0wWJNenTpBeqVWDa1JvJ6W+NJdjxlPpRq5pFM51aa+yz87Y
wc47IrGrF/Pkj060J92cFKWAEr+hNKxsa/klIua1SzzhUTWrG/0lq9C06n2Tx8h7
aeHMeriLtmVUipZp7uIJzIG2N7OQb3i2HjgUDhTaezRMdj1dP4QkH2L3iCpBLg7K
zYLrwXVu2CmqoSAl+u4NWd1Qur39TTrokS3Cqwq7VrJyOulsrdOMxCf7l4J6mAVj
J93I7gnSYM4bA428DJMOgswTSkKPGMCT5tr0/Y68EVz4wPbCUHDhcgHoXOix/vqU
9ndKoX2jF00Zlp7W7PtVBJPQTLJfrQRKkeWQHJhPGWFbgbuj4ZaOgj9w/yqxULs5
btAvF3pPt8XHEoZCovKyBDVCUnRJbig1wT063xL14zhFGs5Wn75ab8tcEAzgIQS+
2rAyFjdPkkMVy4Rf5TZmoZ8sZMB1Vl7aoaSLywVT6mpoE/soyPV9fR/RfVGfVSnz
h3nv3Cmloyaf6BjsECgqCdDYCn62Lb7tlFQXFTbw2P0JpQU21u/EH7v2/IDsT2EJ
hCAD9BazvVVCEEynUImK7tXkvPsinT0XdEEZs66fo7YUM+gumv4Q05ClVMGzfHRA
/a17LgHa9dRzZL6e5Ryi7bWJF+ET64blnFWwnGFUcbm0lk8oNZBK4vHqZvw1d6Pu
ZfCoSElVVuf6yqdGQGt4UTq3CvwI5Hx2G6zltJAFAkgkVKFPrKLpRJMeEgtsEhVF
kqQWJhV4xaa28bWG1OA+s4uS09UIvQJRKBpvYPjEMN9ucGSlkJ/9yj1X1zXfHIzp
SgkiEBLa61mRJYfoPXrefKGJJj+hBawWitAW09nPCNU5Tw63pbxcCupDgKXix+ni
+WCmdKXzS8uCZjS5RA/Zy+l1ERu46bjjArz6x061HuAayPHDuWz9wL+SuzTTvZdf
obvCfO5gUHJ3noNHa1QLgKBX9nO8N8O4GGG54sYCvpkP2YkS8Pkt1W78/gWRCVOn
It81M9wAeO1Wpcn/onrCOdQP70LfVFZxP/xo4mQlknn173bS244HCNzTdyN0MLA+
cAY8HXTaTNqpZc5zNjT1JOe2WeO05ROfD/8f/jJgsO5CbF1NN59uNWLtc6eQIxsV
Q0HH49+8JCenHW1d3e4+8bZ5qGXtshuNBmq92NgTXQUcPxEJsAipR5pTuTZHUEyB
UCANR/ejf55SvKFYRbdWvrtp4IE39NbkVXa8vpyo2IhPcaKK9nylInq3C++V5TTY
oahjCc6z1dWNscbN1BCEb+OsBtp1OaF0A6baCdUoksh+l70IUpElmWaDTBGwH1t9
rCAtTX1zA8ZPeE9Q9mjgEVIxSUJo9iK+TWWfRD5Pi02tF6QlLauWm6PvD0S5X5he
Lvq6GEUVromNsVitUIZBAEaFsmyRb4QiRf91290fqN+DZ5FS5QGXWj4rcW/GxzN7
+MqIDivTFcW43fd+r9oQgKtRsQR97PHYhyUNbwYvFJMqFoo/J8ZgwOU7vPOJxhlh
wTJkZnZu7DTGFRUPJX7yTWja3KrVWRBpr99SnKsIDZMt3j8dPq4rx3WX5MRl7R+y
86ZtV6/RYfH9vpSgVMu8CbsIqfgpzn1ajNtaECvubXS5hYjHigWxlaMPr0MYML9d
Uglu6u5KYl2WK6gGBWig20VOhee/X2sauTLSX+r2E7XlfbX+8hJVN1f2nxdafwaQ
YohkXBcq5iR1CcP7XRm23XUn9YN0KTx6gd5lBHfVrz/wJqgH1biNUTT6aA38wUWZ
iVwNnK+fF3tQ3RLPkYRkp53O2/xOrV6+eoDLRt1H0Fj6wBlhaTpY6z1AX8fGARJn
VVFgDqGPByhwztGA+wMDgwsw5fPBZ7GQOT003Jws9c6zI31sVkY+ZwyukmN0hKO1
l9YTkDT4MbeInlDGjuR6RrQInqrVWRMaKPG506Xc8d8zRgyVQsFLR1G74QABVTkP
A9lsovBN/PbPNzUv7lSUhV+H5ZqMPGW4B7DqkqVx/IojUQ01XXw6ccqZOvo5egHY
Uzg9lzGOa6YtXveNG/5jKVmpWCC+03UbTa5Eg+2PRgCUZbx4guYxKyDELng1U+fi
25fT+IFNREyswgWxOLHCFjrDVb7igSj5RADI9p6OJk43ApG4hOls1f6GxhCdhAPC
Vq6wSopZirdwDjfQ/1Yu536g2z+FzgTD2Uv/to9ufQ0kIxl7OVzbMNfUBFGXJ512
q8fk43zRgq8IAQ8btBLV+ofpevjMZ8b3kJj6U7+D8OYgBQuScDEY00ByoyIiq8lu
tXSewgr7+3H51qnwmqIVaBXqEvmbdEid2hccgU15NYquPdT2zqd5cOjiB85fp+Yk
9ScfcSeTt1pqDXJvyk0Cu7ZUAdexyAAAwmcsc2YxSfiaDmToTnHwle+IDwm2G80H
UEb8JS9BhwzVLpsGzFaFwnRuGt1lk65fHdIhSE6ZtAMiqBfEKiYPBR6fdmW5N62Z
iIE1dshRsE8QOAEroPbIln88r2IjG6ojTLjiv7iLUpC2ps5Eg40R8nHZJ9oLZjug
39LWJCNx/PNXVXscLllFtgBc+FIK0cx8tly7i6ExrrPezp//htEstHMivq4i6zFZ
BoFFGsMM+aUGqWf9x/cTGIGI9QpNytkqLRcWRi4kZdEQ+2zfDGxrAQsuCuym4Ewa
k+FqZNQIgSmj+8KjnW1RcbPAoQkiwAamCvS88Jl7avVr14XMUvOhzJB+IG3C7UcA
nfWFP4b+dJSifin+jujomoU5x6pL4lc3hl1IaWhotAKiQiV58YbaHQXbqeGazaNU
PS/bE4T40q8o6nKxTRegAOtyKPy/LUnehj2Gp9kUo+fWiz6++FUbXRMavxEBtoAn
NlVpVmmQHYPwaVTziB7NSdlz+ZJVDFtjJBJuB5xCHmZ19HMsizrzoHnbG0stoJgK
Ri97gPxR1VGY7Cg9oF68GX/cc9IRa7Y6j5ZmIRlzHeBMkHQl8D2Tc75AyN3ZlNIz
gLaR/aMsmzSLiribQhJdv/wi7VRfl1CKaKcVbA4h3ZDL+zZ1wz1KJ0fnYQkoBwJO
7+JflFfhUB9Uf8A2hEsvZ/RMCLs1fG2tYUVl7KrzoBsIy3FUub6WGaXMTpsVig8u
p6Sh6lSFAewadnDdIVqlCdet2tRY0qWS5HgOU1fbiC+KgKwkEy2B0G8Y3sWbrUAK
03zHUfK9r+HJmm+DjKt0PC10jeVPwMQp8+nmY70iHegRjTv6rl6WXA5ETcNojFlj
yY3QuPh7/tLOSwkmsi55Bke18sl/6nCtNkUO6r72UoXoNF/dZyMublZ2KsWsHVlV
BytXIDKhp90IQ9h5+E0HTL7qI8viyKcu3VbwgUbLdbKyjn44hQXathDQH2IUVtSY
+/Bdo5Ft5zlERsUNZTfIwv0PJ2KSAeT5oKFy9FaVtB74EUKe9Q75LBWL99hGKJvh
fMoQQ9eUv46HNM5C+8y5s2D+hr7mw9SLP2Qj0QE5AOrN1lP2KHOsV/osxXCsKE/X
1W6Wih+eAbaqUqDahY9EHZ8wjrldBfVKs3KP+ofgJ/LUkZEiu6vZ4SvA4hRw8ahT
HdWS1h3cZPYpv7HL5Xavr+2Mt+wolOgPShTayt78DlY77PP+h1JvN9ZGaaaPn2qq
Ai/euhOrVuLceZBnjnuFPEHWC7lZD4lnsi+5lxTpSJz390nqpmmSAH5h1k33wlji
/Nh/E3I1rEIR+Fz1lcvRfrlaKKR+eOT9P10FUsTriMJd4+/bXRMr9hJwj1JsbyzD
wUZSQxBEv7F27HA6yqY9qCrBrchicGsie6vT2Bd0bpCweYQfoci7ZBiboP1RZd7y
EfKRupSXOf08TzjDpgh8kGhqZZonmedNQUH/YfxQZ3b9pqOKewvSogcJhycknylH
h/vcl/4hEAI4zwWAOroAh3TboCAxUVZHe/TkInDDlOr14GMCXqq9fgL5WQmsOxUC
NDDSNcrFoza/XcJT+vCCvhFazE9Qn39LnaSi8fBuNyZCSSdWIft90psU3xKvk9Us
9Y81NXsvn6piT7rRyE1wrC6rj3037ECpVrDCu2HWqPZnMtI7rT1YcJype9pDRcwH
Ra2DuMANntFC4/zjeUo7/ufJbtyG4OATQsaMokZ4Fnaa/r45N4CuA1+uWExvhwGs
82mr1urXSTedK7QC9Goo8i9eyh3rolvaHtkJc6HBG26RB5lnZzHxDM0tX6tnDWx0
E5mMrdvhHtVOlxiIN6Sgz2lixgD6uFo5bgF++1hczzTPe74eFeYksAnzgjvKvhyK
30Odg1v/tb4nfemRh1hH2RKP3z2X3B0Z/kDYU3ANSe/6lErXYZ3LQoWQbTr/Yikx
asFxXteVkgacmP2zTwcEWaTi/sZHTq5XNMwJm9eSpth874GUT2LnWZcSNUq4LRGQ
t94V8V8kpSiWvimAQK8AthRkfLniT5oENQKBLKRtn3+sheXCUuddA04VRK7WuyyP
2zRST1vP/ZWSy9nNfUdp9bVJVFf5mS1SEdZ6BbiFYa5FZP1c9Tr1GfO5ODkfDO77
pbL987x25vat6HQI6xwLZqK9sTQB3CvCPVvC/9O8PexPrVVEjP1/Gr20EaOTboxz
qVM8Y7Di3QdpNiH/n6CPUPJbJ761wHuQHY2dvPS5xrKMDSe9GOrKsQI7Pkyzy7hY
bHJIdVcupOZngYtYWZaiVEF8DMuZGa89Uw18/LZ4CwrW/97AloFh52c7PTh6Pc9C
CpGZQOcPjxDQ6Ae152ktmoAGlAcDeawelG1MlsUCu9PQSdnvN8OxiAcnkAebEkQJ
8NK2j1VCz0ZIeAPFIi/nD4U3vvto511TXijdHCMm69ga9Cgpr0tHmKn0HmLm0K1x
jb5BOzS7xDi6haXGYJGbl+sXf8EZwDbAV0HOt5GQYb8qGt7P58wyFDYqt8cF+32y
3PRjPUQUhkQrFgUsCwyNVKftdrwXxMCFaNQKOr7H+Bz48cJyyxHTe2q6kj8fijxw
FNWrrPrDkM4nd9pOQG5co0TXguBYGfPnWoYFBY230LPGjD9M4+Qrzpumd8O1VzIS
vELxcCZUr+GeljGocFY7UnYWFIdipwA3N/vH84GHl9z2eGv2fUyeTZDcTvyMc6BH
ZIJDJ4T3ZSu5nuvhoYYBwBnqXiCibYKITX0QBeAdseJ6PHBrl598JN+BReHCK35o
40mj/Ukue5wLk9HtPkVCzmWORH9EF0z4IKqSDTwyRPxmneE/ypDOoVxZlpplgY++
vi20tPUPjf0OfwOPdTeaLquit3GpmyaeOlLI49L8mCZYHCXRJgzqwsk4ztKVCsqv
qQBgejWl43uNYl1kCbOpFN1nvH5PB5nMx5WbYTmrtQFqA1kz43aXkJ6JRkwjNiSf
9hLfpfnjsMtjqB/lxNT/Hjf79hPlVFe69GMIRjwBwiBpf5JS5BZsOEnMqtjL+DH1
0aE/qyWgC30UTWI+H1G6tudmYZnnSE7BaU4+1PzBgC7Aid6hjAeb2uaf8YUhrkSt
PiWTZd56rCD7vDn86UwVqwbuEgSM5tnwO9fe+DxdSp93K5u9rQ/Ww+kkLuM8dXe1
cTaaAiwVuGg2AzVE7P/+FK0HvBfMdtv7ULVtE0yc5Wy4E45IVPcF87JyVMEW7bI8
TWkS3Sh6Fse6PQObCgCCo84J77ATllmYAJkai2mvqHL7jRQQ3EmND+bo7NrUuuvI
AWsGL41HS54kuXkHG+ti+6ke/hJgyDoZPIO3bXdNvmkKv1n1cg5vcLEtiMombKQs
rYtUg64aoClo8KMUoF/9JPGssTxpOf7CeoG/enPBYR9vK5aEVbQh3e2amV8soDft
HGWa4vxdoWCSbWwQgfbBAtA/q5eIWIBl+6eHvlrqC6Nd6hujp1Mzg6RIu97qqQF0
lQ8OiTFAEB+FRfNDW8ChI8o8Cn0m1NPn+GcRKCkc/AUyp3wMKfbRjfKadnvFIxh+
ZUzF81SZbOSjnaL54LB1VlpOV5K30g3IG7GInw8wcsUtAb/FbJZax7BoZQpc2que
D7KEDje72SYcMpzeoORmTqPp+1pP3BCPTncQBYAdIR7l1rI6mlW2MjVkdT9OlMq8
l+nutW2HCREiY/e+NBsXuThhA4goAOebm2ixyn9nfFzeTfrDq6WL6E4cuZDIqc9B
Y87BXIHrEMB0n+ut08Lr24Mi2+wts/OrXYwBeOPgKCb5u9qkjpW/T1ht9/j1zR4F
t5zVsoXzjw0mySvVEju7xWBriFtqgzXHKaZ4zUdTsznxs2FVWHVDXQFycflhL9y4
zefK0hPRorrbtlRzeNmFPqe/tnukZb2EMFrQcT3DgPWwEWGLca8m3yA+F7tQX6a0
tRDag/Dy9VFH3BgBQ/fAnPk2Eqk3Dd25EMTEN8IN3FZfS0mk6a8s7nufJC0TktX6
MiAXch3zueA2q3y9euhcMzft6igmq2XuW6SeQJLbBahE1q1fxjbJV5KRno5ff/As
U11RxC2LpQ5Ga7rLbSjzn1Ckqx1tOCfab2ECBpxwnAWN6726Cth6b9gsNXA8thn/
OQ+M66Ndysc69cVmLQB3XBuSlCzEE0fEin9Bn/KrpdBC8Owuc614h+w6apc3i5qy
WM3bLI8L/hEJRpdMNgJMZ2qdnUuCShib8/Nap8CaF5qDFNWvJv3PNWpcyB9db587
AXgZ4YhoZg1TLvOJGOq+nn/nMoP59cR/uMC5LS6n0mAdYutj+Ks5apWgxfjsDTVE
L8ZhOi53eE+3h8FO2D4wPZ43fRfSSE8eq8+kTW2VYj7frT83ctfKDeZA3oN9shlZ
Z+ER0pLJv/wjJyXIqrwDwKn/+9LC7mgYh4CzSakxxVlQYAJ1CBVYkoZYW9tOmiC1
dPyXg06ha5Jzkaw/TWX7KyFxSRNql1vN/NaKSe1R4yAoReYHTaWQepurIDsq/34I
9oI+sG6BDDMhewK32LRrmaeh+iGhzyq287s/OioO5ccZlPyxLzehcw+tQaEnRKl/
Lev8Ek3uJhzmfldmOsa9gZAPGwYGEmnhFjGBI94F7NymLuXl4E/3G1uTKgIMx1Iw
9BHTobXvErfx9PHnQBwXvlUQFKB8sgKtT9qZbpXIJ5UQL1CfqX+zzZG2p/kzgyBy
dXZiL8SJjhz2lJGtjJQZxUJtgU3cTvI1nCFIckMnnlDVdm2wwQ95MosN0EKvl662
p9MCgDyYw4hqdFdb9uw+Y3exaVtDsOgyMlrI1xQ3x+CWXAWzc3Ixy/82RywB2UH4
1xxJeWzE3kM1hsI6aPloJUyCUE1FtKXIIdUIh8OZYZ5OubbfMJOvQaj6VY+dLvXw
ZUS5jgkah3ZQKrdZF1D6wFErOcvMHKC7t7zccRGz/bcwBiQuN2we5y9fy+qIReHC
G66Ksr5H0bhpPUucWN4Iyajcb4C9XQyt90MKCSOG43OgjMRPS78An/9a06aKCBr7
xPwsxsi997ZrMC9Si9t2dAIWkkTzkYZIw2A4b3h8KZxtefdN19qgveK1tCqG3Zy8
G1TkIhi3+wXI2TthdV9yT+EFdhDM654iDP/zVPyLI4d1HdaWyzqVysweFs5b+TQM
4uoDDezyaKNAjFSHSkfadN8+d/H3bhQGv5up017IDJ35a4eg8MzTcNDkXN0Tdm2n
oa8+6ShAcHAxmsRdw2HduD0QSYNkySmvSlQoYZtRPSxFLktaGkeJaUUtuTxvP4kk
W5dHBnrFbIDtf1CMSsS5HB1Jj/fboAJF5psslGNgJ1tRfhBm7YcbmSbjuUmdb3qw
MwsOS6QOaXjIeIQDpDCPlBdYZRAdsRsvdUGwMLkaIzrokF8bpn5h9loig/n8s2LH
Hid+bckwRHRZTpscgZvAFOsG6pZmwDZELrdROOhwbyUbYJTktvP8Lt976BGR999N
3kRexCIQpAOvcYTgRXzpPXm72wWLfZL3ABZ2ojL4DUgHaLGqhy2rczTL7CZIvXL2
Ce4oK4Tp8mcDG3ekvyLvlADuZkj02xFMiJa9ETQHxhx0ZRlBMSx4y1FDwxYN6jQ4
u9VV1skcMhjQvgP2aFNb9aa/TC5hgnXiX71o4Pb0Ikb2H3aFxy2rLnH7ce0QvCP5
s8Ng2tulFPwkgk3SMEuQP/b9K+FD2TPrLQE5ZBe0Wec4aUtIixS0wX/SncgoR14a
3ljjCo/xo3R6Epk70bjv/WMoeXBNt9aD63HzMS3TtH7Hm7j2mlU2Mnr4C5i+oAQL
iLRthh+tnIKJ3u5mt6dNIS7d2bd2HoUCD/pHvd7zCgfsINe6jTCmAC29Hxc91+fs
gRXJYzSF7JuFyd4hE8ot25+tlEO9SNQiLsMhnkGfyP+fXJmNPToT+7FO73qjIFGm
ASUxkZNEXjJ2Kc++ifNK33kz8LxWBWq0IUdrVs9LPCEG7EBv3dZWvXFTquxXMk7r
RPvXtD/VnVuEZdcEOWNSyfkoTCgfYeWzofRy9etH7FtvAUB7Br3KqoEJLKA/oJMU
92BI0DosQAGM5qFpZRkltPfmkX4VxToVYLlpOGmMII0sIg9s4Aruv/K3tNdhra0N
+yT3Zj1iIrcubTULCKi6SBkVhjNHHSECvEdSqzQoM33jj6+UVGnrIl2Do8wmuIEp
l6U9VunBfaAgquwlvDgAC4rLB1bhRQ+sLrogTiX3K3QyFN7dS5iAGL9qgUFwDE3v
yPenaTxEhDgArmw3N1IRbJKBFPs1XuclvZKBzph2EevXIVwsUPWT/8bSnNWUBOBR
L+mSTdtcpv9781otAnchuGmbVLVPH9PB4sFGj2yoSAYbV48K56x8cOLAqaIdL5Sj
8X+yF7nTsgDlb0wEenf1gqMwplwT36J9o1qVDaJOtzmG1E70Rgt6JlU93o+wJXmj
KLNf81fSs5XGd4U8dw72+0wldMTilbPk/dsQ/j+xfDX0V3YzlmeoDaIgZeqir0P/
2CSZXauIZ7FYylSOFvA1ATVPBz5N6vKBc4OwhHXT2sMWEaCcjZBv2IXwlD4Ylzo+
r6y6f4zo78pvmEJm/9qBP0AFdTpZaOLSDHMg2NUKcU1YIvJLypTcl/sjWwqaOEB1
+rhV6sTGRT6mMjfdWKbxzDLXvyFw5mLZ60KcRA8bACNXqqva35CtOrK78IFVbi37
NhmndtgldwR9ATT02HbhYn+NEpukRMwEatI44VrZLVRuxSN9fC25B82FeQQmuIKf
DEQo1ZJH1H7WSTgPQfhBML45iCPbZD5oxS9EEAzzBvBc9mxl/zcjGVsWKhPE+1B8
OWqwCqYXYTNoQdud//jnNttWILEcY24Ss3IOIPJT+hhqM7bpM9pq+SvddUtOV4J1
dAf7TKu57wC7Rg4saFVgIg0VFm84je5Zcx2bgMASgVLgzxUOLYDAO1hhiDhYR6KL
fBTkZy4SpbhEFqx3M8bZVHV34HhX9qdBwiDxNBQd/mS0Ehx52NYx7zmjnst1tbNh
Sg7O9GPhZ0ZSVraeFC9i0kXtMAeqsU4jFL21IzQgjSc4YYFxiP8gYQfEAa/2sXPu
jQ/3htPteaKL8q8GVIagRhZa8ys6un2OjHOM7syC3eKuZ/b5TGVJcsRQPK/pdQdy
IBhNznQmMwlnTZP+zg4nHoXCXj2V3lG3g2VhazEuBnaUuM5d2VJDOWDjl7KMkcz+
scVNMRX76XjNu3tocKX80Kxsfdtu2e597pV0ZfRkw478CVhZv6prfXaCEFL7tOpL
YG7HIpaJ0f6O5udyix8VdOmZBI6500GdnYUqfr0Bdrs+5sWMsZ0pGn+z5mEPi1tY
CSU1VIk5VSJERJIhQEele3Gm0UimMmW0/Ax4dU54t71K26nIhNdfz6TBwtEk6ZQK
qul81VQYAQjdMZVC2CGmfyp+pgcsHApPyhfZkm6H5U0cyPv3pBbqKjASxqY9kpTW
Zy341muI1NQRZQGJChH624daZioZ3w9VGF3pRj8/GEcxcieELuZRUl9vxjVjOpoX
VCS1mWgBzIMF7RPgpjBSHjFmo7QMpXdZdF8CP0fQwx/NOJB8DmCokkLZSiqYjRSx
NtIFy7v2m2TSj1JCgyQJyy/Adk3O3SIwIDCpo9HHjeiN4PuTWx0yki7LGgKVxK5Z
9+6KmfFRxVd5XjUYSYDIeKdCAY8e11dsn8g+KRnVi2ntJ/n/znRkXN6omUJS4vmq
S0p0iY+rnhalM+Q1G9wMw2Dmf+6pqvWco3U/HPIlqAfLRNtne3xC8BI79BunDNH2
AEAWK8fmc3sQFeujl+X1PhblaWaaG6FcRbo7WvRhOD1rLn0DsZBHVJTPP3zYBZQR
olC1mSz42w5O92YgpT3HJhW6ExibuZACaS4gSKxAwFRDBqsYD7wKIdfBrZ257zxM
hayimZ7OFSVxsAAhzzUtjBRrmXZEpFpQqttVk8EwuTohvAhcBVKr6H+KlGQ4JSKa
oEG+NmOcNjTqRjM9Yi1dfSb4FHKFPk9KKTsZVb8q2GYfT7BylsSc5yODzdac/YA/
Ep9tqNN2ap+kQcVGCLPT3jRvZyLrtbYChjyf1nqvt1E7sM0lodqxAdBaa5vOhvFH
QKvq9ifu+NErXMclsOtUBcX2WZKDbS9nKLHYTokcP/eQkL0Nguoln729vtLYOZL4
ednnFykqb5hnEdA1HI6aZyI2Wutl219SxGP94Gr/SzQyulBzHJqdU4n/Oxj7kSZ8
PaIQFAaa80D67jHtyr5GXaMKBj90QvFzNQHhKBIzEWDiNVFZOJWXXYxYAsV2mW6h
9BGpsUDCs0gJ8OAH5inHQnd33yET42OdCpNxWzYaGv/IQ+SvvACXOTnOZJly5iey
6P2IRuGkX/2YuW+XweSBvaXsJ28Z07i+kWGvGOiHuTm4EixgW7KemlBhW4UZ/dUO
F53tAtJ5FqVbgcUPbBRXQr5fxolZOu5jDc8JV+nQVep2lLxzJSQmpTZtM38sUWEl
ouEkNM81XQBnrZ2u67cm7j/UsL4RlE7MIdqSHoxokx2sNwdRYxSeVDy7+xsQQNrJ
Bi/bzRYYEdtzLHlmjxRqkQOuDdOPs/W9wVhOBLXIeycoVSpO04kR6SR/oGvTYucb
IUb4gl4b7D+3CjU+i/bWJk13Y4FRI2+duPJTkAk4f7nZbzS2WV/ftUrxsbKlAe9g
BvqIQALgoMQxq2KFUFTNIKrWPb6OeLjI1f94uCgxBxgkSfOthwoylYQc7363Q297
9Jp9TomKrAsCkKxYGNHWQKuRdaejHtFxh7mvvCVgMHHTYRnCJYA4Jr9XdMJzCjZL
ApWsjEER5L670SEEVdY+K6mFsLaxsw4NIg3QIfIW7qZr8/aL57JYQHHKnqxQrrma
Xk64Yt8FHPsJbuteFqiJdhWC7rmeYzl5WWMT0XVqr2/YkME4A3ZcwYPYwzkiXGFd
vF44r5zElr+g6pPsMt3caY2viRxQeddqXAekRmI6TYztijq2FmTaas4yqqs80J7e
+nlX7Jm7FPtqemjZSBQOSgEwSPWXbKINdeobQpvk1FV274p1r9QIfZbW/U29pckS
hMdMe8i6hnUQOLk5F0QNMOjY+Gqv1UvxrrsmdPR+yfVUqSHt37tjbwwpdLDWHUft
f3SB7QxBUqHHCDfcUqlr3rgNfsGuC8sqNp/jph8if05/VdtlqngV6iqvcYtTpcj2
PLN6mpTwRED4xfeTEivygJ/nuJ7mdfscDfn6RAt8ocWPaiHGtuTj2kgcczMV4QVw
hp0XmxFNGLhzDzAsR6vKRKBLcU5bVOQby4co/FXxt4jgfm5v+Hs2hFpeYJLZnbdn
OzlGzffmbGK1N0HK2prs4RpD9eFwp/BJtTOvMpdz89TeYM9JU3+J20vN48p+MvLM
LACOnRS6Nh9oyu0Ih4+A/LQ8Qq8ZXD8Fy2TdIiMMoxdatt+jUlFUTColEeOkYqsg
rHF68ARscUUtWx1+Ts1g4xoSZS1Ke2wlWWctKnwyy9tE+EcQicU03MoHwunFR5X0
K876csAm01n0GsoA7Zymz/oz25OyoP57/dvGuCIK7EXP5XhDfwz/D0tYEute8CeL
NP+9X+g46VuuoSBbLBlDQWD3dDa6LyVyUHxeDh3TZzewTcswMCIbbqx6mkejYmB0
Ih4oxmNsK5lofE4mFSO7N0yElzjfJIPcpFUs//gESvMLf4nDcsyrhthw32KSSz1Q
5URQnBfKxijw2Vvvbv+/iAKOYV0XYw6fMKquRzs2NsXo5K9JsGSO4wL38/UEky7q
OavII9WDXxfiGf38XxQfWXw+GpmExtf/2F2aow5lTX3AQPsi5t6SepK2vwbw0kzI
Rhsh2oLoycKyGUtfHDbLmagyUC7uDpYwbcQqE3OIpmlKvjvRSDpw5N+Yw7pw+H7l
rwr3kryRyvRDQcnCSH3jVwLuUBGEWXFVBzrRDAl5U8kHuxa07DisHyvTwn/7Fq2c
L1zkVKu6FqZynNLzSxe3+L6G6EAlrKjKXfyYeQHsaEMlAG9BNGeAigZYPozh6e72
IQi4grAeYwFVUz/yL87RgVdVu2OH47gpDqF42YQ4kw+XGmH+9J24Ey6qfP6PFDhn
mRj0KtjwF7BgLyIOjfZvLq1HV9823/jKq66VZ0TwYzVwyua5UGlmUYEoYndcZaLg
/J/5Zq/xay5krKa4cUw9k6yfINdtpJcsj2if8NQNqjtemERnlNs9lNI7Zw4EcDYd
NRu7zXJt4OhcJ+WsHqDiBhDJ3OKMdRNPba+aQGZYtO4EIfHRBEKvgg4Qwx2r17mE
GJ0WKEw3D2/6e1I5JNNbKYrpbIWXVXiSa0BkAjEBdJxocEUG7/X170zbMBGvt6vW
dpo0oUxVqlturj7ucggI82/sEtI4he+Z5amyqyhhznk6gN2EroIOqvRqht5Le/ck
Wr8+s2qencgONQchzmLaK06yEghPhPp5fAlB3aZU0E8NoUxp/E1+zoHiI2RjB7mC
4eILx/1oBAbQ7lhRY6kjSkizRz8kjwPFaTYQlf1C1+xb792x3ihqGNxJ2ByqR2Lw
KHeI8WUvoJlAkpNwes03yPLUHKUx8zAq/sFVr34EJfk187Xz2walq0sXB972/oyi
vDvzftVuEqrzsAg9LhIWIUXivFS1zRRKG2FmUR2K9jgEUPSL0lLnkK5FlU/ZXkKn
zwNfHMqKkT7c6pYQ/NIdIdk4nFAvMrgifuuCHuu2NBnwCHWjWTtUrUHShd9cXBfi
HjWUu+wXeNyOvF8fwplJbDI9I1MRVDa+tGPVe1fFRTY7N3JDkZNt4tvps/l+PTmB
ZdWsbMNd6uvC1UAb579bSDDP1f2UeuKhz5VAlFYBWcPJagjbg7KJEJ45UwKstjbW
QumxCEhFJbBfvWh1ESUw77OGmGP1AGn3pE7l8VJYtvnqHtOPmRpyWxsRZZYKzax2
yMyqwdkiL51koNB2eGZ8WqqTVjY7JQ2l71YUV0IEO2wvBk7pFtUi4ZnkebVQ7W7n
JM6a7EXM1XGPKIG244ha52whgR2nz12wfiIdh6zzevz4RaWZ4KBmfCk7DwyjVQx9
5+P6dlv/S6eStTTJd8Go2BKWET1hB/5O3XDoOIbg5JEDqV2byULsa3PxtOXGapBO
x2cb94jWCBhpuDBIHGFSvd0Lu+ehNNo4rjsRmGl/TtizOuiY8/m2x8lXAyxldyXj
zhsLbyvLsRDYgjImj2EaP1o3J6kUdB4/JUp8e/MfdftSyJbs2IuLs9MY1MShqzgF
xG/cVyM3YDcWtz3SVLSY9eYlVujpLhNW/oSKih9fpmZpQzRHHv7rcsMknFSAWDf7
X/VTOHHaJTG/+7wFwhaOnlBLxb7Nk+FUKh9T32qM+qByuz5KPLtu/mUVLQEwFjLE
0p/zVmaFlMCiAKdrn9pEHgg8j0xJEyBDs/3bxqS/FUXbirJhGid+13TWRnVkEPDC
yxTDDihYPMXAAouCBlulXf/xeId6LwudSOf7m59yLeo4TE276Ui+mgGFi6MkuSH0
l86bZUsMoAwgOZO1Jnqo6QGTzIfbenvSx7W8Qeh76cpNgPT04cFBQ6g2V6H4YDAB
8qdMC5ziSvIQNty8hK+/c6XG8KsaNUs9C4lh93786aqJ8+hEaFbxrJgIF6qA68Va
0XIFmwyPLkCa3ZonRHA09eWj/c9FATqc9QIFmMmhYB4B+JQPaQUj5uiFnR7yXUGU
8rZxdZPfzytB4urNNg/ybLPWzy4laEpjrkUr0tPiyN5GBkx53N9h0cCKN0PwQU72
pAEzQy6oQum5wgSqqUlR26sQCK2JsrdFQv7iJmVbD0juR7x5V2yQCTIv2fPYaBbN
R06ouTnPFnicKvp+mBSsO0yJezVYFlIglkq52U8zxCCf/SoreMOtrLf7+oWUYpQ1
9Wp2EvCTTbHVA+0XIr+X56px/16d4ljenfXbfSTOj2H50Sfaaz9QQisR/YsJn79Z
t4Ni9/ubL3IDtdyhkL7B/8+o/H9/gwwD1gDoj3KZUn3UkHGVd6Dh2LwOQhpOolJN
poYHQdx/tK5vmugUpng+TknQIMCZJVBS7IDWPN0Sc6/Y6D+padrau6q1q0+FRvf1
2ksC+PFniuDlwQkV1nRat2pIB/Ep5ILho9wm9qhnAomNBa5l2g5+cGF8qLfxSxLu
YxKDZ6pGg607giZweOYnfm+7StI+4R6/bGAPEBCTHnxFzAkYSRNKI5mzITXb3+pS
GGWf2C2ALLJfhHLqGWYbp7PJp06tRdqbjJsk/xxQyER1jjyQnqyb0JilGM1YUulD
29hINUSc2G5kNdUfhF8wGC8u7rS2uADZKbYsg9VP8XRWLzTqUga63E97uK/BWlbh
q0Ydmqzw9nhfKtQKBp9ijglsuEf0tQP6JKN0VmZbdEKWQq/2i+Bxorh/VffMGiUg
Rn2ygaGv3cWdzBX7iX1pNG5jQK0FGrshdX0bjL+iJdglaYZiH6RpBVrHs8za8qHo
e7kjL+P7Xjd2CN6toWQCuQndpcXtoOTP2Gdhr0Gj15BtB1QL6EnFtgWXe4WM1VXH
EhAmK4+MGLRoB0oL6lg33j8pz0X9xahJ0Y2jRBf1phjYm0WbkCE68goZCXAgO/yr
T+hIa+jJPElw4zB7YY+7DcgLZHdtpnFhQdLWUxOFb9pwHsvMdCrKgbO6ajdYc7cl
9K2rsBMK+GBX+zRJT0kpSJcbF4c0JrVyAyVTDothINkXaAF0JVBV+dby0R7ZS/4y
4jRF+2VVWNpDOSSbBNpRITd82BoNjrVW7nZof4PECpZBuM8k0aUPKTaY+5F8RSqA
Rcli+ZLnsA7QuYqV5PPJbtch5FrsH+BxfSf5YUtfUr+5ZF9VHmW2Mjt3pxxpH8qm
jHJDvepgTe3UQ45e3I4OceGLFmUroi9O0wPvtXQVWlSX2aBFzbZ7vsQQS72Zytt3
aYcs3s9VziFQx8x6S8WmfBwcgDkknmlQ4PqcoEZrhjiX1Oxdme8cGmqRXInPRAv/
xNW+Tv3mII+w0EL1XdPD2OsbAnlIQe4RhvZQ2qi40MVUFMjruuCOqGInYQsjtRd4
4SpHayCLxqI/SWJwuOdxXFhNyZmGdGy2xdAbJ740NLJUdwXShJxv8vdxyRXx8/Uf
p4EonwCU7/7Tq66D3z8IGtYTJTzzy5yKqAzGULMpUFHyVkkov9ymJrJvAyqffzgX
x8Uv4LaTWXxJtgpRuWdq1u/qJE6iKP8egtGOIwPjwFvOHWpfG8UFwacSOeL+zbZ+
XJDqU1bXFw+yRfZsRAekkU3Ypsc0cvPXlKDivXvn9DCfitpMS5uKlfk/xK9HC1uW
0BglmHy8KuZ96uqhSwAz7ApivMyVsI+9H7vCl9S4PMIRgFa39T1BhzmX2Wu2pmzN
pWrVAW3kBpCjbm6DO4yqVyEZ3lZvj5PohS34tfGGo0JMnd+bIbbtqZPXgGDcCqyA
iEEb/idVwNDNAY/fNzLN1DoKyyw1kTVw4SF83stVpgtGcoyioEVIjHfAPAHRTOFv
uJ1HfIxBowu0RP3J/Q9uCTBMenrLmL6wpqXeQY0MUE2M1Phmhq2iIs551GsR0xCw
EXfEsN02W1S30EPLwuWbpu0bD3q6XI/wxwkv/F5Yn7XT9ZkRjsomcat7cqMXuRsh
V/EKhwSsvDGU4+Wngo2JC+3WfPeHpkQuIPo31TjKoLMHmXp716p4Vd3vdQvQdZln
DnaVRiDg1KJfo2qSORFcZUXadGH/fAmjW5mFqtshX9oUWLhBHRpWXe4THRVZNm4k
zNMlbe5YT2jhL3+bJN5pVtIu3mYe3ct7yOZTloLhwPihRDOSQcSogEhoQm8Id3pT
4HFzIdsjMXdvPywpGD8SLx9NdRg0XuH+trakDzwkZIlpRs7XkCjYNByMuTMQpkSv
lom4SCm8fD8RM0nSboHGE+dD3I8eyX+1MwG4siWwwQA5n7d5wihu8nIhdajaCFI6
1piTtbp77mdraSnmsmeU2phtwK+IyU1rZWx15Gud4u6j2Nw7jADJUsqU2xVwjuCW
UDTk0zI5cImz+ZSOYoEbJSt0tl5b6dZo2nZouMBwxiBNJBJxJyjL9RPUrML/Y14H
OJkOgp2Qyz2Db6X0G4Z5ZlMCEMciMVvu7++IDF4MPoznyjbUWDnV1thYLNwdk2iq
B41LNkatYUiGS3VPpTSMGuVJOghleAO7At3KpUUxaB3kKuHIgL2A4pZoCTeFPrjW
x6/4TKBmsYWqETNH0OSH/DLJg118QXPI8w5zDlx3QqNa+Yw5gYMjeCvnY6jTgo/3
iQ6P7xQCDZIxady81vOq/aa9wgYrZP5FLiTVGCjvg8oPdmF1z3UfD1n0IL2FLqpg
4n+coUhKz5ohXg+VX1dLDUi3cWUZJUVPZuDVJyGey0ZoZlgcOuqWR+F4o3hkIIAk
4/XXJ/0LZuO/pQoDuIZLbpVG09hEiwWVbin+DsJNr/zMH2G8Ggd50FjmJi86tFxP
n1PmAC70W5Ju+YvI7/iB0K2SKgmSOafZjbj8CWHfbCEEDax/5l3hIEmMZoxCEUpF
XQ052xy1ZV664fYHmBsxhseU6hhDyPSaqy+L/6uR8z0nDhyICnd9gTybAo6iqDG4
EXrFpPeuWVj7EgZnRybzBcqti3R0ITc9Q2TYvPmqKIdf83zAgPsmPC0QA8V2lRot
UzXssS04OJDTdMHUe9LQTnD6Vv5n1Zt9sNAIdixxpGp/CaRW2ftwCeGOVAs+KC6X
2ho+mGfLFDQuBKGTlPAxieDMP684sru1rqpP1UGNqRZ2ZWFo81VnsxpUaX3T5e1/
rBn05JQ9FyoT4sh0X7wbglouZetIZUEK7poKkDNSbK3vG5iYr/AXvOwiZxzovsbo
PZh01iDfwnzYdwVZ6RA27GV6k0ptt3Ck99JhxPhfplgxMfwpyO2/PhlRwgUQ7Svu
t+ARHeT6ZjGQVTVZDy+ts0OXIWp2oyPTnVJCQ1unrN34r60UmN5y7jh5OWufLKS+
KtC2n4KUXyZGlRjOExKr5Ha533vST5F+Gmx5TL+koIzwO5J2zXPERVXomiQcIupK
5WUig+UiV3Gxm9wURzxUoZNGqiS+TEFFBPWrtaY7WSAsGHf580Z/vLW6cQ54Ps6r
Maguy1fQzvUVpA+UILbCEj6Dg3UJWL2cZXSonX1PAKEru4845CEGPE3Q+FGpXzsd
9PFmS2pIi7+2gshH/YjDVWqy5FrkCZzTNoXt2p4ZOEBbM61YhAetCcVP8qzV6Hdh
lbxKL2GzZgBQLrRIVr+892lU8pqQpwOws6j9/tktvPd/36KdDbL1WcNShSU2qQQC
gYSA+Gy1H944Z48So6iMC1dRIl3a/GZZ2rzbdXKdWmtAnK9GwSC4PHMBnGCw+G6+
+XrJCa9hoWgY5y78yXoMk2SXDnaWba1PzdNy6jq+746lgg9ldSJRsdXNoEb7gzCD
pfBtzXcfC3rX8DHH5zA8yqNetTRAlys6qPRI1+a0MG3NH9daAb45LBZsaUzSPl8l
tkfOS+L9sPQ8f7sDrZu7GwsXiubGiyfItdOWHtMrjPedrNJtyW75/23AHA9DSFTa
d6/T81Bui0kP9MpScXLDQ+pcRdhAbgvuOJPC5wp56I9+Y6QRQKrGUPArTCb7GH98
Qoe7CpnKsZr+BSEBDrT83gOL/Tuo3eVCErG9VDqyR84H5VgfKHKM6KVh6VNaBaHQ
RYEnDKmuBdy9VZVUMUQaaRkanX8MdQQo7mYwabSAKeLVMIqpTmuoHVUUL/hNWa8j
Lfl8Mq8AqiqOEJJn6BM9sWe1yJHlLOP/83YcTWR0WNNzWfhZ+JZ4iQm8yiSRUHW2
ZojZVc4pX8glTJByU9dGW8jSsITF1Fe+iehx9iea1tHZl5TwpWgBTkvA7K3VHYrU
4XNNj0Sm9+3n7n0FoV04FmHiMQS4bJu/6d1PCbPIE8WLveE66J4Y8PuaIkNdUPJa
KTZRjeS6Oy/aF4HZiaGs80pnvmms4PSLiT3w0LFGL97hkG43BE8pfkonMyN8nKe9
K56Q9qxK4H6/NZMkUNmZbPIMxF4cUkRkofUHnXdYpxs9MYU14/ftGXCKRAOGOje3
rlQRxLIFzY06/wvD/pACwxsMzuPd6QOqgb04UXvuurz/zlYjJyMrWm/Ja6Zkd6M8
eEwXVuzMqlx9dO3YkcC56lbC/jyracAeWPhRdizIg0apyLC3hRkCUwwPMTA8wAoL
XDaQmHoFarfHEjsHfa1NDlLBhzTIDKa9evEuau1il3t/HZz/bB2EAtHoIskVkqD3
gqWw8J5u+7qi7ATKzoHxpx3Xwrt0Wt7kzqkKv+/8vEWsBNUzxxtTZQYDOjoui/gu
2tUnsVAwkcxfrqq/nGDyBVs583VoL4ZKmPSKlJYYeS21pkg/6e/+2+12/bSH6VFa
qqf8479p9gJQOBzXzVKLFsjUXTQbjlOanDbE17giTh4bnlvLbLzJg51O9ApQueyq
VaMIghvJoZM0PTJAUZvlml1H3as9EFWTQibhEy7tTyBkJlVuVxI110IYETsTw0aR
DEAQvsZEm5n9W4Et/9LNU7VKXcXx1IrYYCd0aOe8kyXP++ZsgExe9gvWgm9HjitX
kiJZD3K3A50Pe5/dX6MZ/quT3fDjnP8aJf0bCUwZajGNeuf4kaCLj+hWbuNKN4i4
dF9RYWxSTN2TZPKMprK1z9y7ZZMn6WtfunrauDeYkcjY+5Bjte1+pontSuOUHFlL
4dPRGNHDS5Yuf78uz73kPYa8doUQCnG/A3jmMX612ahSGiLmnq2fB5CdohJJOoxp
xFO2uEHvqH6A1G0jfSO/1eDvSTlPGnVtqopXedlCCU5hQw6p+ePD5p1yQ+2wXt+J
6+i49Jdf/OL7cEzUjoB+WpPFsRzfLdSHpS8X/tJN/o38hOeo1FMAuiqDYnL7fi6L
U1812vICpOpt+52YiqJaQvnh+fcZj07v0AzTPGXZOGgt/fm9tpu4Lu4Y9RdFDpEh
i99dVAVWdaDD8J21jZukGSbFD9aXQWz5S50i8mpOUV7Xj8CPhuNJ4JG9O6ROFZoX
CaHGFHESJ179nmhUaNCuKq66fgtV/EpNX+l6A8uVIAcMIMs/tR7kz2IRLzrWc4PU
g3CKOfFN82TxDQ8VPuI10v4TzsMRgkjrsND/Mf1kdJNWZStkK7QmFvKIr1E1EjU0
gyLFu5SZhJEIOz7AnS/+Ktivwfzv+DvDhznVVVkzXVGUQOamqRPvoHHI1L70l4Uz
OpCSdOtmCuuFRq4UoK0ndOUup7d6Z5Fnb1yfOecGqsVKXyUz8YerOTeU4osI6cKi
JfKMjKznmhNoXogs9OhRWRCIFlN0rMCLTJU8dce6Mqcib6Y8rref3oQmZy4agSbQ
RAb6K8+WV+aqPE7uNnn5XMN20sUoDWra4z1sQLgVaFLI2Z/BGwseF6O+/EZE7Viu
52pXwuHY8tfZ5lL1gRNJ1iTFK1ZDkQYZ1hNFwX1E/P8zcs3GEj5XEQKxi/3zNfU7
UIzyIeD4LjNSRVXpnp/yDufBEGH4Cb9BTmTkTUu/ZvE1uGvldSdhcnKkDF1OpbHm
aGZXyUQZ0WPNul0iX+YC4HhNvUBn1Q4UsoDQtZ7NnnC2TxMayfXG9WuVfCElHeVP
USiaYMZi9UkXsHQiOl9EVB7wcwiYCnyr+G6EdOKYjMh++72PcrHHo7HEVjLLg/U3
VfVAZGZn28jvFXY/U9FJl3CaSxL3vdn7lYyHzJ9mjdHBthv9oqdLNrFLC8aKxQKz
kuicMvJ7uYnvtqitiq2DaTWN1AtVE+ufQ9VuX0NerWvzpNJVE83H3iLO22cPm4Gh
yTDx355Tq01eTTETkeAC4EZM4nuNKk11gAkvzX6KpZU6AlQgDjtbEgv6tcocCMnZ
C3klHW3jXPE2YWnZRKyYeDCFROZ3xOoZbsYTmuQsJDIQtVG9+/LVV10cIqlrBE2d
HdAJtpfZVqr68u7800HtYeS934dOmL+ig+NVLN/Y90lYTnZ7Pe7noGRbpv7Q4sa9
Q5YzISGrMmBdzCEO1HQ/z4hbc8KbfHL486PfsRACc6g0MaaiP0Jqr3wr0LpTioTb
h4gFKp/FcjRocVXGqfy2qzv/I6KBaO5IDDml7XETB9LWvs2u/XvJ5FDmN/27M5Tq
7AQCv/7DWN4k6DPyScYk+KL1q7oUZVzNdY1ee+eRnv6Kq8Ke49manw20GjKHri7s
X8j20keR1Wuq02TDVKCwl87AK8Tx2EQtszIPx6qko+QbTVFn6F7zlcmdmeqVTaLf
ovTsahg15lWao/92RZYf8BSp9pAPuQN9PQAoGQ+X9ALms9ttbMowqs0IZ5/kSu/Z
BPeupf7xpaSbajxnpXUKRc1xTXW0Iw1KCZ39bG4V5nHlVrG3/KKCg2GyenE9LnSF
rmiUeFju5ZFQcKItWbodGxnQSvfLMjFrnn1BRycYOyAqnKlQ28JHcLyvr2Nt5bIB
8tgDHfAj1SOkQj7sZ7TUuAtxSs4vGv0eZak7lQb7r+2hDl753a32mOisACQTg2vw
cyKJTWgTB9avV3ZQ86HissEIFWuzI0WYq2fndwRkCwvUjDc6xm4nzWlAr5By51GO
x6yCNEr7vxCcy/wJ6wFbeOgNAI3Vz9opHzH7Eaj6PKBYN99FDIhuCm68gq++YoMi
FLu+rP2AhTlGk7OTXqAXjaU7YlwfTuNqdHRVrGEZwxVzJEhQi8yA0rGUrehoH6/T
JcO6JaGUvcHbGgur+1iW8Mlu3XJEImIk16nHnEmMKAxvYvpFW6naAids9AeKBl8w
VH9cfVUobhn6LAtZUr4zhPbSpB1VzOW2mkCff58AQOrHaIQPYUSRXzBorvJW17z0
0CI+vayGxpxen8yX1ywo+BcyJSxa1yFOyr4WWbp+G5cyLb2pnSpkCd2ky6eSVsL8
CvX12k2k5z266bDTQTXk1DvDPeE4W5WNYBwJk8d6LrKJfZEnjFgXmltF8Tf0Qqc+
U5mf9jBRK8rdzut/8Z2rad5frAV0OIcZtCah/p5S/IUomuGOWw/C6VIbnzmhaY4s
EmFb+uIYlhMabdoJysSE0Guv89qEG01KzCFzY4Cvg0YQKXgldEXXWzvKYsrd23qR
+DXxtgKoriqxY1DMe+TD2QGDabwnMqcVpIfM1RUonNqH/oxyB0leFUudd2xk8d8c
MzHILg5TxD3N1hfc2b7gVEYYVuLoN4UNmjcd5Cz1MnKSwl0/RLl0JJCprqBiCMN6
J6yz6ClvLz2B/2yMn2tfmp1p7GYz66fY10Avv5vrR/fUrD1QdHz6nqdkWYtFffZf
2THMijKFDa1K3MRgBow+BnfEyVOAy94Y5lDes39jxiAWPhMBlsvSOmZCMtGHhoDh
s0PIQpnL4yvc91yf/jbKyKI+yGXPy7JlSbvXW6OCdO3dU/F9iiBqGH8ncpShwbCo
60B22X2fB/alXPrWITR4R+Z5mA02EdzVZMNdOTbxnhZNORkgaGW6j6USCMi0TGch
4XU7RdPFeWFwGW/UQPAvRfzHPvxUQGSyVjdqJOg36vuctHbYtGBuIdvFMCk7XCbs
RVbFwtNHzD24PDX2zwLCYQdo8lIE5ZUlZT6M7UcO6ptSAH4uhC3mL6EnwV6bHqdz
JnW0YepO++mAFy8RPFhUIvcVopqoZ/+h+7Y2+xzfJEx7KI9rlb4RMkL4qqLwJwv6
Z8PvVVMM+cT27lnRg9ocW6AeLSi6LgTZawh8uxYxleKQYy25QXQNh5o+s7v692kT
3GiGotMwKLB9RHIlFMOze3FXqu06T0mHMRzkxJUuKF2kjhA+khvOd1aNRAclaxOR
3fWVEAFeL8Bh6lVf/CVFlAZO1iJi8ah1eSgJk5rO1zL24UP8k+E0Aom6RVhAJX23
IxKdwbAbEreg255I7VEOt98ti679MjTvCOY/kGP/VNLTQ4qHd5j/7pouGoP8oEu1
a8uBXdTZi53pSm9bR74UkHgD7SrLuUKkoWHvOXguLJBHvoS+6jFRwPEDymOH3AuA
HLQpH7qr92Obd5x1d1dYJjNE8D1Ec3yFqFVGa8EG9VnICtjoTWiNxzdtDUChzbpG
txXZBIVnqZxaYU9nhOqpMaeq4SJCEfB37S3gSmoXPQJaiZsFxk+21MJ1tbqc7l8G
g1GGfhYOItAbzf5mY9FTdyZg6kIXpR9aViGv/bhVvLkLuCtnAN12xiRJFR9WPm89
7ys45Y93h/KQ6KpGfYxuTFv6FsTyfqe1cFyN6Q7CA68oqNAkIUjVZ6hvTCWvJd4J
YYqHWKVovSGd2t3i1xXiJvn2WM9A/lIAo5OjCoI9unqAp4g0gRYJojV7HHOdZxco
N0LSrXMlpeuqSNe7jS66ZzQPn0LzVE8ZmqcqUpio54eoWOXZW7MlU8gPO/FExJ4v
cCQkcKV6iR2FPLHiUIkuWusGapyxNj/0OSTAzBoKgSyfd6mhD1LiyJzxiaM/P4mX
fItVBZ8tGmmtVm8PHBwfviwgyezAd0UoiPM3t+GkK0kwKGkj2xNTf0JjQ5btOQTq
rltpkPx3X+LkC3gifwq2k0a5biHwYAs86bIEeFHYTHionMzbra/ZTIO/w9/xJ4HF
CJKRXcL5O61beedoucYn/Icc+P0+OE10D5Brt+tVtCsgi7QDFlLw/BEZyEM+BnKW
amj06rVTytMO4PZTIpBQNZj4IjYYCXcIpTdlvjlJEDUdRiVrT1ucrpCPMpmy2wIv
jYNFbzyjVLnm31HmQG1EkDJPw14f/RfghUSOnvQumzPoVCA0XIxe8V9bT8VztP2b
e6qMuj++hPWJkZg9Z1q1SHoSUloew/A68hgFSHdaMO6nsNftb4vtRuu5DV37ROso
4Oz+z4pCaS7QMdNZsxnpuvG9o32ARYxgB22JJ9t0Gn1WZtieZoa26K8P+Ab0HOgQ
1yOLAkONOp8/ZIsFZGPizXMvzW7wokt3takoVS7pjbA8cgBEDD3fn1YHSuRdbxjl
IxW+TtQSoM1QX8Gry3DtghX6+K5MhBFvVGsboMoYYA6LXlzeeytniaAKXQ9QaIci
HnNqvzsZizoeaYMJpCnDE0IVQEbHMIEIwyoIWQJoWmvdOon2Xoqp2jZZUyzwikFe
Mw7in35DEMYGbLJsiouC8f3nFg44x5CES9R6kiwc9R0Hh3et/vc4Pv7M2PyRHDdN
RewsqER2PgUwdDdURuLoZafTU/QzLwq91nMK7Aiybj+wsJIR2+GohEKTW13tP+5R
E0EyNWn99EnxJ+y+s6IUAw9wB8JsZ7roBYQZqy8bOoxmOV9lyDZW57xuGOQYMQIs
YW9RIWnNuetzOWT9lEysq58zvD3m1Y3NPQnZCPiJ7f7r5/QnOiS1c0r9iW01qS3a
DIlq724/s1zF3WkKGlNqFP8chyxemTvmfqgMY9VEID/udb4k70mVWtD1n8KynYyV
TFZex4yyoD9K0W6PMXnfwev5qb3g85whd1D3hwU7IvMZD14n7RO7EY9+G1FZds5s
czk5qZxK2rwBfaDJDqJGwgwbRUarKBMdJRcvwY0OwhGuAQoyRd/z0fDdu+sPbs4Z
HV9HthSaAQMMMHfxD48KzV4FFa48iWBi6wbBw/qyBkXYYM0UjUn75Fvb/m9vtJM5
TYZloHffgYdh4cQWInvRys4iUd4RC/T6SZfIJUyurN75oLCkTVdZsRolNfgQQhwd
tsB1ry7/gaK6gnKLTWbzC59E59vdGMhUvc4zhapOzThEjXG5aKVkx+nb7a1fpbgT
xS7aHAxEH4LScHitMWuz+zxVemXw1FWY+JlAJD1TS+kKrvTsv9oL0DJO2L7iW+5d
UdBTqtASJP5NGigQRmNxbsDIpc49u8d5+ErScbPs6q/3OLg7LS8qj1KKki4GZUfY
1vmx5paF7AI6xLp8L7qmIBvTfKCvVTcTQwmggHuoATbOaUsinQM7Jb5drJ+S8Rkc
1ItUpsHm9wSI9sJY+e2GM1f6QB6+s6RFlUTGvIHkODxxKk0D3y/fC3b57TX8klAV
M8Z53RrUzGl8YiSTRcQpld2wvunpvwUyXDhn8ucizs5iga9BpKwMZMwET/e6Zz4m
6Vdmpoa+DGDWtL1dZ4iSdGqUGCWRDUZkXygk+ayexL8nnZIRcwilMe2uzM7KpmMD
/aoW9UPNPv5zzhEJNcd5/uOF+zk6YLPFIzw7Ujbdp2OcqM84viB8bF202suJY8zv
2XxbEEmadn3cenn9MG7JxKY1wi/pQlV3Y08hsYSBcHGAGrcIVbBn4sXMTtYiDQ00
POXIX/jOtc0kaEU/I+bJ8pegblwCOFbWsv+VPWSEkUwa0AufBDhXbFqd2Q/lT90w
XxrBiJWly0MAKgEjAFg2p/txeTHkM9xlXEN9O/VFGu1JmkSy+AFOAabklzxvTaIR
6f3hBZewyGUv76EM/Wi3QRZzdKCyEY0tY2NvbOagLYP9h03Exfp0w+EhsVkxub6g
URE42RBJP786seEyQa7bG6mMW2BLzlN/TROMHtEUMtTAXAInfhPHqmkON3HrJxQ2
SwpKBvBae3/XdJXXhIqP/HrvZYWTDCjWB2DsYqIvMBFLA5Gteul1SfwQjafQ85Xf
tQSDse/uOm/8cLdkQWmbt97jWAXbbZO6cfiMvgg9r+3DbkxC5PWKtz8U+4pOXOVx
lV4SH9/NsA1qNkX9sXxTAapcIqmaqrkeO6p01Ow2jdblcKmPASCx1547NEibbDRu
WKxCIO7ZiKr1NQVnuR0wj3ILogR8KJbAVzZLFSu17A6N2hlyJYmnO0Ya5vsjCvci
G1YThv0WwIVxAqwrlfPFhG0HrE9Wmlq3xyyvBFaSAfh0LdtIXGDJHcfFFjEqPDqu
N694g2o7wxdEsq4r/HRuyEkAnTiMqkHw8ZD20fwauVJioOeF235gddlmWOl2J+wD
BX5/NJt/ixK0ZyBByZoZ9vG9H3Uz/Ctujq07ubxHk7N0teZkG31gQueIACQhyUWb
AQS7aiAOt2JNI2eBK5Nhn30BmWttfXdMe9SyHr/ReJY8TwzmMQt0ELnawNSUYLAv
Bg1hb+CrZi9xXKUgORvsEJKAi5e3h1SfXyqcmIMdCNfmzVCzEsMs7aJtIVLI6Q8D
3drUR1KGJUTA/bU9KeDhRRKIH5TxSHZ+++iOZ6LosO9bJT+hvnnatDJbehwb2G1C
PFzpS3SWlW5Bbjl/vefW2shIWD7dR99In6LwPr9OZaud60W/XtZCR2eWQfxXif++
ZJRUJZldrc1ikCjqh7ua+BMKZe974A7xafhQBsV8xCqa/Ids9J3Unk5OAGrnrP6t
YF92YJQJjmcOvxynW7FUcc4/CsuHHzyCAZrfKzfLtyEkAxb9y6VBxwaAAxCdAm2t
xB4JDaplx5fh+/viiFqhxBcmxJtdIx0ANjDg1bOv4ax9IkvsA+dDRM8rC/yTvXEM
/6xF3E7TqAkF3sUsw10GoByH+218AD7lOE/Av6WaT69ER1CCmzEYvT+cXo0NYh7V
n/M3m0b9Jlbd9pN0Hv7OE8Wqp+oV6sRew6JKqBh2/mBoNKREeaN9Jnk74SkCIYRh
GxfxdKZHR9uyWZv531t0wzTZTi3uo90nbnbjvo3bVlrCtUvnl0Ppa++YmQsYVR4t
u0kMlYfiKvdbvBVHmTgmU8pXQISyXVwallrZj/MEwV1QdLWa53+pLRQNQVSkzVww
rhp/3/iTDhNt9Vv+aXYWj+XJFnnlr/6S6N850aL4WsuC9E0l5yKcOqCMNF9eZ7aU
PSSpR1OGhK3tkpQBBpNfrixkar2ePV0eilvAZafmx5Iv9+Im8Ih9nWnzyXYWYL1N
LrMVU/AIpKCySiK2nduE0UqtjjcwcHixamgprvmr7z7GhNY7GVgfWNwuZm/qOsL9
kxBD68TvXiy4bFPAOzd2EOxTetE5p6b8iU5G8LNqE29sglus8m45KiNsu6Qj0GNZ
XVKsEfNby+D4Se517bpW2aPBEGPe4mHZst/TqFkkT/1PWKmwDS4AonQm8Ry6bsbp
KMbo3lxtoejzdamrr95cF7YCbDkD8pYqC6AUKIUtLxHlyGp5W0PpWl+h7nF8Fw/m
mCSRhf9epXkxiBNMrv5VysDX92wkrNxJ4BvNlsTZw5Yt4ezcd8ZY5wR7Rufhp/TZ
uFxKe3lppqG+j8+EUcyLeCp3ObBWTIdGaH6fWzMIK8D9lqX6b4SBG/d0/pjlk6xY
ah2JtKa7Au4iIGLgbb5ke0igsFupuzlkeGcUSkqO6/Q/tilZb/Re2BeDcXddu77s
YkKYsDZpGa3hpIbGcZS/XtdvtLH9ggrF62QdL42P5fulusgpFCCQiT65/5IstiOU
BUeAvsfUUmNuxL6fgj6Rx67GV/OjBNGgCf1rS5MQLfECTo+bzbXbT+K/CxRod343
fpArkTiknKCA3PQ7VR6L53EfrLV/2BgnDi87cnoYIx90avl3b1RaTPpUpGs8aqZM
kfcY03zjmDbLGA/dwKaZjGTOPN0lsohYqXYsr9tFKq8q2MO6cpqPi8Bl/mpwbpoC
8bda28kaDEb/QKhfzLfETg+EAL/Caip95LWADAfIteLUoT9mofrXafKWh7YF9DEV
PWVwADQ7SDl2zCe81eXv3pUiwxmwB4RSL21LC3OCFbOqCIoatSStPH6vqX95UvBA
kN92loAQYolEXg6EwVJDy/BxOQDpvyS0P4t3dpHPoh4SeDwJ3JZvnK6Y7npRnk5l
YzqSpewkZBw1DTQ/cB6ajjwT+5NzK0HhxI/WZdGdvmrS8eZqkwJOjL4D4ioZIQkF
NzVd11pFfIUSKZN1NaPN3bmbrvrl++LLA2GBKBwow+fmO2ZHBzlpUeQtXw/ZTWfK
dWYXgrp38+v/zRWmdi7soxhoRSh1ALTphyDCgIjJCMJwbhOxJVv92RlyY3slj7hg
9p3IcrUctNA1QdCLAFUIR37L0Nu5SsmGmH2obDFqavHH2xjSXeb0PW0Af/eBjN6z
zQY8xOUFq6iq8JClD2gb1LhVucZAYgYzBqfXd+P9Cxqp6aYJ+jCTPWSXWSJMp6Mj
omF92D1STs5dt7KiKbIf9LiDGAZFjohOiXiABIzyZNVKkRWqNZpjKMMjZJ411XN4
JUHx7bk7x9poJOrEEUatndJfHfgr5QdWbPoEQEfngQfW/jT1Nu6DmVoARvqJWJLk
etF64G8y5Z1qcbLcooa4+zMV6IK74aaR56cDjVZSUtk3fj/Mkskjx2dgQ296/Ggq
p+TlKYBRiNIIkLYcaAOJQvEA3MG9bwbR6zWKXkVejmsjM6KSCktl8Ga3efYs/ic7
/eBb8b03ToTb5Y2xpWzo7z5ZGGytmajPd5hUtsaFvifL84zXpu68A1GM8h+o/cNt
herFTAS1/Ydsraguw0FTo+6ICIyvsZElBh8qnrONIDAywTMyMfISlpNN8zou/McE
p5vK1FyV9Et5DaPaEfk4lcv/wL9L/oqhPWRE4WmGcDi2QhU820xxGaocgKAfCOCD
7WYeAvJhs+woIfHgT1tbHuYDz2Wz4fh9HBujXADm4+F0kqHDvB0iOQ7Ra88ORIfw
q6Umb6KhipdpO0Nt3F0tKqniKYzXF70cj9XzRITS5slkdFHuO9mZ+GWcA/x8Fq9F
gS87SQ4bcQTZUu/DIE/aD3F7XO2DAhQQsVgI5OwOojssvL3b3dVrk/qmnBIkmQ26
0KHBjIxp+VTdU49fCd+1MMkBckfEF5x2a+6o/It1Dk6xmS5ee58bSAxCwWOx4esz
p14fFXqfP7aPbC0C2DbBVrfg7A4oKpNOB0yTD0B3HATgOEsQr/J+NiXbjP2RRpPu
Bv4oS4SLm6xA+UfQJ4g49s6rqmgMh9XERXn7mjerAcnasSTkaaoB7tzbrxLEeOvD
mGolZwFJU0b56vbuHo0NbG8qv1jPikX6Ev1Uhl/vYutX9Qfr3QBudV//ZDUd1q6M
q7rknyV7+haYa8zyOOGgWi4G90UAbGrYW196qWBTKfNQhNiHS6PyzIsrMcxbp+xZ
eegwgAHxdciOo1IZm+HscyOck7oe5iMZDgJ56hssPd7IcMGkk2wJlVTkZWY44mtM
XZGF7V1/VGHgFmO80X3GPs+Qtp0R2BULntCWID4EDbzDvONlTsRLt6r4UWauWV+f
82KrVGANHlpJwNPdbCk8Syg5I97tpNt4w+9OaU45HhVpk+VXi/+DpsWBfF88Ol7i
8nBA8x2bHiBKYbzJBrsXv1AIFxoQ7H1V4zKLNaoKngORmvMzBOKGvfpt0DocIXo0
jnePwV6V3jhnONCjxwV3GSqBTMFAZ2xa5WwsSD+Iz0jJbsiLpGv//LRgeVePcPuW
gC2w7XXgnKn9097LH1uSU5BhLtlTVOSLpzr5tiQTEAGfpMpMwBJricVzhG7rwU7s
dBzWJ1XeEqkIsIVaMIzhv4+w895cEvn/wRP17gHCvkHnf/7MnQyHdScOglNBlK/Q
laI0PxT3hTmZK8OUSFmINeMjLaTtq4NtorLessQHmj7qZe6ZDF7hBxZ5P8uh82Wp
cHCHFhhoWy7HKJ4KsFPz1ars6BIsX+qpD8RXdVDNx96ElF/xBZdgUyzS6p8q5SKv
/AVB+00o0QDa6JJFez93VNJYlGpcj+1t2m2mfjc4JpiP8YvsNosLWaY79nboRjvG
rPtv7ODwj1NSsbYjlEHCSnE8JR9Wpo5+n2ZX+Qi4H+BT1tS99d2FYZjkRF40glPX
xkwarLJyPGP+U7tR+HHj2kgJYUdndMP4gO3kDJoRKwDmS4WWBsm5YeVIW9ykGXCB
+na7N9sBSNUkFXXrygvCLauva1iUVGJRi7NCr0K5vPAVHvMu4pC/rBekFs8ofVXo
XSmZfrP3sVNh2ITIbDFDqG7brLor4hnU/WB/XAIhppwF87fIq9MPL7vEG1c2+4T6
klgtI+Hx2a3KeDS7kIlIfVHD/Jhjw5Iwt6NFFMNIU/UV4olivJdc2n7Mhd73OO/U
GI/DHAHqd8iDhFg0/RjiUEXAcq/MiUTNWjyf/p3ZTxGql2posRv4ahXJ5lDqXXLD
jYBQQrZ6F3SQNm5gIQvOFWpOw2v7Q8ZB3lXcIAWlq3aZmnQMYltKXiSqkSCz/QKy
YBf6PLiy8MCwhRKlLvdNRqVkXGF9Z0qWELTdv5+dXjPtI35qwMrHKlFqCwYSzU4s
E6mQeoaSBy0lXUVcCf8MFdBI40qSLJM0BlmKzaQXyBHtIdUZsiOTGbKkgXlT9cxs
2wJVXQ2gAL08nuR5sRq2w7mttnDZ46c4LpzYLzm2Pv0jMmRgrKRZeJntCLs0TrJc
KcdjUO9t3M3kJWS0REsVf+6rBC74o79yzTXsM4+A49EUklsbDp84kN748/gFMUej
jlAC9BR+FNy9StsHdF5raJfzxn5+DVGTeZfbj4KEnosTqXrG6m6FlWwmsRvDWckP
JhNQPrdwFnkEz2PWsDsEP1k7gcCkkJxYSW/mDY5uDSHsxlxXAQJqhHJbglVrOg4i
Tzl5YMSt58k2bezQjmiLa/etCAY1y+f5Bgy/EyHrP1bglhVXj4QXDI0+HAuyQkPf
SzjIu6AGPuGfp7vHq1lEYB9Gd5ctU+VjIRQN4KOQsF/Q4VQlJVsjveTzFNaKpmrR
Y5M9iHHM2JwFulClD2bxUmZEndONetLoYA9qhmA/57CD7JSSuvMea/Qhad4CeOJV
G62WvE8Oz/r0JGH/c/+m74d5cD+lWbHxpiMhMoxRgJl0jwhNbWGMLEq7+QhzsKtq
/Dt5tlmfp/huKFsnUwE+p6ryZXOHZVHb0JH6scv8VR/6v14cXeAQqq23pcZJrTNz
uOaHzO4NAyRgG952RUEveb/4T3COZhAOg3SdgmF/kqwGuRTy6z+IGdRCQyPfJ7JJ
9uEJZ+rZIyMzIgDlnoMk/RbAcnSmod9ijNEjhm8KJ6FkIIyDC0ncMWvuLLC16wGP
Q5o3iV268HKnHeUTOmObFSluDH/b9nro4bskTlZ+xUXJgJqyhzFKQazBrJbWd6QL
237lFAZOUSvArRM99asdFTfT5FMUhiFsrLka3A18YA/fCH9qfj8vkoh8+9SRVTQo
D3GBuOdTTNQCQxJhTeg7mNwi4SlhWAtnbE7aR4dbmvA3wan10wN1DPcf3iE92YJ/
0HKERFmHyqdjs74wW8tR9xF65U9Qr48aK5lwLrtQM8EZJQ+KbnDJrsfVwdy2FVDs
9VFgHK8Ik3esbdFKbAMSJCVgZXYbk7ZUcLvNW9yqjHtwwu3dK0Wgmyd/VCPfuebi
C+IkGPgB3VTyFKtwECwrokQEnFdJdwab3rZ4iPvQ5qOjwFxXlyBZmCIIoSK6kCpF
aH58COdsL5kjN5loyYVRiBb3hQV8zOZToolt7AQN+3Pn7HQD0xcdanROCMzza05h
sFx3UmIIMoz95mUDm3gQdMAgrYvGPQsZVPDQKdzFOhDu0h7zoSufuC07DpzNV9Ti
ML/FDGYg+RROb9M2YeKE+sZbNNv91c28pHN17aiauF8WVTvmSAhhiXSu9jIn662W
Vt6F9/IcQX2mdHTgUVzAWVUY8sUcxt7qfErWXbdF2MTJOoylo92p2DsuFEg0NLN0
o3RumQzQStbe2caCXj6MVXEUF/FqzL9s9BKF7cDYeQddHWCCHw9/kF4/DonE0qS2
T6Mte5PnIMcuc3r6GgtPQyFmzxi4qTi24Epn62sKJq8zSbODsKN73v9Z9mZfYXFv
aID2tFESswIpA8jZJULO7vKL6wzxOFa01vSyoD1GXrJZG2FGkEuMDake4E7YgL5T
cvyV/pspQQq69BXEU44BqyTfekck8ZmN0spnsbouqC/Jz7ZUVZmsdC4TZnYU8q8m
sR5IZkaFfytvAGj+K+saNsQEVwgTTg+/0Gx3pg70/+SrGJ4G5nYNh+yV6xdG5Gms
FAA4fL/rhCWON/zqmLe39hVRfcpT1zE8yjgcM3vcTLFLHNkRroLOJpMX8SVY0mnD
iLZLER0n7Ss+EdWS4MvuK7mll90l496t1vz7HAouCmnB7UwMu0y7hO2VRCY0y16A
Vcb0d+trM23fItUpHo9+0orHDXANFA2SgUIYKdE8SY/GQspOcJe2WBtb/D3POpu8
cPs+yB1dU26jqqbxDsFDw+mi4FO2kMU8ZCQSHyOGIP5R3pBcOrFxU0ad+CrgpZG1
/G+aIxOipRJOmx411yL6DOacr2m0Q88lOtit7++qFFaJlvjGMzVEcelvPwUBArF1
5KNZANikuOlTlZvfq7dsCw1/Alp6WxH1SHVBNx0Fx0GZeNK/jS95ag+DXPdSETue
ew5Wvt5W6MebOOgXTbmTVdUbwQOcXOHERmoMFchW9pDEbEMs+Q05yzAIj4O9Gdbq
kw2GGCD1tuf49bpGw74DX78yykj9o0g/EDLgi4DTpj9TIKnFuWJog24n4EvzmAzj
y3bQBIa04R6U3ciIL+CUmBPdZzCUFDaKnoBkoPUY27YC0E0BH+JBVMs5zqXY2xpj
GfXS8TTKSYYrQo0205981KRLf425/gEmO/N2w8n0s3s2fWq+mf/uwatZFq0mutZz
9GsHbcB1Ll6iwGzxx3eJBPMTWbliLzTMCiHT5XWlMgO7pLvkLmjARb4rJG375qvF
H16VIO2W4Xy+xi0Vc5wmNyInVREmD2p4iZIlv917UaR0nsylu1vab1SUFhJ3YFKN
fClUKo/VoJT2JLtVOGrAkXB/6btTEkeepuYVIx7e1jrOMazyHDRIz5lpMzTYLNmb
GGaFX2Q5R91bIAjIni13OM0CnpRIBI+XlfbsKvNkUuz0YAy9/1Fb5iakVvSssUOd
uFY/iI/cUrInRwbBVnM5KPWP53abNQwBiBof9hCjkqsSeJSg3lfgbIASDyJk9fNz
qRpQDUQuoGrL4jw3Is9MWIceDy5jWFA3JkOcsuceLMJrnyvzy10OKS6zw0df6XxL
xRDuMhZI9odFa1zDRY+xquenB5iWfNuuS0fQdaU/vcU93AjR4/SM3OXK9wEYgo8E
tjYQ1zyz+ngtu6ZlwykSAlBCDEJSy3ok/vAqlfizbkMZSOAQHny/b4nKJZbXfDS7
E45ZiXH9VcLPwBp5erJTaPnWyBUHF6PvXfNlZH7666/3WLiEER2MZevyghabN1RB
RoHyZlGBrESZJE1i89KMaW/O4bt6p/KX4sc0jMmIJAsnKBN0E7TkYxjgdifUDTrU
AsWIS/pzMxv+ZWHTx3aibIfo8pTZQ+CAjqPfwpYm3T8SohBsi7sZ/IsPhn86MRG7
fjP4UWP89xzogp9L9jC8x+qRT/CHk+8XUNx5Y0UkP43sOptJO+ly0NR1/Jhjyz7O
C8dfc/Nb+qJia2jOwq+geiUqd1Qj/iEVRaKUaAPkMzMvatPSIL2Vv9vKoQTuqh8g
c0rxcinNHh1Bv7hIxQbSuqIiO3aNwFss48atxoJXGQKN5uqrWoT9fWAXeu116PKt
MAYfa+l4aH7H1CMuGoz7fRBL4hE1J0dIrMm1AOAqi/RnwDjNdueLrzLUsPYHl4Mf
Ok14lwI+bJtTubJA1NQoWAPoqk0KWujOn+i9zO3ibtdsIns7ozA7w+s6Rgvf/JA/
qGVy+JFGw/XVYTVh3zVo/qjRklxfFTDfWnoQY8qHYxx2wQ/X7tluB1GPvnT95e72
KIDpLwfkLH0PEqiJAUOhan4D56VPqQzIC0tJfq1A4Hb8YKI6hIysl5ISXJYCvzE3
OLmz/4H2m12ieIEGo0HqwA2SDPFeZ4uNp2g/8zmKbkyRemK79rLCxvuPlhKAZvq0
Q+ban0nqLLaQHWe5bupZ1vogb5d6RMgN9BF6laWrKA+MHUUUtHJkBGzd9cRIYPeJ
zzDIpsGU1kUHUH18Vn3+fIktkTW2GXcpySdpRz8sUtA3LEPQVgG0YF56qZqQqCxX
dOXqCjAd+6M6PSvrH0thyUUIn/dznj+K8gyD/hdfE6TEGUALOQo9vO4mcMfpXAq4
sJVpPJgFWxRtBEiFhQzpu/0VnYPWBdJVlnB4AmKAWD8Bb37W5kmVzyjbNqlI0E3R
2f9RmSPuYh3PJONDszoZ3LS0keS1+L8S8FIynfeHTf1d3hooefWu1FTbUVqND+rX
WtpeG/MTFQI3HHpNQn6kfQOnyeCCEm25cMnxDUCzr+z0V+SxJ66H9Tbo8Fm6ieph
6/tEpC1/1GLBjKD7gmPRlEQMplnaI/3vbGuusxKaiWcFYm4tSj5LOYUKE4QanI5I
0Vo6TWz8EM7q11GfzutVemlwM2Ww1BL45oerC2Mxltn1ngN3eoy9CGyBUuu39K1m
3lpq+zOh/lFAg0OrZYIqNIYga654sJgsiweuaTAmauU2bsqsaGu2P07ixQFXUiTy
90llso/iteghoL6y6DxIIJsWRuLUmv2+tnS3rXYTX0JNdE5OTNsDhJKoVSSH96dM
ypxfyac6okDXTb27jO6alHU1YPTPUeYtY3pbZxfNrb8dN9vLH55LmskzvxjN737H
9fMHXUgq+8a6TYm7E1tl/csOsiAFTWr9je+vbEzhoSRoHFn+st6FyXyGWkYHeYkg
qeQwvzYzLm6KpWFH2ple8lNTZvSDjsP3ToHMDaz/H/h8sNIJWUtjsyYOMWSl/Ree
mwAUDAk5KPEHIG33fwbfhsA5DUAltzB8+KDqrRVfvnbYxp6IdlwjaZqDWFtYzHYC
BY6pr05oGvLw1WKwa4VpyfAUEvC1BAmOEjzmgB8gL55D4myjw3RPrnGMWca2+Cwk
aVztz0RWG6SJcovWeZxt02Uf9N68wtYT+xIo1P7Xn9nwWpog4CmRM9mZ9JZoLJGp
4u69zVi79z3VaV17IdxYfuKIg5o4TCjf7nAiPTa/Kwg+NOGUWvsuKdEItxvVHUzv
IEAN+c2eJBWTp63H0cIlbVAHqUuiV3g6SZQKzKbxv/Tw2vj9eDBB4yvNdQYl03vR
3m8hytEjEYJS+MBsQvSQoXtZlJ7ijUx4MlFLL1zA2RriYP5yDl80jXiCooO2gYpj
tI2U/GwKRNCKQpzRJHqTzxX4UGRbtjo/cSyTyhpOWtWygAze2dxWfnHin9IXI7jn
V07pCePtuAN1blF3z1iZwpceG2ShO4yFVcEs0qQljF7/hMJMtnb/EUt/DvrafXIx
NZypItK8Wm2y2Xu7C11RtjeProt4jS6g2NdXkC3kvJum6y3jj4h/dMO4PRbnOIak
e0WTSEa+NVzdKLHg1De1HdZkqv5Rmnik4TCvG6nmIPFiiqmBAZ/Mf09I9kBD8bF1
KR2x5yf4PZR2uxFXuozuyWrnSbTtTx9RfSX+mQf/kycpi9/rq9OBNOo0hUUcV3zi
g1eZXgGwohGLgcIH0aKGdyXyDzsWpdgZwAa+boM38jSrpiAM1cUKOvQUSCBhwxR5
KshAzu47d+GIGgGeXPYRo756PiFCR2bcjhVvA8RK4L3Yn1EbLVHEKtCtuKbONpoF
EL+AoY5Yl90rKI5Hhvc04N41gMH0cLiPOh+g2IAMUWf+lbGtjfcOHWY7uOu6SSsP
q+ARsxNTEVFwgBEOZt/fVaGSeXxv0VQof8sg4renoFEDeCE7zL/ZqF7DeFXY+wwR
QXurZuJFiWRXlPXIdfp7tpjElRnMqkOjqKzrES5UqTALLoy5G7T/HAIN13rXMaRs
LadS306i2ZCglt3ROjx4tysMbno9krIhv9yGVB6rGR1KxRtBxPhPZopLM5NC+Kkz
7LUs3xSOi9t53YJWPjw86hNDqQGDZaIaVFNk6bleyO0kbzZR8kikTc9codshfz43
WP8c+H9ZN6b+YVJuMM6gxcijdFY6f316iVBW8XNbcCy5+nckuSsPJQhrZk+7uP3e
mvumA2NekEkEqHXD9eouldaNKZ5u9gRapGd3yDCWeMqNHRtvPAdr6Sxs+qAl38hm
0xguQ+Xo5tEPYvDPRspNXaPK/v+MsEKmS6WxfYk8dxfClvU21vTxT8RMBihlEsLk
Oyym1Fqz07pufZYSIwn+6yBXHsyAlf34rYY2FNabiJfJkogiIdI9qQVFsO/mpwtF
eE53cYsMWcMndH7pmdyqgikBQ7jOnzlRmqcqLCLQPj+WaKpf31OT5hF0N4npKa7h
rew25JmiBbYudb769L4IiWYiHrVhgGVhRGdeyunrL3SSBBpNJXFl8LNQyKHDmjHT
Lrjiijc2Psw97nWvY1ZHzAwmp2chi4wU7tG8w/sm3itq2DZyrH7q1KPdN5cjfzqr
Ewqj7+IziEzgnQf8rlTKs9/W4G0A93KNeLbcYr8AGlbqrEzkJUhmf7DfxgU5+PQt
abgldCcSLCYq4mI3z1blXDO/ESMvhaIEkvfDq96m0L0TfvzlYe8/RZBNUaX2gKte
S1rIZVSgA8hEvc8pb+VAnZ/Sh/ufXn95WTmISyms8A8dJsrPmCaOMaaekUolzxfp
elRC2pRvO53tzA49LT9lVEHcnnvST7ORaVMiEISJv/DU/mTOgs33yMZe2pzmYru6
i5g0xt0G9CPlp1kwPTp9Esg9iPWYFDCXegTJeF7ML9ZoBPyXngUgyDJTkVc5J62g
pItvu1zVTLh9wLja63QJ3IPWcoRWpGzQb26pOiP0f6dQmWGmSjRsk5EjvImNkLTZ
SvhjaPYboHTNCQVbTBzOSKbGzfxfrkRlIggJhRtA/RsGoqwObUNYc9AoPQcl8jGm
xTzu+wJgO2jN7JyYk9VAlHWnGR/CTtDNAh6UhPRbLeWidLE/Ht+KbGwrvFzPk9TL
Lx5JDs7iuzPYeUFnvTYXWJrz1SEfl9Ggad7hgcZOwP0cLqRDR+GAlCDLChtzEoS1
Kl05IPLyw6bU1/BzKkWhn1R7hi5UzvQU8jSRAdvRPsj9fQMcisFXTr2sOb2BHFrY
a8/98T/ylMhAkCtQ/3akUzkTg4it1grnXAgrqcGOHVCfB6uWbDC2DnhlOTsWp8f4
9LYdMhGc3UuCgiyBZwv6TtJ2T41LU9yCsM6EZoC9yASM7fVbzdkbBM4aWjM+jpcm
pd144Zrnhy5cHuSSE3NDBDLMZMfLwtptROR3q1tAF/Y1oWdSIuZdAtf8jsZY/CiV
yEke6HEOaVAx85/y1qErqZgA6/97kbLZcujPk8yhvj2RRUxtMWM2Uj/OcozlggJY
+i5mYbLT9RIIZksY43Cso0Icx+PJIiDTzuY6kzQRNm9D+UEu0OjQQqaxMu9J3Kg0
L1MT5aUDW64eaXpcEn8AcY7P83qvjoO77WZH9NpW6i3lJMY9dgxkTt1hgtVZ134D
a4iGrGWfcAbDRY0vS+9fdwdyOYWTEKjMTmOh0hYcZIPRc4I/XD0f1w6nlY5Hzzaz
7pbcYdj/i4m9NJ1WTUbdyGK+ZsiIGFltjbRX1Lhzy2OB5HjPXGkqnVOsgTtgLR8U
hEJpZuuEQZ6xsjwbAtIInR/1gQZK703rf8RSQhvNj0urwQ/RqvaLxAU0hVz1vvRN
MXN3lD0nB8k0ypwoEoszUkcIXc5EPno4CdqQxmEc+d9g3L4Vh65XgbZ5sk7aRYjv
K7/wC3vYV815XN2RdODuDsFZrjuP+PkWfgCEBINMctQ4Qm2jyJd0MYfgs9JSUVry
Xa5vO2q88TKBzykA+N78kcVtK9E4K1iwS60OzGjWDKwfKIbgBOg50zoCWmEOqQmG
6q+Wwr8wqVdaejVkL7hq7TR1iXYPA/voS/XaKEKzl7o8/yH+envAi3rO2IzuOxq3
hk78cbQM105rEcvVUuoY6iy6UBFv736F+5qy7BoYaVKLo9CJT7C1CdstrLr0hiTR
GazCPrIKCq1irxKqYaARC6PjN+845ycZHjT+oXy9pWP2lqMYO4xvGHLK3UEmjH4T
JjXijSsnw25ryRS6DtdqwT04+Oj3pCmcYiXbnhQT5lX+s9Q1qi0Kr6Un7gkO+KPm
tj+a9vQcZGcUDXVt44JbZ8wbqKTJM9Rh89jc56vi2EjTFjZOb8/AVONPyr4eNMRS
XrLEGoy0vcJnXGOlvkf/WwzjQ4KRnHx8vH/YBmGGJqa9GPB5iJy2nSHSsOJqBYQL
mTa+aFdVhIKUHhWJP5UZFLrjfmCqt7akMPBUSEPXLSogH0fu9NzAq6+5u0eHhHad
sHhUoxCQp0o8RAyZHpgvXQfQ3oIJzZHqCnA7zFx1BBOCrZhW8u4c3kt1oHnt+H7X
MyUJXx3TiXRd2ylvsGIABL6wn6FvNfsUnx0S/VfCqDNFsec2/igow5dD0eEcEAVS
6/6zfUKMkkEw7YOoAwtMgKygTgTPUBL4NelkNG2NG8lZ+JJsoVi0ENOte3jN3tl/
gdOW5XBif7iIKpvPNEFpC/77qc8QNJ0hkWVOW+GAGChzklrHqWrtvuMCgXMSIqFa
EEf6hkqkEri8FDGGvW2X6UiTeNp4VnwSayOlv0WQqbyYFnM6M0HRTO4Ew02mB3Jp
qrqDANYdIzvkVXldohVWmjicjS/EKLFUA7p83fNx7z/uJ/4sQDHlF8/sMzmjwmh9
ZF/n1NQesiB7wreT7lUXmVIR/UaWpQ2BFgpgAFin/5aTkjH6GyeUkqkO5Ooidkgz
I5sDVa6K5omard++h7apNuNXPzKvfDaLlHCCtfqH0tzx6N4yzwg+gBB97KzkSPYj
2TqbEQmK3cop2UhhuRRXMvZPeXsMhrQNXuNygKde+wrJSOCGfwkZ5Nv0o5a/g0TS
oT2scq5vItYlQLxGuSEChEn3KLCNH7iErNGLguGz9awMoEMKXLbhZ+NWMz178f+x
x5H5WUg4e8C51RPeQdzGmFfOCTipBa9tZcRdGgSgak3WgH83Vty5CXoPbdpSQ9dj
/1a1zWlk4jY5mSxPp8CxcLEzvAJjYOU6ycgL/zSg28zKjpD9AXarmygCrqsV0jzC
D8MyKtP01FJ1hYOolri7Q21eycSYaApTzGLIJUbmuywwahAREdzbVjrIpyo54Isp
sC3E+vD72t2L+EOl6wIQvJcbtIwHh+AuaniGO0NH/bK3HDyhRNMxbSW7iQjtqw1W
+EfENWGpSyqtyS+PW1O6ONSpRO0mpYZ+IZepdFqemb8c+LrP55YnEsY2ATuABH7j
tfGtxbROZY/dB6KVjXkevXGgSddgi8ry3orXROEZuk5Btk1AVPyFJy+GJX7UHoVS
IBqV7hFWiwNKpYnDDwPBbY85JW3WkzL+O2puexdSxuvfQUEP4XtpoAfS+kyvnTVt
aCDJhYSpN43D6VaPdrWoO9xBPHhHBcn9zK6EsGX3WFZ9ieqrkgHysfcg7j7l5TS5
Y2g5cri4JfuY5Q6wvzBJwnzj9gkmxUzDBbkey2S3j+YyjZsg1nl7Fxc8O3dguxkW
dOULc8t+MKOAAK59lUP8uZU6i+SdwJO1ejS1g9ReHfV8sXKJVINdf1MwIx8ZuRIR
h8dLVNL1pR+CkRxnst280ZVV92WnIKZTJLd1Cy1J/qJvdYVtao4ZtQ+/Q11vnh0r
S75oisyJucok7qNA+hVkPXWyDJTsFuxkvYzU+NB9gHg13SPO/Z2D5EIYsxlwEfjJ
NQw0fSGaNkZu59nW0LxZ11cGW05R63649PJ5jwIQ/mfxiYEDINgiartzYeeW5f3j
+QWRvq7eg58zV0Xle8jnswbhISXnmblNxsrqANJc/jXmVID89kL8XzABD6w0HI5g
sX2EJ6gsq53YzN6Mx84ynKvGjRoP67fU3pxVodwjeRXlTpRGEC7HCgPoFx7ldCnw
seKxZjP0uclqeVeZeKC+H6JAdd0CHSMy+EMtFXXEH7jdHJTME7kZLC9dGdWlOKT/
w9+0E0w2xCB+ZarvRuiFmHa/eW2O6vgyqflYfes8ZKWT2vj1h76vF2f66eOfL48Y
+H97bJpZqKLBn2jkNPpr5RCmxSqsLvREGmLhinfUygm8h5kXEJg7GclI7tbC/qyl
ddi9rXiml6YavaMcJui+xcEPgJ1GQAs6eTGEjIB13NEBgwGFDquAYEKwsJFK14tB
xLZlsDlweHrOV8oIUTz66sPtn8+jbU47Nz27G8W6xeXLE9mImRNS9QWSELaQrI3t
HCgsJQ2TPSUHF6n6l322DTKDSEAYD46y5h9l1I8f4R7QHDBan/lRJlS64O+DHZ2F
Q2INu+oqZsbzdnDDiVEzOZvVS0gfwju4bDbrscoUK+I75wyk0drMB4nnkzgtkyFw
dLclKU5LkcVp5n1IJrGBXf+12T9r54BUjhbYvP+jpnN+zF5Juk7jBE4pODIrA7z/
EEVkqkYzuq++l72JGO9siiR2wqeccqB4A/q+vE1cUajXMxatkKlxMv2P1WAoCvXX
5OfJUUNu/YotTLTfNn8antLS3Pp/d12OQBduCu+TIyqhsgqYW70bVtaTyEI+ecgV
GuNeRdU8k1A1rYFhHVexsSQhpEJm/3zcgDeNz96WXMnyfuyWBac84Hi5Hy3DN7ml
KZ0m+VPARZ5gA356GSLvL25gN3Ts9mMX5Cggzf66Ks50kJm85TD7PoaSyU+UaSKw
AHxufT640YveqM5A0HoK5qCkassKtrEorbGUKxdk+LMnrtmj9VDBPuvZdx6VLrTE
mVeOlG27XgSXK6vELKCLk7fP/dchJaPlkuD8rGd2kV6Nsws1mf8AhMcs7OvZ+EYa
ucQD6Yr3bFWvLRpoiqH9ew27e3JaHAJCaj28Knfqjw2DW2WFamaWtvuX8nEes/AS
JHlkh9+jPYpAAd/IeezAOszwWXrTGbkWctGSaEkv3P8t3D6I3cbORjQfJb5cZc4D
2o6n/jqyg7BouQuCAUBiHePP62HMPaznGnHWxEnGgGqXbNpmWE1oqsLlbxJs+ocm
1YiM/wSmSTTN4hA5gbS/WxfboRNJ8Nd+o2FCAtoic+VDZ6qkAygywm2BGg52k37D
bUhajy7jJ1way4UnzqA52aukS4+4EgBLhTVNtuG8F4jBER1+5OlmqzkSy5bKudIg
5PD3Jq0wSaNKWuZVwYCSPr+yynnAmU3jPqERNFpUapv69/EG95/gpFcnYwyQukeg
aWjfJS9DQsJCGVdr4jcJgV+Il31W4gZj9U7XXllVU5eRWSTHSakk6EUpaTZZOSw3
4e/AeKQE6nGEG966wiCSvhrUaeVQESxDawpIi2N/mnmD99dawM3yowA/HC15pZT+
GwMprJo5Qi/aN78G0nSRGBnY1JfLQcBGjECYg48NgZ7UsEKykULqssrGvfYkVMfT
Mfxi20I9nlkAf6Fpnnof3LuZcogg5ixrqXlrriK+zc8MdPZ4Y97/YcwyJBuhssjC
kmNLAALsx3n03JnmsgFxTZqkcvkIX8373JH9d5SECNhFt9zDP936TQyCNtHQMDFn
ShtHJO4u0w9St3cbzFu+gDm7Vas+xe5a8s/V9YeEdcA07eZSUZr3mioEqCsuySas
q1To+RPeQscCv553+fmT61QizGkisDB2eqaKLSoV8mR81krUfiUTYh56mk15MI1c
n5Lydh/yLRGCRM8GoYBmhNErQL4deNocrI6vvCeX56XzL+qhbnYYaRqYZsCPcQ0B
8Rx9uDzAORdFZpYToNCKRPrNMUuwE+xymwjx/2z1MCMGvpPzWMi1ndn/AW2IkL8l
YAYqPWapJ5DMt2imD2tJWBANToTQaPN5MTHH8WC2q19iiu0Y64YoGHE0vK18Ifkg
BeqMu14EHT3w2FX6U8rL/4z9ZTRbelQIcJZ77HBmLyzrR875a5ILiKyDxtpnve6o
xnmifw4c9R7qNDJy7RXN4C5FZZpt2ovvXa5fzekA0iW5zfPNtGARvgOEA6oc0HW4
vFNY1d6pPyzoIPt5Ot3c70SOI6IQAbL0JI+1T6OzxVb+m8MT47JHsNVaU3ebX92A
C9KpHAhguhTwRWOjz7zWT0f4lJi5XiZvEmXEeG4ycYhw8LJq1d6W21US5EGwVoGy
6aio2ij4NYRxBHeGvx3B/AJRhibh9mbAQgclo7oIBe11HiPPJ9k8DGb/4TH0LdSd
9bH3Ow/JOIfiCkOOEoL4giixPTfx0PvEpuBuSwB/7L7t1NtULHXB2ZufUmxyTSUK
I8UtqX7cc+o9kGxorj8zGqBA2ViXfYRyZbsQhZ6avyNCUuab8ZEFkA/WEquhyl/v
4f00h21ykicuzm3uXa3zknoHBJ5ZNYqOyPiUtd1FkmtjdVmpm2j3EIeifWxyQjx3
LSX2cdfcLkeKbl3KDAxI6rD2SEBwmHFKVMPbYVijmg+Un9mSPJ7YwQ9GNmzM8lWM
5hGMcdtEsSQE+zc/u1GscAWuVcIKymi+ICc8aMjq3uy/dknUHDJ4Xxzvx5AkOyRu
atau8CqXp5QvGqpyJ4Rh/kA2SCT97nijG3G5p8cImeTz8RhN/aECoMJbSHUDAM+l
hGD+23/gcKL9ll+5VOGYU5AN972TD/smXtlRs18nnp+K/MB9qcWhZ/Pag0U/qr6J
XpbBt5t18pG7xONjRoFGvTV9K3o4vbg9ZUb5hKdbW0hIy9J8k3Top0uStJXPCZ8b
RFZQJTHvj8PJwx+yD7JaygFmlQeTS20+ow9x8K2lJFeNucSVUR8uJg7abt2/uagi
ZPZA/IZf51galX6hfXURjQ4K/KMIYvar5gl2wwbMYmxzJ+99Nxq+bNmv9egJEw61
DtkXCT5ucorOos5cbVuX5D5t3ivtvaj6GjwLsfBEKtj0uboib72USfiIJCKuLM+l
4jF6DCd3+ClAWwwsxb4vBQWgg3Qv63AsAdDRJhObCUaUDOjFG/rr2LGoULCAhqJS
K15tmMGNxDDJ1mkHUzgXcxa+fdOOA4sX+wxhKxmc2eSOWCnNO1K1mGgDPMfT0zoL
kSQmc9qFFvfNpqzOi/S7RA/RbhtsyAZNDLy6+pcPFjINQAV+c4dfwjweC6uUB2lF
XkdB70VxT+Fs7ydZbKjLa6V32WBvyezd6T0pB/inTlsTzsOb2L1335Ku4wK++cbA
xnZt5ksXgI6jUanarQqomLI2udW2v+/YdFv78Yts98VNoHow3l6yEDyJywbCHXyW
Xmph8i51cmOVKAC0diuxP55vf7oJa84yxVCFvUwDcqWWu+5fGlrYrtfxQC1qvUg9
LsAXMjuP6qAdvbxScm60J31qD8mnM7wf0iMrHmRVyQM0+jmQowGDHdtjfXsADG+a
c4o5o4EUciZvBzs3UkpIOBv0cHCk5MV6T2fIlhuUFPDEAWuBAPru6nuDtiCGVf7R
emBwL4WwVzeDPvBxZ7oErYV/SyMyNVzoqWGsXQWd6H6rDiXPuKO4lYiW1rwAfHSl
KsSmp723D1EZhpzVZICl81L580GdWGbJgrnZXo9DTO5pr30BkSzUAA26nC0Sdwba
G914mr4Tx4oBDkZmjjgsYAgoZGlqEHE+40xeK4NzLAq5vDSZ6T+aXFohYKW1h2oe
vs8O56H1pfk55qT0LIJZAIIcLKZo7hOa99IOMBsiyN+6x52CeW0cgaWu848VG521
tZuZ6bVmN0m3WPmiCOI77aL/D8yRQMDCsQkf09wo3zFBp/Y+ZgwMkT+YSREr9UlN
P+iVuIZC9PMaRxCLqRA9+dtPkMHPwxypCPv7j/P5iJuW3W1uM01NG0mtrJyID5+/
s+dLON34vwi86POwczIDMdtYaOECU7dn77Hc0CrYAGgD0DKuRlsIg5y9DwOBemNm
kb9rYww7tu/m4BbpioxKwaPa7qBZr7vqBCqq5Y+4PAOHeubHJ2tqQCQ+dgaAav9T
XNso93LeC5b/ECm0CGGFD9JRRYNM7Nw+lAdKlgEkRLXHftvX0ygqDaW5VnGVcbAZ
AfCm/WuYej2/XDYH8jHlV2wtPZj3mZfA66RKr3cEPv5n3rWPsx+MtYvOZM7pDlBD
0IBfhxxsr+XSt4kcUBfl+CCUTNDKs2vmchI7riZl8NTv2EWKAzIfRRlxzxRRdEHa
/WFwMlGf5LOv5JYpTmRJNv0dW+vFmrNiMZgKb81uNUj4X41yQ2B0RILxBL9KDHRw
o/4NMDPQJgNXnL8LLiGsNCBc+XwyXzAV4sNAoorClezuVD9n85vKBrRyWtbnqw39
aT6noxR1iYwY23JZctWGr6Mtwf6cVnUwq9gr9OultDXsGgdKT/kTXPKEm7FPbUXO
VQZmZVyAwSqPuR2B3xdFD3p6JLPpt9aReqJtf+imZrLH0TlOUc29m2r08qwyD8Wr
0MNQMRsmMC2SGMEJfpnl1o5ozPBsmqA3Y9iUTRum7qBdtIy2+Sc71vIn/yzJe8Yh
SI8h1b8lqXDh/ra3jlECyMUrJ4dm3we+Tbarj2asTZ20nJ8Z4VWytqpYu78sa5IU
26Miwa/riugUoCagfsQFN2L1gMmmIX4mo8MLqN+mYlpwhg97cg6UwHFawhTaWQI4
oJXDgsPZ0yAoo8fQCrmX95rpLGTTxQ7aZWv4c/demmqZHp8hlchpOFEnSdutvJv2
H0BlySnr3U6SnSIhq5w1VkejnQdPCdaaha3GxMHwruAJBiek+XXYNolWVGrRhnIf
m0DaijaHPft9zKFdNL420EEWlT0oVaZn1BsZKi5pFBJ4YVlwOXW+DuPFHTvlOg2b
S1pcFdMR7OTjxk64+AnpSHVy9sfarNsd6jmwyBXjQHM8VCBEOiWYAJ2xw+PVBWD2
WFgJbK91HqtG48AXDN651XrAz3m6nDNcVMNs2skGCY0D0fkbGWkYDbQNzOVcLE8D
QghbltQMHk1BAd6gVAXhTjFUTzX3XkNvDEL77bHXVS1xxYF7h1xcxrC4CdUY5fFh
SBZmBEgS8OhFidesP7Yoa8CTtDjFD4JFFxmfzHq9HCE8/oYdCNvuyoM6Vit5AYKN
z8lCSQGNpulDNUHgJUEOA+DNBX18EWyj+He4DiksfRyecAB5lKowEfI+ZITuaZu2
WGzscwosak4VwKz1TcL6EWEA2i/I6APe5yyMsPwvdnAQb8IZ4yBk/3bRrwWqAZP6
6eLRH6oijminN5TvcQeaJzghqNLSZUnILSJliRtcJJ/aHOGvxg4K5uKtW64Bbwpf
wGyagu23EjCnU3tGmElh9cRt6lZcfOIDIkaoUzXihYrO7q5yifm/Bpvr+MjO6u1y
Hq7EuHH95SrmE6ZHcM+X8sW0EoqiCLVQe5w5JSDqlD2U78qSYxmzyTE/ZTnvf14R
eBURoOS9BqRZtW3yV5b314Lzqh5dZikraScolPk8fJcbyMXfjlgawVkvmAHnpE1O
/W1Dxz1ega4r6eHTnoEfNSWyRsjWmHrzPM3ICVdTpw4PZCnp87QgbDsApkcYya3K
WWruUBbE30mfAm/dgdKT0UA8bNA8e3VTpyu7V95/mSKd+1VLnIiTdVNjD6KqRn03
vu8pJpXhodNyUPrChnFW9GH8TsvLh9z6tDJaFGn8hU8F4A9tebBBxRyM+G+ZHLhG
XCk+gS82zu31HT3O0dSfEE/3uWaRpFuO1vYfYtYO2h6GLDBH8/YVdpxzr1tzTkoV
yFchb/DjhiSN//im60SCB0gOYMMi9uJF6S5zd03tP134Ca7pL/0ueMz7haq6Ik6E
SRmt+oDNyBDyUlaTVKHsHy2VnJiGTif9R8a5N8Jq5XY3vX/vgubthJwCKSB0U4nU
sI9Jb2n/SIKBQeWsPMM56+wDvD8BXvrTb5Qp7Vz8oAXs7k4RpPu5B4w6pc2NpA1s
V2jdrtwRTAAcHdCup2EwAKPOVcYNmceENg8racHIkWWhClA2V3NypLkUJ+OeHLl+
EAWOVE+yPbEsQpNmQUkpjQtEhzXkuaUfr35AbjtN/H8g49F5BQ3tDAMEw0kpTs+q
1J8w/ndRmdSgcRGRq2PpGijFgBk8JY5/4uQe2Wl4i9z/DYgJjxLIVK3Nl3cPA25l
vTqwhGTBnEgAXEPfv0ilzfSfM0T4faRUAtb8SSb8zfAWMMw5bJ6WXp3WUwc/27OH
/zhiVQ3YPWAxT+2F334N/qaShD62UC6vuoqtGgZ5URwtKxJ6KqE0GUVsz2+ixA+y
+YZcH2mQRyaW1Ieu7HUOCWIbKwjqV7A5V4y3vfqAtbvnmySAumW6S7U3Tbx3lVWQ
z1d9Dt5OKNKclR57jIl7qbPXfRqt9kWc5Q3uw9dy3aEU4R2IOpqPh8UxI3HbdQHA
uQuVYBtcxyITdbF4QeJBsD9xx7XiBRIdZm2UJ2YiAgGaLnmVO/k9AvX7WflQZQZu
RILQPluYKMSu4tcTOl7nj+ewWomBNg0EQs6nsxfUuK+VfEoGnmzYQ2vkJAQYszrM
TZrn6ploLE8O/tU9jKT6W17q6EBsZT5Hnj0qUVauWcTP0+rte9x0Nap5UDnpgdiX
TH0jUKhcFPhDZUDK+fvmvfMzMN5ZyH8jxDjg+2ChAoFzUeMRKwLAfb94hdYGtM3c
d/XKcL2lLKS3dfr+GlOoiICF1wLiBZZZ0n/xLEbiI8oFlG4AuaC/Wj7F0NNx+1z/
s69QcWNzrHjRoqjsGpfsoo999lfAhflXdQEHAq/tHBnirdgGYRz4iErUxSaQaUV0
B1tW1nL0HD8xzMT97wR6ajzeGfq2meVvuOHQduxN9+IZXOqVyKbnVT22h8oJxe/r
0DlvwXWQ2W+0pPiK21SGQGTbjV4jVO6sE1RLaaYZGXricjN+uv4SO5yw8g0e0zsB
GiEbOC8WfZRzeRze1UwSFozUzFRnGdX6VPg/lBFnpvsZpoui94tE7eX/dGPP5mV8
V+rU37LGCBgWEKjLdlMgHe3bjZUCJOd+i1o/R7Hj6HOdiRwJtc3Le+C365Dt7Brq
RXMnhIPYzcwezWnibKLxleRfIPac01T7blfcKBXsVgZ0CbJ8+K3S3kCGDofFCLlY
UOe6P/I1+XG0q1rB7lagnKWFImnwwZtyduv6Cgnut5wlGoEY/BYHtJw2eBtdf15p
TfuWbhMYKWnnU2+GBaU+0pGo/YIo7UncWs2UvUCvRQWvsKxnAB8e2LiFBfRTpMdx
S5o0+7g19h3jQOS1lgmaZbYohrKYHoZJ+haDUjRKehXcs/gykiUmimrA+PrO38G4
7sJAPuQEFETlI9kFpNHilKINz+YJZqswIFjZWX1iO3d+D0TeJp/e3q1x8EDq81ki
13N4BYFNCS2g0qG5KYs6UPm5VM5D7/urrYh9atmDMCwEL88BpVdY587a5s2OILcb
9gjCKnMPaloNrjbgfp836wCPg6Wd056emwTP4ytMFpHWJqO2ly/ENkogMtnjzesj
NVL95qGrJbywt3TfpblcKgpg6SKa5sTWXL24pZthYvLwYUM5f3dhCJ8VGI6hjb8k
z0L/HIySd9tVf1ujbejsWGatfRRQKf6AXUVXU78nlykowp1qJ3N6BSNNVSyHete6
eTNHcAYY//sbfPeeV9Ze99hdtJSKnOs8Jec9P8g4QY4qsQhX9RtTkrp1elY/TYAs
fCdRt5Hmbq7lDrXZMx6vlkeS31Oaeg3YJUVgDDCPGGm9HpJhWWOeB3Os+WwMWrNb
9Jz4RJLkBmEQl3KodFbfrLVFzatcjDZDehMwQAMmavjgW7XupPyEOBtUG7NbnZqG
8ob8aQGklw2qvQMsmYs+nsNebio5Kj14WPQrqhqCwXREWuG1NAuz4seUugb9FGaY
29KMxT28CK/QoTBx67f55k7Vu3NazvRrFVammVVK/WZiSsXCbnOzhD2sl9T5lol3
0YRMEjr0B0KHOFBs2ybBJ8WjjrMpahZLU2u4glrYPGFtFZK4LFzx+f8iHWdhAhQC
ikFV21KEUwsc98DU5ZprQzF8XLorx3OtONWPz3tRv2nUT1UYzy9G5RSO1eSLFVor
JA3fmqrsKbOgGsH/GXn4Gz/j90qnOYptxtU/xXV2OGRzJvslFXutW/gOCX27gRcv
kN6n8mHZQJEr0IJvmvOsNa2uuw3UOuh/vxhB2F17vZyRovApQZ2k11r0e5VsEljG
TgVJL09NT02ZzFj807zPdHMGhYrXPjNdAmfy/qIlcjkVv4PkyOhHVqj1oebt7AIh
mIQtXc0uYzDvtEIatAMH3KWc3w3L4GEv6U8PyZQzYAU9md8fBLlEHPDcf08+9el5
2t8XXfj0NID40GNZTNCJA0z0Bw1PS1oCtJKgKxXmQ2XH8wHwFiTWqZC7sj/Tihs7
Oy4dNWFb7wrH7Kb8fuQWDxCgv6dQnd3221QmSOUGxkLvX5Fuc9C+DsOJzjkV5Ov0
dH8UawhrmGxP0pTjfzen/vn3kFSGJRzEMxaL4wyhjDXnjV7RJfwBemQIFmPDIQyY
hpa3kflBUzCq1q2T7EkHSJt9FbCPQZDQxDJYbib21nitp/4pezLS2Ghx5jlCcCyE
2yDDG71gW7UZl2vU9YlMn/nbXqlmOdnkcXryb7j5TkO7VkHj+Rvr7oWJE/A5oM0Z
m2T4dsZ7axap0ydd7CMlY8sFxyZjg3/t01YcM/r6loLHUOcnC9f5XVLk73d+y5z0
5Qxg0ZTWsaiqBnajEAQ0jPrfUyQfJHq+Z2eUifMOiHZXHCi8JSYSDr4XQjQ1iOiI
TfIv9HvFjHKUIE1TGMTZtcHx6+huUg949nHgWn66IU86TmvsfHuFJPLL5CQ1mDQh
T3kzkyT7nkxJRP0gWKpSIR8lrGwT6Xu566MRXlMT8EuTv5QIJKZjX/b3fAMWy+5p
q+CwiXVrVK8FbJgoa3bezjn5mu56byFqcv/vmW+IjL5L/rtCK9wX9drlDNvXm/mK
8Gj4KPdL1nG8iKeYF3CHqq1hp47Ax3vfUVOGxwTScNT7zd3V76LITbJwciLLWfTl
12aqIgx4Jym+D2M6f2xGhHhwCPlnU/2+LjCebVfzFi1xG1/7h2HB2lkbcPfUfwIn
ojnTg/WhhhQgdQhIQMpyamitVWKQ8jRxGVZxZt/3PXPeo3KhGGHEcQFfZ7IwH0w8
1ObUeWAGMFxSIq1wWb++f0eqyE8hjuu2gzixCjb6Z/K8sgwAl1cmLq70bHsvOEav
gVkpUfrPZ/Jvpy3bbjc8hAE0aBfnsRStVu3cTgp4dMw+G3AN5uNwGkTyPnHKHzSa
kum3s5ZQ1zVmPsbh/SZH7dfQwa6k0/tL/lU5cnWaMaURzqA5rOEKon/9sdZO1Ut7
secbQNvHyliHDk+nd2MyZJxJqhJuRQM7JhTZ7D9odUwv2vzhj8UDAd5ZRAq+rQuS
Vzi/lL9skZx97AYdKjvbA3lzgBtj85MDPJ/lhe7tp0ZfvM/j8h1Qs/COzqEI9gJg
uMGm+5mxQpS2S/rA+aOQMuaz/jl8e18MV1PpFLcM+d1qLVNs5rBZkgDwN45Z7kZV
CaY/MCVvI395vKjn0T6IMEdzRrJ8PpK1SsjdRoOa2clXXnF+/DKZs6GQJg/X33jR
l0uNd/VtiZxcnSGWeoJS2d8CHL4JcZhU2geZl1ibx60TUEPfSHhX1UTOFYXydHzx
3RH6CZRgFZPok/50W9wBJaNsC/k8h4Eq0/gQ9j9neCdeyZ6zJEZC43O+EbfnJjxe
tkUvf5sbILllpxchR4m1Sb4fWN+RoqfmOoy0tLYhNE0xCG+rhox/yhyAwBPsqQyz
Z5A5digiPQVUTY02fVrjfnBrCzXt9ecM4ybw5Urbl/COsWziLb6knW9SyCuFzeIu
tib8EM3SJv6sFIS7/9PNMi3SfVakVH8QDpUJ6dhQ3E0EHy/qVwgOO10XvQf/f4Op
L0lQzHwUN7BTTnGUpATsWLOnvh4/+FwrTTkAmyQSsP/p6gxCx1S+2mmRTICfSkxX
Cax1eSSDtuzYM0vDGeZ1o1Z5ziSaosPhlfiAwikiOh0x5cvtKxJPIzOrBKoloYvM
5nzGhwFaEvKmezrQ9gNJG7luyT3s5lKhKrzdX6ZbQYh4D3LosVgOxrnYiLorztuy
OuG6+lpgiKHtJHYIDtAFBpudXuYVBJbQZ9uIBBq4wUttZvGSBfy02ED2mT8E6XIh
qkr4nHaIcr8GxiRsg6pB/w8flWQYKlAk5RdHkvD4OXXLJvqdY64XM2vlBc8mjRk8
yI+Ycun5LeiCpuLG+0AJrBo5NCV2W0zhzCk7jVs0aOHONkJA0vwlcnHj5QNzeObk
4SgtaxtBs2QWdnli6ZR+Gbfb0BHzFvtC5tWtcSLWk8d/H4S4vXVV3BRjVkt/RGKK
19RGtNZiHiWqG5E89ICGt6fpbU9c9lQ1OJ83R5m5Ou8mzX57kZWOJBIY6lZ4BZGW
HNFz73o9VIg4BlF5dIKrwjfNq2TskzUMlyEIEwuX5KYbl0h9KR0W0QyBLV7xmp4T
YtzJ50wA24AD8lMP+bxpgcSJffhL7vSPXj+4OQcwq22ADG6Y8sBasgMPhdHCzlAm
y/l6tlrXZltN/IjPP9gJWRmaQAhjdduybW7W+TzDAMPmddInq+LgbZz2ok7pMQBg
yuZ9vOyDHNmmqdmvhLhvBn4NSNrWUY114ZO/A8tu1q0T7g+5DkEfPScExe4dl6pV
R+fz9F/UHqcPG+WR1lU3NRy4U/J1uDvliF55nyfsps8EmDvpWpIVIBHXMyIYxRAj
7egzDDYviXO1ZxVVF32dEOd8gxRgS6vklfj242yEtAKZRGICVG4E5dg2jZzd7xaM
OXXTo7tGXh8re4NQQz/GUulNy4w1pZBRrQA2rdo6FTII3+R2s7uWBL60AmUV9R42
J89wfHljMXo7n6MZbGWWeo1z1Sph14V2TbpqVFrxt7evkcAYMJL7FGNoro4GuITp
Gx9Qosf/jXvuQNfpttiWKljl0gAtMn2JmMXeIfXoBKY3JP0RnQnOJ1V9O/IEver6
+zt+Lfl/o8l0xWLPRpnzJP+rU45DkHk/ou3Sm7Kdv+msjPQ1ScDX3J73ugMKuukb
ysZQLHDYz66xbQseE++Zu5eF98LCiLdEuYgsA+vxvRmh0yTg8T7rJYTRwK2w6ACw
+TvGVk/HJA4+m99TKmPzVGerCFab/3L1COF3rspDLcqaa9zfyazAOIQxigtOz8Kp
B3O4C6vguY1UjHvyFgw7LvFT1iK+wt/AeggXOjPURAyZUgYA9grabZ1/lmV7lmw9
L03HuHd3syK7AMUScA2PLknN9R5qi4sqqmug6I5Ic2RRIYtVQw1ppSogqFMUsDkp
XS3HHbA1i0xHcOuRJXEAz74NviI54ga0HZdgh8QlqdT7orjRiuyInnl+ouZq/wdc
gQpXED3y9rLYPLnpJynTWi7N0Rwv8PLczchnlg5o0OEZyBJD6c8yVqM0sPDLq7Qb
7O5oWGpqXRRdTTJPUPuImnYBW+wDgh1cRrJttY2487JJ/g7brmifPfrmj8w3jqA2
tHYT+z+AI9pP+Oa0BnSE287DGqPUGVdAoKlxkyheDAFN0I94KLPs4yVK596Wpr08
FF7BQqTlltMPWNxzUCM9Ogsh+5Xm0SyVNmSmqNv6/Vk4lXFZmiQ+lR0oDBcIf6qQ
hXp4iA/z91EqKO80b/jH8AuFqclPZgRVQhatRW9jA3HXS4gwu6Md+geP/hP2drpW
BU/M0GgaaQVIfx36PyT24zHsqm11tECmKaf5jORlBMnkUyuL/dg86HdF3Gk0lFjd
JIr6T13IWs8MHPjieswwtewCxPNWxhX7+5s5YRZiQBiuTL6x6l2L3LDHoASNXkBq
sDz4XskK/PMOW1ukBCyFJxdw8BqDj4AhtDmZ5GEptzqP9ushEpFXOh7f/hyBs0ZJ
B65K9m65BbS2b0PTWqzoa/Aq801oYcKB9F7k87zBXhCBkUIvSYmlBGTFr+CntbIy
+jQ1CHcpthCzgGcduDNDR0pxkY5ubBkih8uc9OAdWg4cgWTtJJhkZN+NZCBC1Zl4
Wzf4kO6HqjGe7X7y98X1jOF+V9zX2NPQ7FH7ai+W0LZ62FX//XZbx8mFe0cG61Xp
s2du3NSq6X3WxK1ZurkR9nGE44fTRWtVs4m5RN2oV5yQqec0/TBqhloLLrZKKKEu
Lax74X91EWJqcrQq4hR2CUDvp2FDZY/FYlWFP711RHgQPifxx/2iw9pOtc3imb7t
oTTcD80wu9J32dBot520WqmtS+8TckdAfAebB9CABN+jQOE9rjPqahpdQyFOqCQn
+UEoLr7uWruhXS9tC9rkIht6aN2+fMLxEQ76rgbb+yyBLUa3BtxPJyJeyaKTGp+f
UdmZJxk+HbkvOXxIKefz+p5zqJv8x4O07tKauj6ibR0oyUpitTkTSMgaksEaGhsA
2hoqZC8kAYGyd4XJN1NexevKKxVTHAROX+TvjZlOD974VPBhH0HqPP3kRhAcIwFJ
ElTFX8xyWfzalYAWV2U3Jy6Xsc+4G1p/qCqzG3UOKtATl3sN1sQCMvG5lvl7c67W
GqfseeKGI8VEh7sKtcRyndaA7eH5GmdPIZUzsmmS3xB6ij5OTc4/Bd20X86Xy4Sn
kLUB2IQ7ITT0sllp+Mz/p5spMNwLCoFBd7+aP8hyDWUgUdw3IGXqZMY6ZgMw6odw
ogRuK5x8o77nIqDhdGB19WQJ5JcrI8pA8usvV6FeCubZRlvkxkzASiIML9JhyseM
q2T9gwnbUDUwA1F1BWYyGW4fAmyGQGxXX+soIZHnPGGap9C8zqJQe61lyL9DI85d
C39WRvJ4xa6xhPWT+exUz9O+/133WwxmQOl87FqqMfzpaDt7IWTbBT/Dq6yS2LJw
RvouAOhAwdJZMFgqdgzijSnO7BBKFJw8caoXDJmlqu3N21pXohyOLunC8lJyW+pv
qWUF8h3r/4aKliYYX5VKQYmBFaKIjlVOPW531alDc6y0t7K8n/CNF7hMWdUZy1oe
3O8j7LbgWF7cpb2i4vNQ36tu9qqO2+/1wS5VLGu+2dmBUbs1OQYIDMV1b41XUX2L
BM/44sQ43+Thz47X25CQGedp6IZaqQtEJkrnTeJdX1/rR0pV0BpRbmqNV0gSAdzG
nveuKkA1iJCldA+bGwMHKHTYuX9n72JzFLu0hbeuECfodmXwQWcYNpRw8q7bl8JH
TS5PqUoxNxWCBFw5DRQwaZqhY0g2YTlXBLBnNgFC5mbjUTlRFkK+BR9hzNFnE+Cj
+kFvrgKOVUzPOA7maK4rSDV6lpBXluXYYd1sVg5FMWX+h/0bgfFoDxNestw8eIHm
epnHr5Z9ZIICg28Wbb3ZSG6iTkbdDHm4eSIyuyNMbHBp604Ff5yrztQkHGpJCbLa
PV2Om40v1zeOWxJkV4GuP4zRLSoCqQMjDFdi/xywjEH7EMuYBhcvqmB2Iehf2Lr6
m8wqgZ3bTsEqeM7YUq8X87uTmFygXatEzvTkWuOPjYETrObHHJ1kCgTF8bccvL8Z
b93VXWiytnZzhomgUqQA4Lx8wNTXrqiQpwFysM3L28vEpGiqmAF3vHhgSSTlUaeV
b2cuASFGX+zYm8Ea0FkjrdTSCGM2s3gc9kAlweZqJKeeDK9NJox1QWLgCEfoB53e
dYyLnjB99VaFgktRMV0Ia5d4MBfsnQda6JinnyElsRmco+vp90Bsb5Y/mbdC7VVF
hy78eAlCmurB77c9wlhFaPYEe+7WxyIWuW2G0csNoRCowGcAzCIVkjxQgBWyf5Xj
FtbblSkuqjKHzzC0wgWpQVnpYjT5CuOy7lZ8mpnHrG+1CZzys/RKiA+2/nqwRKUS
uQ5/S9vplIioULjdu+er+7PDlwjhF/4f2JdIXFHKy2VPBa/BuzweA91islnE513r
DhNcpPUHx/MgLkLwTb6xQ2HtD7pM/eB4+ZChAy0QkSIija16acjyAxJ2jTMCeeEA
YEqv3HWs0p39CDmb1r6w1ezvIJkrmRF26Dt2m/oeTqRza4bmiZsZbFBtRKGetiwz
HRlOMfblX98hhMaGvXURO4mFjz567ZNjtEvjhDVlIf0EZjcDClGkHx/QZ6mUMmJC
kTFPpCZTaJuUSf347Xxwte9THFXLa7R1Vrco/Avu72aMMfGoiID0Yq+kW/ykV1B0
ihRlv2rzD+T0yYwrh5qjSZJs+klGdGZ45ZefvYLYKDwusKpNN7RxtzpdoRTM7pHL
FnNuadfwiy4O2zLkWFbcr4Q56d1AZ2QNPBJOIxQgniIAmeBjs9rXK6bMCtmx+Y5O
PsJLsNkzJp56CiI5YHswkp8g+1YrKILRqLV5fhvbLcRrJzdwhukOwuFfoqdhqnNB
E/4WPZy6v90ZRDxbheuYgx3euBRslinwQlODVuNrev+NSjVwsmQ/v4xUrM6vbRVn
1pWoNvMhFjh8Tc6NV5cmoPmcvEP+/BN7pkyEKz9B8QyBBeZnZgZo/x3PNVcdNTeC
wE0+9s3D+kjqj7UjJBiu6tkMONcNmc0dH7BgPgCfPgmH1XX8qx36tGsJUWmsaeRO
vPKmiB6xiCX3qyDIRxWQ5W5I4j6cPQZXkUNtIZhfpGsMSfLeuGs9MlyxMTPWmGQ2
5lU4Ufoo0tvLdycaCfosblmqI5qhh9G6cHXB/7Uo5MZO6LaKRF607vMcbZO3r/4s
CKdh0dar3UY3a84jcK/7xlpZqE/xBqiR/v7yoTPSCNDBDDQOtPRM1uxuJdalMKqx
3nznlK8iFiSYTj9x7JDChTbcLDViCUf193moDEmHgV/3DLTNvDd/4mA7jIpcBlqq
meFxtW1Aq3E3TB4GMO/f7vjnBUmpHPNotuRnfPA5Czsm0YLWeFNBwAf3QXS/lfIf
c0q5iL38Ams7lcXJMOqQ6BjQTKcA80LLlYDYTlLl076Ry3vmIL7ublBTMi1/kbpK
73VpKcUJ7taHlnpW4junji6apIkPkqiADjITkGPEAsnWIp5tpXAH422WmzLKwCmU
XlQ4q0RDekXtEWCwMeIOc1NsDu/xLaR0etJ/8q6415DVGPmaQjAX6+9YmAt5eAkU
vgpjadt0i/Wvj26DfQAaDdkTFHMqp8JFZSid69ujjP1nhfghGhOa9JdN80TvAsXD
BfeLK9H1SRDd7F6UygqHZ0+pijgk3StTtaW+DI7nQfh0eWAn/KtHaZ1EsqdCdEhY
kMM7vWTIET8rynrYP1glJaereZigfn1Oa9BsSh240GezxKf0J/xwcA6Q+hMJFiBt
jpI11K9P0iLCvsPgLrKoy5EA0rjly0XiDRog2gwDYffKcLmqiFCIcTiXQ8Lx7EVi
oM2xG8vhZfD7ttRdPTDn52Jl/Tg4k8vFJaLXAYSqgJMM+/8TkT0ZLKyvoT5SEh6J
VWCNAfc5MnQr2oGnpZt1jOy5N0kRAl7jykQoUuE1L+lgQ7xPVqT3TKwveuZN3gR0
CAiYOQfQcEB4Y4jjbM0esnl0LHKK2Ez+q/Tm+FCw50e8c5ZGcZ/DNCEzlWNnl+Q9
uln93+fGgA9K8wzFE/xf6VLhI/Nh9ULO4tzrCe+PdAagO0SpVxpH0xLXo67OGgmh
NMK4dWoIyTBYzusZ/rAktg6qFoBxMKdjArWZlHSRkLlBnETXkCBGiFQxkg+HTwZL
8Jxjw1LIYW4H3usveDMcCppfCN3vkUPqVDhBrE0zmAz1+QFliB62+2qCSNSr9uFg
nq4cevlgJsuzxhe29JijOTWsVXMzJ4Lk5U+nafowihYd26kseCfqQG1pQ+1zqQZY
ofGRYC/XFftpgrgHNivJYDWw5/XPxe11idicPL444cKKT9SX6Z0onbEmsDApkXcx
Ew59CSpAZx7ylQCa3ZLshmd3enk/MIn4xlRoON2+2ubVXJQKRIJ/Y2zEnCQPeJ0i
o3rpdwQlwQlxgxtZhvIzBlsvPKZ3PM2a9+ygClK2dE7damJD+GZ7OpX6ecn/k8+Z
GOt18Do+CoxrhILU/BtWvgrVpEFvDt8KSsA00trs9wT9gTPMfM+wmcxf5tOvAek5
3G8ILrXRdlvINBCxwuxwhyRrSw3bvfdhWSAaKxDHR3cVB0XvqSVQn9pMJdrwNnI1
MW2Jg7LAOh4GZWrqYjSvI2XESOJ16LWcSDi5Q9G0FezrMgmj3z8Rt6Hf3A5FH02d
VFnVvD0Hwyw1vJwst4sxMOpe+WE37ylRgFeMFwUP1fNRQzaFIjdqzAbNkN3yb90E
jnHZnXUp29BW15z5CbzYNLhnKP/8LAOTiHrL6FFFD3m+DrAt5kfOveMBA3Xk84hE
GbOWhzj2cadQ04L4riDWMhBimoxgD8NPli+UShd2vVoxRNIru4WpVu+Ep+guq3rR
qdkUyUBFNN3wQ2dXvusQSpHysVMM4f1fVnpCnOaZeIpNAzuXkSyz4gig7yE5/o2w
5Q/cDgjsm2fKfcbNEF/0Ei/+vim6Ko9D5JioJFq/QeaYO+NOJqclDoPeLnS7PG4N
vqhur5MxdwdiEe4LE1Om0t/yBDiV+GIOqckqKikc4mvUGe0k7oiTpc/sO1dcEt1u
oz0nO7WK1pYvE0gHlxHfHkjuHHe68VHrCiWkOCF3PldgRv+Hu7NhtFcDwAi0sGYY
mfctZSyBz8DdJzmUIC+8z8VZFPxtpTO3B1pFC/RNuDRhQltAs28cH7CcBRvj0dzo
/qBwqQHIG+kCe4TfCD3BQUq2pE11tY9lzycEb8ZT2qP3/Iz2SIxVn0ug18YpZ9lN
cIBm9F4Udlj+noNsTbSUhlgW1GxgzvEwrSp32uuTsLYEeiYdWFALwy6yOK4g7xX+
a+j0bDJ++9N/H/LDdOtJEjgznL6hIR78gB5Wq9UpDbRBLZy8kUjCQR9S6MeRVZXy
PtdZkrgEQve0Npky8vnfn0EfY7o5ia9TX83jg8UIpftZ6gwGEh+sA5Q3BEUQ2swp
DpIfZMMeNzcjMBOt0h2I/myUJCQZT+rzVwLOqH0aIYICPlVSprcqcYQm1nWfVEWg
VOhlcVulhRjdYgI3+5oOVs9LkUR/+fxuZSoBlPBG4mm1bUU4j5fzNZ762w2Pldzo
rrP0GoMwqr3uPiys7LQd1NvBJWqDObVIW51AMeViNJC0cEbmLXB3EY80z+Nv6RFR
PMg/CRYRzr8MjTSNrgF2Nc5jw0xJWEsy0XUfCo9nsTXDgjIx7sUnz26FWL1KKX98
qTjw7nb05SPoprZZGNhf/cDoU8JavxBBwPNQXJ/3MWsTi/3qd4+IXJT8Vt3LzYus
zOmBIvWKdsDwbbYHBkRbsMGxQeuK5CiBHh2j9B3ZGKWTKEjNP6w96MH428LuopZF
t1yoZugT4LWav6lcnwt4gA8zJFxo388bukfBn2Twt/1FQ4ww/BZY2eGJP1QVZr4+
MoCKUO3dxhkfWrXhSuUeLbe3epBBjBkPk2Pd+f1XxQwgtV/hp5Pr62UaISl4eZ5u
0ACyF/TbDq7ZtSovN0fPT2IpYzQiVj7O6D5ATpe6mqmF+usdYjAmw/TiPjFKUIxo
bT5Chy4f/uK/GjQjKHjCw2MS4aYqtKD3nnq0gocJhu0fg6EqoCB5iYd8LWvkhZaN
h+g5s71RbKNx2E9l2m6jtO3szhP+7O5uVkeJ7ZsgQHp2WUsLRWlLj5XDyFn+jlSh
DF/7dQVKN0Vt13nVdvb8hbERwBrbD9WR/M8HoO3M0nXOfuH9NbLJS7LVuhcupobS
L0y+BHxsT20Yweoit5kCwykD8p9/XmzGB/pL8MHnYUQIsfgMI2s+SwfsTrEpzCYY
KgIzPH+uF7dzs81uKcNZib+CRVl+C9MfQQM241kTmW1TVNxovQ2zt7XJ/2Jd0mS0
8MiN4vhcfyijXYiC1v4q3jFsmHcSIXmb/1eFe92fSRKl9eUn00eTHW86Kg8C9pDF
GkZU8zjUzPiaUZTWTjab36J7ZqpYvtC1Wk+rjhpym6vb9DtAArFNuioJcZGCmeyA
p1O5O6jezTlBc5/OHgdDchKjEtaXlYj/vZnQtVRPgYpqF0PzRa7+QUocMcu+7NK/
is8W0vN4XTbcaJ6e0f5xW5VWNy7uXmkUBL0WgtgU0X7eUr+BslEEuxsg/8RCgGVA
k5TxHUUjuUjqpyh5936Uy3t3w7hqRQRXPHtD8Jd01wFPvM1Bhk9NFKcdIV7Rk1pJ
iki/Xg5RaGPY68o166uKD4pNR3ppBRHyijVzfM/8qBDSddkLNV/vKbwDH3L9W0uG
1HCisieOHH9WzMPC/mb0me99+rNe0NxHgyTPSAR+44Zb9eil1ppUYOs68WTEiIfY
HR5x1FC5IQIDIygd1R3IrFZscV94L5+iwfp7+evxi8LfSZplZ+GGgym563+AxcHd
mQOBFcAugAaUz0LzzT6a/mC9pv+q101niqDaqp88FfTGOsW1P3QqoS9IGSrpMf4V
XiLxSsz0wg2AYzspVYHu+a0RJPm9fYRyDoZ8AVbRUm48aqr97SXJXferQtd/BQGb
9tT8U5aJYYmQeW6G7+OhH3l3dV+qrVOOQPqD05chMXL2fk+n5yNoqPoONR6M+whp
MdbxIglI/6cBG6gGK3RGbn7ftcOHEkHwt9486ufit8Fs+aKdrT5oVXZRoThZCIbG
PRIYbPnp3PNBU2ifUoSj/CMHsNrn40PCfDQeJ9z6BBBVi1hjhN38tR8YjVhhBqEr
zhr+Vkw3D7QWmmcnCi7H9szgQe1GeHtJQlgON4sCXfZUuFFlw7zLq5YL+UpKfATg
8oT1C1d2QJd2WVa6yUJUwgSbUdsx0D+V0yErEd0yN6pUCZbQhLVoz8mfGPJjRU+z
NlurdXMKxG4N5Rs+oO7Relsq5CLbE/uRID4XfOEVib4G/ngjvNlChzSRI6mfsok0
1KfSYGZJYTwV413Zqsy7o8bw0uLRMbZoPAvdN/AHH9BxSS8hbWSqh8wr+J83KT+E
nWsnne/THk7LstHQkUERzdQ75QOflqbcg0t1XL4pthIyU5hfsFnb6/GVgij2iYdw
95/mXgHMLP0Tc2qozDnZnM/uaaCBrFUpf6vh099LTi9sOAiE0YWiRWgI1ck59dHU
ckoSIp0+SWc3FSS1GctSVJaGPjaih1vdrQItLLG1HK7UgiE4SrogMX29xDJP4y3X
u2nNyKlz8FQ0GHqgyMkX4c/it4vTFXfTXYy0pnkQf8Z7Ry4PWm129JVIaiwTgCpZ
0ewiW/6oSMVHRFsSdE2zVtQdsVO0UnhX48FoQWAzx8o5NJSpW41Yqfk3x0AGmCuw
4/Zmi3O/Ivyy/zcFNbWrzkHCyTE/EAEz7x6NwM+1hG3vbVKnJm4BjpHkFHmLWUv6
tGTmdM8MV3WC1ekUoKkEKDt5StFrkYsrexCjclZu0X4RnQWL/CPAkqjVnAEgrfPs
C570X6tctGtkPVHP1X+jC1lkmXGDW49Ms+XWpUcXWdCt6NCwlLlY1oBnyYMqmVvR
yCzaDIVNXB58IXQU9pYoRoHDIY2iNdo3GRnqcMK34q7Nto3sYQLHFbDrTEXQbLTU
8KSnJjjpUtlIJBzH9ehO/r23vpMR9w1ez0Fm0cutf3AJiiOtu1lWN7AUvm0HGUJr
T/sZlOwBpxjZ9XFK2gAqZg38XDwribUAZniRHQ+sZ12KlFXgr/3dBrPti45d5A49
wXfQaPlmlUwFap7czWYUAQzQWVsRdbPH83VrkaEv0N8vHBcCnRL2/rFAPnsuN1hS
C7dOyJD36gSGBHAYIHT26OJgzN+t8/z/mm5sXWqyTwbt5VcmlbbaV3+NWL7wrQkE
O6hrUWwbt2zOPDiLFTmkpfbZbuLBzI87kb40X9r/6ViFGjTl/GcQo2GG4+LcnMSY
xkdauy3z3H9mF0L4QypHvg5MfAM0RGrnwrMSjqBB86t1Afd7+alWGgrsqPsIaBku
/xNgE40PZASXUpHRBQh1bCVvqwqgkhNJemSsGFvvfxUh/NrjZVgUP8YIsJbufkYy
pZhM7SfAE5g8T1+VHtwb1UM+qUh05xNlbCSFSG/PI3eEuSGSyI5f/zouqiRBzjgM
eBXK12vwfwhUYXcRGpiIRhKo3uODs7uhqrnkHUXJwPXji+2J58I21xnwHe8jmmFW
L/URYZZ2aW09zzPwaqHj5rwM5BQUYJ5fPAE4ehXnifz8quMhQSkni6R7Y0hpQt+1
IrQdCeFLpl6s78vUOa35AJJNivFT85znmz+PzIWwjy0H+WFTVYQkz0Rx/VcF0N9L
5fV90qeqphnojnVW51lWl6/3eitahGE/YZZ0XewlNC3DZxnHtibZmULYWOUXm060
0qf/KHNb3q71GOVmeBe/A7DNHUJXoFgn0UwACrrtkcpvB1j0AG4+nWLo0byT0MZM
3DF2IJL7bXteeS7Rtf87kXtE2h76DzPxr/z3UxEfKSXaf6zZ+iyvmf4fIpsw0TRO
ksVhcRPmQyOjV1BLixA2djByv6LB03HtENdakz/P8htgldQp7l4+2zEt3n/9wKZO
BArwc4dwKmJEIwm7uqGCwCETu8pI6aRxSNQxwrSbGnjgAJHT4RVagAPqpkFHvmhg
SahaClTSP3FxAnSLZ5NoNc98xtEi951di9oQn96UD7xttPCmawiQIoOSAnjCWWYh
uDFnZHloS/Ol/V1gpvHakPTIUtl+htnEIWIsL/S1wSt7iIWxb+wbxbpQBw4J84HO
kP3JDWeQs8OitnEsAH1Vktyr5X897hs8XbWQj7di9p5Ob9kkO1CVESZiiPFgWENh
U/anpzf2QzjUx4Zo5mST9Qu4CODMU2f9gO81ORYgQqY8yOHMUiIfCkSPBJGmEMhG
02EabS+LuSrYE0xNMKfqDcV5gGwx6qy84KTUV7POgTLJMVnBxVlhym+I7257biYP
gudUmurvja2s2SDWVpy+JcBJthR8GUq6XHyxNoZqGXHq5pWQtRsR7N6ki0tjbWae
yi3sBrO8jf1avatE3s7t1sp+P+eyyYLoQvK5feleGS3KyDbz5QnUesrMMZGO6hBy
1zQFN4zxR6TyyIaAcdcMymzvVewlVQI/7b7LclexYUabJnlcCZfMNaD+/vuOMZ7g
CVHuExJ3OJHin1Fqv+aQR0H6jhegYvVx0GifMjXvaTNSyu1If4ydWsYTHBLFvnqO
MZV3vubK4hdHS88SpEmcv5cy/xPo3PHfUvhYUAeC+/OAoylZUnnh4ObGw5HP18Q6
JrYSVHjuEzH5SjL2lAksOxlkn9+SgDn2+dS9uqvFc8hcLZuXuicF/0MQPx/K/qn3
Q8sh6sLLZap2JZh2FjZT6EPAuD/+H0rs1GDugmSgIjN0KGd3yIi3BrcqUgf16+vw
2ZrJ6u0dl79WiAg25+oWcowqQdQJfomEOFucBDPTqe6Cbr5oaJervDqeFbblRSIK
Rp9ONByWiDQswIb6321e18S7GUf6hVRtKUsUpufmhg9Q6Xpb4eHH6tZ1Fxvxu9MB
vNycRXxnZAm9EUECrjwfHV5DSGrxRsyG1IrL6hgaAT395vEDq70f5p+gwysAXC6v
psRk97WH8N4Wli+Zek2Gx7SFq9hgANue9cW1tJ3Ib89fRsgEeFbqups33dT0jPIt
Y0z5mLi+NZV0fML5fHjgZqcAr8OMZ3eWDLHgzNiTdbhyN/rXvDGMXehlv0dTEiCg
kJ25jYn4UsbB3b/JlH+JMYcnYSsQbv+JDDETeO7LM7gt1voJlPLnUOTqe+/bmQli
w8YaCmpgzvPgGIGVUQHLKYZH0GdUwiDocL8gUMYNTWWVOeXlCGltXTwd6CmoUV80
yUQCIjjm2cjzYweyLzUw3XjkqOqoFOmwzvblVVgAjn/AmTlg+Omr/Lir1akC8E7R
dlliri+8wXT3H+6b/468YCG2BeXMEAkU0YyKScF6PjyaKKuryDN4STs9cMNsd4RV
nRVpKrHJMOnIIhle+rruAMBtxnt6KNNYWUAMntH5cbrk6w57zzj6xqX6hS7sGSRL
t+LGEEKeUPrq1PBRlzPK7tfFxv1XTOq8vrOsLJF7W6Yz5X+lVaKn4W5WuwCB1T58
/3OYvGtfh+PydNCgjvs5ydmT20j5bcDtdmKSuxA5TRfJalybL9c+W0+9X2vrKUuo
f7cz/Y++jxWqffi5ly8mJC0jwcTj/8Wci8JYiEg/ccsG9hpfHEED5LuQa+58Iopm
e/kVAvjR2oF4W5LMdRUaTrSxv8h727lM5mi4lTUfhSyZJwHFNRk1z9yFEBJsEO1y
TqhDy1ocuMY3FgHh2M/W9qg3EevY0F5MGgRwD9+p0cKtGANhMRCGIhhdZ9tnwyJt
cInPjwXeWXS6vxGl4w7UbDjJw7rF99xlrFczzzXrqEdBAX8Qw9knuW7+o8ID1HWJ
PQ3vrJ0/bEoaB4mM55faTctj4ufaRxiQGkSaeUlxAQQf894L5HwwaNXeRe5neGGD
eGDq7ERafFGN0ZQdfBWwHNCpZhsI+3J4zmpcVipu3BIYn56i06rufiRu/R8FOvkd
81p2IBV1w6CLAnc8a4AALMbJnFTnly6mM5uDX23LeyouTIBocuCIrnz0HdRT/aGg
jkdbbO59ZafmJsixzScY0OoaWLk34atnKWRwHpuqolTI6tmTDu2yDwebgBWg71nY
QpkUNfMaTE+BzHVDVEH04DQ7FuWZFT0v8MTMN7OwYmtSZbCgrrGmyDm6/ucsJn7d
MgdrlbZ6hGS/FHGrFpf/4Knwj2sFcpQj6lQCYnjgfBoWBAwKD6RZg9lx0agy/nl1
5hGs62k6dnQ8n1eAAr5hqKxZzll56p0IoiDPxOKAilfkjOwez/VGdhq0q+wiYh7s
NJkal6k0Yr/cKqK5/iItwX6B5Gvlfv03OzckBDB5tzJ/OxKRDcBrJY7Qc3Kto1EG
TQawjdgFdl6aMlN+dWQOCJD42rIgExHHmvfWxJxObviPHs/VcD9LKv38LayTWIJP
i6NMmCB7h4OkW58bDOtduKyGJfI8MEeMVGXtEh0fkC71QtAsuZIcb3BRFG44sX9Q
NM/hu3Op9NprprzCfDm80d3HLZ3z4+vfBNHveGZQu0K4DZMxcxc7JwM/KFqW5ayA
0T032CPoCdshL8tJG5ir0RH12MXmKwAZPvWjSB0p1zxwhk/flLsvWo4qi8B08Noa
OPy2BCmI+D1u+JQUhGpx6v/w8R3dQnW3qllGRIOzUmfmGJLRMsxgnSc4Qn/eCZ2z
94doNXbIa0vXrcydyBqjNKizB+100Eqe5V+78q5OIWXuImZ9QUZuXpCfu7Gkt4pV
aJIptuf7K+kFTRj/yQwOvkqzFGYAAzNjSSCcYXtlnu6vxqniPT+uDU9pCHFgnSHn
SwV1hIKTnUFlTRUclZmCDK6vAKJJe4kyr/PLtk0EhPnqNYyXLfzKIjUS7DeG4Qyf
lk6wlnjqAF+Q6Rnhui7ZE34gk05VpmD81ARLNsYKJcEj89tEMhWOsYBQ/MXiLsfK
nNq7LacXSE0/UiC3N3me0h71wNYo4xm/ZEhs92WEV/3NwmwZJOk/EL4jmSZXeI4c
1HLHkPH0zPvmKlSPThi/MCXqUIGX22VM4QWbSCQ/D26SayPTtLMGojfPxt2yt4Be
YVH1WSv5I/bJJDTfg6+zrjUenC++2cRSMgCdYcKTXqfQqE0WG+hqBr/HZTqGt4hK
2PRwXmuTcJPmiSJOzZ3mzhe2CF2mdOVG//0U9ZBJPSBAyk+3NDC6LAcr/+gqgMey
0igV+e/Shse4WRaUeX+Xq/5sNzPz429wKvl6Zpkr1C62PsKyEQmlTRS/pYn72H7x
P68BQRuxkFu4XCMCnCTEvk2guPDBl2WcJuwD0D5PQf5RtrvjGXf5O7SvyJ2Gkrto
Tzrady9tV/WX1bz7KfDqISz/YXAYQ11iw7dpV9cIYPfGWIkFhZYV69/kLaIblu4Q
dc/zc8JQSea+Bpk6Y9Ch/EoLBZIDSDSELQ2O8llRrTm1hFmsn96dc+brbVdTZs1O
hcHf4dz0ggB4pYxGr+tnLJ+A/jeRddfi6dvEyvrPTgTcb6fBG7co/iiZdm5VgQxn
lR6Djby7zafGKtvev+OFiX83zlNY5ybTjkOx+DMA28OOL8nUFzHLqyMZF3ulOZJG
ubjFKq+3ao1FEALV4t/zpI03BTyF3022V53wuVQnK2341k6r6CsfnzLVx67p6qf4
riynqk4w8kKO3a13ay1XXzxDTriJubUe/qBiTw9OBSQPzE5356V2mgpgl75zEvau
ug+cILP6Ls+1DsNxEAcyNJuf4PVPGYoD9cvRzfxDN9abi8x56OXZxktB7CTWthLl
maqzGIN4FRkYht8GkeftkmyU0CZshrt6cR9c6N+Zj3jGJgOrk3FFyDCTWL0RONNj
/dArTYAY6Rc+4kuCRz7kyJ1I2uIjen/GdZtf0MYkrOSINENgulhUMkEbaQ2Aw7D7
WDRsDrrKR80rL/Zu5p38A7mlWEz0U+aGghmgOfkw3fYYhfFs/4nA4ZciR1Khk/bc
Rd/wVEdWmZxlWG2FMrx0h0Qj+2LXK0cACfAbGLXbXRTjw6hCyijJlwi9niNvZobK
tWtFFGfBfLi95n1Hc9rkAJxZSpwDksxfgySwprYhS55AtJ46g5HqoYIzEXOrETPa
8S7djny6beI2RIbs1a7pSOgiPWsovgtBM2bxjH7LpqQHyei0dIibBNFYBOoqBWMr
aUM71IJT/d8VovjhOn+d3hWp27X4QQj1OnXg3kckflAjzE5p88LRRzmjXtrVzfMk
JJzQdMZg7W/QR1Sg7vJXqpl3Pig8D8YorgWKCjg6FHiCXPKQbqmLmz7W1PBM3Dk8
etZL2fHMyr1YRM+UztxehLQ58QHdKwaPiMurUs8uKHMq1dWbOb5FQK36yaBR0vk3
KxfVoLUDqfXOpXDiHxjtSn7u811C+VH89Smpqur/nOdBN8die2d+c7E08XhuW2fo
OtfAedXn1NdoniSm4brGhtlX4RR8nuf5NI/tl7J8YYXZRCdhE4fTXasD7WzDObgg
ScmwleYRKw0LL7bqkcZoplf0Ej1ycKnu+ro6Kda6W0xlpTGwVdvRg+Dpnkwx+KiK
TsasXkT/TSZsqKljLv83HwtMbez4gY5aSGNlHyWJ4ORtSPLi3mExr1HPPYhZuoMr
xZBNoWGtqrGkC9hSXLvBFBpTqOqkvuM1oPg1CjfI2R6VHNc4sHpGe/boQmrpQJmh
XBlT2O4GKY2IFtRBxo4kNJnhJ/3S7G5UqXWjHqLpdKpLkzscgaJPQD+cbAFIcN3a
3H1Gz1/IG1/zn1MvMXxJ//HXMUMjgo8DtW5qU8wln2ckvkSY1jDWDQN4AD3LYoFk
9DIE03wKCzA98HScIhL/fw8ZWuU44npGe28si5tG3CY0xqqvk4lCY6t/wD3C2a1g
bLqo08Agt/OjgyZj6e7qQvrCVmBw/Aozqn3E//l0AxrqvmACKek3fHgL6f3/pwX3
Fw5EI0KKd4JaLtKzblkXSz3gSt3B/jKHENjTW3/HiQ7ZGQEH/PsxSO9i9Mky15WN
bZY74xidFQsZ7DWZ0+Jkggk5JCU/bWWDOlwhiBOCIhbeapq7BMlJ0l45hf1kzuH9
Q4+NQkE43CfUBl7b2JYKtgROsBZcm6jqC4sRsbdU2+dbc8CoUeKj/T04yKHtlEHl
p4JverPVlPFDxzQ3qg9V/L+mUrVnxaqTV0eQdOuDWV/h77DzKTpOcM2N6nv+tBD/
7+RoB1ayzs0fkvu0RTrPTq4VbFaOIZ2IlIGeKljp5/vLvNnEvR0ZYkFRWMoGnnsy
EEtI7OCpkTgYkVDVLj1Gb4KpIREEoxjpY5n2jyNkvR+VlRvfG7BQRG+aV+ix0SYj
ML6HBwY1f/A7UE5U4H6viwbNr2dbpE/ACss6A2dzWjxpAyRfqlSUoZF5+cpLT8FV
6Sg9caK8XrD6PMjcoUoZWMD2EZqj0ObnnLXaMHECAxUOyyVIKqsGyFf1RnFKN3RR
6xWtel2vWEfglwXvxzybSdwcc6ErB4lGTDrkPMapuL8r7tYhSX3HZTT5cd6em5pJ
7eXMwvx9BJveCBfad42a1jKZMpppyiryXWLr1Icpz0bDgkZ+jSzq5+fEaflANy41
8OuKt7fSVQB6BdYJjMFmJSt7pHF3JDU5DZOv9/zsVjCaVba7HCi7pg7DiVj4VtSA
UakeMzXSSmSo9MfcmSlpK7ueIDrc3wFfdRBGKz01HeYBgavGTNvhI/fuKD6iazln
pcOLrTBbGMl4oXRZYWHhVUH6wHoUAcWRnFb5h9BN9aBu26OxW86/cWVOJnBFuIzA
Bg0NzeOaqEc/8kzzuzc1fxS16JAlzG0btb/obTiuZa1leIY26t6wfQnYCaZGNao9
WzVpVTNwFIqtxxAed6/LKkIZY45fgSZHNqQziRQkIYPLjgbW804NxoaiFrz1fbPQ
wPuqa3AUpPLXik5wDb/zxjDrHfvCAj8Dgnv20eHRv5zkGi79NJWJsFSBGWybHDRi
2Q9eGEg0+iARUfyN+itD+KDYB/d47ZiUW7mufptiyhGbIR3CG0pPqLmhEQKeKNIE
7zNjDqAoyqm+YQuGSL+qSfz/HRsqhQdyWsbzLrECuTiEJCnyOVsyHSQ5YyUkFXuP
p4YmJIyRam4JSoULzNAsRPlzbtpXLn95tnyT9BUzMRRDV0dP3GQjneR0YlzZpArY
PgKHqOwGor2y2IqYDgidttuk5ubaS+fx+pfyfkThsVmsLFcev0s5KP3TOlVhEciI
8PvIh9qxziznW67VEId806TvKdYJc7dR6m6GdXqXZ/4F0mvXz8rdOVUZcMtrRvia
kwJdDA7voKPYLH8GcuPQLb64ipTNJDhJ/48j3F0tORnIzT09/RWMgp9fHacPFwLj
f+sfMQn7FiSjaCDkY6z6HUBZB9L/HE9aCuLeGfiXjAPCbX4zfyRxmR4X7fP/LQwu
jP50rtdSxWygrFtIQXcEm6PVr9gwBlmEK+xK82xztE+epGTxbqCg4EUFCc/LjMjj
U4vXUQdKpo6FJHHAGgn1oHfN7Rtr/02xsaJIAcs0qt5uE27BaohSuTAhlivD5Jy5
lWFDdKlkC/ad1x/6wL60iSBZreMzmfVzdHNSiS79XNy6b1nTVNX5of/9wbqIvKrt
WvLuohvztN6xsKrkMjb5SvY6e5RtyzUvDuQrlBbmJccPtbKmABDjm8R7gahBWRNd
fKRPiwUIdhgvWAE9ZFnghpEApcpgq7eGS4UKxh1pZ1WLFOc/2u8jRUtqe0xD8/ww
69NKQGVZLQv4Dv+UODmBR1ZnKHCryuSyJ+f5yGYsMhXMO8bOlmx5GGh7x+JDsTyq
4wcusxCczWSEzTMbImEtjkneGUbIipa3+DDpjOPUwUypVZNXPMy91Re7sot42esc
d1r36jfkUInZJR1xq1a6grma6J/kEpWufjjKtAPKSGWwGhAbAdb7xow5zq1pDoKH
2U+Nl/PjdbWV5vyqjyag7rLU97TEZFRvL+UKA5bTUoh6ExU+8dXTVPbgHjYjY1FN
vAMNYy07041IvBg5Uagpkl1GZDEKPEg97g/5QA98l2STomWI3s6x/FydngUjzNb2
bWcgGuCQam05gw3e7SDxcvD5bABWWS4OILZI+vkyOWWXN/+N0zNo8H8DRbx+nbDt
bLUgGa1oR4D2cB/vCkPJdCDDyTDKiNiB+DZjDds8AqiyB9WR3d775hMPzourwQjH
OWqYVX+YueYEaPSBD0AJIGhNQsJPvDFGM8U7Q5FYTWtcXkb7eoQtdBhR+R0L9QE2
SFO5a5moD2k3yipVz6eqJhV5FF4bgwcE1JC9YEXPprnDDAJXUJ8lBxtt7I2jrB+a
S38IsQUFLYFvo27A9Aadq2zmem12xavVLSMXApxVR57JEuw4804osT23G3xayBfP
K+YcmwQHIuWaDvm41231uDbRR9YpyKfuRv4weedopR2oKDcyztWNb+wwL8PUq74h
vY0wB+TtulPPPPsYYkojsnE0V82kxu47QgphbKDE9e/E4Oo82P45M3AZe28ZKYrN
r7wSOrB2SHozgn8iVcrR/wjhuY9UlWqfCmzttQwkBM6FbK7CWDNm8lxDMHE+WSXh
4VY4zLnXkof40Qxt6HYh5++mVm4HsERntm5ws2v/xGdJJ0QVGgec2K33/hRZ34/b
I3PooVPLQJFkZiVmUdI63VR3Dl8/9QUtDvQBiGDXbitbqLfTZgJfRVk93bf8Yz+p
0UYyF6iGTCIU45JzzPXCUhV04mGUQ+4ryFSMc+YElq6Mv2igZRm6KQdESAaPZEg6
S+sfn1pzKz/MGndx64BYKv90WQNtboIs3FRo0sCk+27kJrYWz4N4Dk/ixCe38ucH
RjxsVDuuDdAtymNvdJtsqENLY4+EtKlmXQV2FUyaDu7UiXlTwDOlfGosn6n6ny23
2aWhj5mGOAvGvsEcfdIKyOn69lQ75NuXeU+toHh7PWIEQTS761M33AQ6WF82h/EY
9deC1SoLiI9gObxKNds6kdhhaEAoxCPw3hiLnH2uH4UdwW4UDbt6iEEk2iYsfdZQ
Qim0pVHTdoUBQB9/jTEwrMwLmkRRuSiqTSxHueRF7QELi0KbfXFBlVv7ovuvWfQp
KXOn8AyDgL9I4AeGiTKz3FdfWZdALsBhA8X6MthyttZyf2ORzo3XvW7qjbwnfJ5o
bdWsGUySN7iGdRW8T/XVCB0nEINxqDx4ptesp/drhiR7Ol6v4wE4YK4nvIWNSlmz
MfOjs5VHC38FnOqwF3h8KBV25DlNJx/3n9t4NY5JsDHDidYfNWrwXUXjip/1LYFz
lju7i/Mg9SPoFyOcMtnBRLKoxj1PlaleGs8dAn+cETZ/aYbhfRcqX2h2TAWP3GTC
Zzli1XmcZWn5HWvlkLFrlGSY71ViF6Vu0JUsf7pMKLX6NruBlkd6fO+VzLUzNfEh
Tf3plMcJ3E8mUX0zDdCjAGNkNT98gmzQFMq0qmvi9SNRXGGEFx6rbbP6B8miG2NG
i3zyQIuUaEBrbDGwqQTUtcEq3pZ1zc9Q51cC1LbLeNyXQikY8oAHyC4wjhQzYC4N
kTu/cmSieYVGuwJJTo5ysRygfkPo/MM4av0sluOpoH/eyjDCcU7qFo+N6WhlUW/v
s5cAtCcvjb8PvmPycfflCKNmGhlawJve1F2mNoU1lPQZHaXF3QeingMvkReA3nV5
Vhb9/Y0NNromggl2LIERvcUYJwdHuQ874MnuvvSbt4Qq2lIBcd7qXRaHnyXa9TDB
BpFQc++I5qAM7NtyBLrLaTAsejB5uHNUFhKmm8vCYzaG7jsu485bl8WtHFVc1P5o
cZd+F8masBLx4SdY3Th24NUTyyH2VltFS096DhyN/jwg39sTkCEnPGDvPEaFVgdY
0SClBJAjhjrw5Beg2b/YzMAS9jrzIbsSS7YKP1slP2OlDro2FsVPcRrW2h98Hgjv
6Du/LbXdYjvaGSqhW/ZTGjGQ8RgMo9FozE7jcFE7vazIdIKyiFKIdXB7NiOpJqMf
3oknMg1CXzkVSuzPaXCqsl2JalTB63GrqMa61NQXXcwqkXTDYZIAZkBU/WUAYLv2
3hKkjlIiYOtBbqv6VnikQWYYHGqsuvAOiLkm8amBh96F91hkqHeTKZPZzv5Klnsv
MwTafAD9x33SdNOSsw6E0pSysaYTbyewcQBm1N9aICsPoO8uoiRbOBNvU8UVahXb
+6Q1ebWilS9PoJ8MbDsaitDXThRM9yCAk86tQWWRUETpP+nga6jEEGx1jomzCmoF
4CcBYQQfLE1CovKsubCff3MoIt7xM82QSPpSt+IhR3Nr7FniNKHnyR5RN6QUgU69
WRHst/KfBg5otuaHliMYaQ8ghdNBBZcqFbDRT+UhySo/lxgkqwcVwNQZOdpQ8RVI
04XvzwHadEGy1aN2T1wUTcgey/kFmpoPVo7/cDLE6+47Sx8oRAWQ+23Xz06T1B3v
hZ2eWcQ501Jcf2Aql2wVTnsz+n+tZ89q9wvBDoZLIuU7vEvARyqmkNMASKDCb/zh
X45WBpCMISb94Pl2rRlFSNhs/z7Ljm9h58bMIDL4is36IpahuW5g/42xF9VHqWmd
tIe6aO8rVTxGrU6bjiG09EVn3++AVYYyHeijB6YTxOCF2QLxDJwq/pE9pxIlGhXj
i9IuX4/nB1aG0qsmzsADFUbLQa20zuo+RCZEn4bEh3tNUybduoBvyH2MMf8LZpjQ
WGizrTM88PuGjiZCltUv2QIGRWmVX7KGyA/MFTF63WNWv8tl1PBpOUI4I+znvVAi
n6Vvh0vp87APo+i9Mg+7feuM5LRX6R6tRu6fmpLl9r/uBRab4LlMaU1JY+KnggAm
GyTkjo6en3YIbTS3aqO7iQqtTkCorSwdwh6iSoH1t5VaGIHrxbiDXhSY+kI6cA4g
+YDqvLx1FuifpGvscSkFEOEA/Z1cmAnmqb+ldaLiCGILY7rd4REkLO/erkGY2BSu
wKGbBD4SRA+f1WGXRnjrbPAn7/28g9oBKj0pUEMgpvRzohbgm4tLCWuVkctZ6SCE
qI29oiwv4BdXnZmaFLrq2qQxMDF11COc71XaaD/aFaXx7SL+R+u+bWln2VQI9nHb
zHTT+vaRCwTII0x6aLr0EhQa0D4QvvDxMuXZwB0svhPiydhGZYImdiKSPTZTz5vJ
p/qsFnNW59kJPoSXk3cXbD9r0kTOJ5m/9HDQCzXVfNoB6BF+st926Clzbf4A8AJp
qMmOlHcbx8s4il1r9qpHa1CR1T+DT3Dy+nrnFooozL8FARvwz8zqacCctmkJRWlC
OG/MhWz38zkx3flEwXhabC69ftwS54naLTILfySEXqqlgadZKeyZfZaFJ9ERplIz
vyT0Q8pxlPUhDn9m6BmxW7N5nmNPNVhrVOg79krzY8vyeWtxyKlmoh1FqTEpuRvc
dWGVpFaK5+lUXYBRIyfkktCOSRckXBiJMXzp/UJba4yFwVbvymV8Wy+k7raSeusx
6K+BHR3k3MMGjb04UNufrZcfYp12w7XdLFSKf98wFgcoNSPtVdxnBYwV7fjsJock
GEoJ/j7EIZutfHgFhTP3ORFs/GW/wYHhEceIJt1ORfyiJDHdyg0LF6EwTYMAyo4V
WqQTdQ9XtjQ8hlf1/StRRkx4/eYw5N23FHVZHxU02IpcCaC0o3psb2BJa0CdSAao
qvR3N3aBL+8DVaLhIPsJDZA+jGbRKsnAMmQe2tD1+BspU9oE130v6vxk1Vnc0oGD
hA84jPhtcDJTwooYEYHtVLq9UPFadx9Fl/rpyF/oUACSnjJiS4E40x+pnAwmYApd
IqquwX7XtncOxa2VkT2LjvHi2Isf0L8zMzXqUWZ9UsMKeZj+lox8+cl6/j8SG3Lp
h2BKEu3Zx1oRUS+fo3qbzLrJ/NtLKkA1dsC1ocMHjlddo/LWovvAb8CWBXgfTeic
dgtDH10VhcdZBKbeyt7/OOU00d7F9Hyeaqf8weZrkeZXNSMnACEdoI2mX7WNIpQY
P1/5AO1ZXdvTlZzQgMRbOQoWj5J9Z677rOdts0tJY1K9+/nDvRzQe5hTBwmp6trp
J+3LxTyxgyCkriQ0nEvzN4fzkj4RUkUeWpDDgIUkJpS4BvEfzgGKySIT+YWRU9GM
ul/uu0QfsJ52Ut/Jcckh3O8ycZFMv7vDi3+ZQp0BM2AvQ4ob19fGTcH6vkPA4lxp
BGNXd5PY9hRS5i5hkVSN8rhirz/VxCWSywvOcIbdn7Eq0oG1ipEF9FhRaapoanoj
JZbAR3QnNkIY59U9+ZxU5lxfYtjXKdqmd+XfIoPLG1cowm4TYe5VsW+hdoSw4MNN
D4109XQcxP1B75L7OEtPCAWbZrbNw28RjnqlqPngMNbGN+CnPBj4jTUvWesNkldE
hFqPpe7TfMPJHp1E7EQoYXfHhwz1yWIitCktOAi4HLnRD+32X9oz0YvtcctRzpe2
OBHHheptej9zqjFZPrszQjrRCsMVWQW6ogVva33apA2GkSSDjvvWxAwg5ETrZmkp
4h6PZ2CE2rvmUYzai1GB6FTZN6pAl+J4jvnuBY6AvItBtBhKSNlnZep1eERBh0XU
NTPZX9IqgKetsVHJcIXEcvciMFN4stCEKGCin4UV5FzIeNerwmbdscg3C+gmvH31
kcSPgXD/yqplB1cTDgOtwYgvf3nhn+XP/tMY3Of9r+wLVyxmMFWk51TXhrQzV3Cc
vKLnderBZuBEj2BDIDFhJH/bvnJmYg4y0mOPUXx7tpKlIMJ+BffcyqDKgPVhez9e
z7fmyqlsNSqZuDNbgK7cp32b4DRL5nL8EWfFf1G2zqwvfyKJJM8KDdEQVaUY0ze4
MQOzCOl4geSVA3cH0VGNrGW+KUzASAWGvYP3i5lQHKssNrx2pfEOaOI90eCfRAeb
wx6MahoDD1J7VJ9kM8WPvqQtrvVL9ZU18oFw6ehjAHV5XuIqHt+n+j+OlJTT+8xr
FpeAIJd0iwe5wP/H1W5zdMGveG1hy3dVE2m5Yi5XmzszKPHht273fUnjSa1Bsg7E
yz9VihBKG/u0zybwObYS2XGZz0RAIkvqORfJdSw0o0hn95ISeDccP52BzrnmS/Dg
lGiNZ7G6/2VQZtQ/viGbKg28AxUcJKsX0tIRIEjzVnCGrUYHMrKpfzBD+kbq4Lfg
UJMwii+H787jRXFcMQ6vMrZiKwfu6iipyyg+eVibvGFCpZe5z5JfqlO9DInr1gCL
ZKZihwKG4VPS/Je7OC6zzbi0vz+UjRJ1J5vHlHdu3Mb6U+QOZA7nk0wPDERzmJJ4
6u+9vL5/HqmdBFHILNNzKRKYbdz1NA0TrPPnnW+FVKP9sZf4aRnDcQDilHHRjipe
rhsu22vzl3reorUVF4+emoKJzaPiJ5Eto9luocnEPpRVTAhQJfaxOQgE8CrkpCB0
bwILgHMHQfzdBY3a2jCJekl+vZaxCKVDueCM8hR18pXNZQVxVYLmJ9Y94myGwUd8
h0SfDTfLMTZbu36haCyHrqaA7GK/HR5uDXtUhLk9Bg7J0qi0cTZwv7aE0IeKzwAq
B6YOvGpD7RT4l0AL2fHbMYSFq8hUi4+/0OWuwC653/yCT+agQAvgmUXULugn8Qdj
V3g3sFXj7KUGaej5BxaSQllLt1VKaRGZ+UIE5bhpLKSc7MhMTlAs1MP2KZ2rxBYH
8Fu+bPqgSWrHVmRsBHHvxAVz5LBRVA6toGB5GpYxmp469EejxvHqzzoLAs7dQUoI
Bu2VW2nOSsij6Dk6JwuH6jgY4SwqiCPqDZddws+EZavm0BEsFRKhMjPCaKXNNY1e
dtBcLgtCy/o7cfu6XJR68EEJXNpSymsw3ieK/1fpjgG5omjEjuUuPd6Odczcms2q
tcestVi1eAZDKxByE7dErYLqoh8ZMzcwMXzhKLO41NXXzyKeUqy16wMeYpX7hlnx
QilkZT4IJq0QuSGKypnea4bro0CMkQJdrwEH7WUxgcL8L+E/X/reBmqlJP6U5LsG
3qX+MVY4roMSzz7VP2PuCxYq0AzHZJbSYy/JNM1lB1eAAAdKB3OA3biVGzhSya80
wJlaIiuQsXomVVUF6yxlwPapLzGWSoNX6yevWZiz8FMLldUYULlaZ86ApxI5bzB1
Ahl9M6d0DdxPZHAui2VxfMQ3R82G7TXIicrfWnj/6M6urIDm3uGtjlLV7fkX/xci
L9Bg69wRURlXEIvLrZ7WgVN820nyFVzkb4WA+4BsRf+upLstMONFJzx1/VuaoJwq
zU2xBDGuOEeE8+1nTJZyBGliNKZN9KeN/mYCjOJljldydcfn4IGDk7IewhHoNGBu
KJPWbb3TgHoTftWCD4eKuiP4rc8HAet/0W9XYng90nQSJ/AD/53JRGFWm9NizMZR
ioGM6Fm8s9FvmAmssrasQBUBF8Jwt+Eq/qOuk/MFe4Tcejg7cTswL3ZaZ5XOBk72
Iy64xjn1SF4hkI0cSbbJDNuLOXTEVQ4sqPRlKvsSdFIQuFxc09CzVHZhDfRcMfGq
689/R+7gwAjQhdB+Pqdu8eNBKbzKK5YBhL1yB3cvWeaAkLjnghd+Y+9JA8uUFSj9
xqOVFAN8wNrAj0LC68Y9qCSDU06jefQRwNZ9hwla4urGm8309Jsi4PJg6StAy3E8
TXcvM5YYJIoX8PpT0+X2h7v+gZbxBWuV30X1o+PUgbsWNjNMSxrqX7vup/2PeRCt
oFslLvKNZppx5YkZvfqoISyilDLXDGDbdYQtM9n1RpmnInIsEfeQeiewjcsFrotn
YuruM73v9Up6344Bj8FLw5hoA7pqV1nLL63P4EV8RSjrttCuLsSUYV3Tacsca9p5
yJKQ5tI+/M5Lt++LLS2m8IB+0tGVEHcyp+1LszXdDGE/9G0dBgPyzCXp6PE/xB32
CsA9C/RJ6yQzLa551dQ1+OdiTWb6gxG2HZX7FFcW2g8+7OJAWqVccT92iBFYEHla
8fcvmS9GM92M6Cz3ADi9EXfPWmy0RPHFMrcxhSwsMj4/V27i0eipH4bdEIE5AE+X
qarQO6QZwNvax94dGftt7DM/8KNGMQTPJwA/1BCsby6pkdeOPtecuC7ORiZij1R0
IZ+KbGLJOb//BLiuRlIiPSAN1mV5+sii9F+ktEmarNoOI/xEtUIodz2MQFOE1qLF
IStr4IPIXBtTV7ujueTevzmeBfP48oy0yxciVesOp0T6AYp4dGUGcEuYUuD0c49B
i9BwkUMpJAHSgaf6ebun28oWcEZGELCsiJ9E3DvucRdo1pcx54Vi7fJ2idXDeC81
ZRMEsKCowxxAvp1xN9Ssw1Yge7TJRU4HPC3PMYvrhyIPOx/3QpfrxClT+fIoeltb
cB69R0xwrvcpZK2zFaHhabPtYJ4FaY2jjjBYMDmFsSV5HQu2SZ4oY1R71hiGO8c8
VmWGRPD4Ca3cjDWWAcy9jaZwh3V8Du/+t43wQCTi2RPB7vNWZwAg0FK3RIbOh61R
7qixTbZb3SJINB2wcg7LoOmHx3+OWOaK7lgbi+3vY7pLnwgMxDR6GFqWoImBd70s
HsOjqFjkBycYOiM0A1eCqajiw7YrW1F0Ps/OBfFeHEil9PHtdccWK2iGnHbf+bhW
01AUEW/UDm/39/gPHeycA2e40BMm/JuazReHFIQuOrhQcRR/6xbwPtcpIcRx4YkM
TDTWmR6BnKr+4muQ35anwS1XTrX6o9QOFujAIjXWOJl4VHU244LgxCqevUv2rVx7
vbIBStCFklZ83ZOmoFJUdgUSwQS5G99YPwOWtRgp4sOXbJeYUpkzMSdy1AFLnlUQ
a0gAhgL8oBYmggxQF36WAz6sLRsBNYkQATtEGW3HTyu0PXZ4tjKTheNGlaK2c7NH
YeIpna2VcDuqn0yvFOHMD59y9M2GXkDQbWCOoc5JtQtJ/VL1Rvh1xZ+y56Pnf3Ae
z/kOwlvdntXwBPnvDK90HTirwFwWzYXhYp1gjwhSVBVLiCm2v+30d7Tmr622Aw6I
lRu4cXm2zCrCGb9PGtKCMETjyqZ2QGS3JPgwPCId+CakOIloC20kakCu92owc7bP
K8+BOswz0nz0TajO96x1HK1CKRQgb0MPnGblKMrslhgEcKb7QrRWRu3gM1Xu+QeI
MiJVOI+6lPIQQ4xl60gNXNbaJ9bMZo/wlUDFzSm2N9FLKNfnOvBJ1xm7JKYUr0ea
/UUTg0IPy1zjEJOelqH2Y5WLpcABUWR0g3TjBiFDkhJyZsEBBkXPcUolqfKXk944
DkjEny4PQC8pqTZd1nQsMU8nfPYSS680FTezK3EnW8oOyAI9abFuUjp1qVJTpls7
WbBW5MmXc5S4O6F/tJA7hvAHcoVCGCKQk8s+jlkfFTQUwi21lYr4z5ybT4g5rGIH
X9JezS/oousDZ96u2K+1P3u9gX2K1rFZESJAhsBRWeB8OEjknULuEFVASfMByki5
etW4sPSBigV6bAOEQEa7mUzX+HV3YJlImAYdgpjpWSix4TuMWmLugBRQte8mFOyG
mIywL46rdtOkT8qUcXmrj2T5r78rCiWW3PMOerkmVDc4yir5q3+Kxc79e4W5FDy7
Cl1wtjJe1i2MU4TlI40Vh7cKzqt4R4U8r/yE9o7huAVWiEB85nWVxvRo7AWb2AB+
/0/0sf58+feyVtXvDD8hmERPaQO86rppS+4qUMCJZVbLuQmwdDvbqXCgEUnzy0Dq
GWng8tYMl+Jx1JhFjeHz+91L1479x2OXpdh46Y63qQ4VMh8QNod77MRwsa/ImVls
hf+nZnjzJ1xppSr+UryK5N3cV+QL+vnpV9NBSZmY3D/Dmo+FrOvRPwkSd+c2dieC
W6l0FpHq+Iub/fX8wBpw8Bcln+96OsEb6EoNnTWAStmlSrxVLRYww6lOZH69ZXZj
H+P3moerGLNgHNbsSnrlKENvTR+tmH9yCK36EiwTD70FFbzA9A0DkMOjzo9Ib0Hz
vl8s/a4m6P/Qh6O+KIivp1oA9MWwe07qP01QxKCANhiQbjCStBl1jVeZkC/68V0H
oFfZZ0YR8LEsLAsSEXkanqJ/NXulnefDjzKGNkqam/v9PnRLOUrr66qWgRwNeviO
tjugeMv3mG4xos2JOz/MEBTP7o55EnPU0WYjOopzakg1U61NEkn4fr/cSm5h14Ur
IkXuPjfL/GzelTk/RwsfqrDE9ailqM72c5P97elOaENv2YzK7RqcdN3DDs4BtDPk
U/TTQCOqB+u83UdVdDQbstjBfJPqW9AvzW8vnvsI5Wig2zWoAwTav6L7PKzABFbU
tNU+MoZeaTBKWLWfjDShjz8iYj8gmyL44Q7Vq3tmaPadKl9T87OfT6zrpCw0kA9M
8x311VLI+lRTc/WK18UEW1bimUzRZNpxfZSRieyKNT83pdMSC4ANnXxQ6MTW7hpP
d7wc0q92LdwXTtXt+wgBuHbJ8MDq3FDwtaz4rg050NwU+xVIa8t+Z4D9we8fAXe6
q4ztQ3MS8Xt5PSkU8vDPJG2QrJFRba3d0lx0UWJMhBwmhYb8CnAmHZ/SIJglV0n+
hatgDz6slwZ4+MKl0Ck5W80gtkaN3pIUb7C+1+UjhATgp8nPylrSQ2jONbIbTumz
XtJiz4UFCeH3heatn8TE0Y+XRJnuk79JwZt4s0TnqMRsswDZR+td/NAdQ093PdKf
5RyjT00WzuM49sW/G6MC4Ygc6XtpFloTkLo3HengZyb0Aa4qXVo6tJXCawEvsX4D
w3FEl3y6TXbPPwmVFrQazYvbZ1Cf5zjBFM4wueOIrc2JV/+873ivOePGmPZ/43Ty
sS3PAy3Name5bAAyfhazwTRtW4bE9RnuyIHKAQ1rKd7Wm34+vnh0ygKztwMRgi8z
FiKKNHz3eL76+ZGiN/fLODYwUOSDcdAcYihrqCH0IrT/aNJsIypo0Nq+ODUQ0su3
LB8HSEEfpw5XQVrgbLiPATnk4RUGFxfK1S5UPRz45CWoF0AsARkeSOLiiHJBz1jX
GgjsuyqmjSnMdWakMsPACA2yM9xKjD2SpWRMpGdd6r6dGkiyvmIJR4F8Zr/9O4bQ
wXJhkwnTHM3rp7cp77oJUC1DLdaItaR/4xKJiX0Du6QYn1PXfFv3tbGLJgjiDOwV
GNcAJNsidmdw2CmwB9prmxOlsFIrt8tzSzBazLQs95Jc7G0mZyTAcGNn7tWJ4XrS
OO/b0Rk09JrcKrV08QioKN2ur6dNNEmeu6ToajE3PLSqgV1c20UX9X2QbSrHEE+3
7MtUZGYnjI6ktxFCNGYSIDFfyKn1oKmNzQxvQ8o2VRBSdXnlXqMBFq7DPrGzeP9f
HX6oRVVTW8i11ZBwfWuS7pARFEYbBb25R6CJRiAb9plz7vUhrzp9b09r/C+hm1Cs
tTkSYQppZ0YLILhZ5c2a9xMG9op+mNvytALIeJWYjRoCdJX7/qURv2k+i0TrwtTp
Hf1rb13gvlRfjp/QboeaKHQSz9x/rwOzM8TVIufHmVroT2gNU7LDKQoTujI2G9QV
QeWVriZ7N1antgKrFgNLq+W4EBd4VRXqUD26f8sCGXHbNLEWzIDYoZ4Vv5rcsYtX
6AvN7V37z4GaWpYp8VpQSS3V8SAX4U251rjvKJT2LmjStFVwpR9yfm17Ezsy07ym
osAFV10IVvHjOd7Il2AIeT0Yp1I7TSOEJiXU7bEwKpWpVEE+15Z8N86u5VJUO8v7
02LA99r1eicIAKBkcAqtkGE3wONhmZQ6+HLoSsZ3Z9sJcqbZL5etJ+K9/yW1a9o9
t0nFYKc62btmbaONfZMam+MjEhjpmRMQ09AMfFKuKi1OgfGCWBFolS1JdWBX/u55
kRAp3dQNrs+3M9944s7eaceAz09uZBWXbGY2VYvhEJ3YWTmPc8x5KXYT5hfHRgVE
DViC+qY/aTR6hig5vUG6s+qWL3y7kn8VI1ZNURtbv5pTAs8V8O7lB3r1Yo8i47Le
dr7u786SNzwC1lVU057n8nGAkysHFJR6sXWlq2j1fzT16Vvu0Qk7C/NsxwNTspim
aLtkSPjF0GMC0LWRciVLqB7PXqVkrG/A5jz6ClX+a8ki5N01wwSiPPZ4tBU5Kyf9
QdEbWl55KjkgGrsyn/NGH0N162XCaPiiz0NXj1Fmdifk7uiBWTndSuKMrcG+Csmk
4GuhDPE4Mr5PvJFFKb97o33ECI3L5ijgcLqKTjGplr6nCIlva0zMafoUcKPhrmQw
FM7lpXa82Ja+sS2TloqXibx8akmx0sFA31ajBIC8U8356t4LtQpSQrSbo1e0h4lQ
4JG5cmHBRL86AbYkgAUi7mPCp1XkbuTKPA7GXTLuuJETbGwpq+63J/pO+DkFuLUU
bYgu9WxcAOEOQk3Y/q+WzpQlimGAgU/E39+vc8pqY7rWD0jbYKUIp5SwBfPX03KT
zCzpwGTBdRNHXCWwFo4fTnazhHUONdvYCDHH/jP5U6/sJjY0c8Ky1rcX2ZbIw2zs
OfgEy9Xv8Mv22bAAdAv2bhu/+s2pndRkGoUyJvo4D4s1KRmbbciOLHoTfsMWhf4M
NdKfdW3DQtyNp8Qe7xHaAAO3L+yUNDjjCiG3x+wKeoWiiQuyUUpXGgZS8Hit7BHM
Xzt2HP6V3fqs4s6Hlbjp4pG+ClhzYUzw2SU/BQ71pRicJPOpzw6IkXcIztvlc28O
FVXNtAWjIliJGwB5D9VegYvQKC9iFsyxN+S4RnH8kPI2vz8OU/tWGC90sh9pj5Oj
z3soQYQjZlZ3oVvYGCwsIwJuNM0t9X3D5rXCUbXwxBmR1MnDttQ3y49CAmryO/PD
CRFZi+stBuSbRVEyqgOI2Ugz/TKG2fz6dcbKyaiBbVpOBF6Ac9Bf0CWKmDJ4Y28Z
/415YmF40AgiA7dy0dWK75MAErD3Vin0NFAY/OFwsMOEtBNb42M6Rx9aOMHv7PNp
0HreU71gFiLJMfPCu43EN04/reYYvjzu6x4dn0BqOvopffS94C7DUSPZbX+fF78d
DsfW7thKLPiKm2O7KbKaDwAzFv8JlGgDeOz8ObTlBK0MqGtkBLSu4CtmwuKvAwYi
aTaSOFmKR1ltR1DYjAhoK0puoLcg7/4p94qnnZquG/Dxk/SRHWy9zfIU3zuRsKEt
XVyS4Jqxqy1i5n1Sw9eu2OoiWm1QdyDrPJufrgV+u/nYUMoNHuB5MXwmGnwVmx+F
jM1Gyq3I+O70TJD3ENry9EFT84bRaY//9A9GWQXcGuCCZfNJEM3jM+N4RoyexGoT
gN0VwlofrBKo4UAD/DyISaQdWdxR7qlSbeWKNnNjk3M5sgmWqmHKX5+EF4hG0gWf
pVTEeACaF9J7JWasWMzSTzeBTG7KDm2gvea9nG2iWJpi+mA9kx4XmbHKq7CFY0/7
PLFBWBnklRITVZDiYr5fWlCTyflVCLzVu9iJ8ZEXyZRKyaOm2OgDejoRTF1OXXOF
iLLqBz9OMq1Gq4iIyllPGO72eyfnbASKZxrhwcgBe9j2AElTsgUstNe3AOUppKE0
K8AqyX4AYMArv55mj2x915TTfJ/lVY/tSbS2Ol3ZxUzSGcYfn3VgKUo7ktaEfEW0
l97/DG4uIgMeP3id14eJLmTAFibAuAIFAlq9iOh4grMgJFQzcKtI+K/cEni+aRt0
vZMRCAZfsM6luHccxWSwVJPsH2AV9PRqCBxK6QkF/7COjhsJj+AKe2zzjD5gCUKR
qQB2H1+7r3t8wr1jdC/emCWYI22WUYRWIvBY/6DVxIw5su9miQ7OqO3nfSAtHKbM
CJQJ3WEX7gCSfsKmJvAFfU/7Wi7uD5oN0rq6bHKiLsJFV7FVUJf+IqlZN45fGo08
Ry6tcqwJjklf2lpCJj/WGV5SHOgK8wzkdaUGw4wOfoLRpV3OkO3+bBGJIKcvsHzX
BYZtkeTGJTbT7c0y/HAtoRottfSazvQ4nLSGsgfjrR07th596QNp5FfJTADiqEhL
szuk87FbqTEqCxk0L2qhIQQ7IYagRKYrkjRy7cr1JoUkpa9oelQumhBC0+oMKHIq
j7p8u6UlKXLVxyQvvHZKdwvjxjSV826E8a+6iPaGiAr8SwvoWshjTGt96QqSajUv
cVEBNohS3r1AguoL+QcID50ECdWFomlUCOouGzirUW756QTH2WaFmJD4gcJqwotQ
Gh0aY0hr/9h50mtNNwc+3XMBk8S/Fu3kdrjsfpwn6ahuLS6HXi4IVw5DrKM3LtK5
lBze5f/cjQ8U9FRanTF6CJ2wL6MZwyXZGHuY0cfG5TZlv7XNE7qeKI7ulaDlVrbU
brAKaVB+nWMcJMOPpZDrJ+g+Jbv+cZulhlQqqqh7rZLcIxOw2KGEtYw5+xybG5ad
zJGnHYJhFoX8LDZtOR3BpOVVa79QrA8hJ37NeRwbDIaquRAqtvplU+JohHuMRFvJ
v98gb0NX3xIwT9oALAa5VHD4+K69kV1oL1elWgyAFtIo2sffGv88VKyuDxXylsuP
S0qfVGaEuRCLBgfc+SJi+Ogou9LT/eQYhnTKYydERNdxooDlLTPTHQAXRCI2uru5
/894XEFNZFDbah50ZXMZj10ujICPeW1Y5XOB3XlOJDdptUygbu9RWzzdHVqvxWzM
rz4nPbR65J5A5xO/Iyx+H41hFNjQxtgkyqphE//Q/WFdF9qJc906/t5BhLNY51HI
en5jrdFgpwg4Zxfzgf+sd1OBeVNfdGoUqfr0EPcc8NOutJDP4GFXrqFdGl7CK90R
jRTzBJCzywZXE9Bn6paaIl20HAiNHbOmT2/cK3T1pPz5BUITUlLYZ969LC/cyTfa
JWJxnlV5HB3NGZ7kQitjhgZXEE+BCe7F5j26AItJtlCfjcn4d1vb73d33qdzDiD6
vfOH/Sx0gbVNBZ5komZaEKyipJCPkvX99M2RAy7Y5IB7gtsC2fNB+E7ij1wL39Cg
gSufk8AC9VN00kfhskN+dkXRsCPN5NT3YCxxJwGxTla9zmZloZJBLUUqM9Qoywgp
RmwJn6LsktMB4XX67xPGCXgjN51dWQ/OQrRYlzbK4sq3QAfyZSe3FFL4y/ZeMfSy
WX7gtwHulyLmhluKSjldA65o2q7v9JO6NJsHCtfHE0LJXgvIWoVbfJZ2Z4qfSiWM
IhPTkQbi/ooE0L6u0fCKUnjBA+OWoP4RZb0PHDBI/6Vqr3anuSZwWbV5glShA0f+
XU0Hmg+MNHp0R1qP292wmMNm+N85RHGBqbyKmujM78KY+jhvyiZakrgF24nEGIS9
7t+mYZBSsFap1HSnTLO51hsY3HLuRTrxtSHbZ7e++vbR5a7blBH8+XkxmPRCEahb
ZDE/7xLvhil+FJhRvaIiVfKbuqujJnSb9fcDDkjrBlq6KOP2hcqLYCY9UDjdwREm
19NHl/MhMKTzRC48VTyf52JAJLoM+gvd7fdzWm04p4R8e9WhsHq+zPuVAdoB1jm3
ncFGbpNteaBoB7RrAxQepw6NPr5xE9IpDitGoYDQbHMsvXcfkSwJJB1IRVGYEDtj
huXqN2KQiHaJ9g0Ln89W8/YC+0IJL0rgqdaQEi1z3D5QcC3lmu8Kj66VospSQHcO
JLgZks6Q69Lyg4XM429SCXHsY2tRK7lz4HNz8WUjaMoGZFQoLTdobfE1drL3tAMe
iPmrKR2UWF24VAfXE9WZdrAmrr9pm8niVGWgT1su+Jgz/u5NDR8U8uI8xu/wfVjp
DkPsOAJPggSS/xqERPtLtNTyXh/2XqmYOUKUIf88LgbYUAAFgnQKbFjpDs3vKrpB
rKwx0EllzaLtN3HnYICnUsoGryTJazYIWNYmOvulxoBqpMYdKD62ThTlBqVCCaZl
UPWiMEjn+dAULiiQSdx194lmOdoq9QUl7wAFFKyyiSGTYNH695knDl0jFJ3eBDgD
6RGkGBfAu3jpz0uHM/YE28Ss4YttTwMM77y3gGAn2n8FuzaqtqGuoIBcOYF+tRLb
Ydeb5hti++H0nLImzhH1dRnv6FecIpjnb3kxn59ls8IgsftJx801Xw0A4TYzuAyT
esG4f7PA+NNz/7DqofIwl3xAuCBLtJNSgFSyJFxuknXiMlSunbssY7hb/3pifZcv
RBWGWBmeVT5RHpPqH/Ka6LiLWH3WzXb7f48axty/YlsPcGOfJfbFz4P2dYikOfBV
A0Lho9qyjwH6cntW7r3nS68VQP/jta60So7+t6qc3QfufFl6YHXvqA61BqT0/ce1
v+QzRg9Z1clM7sTf1N9upXT/3tdPhuVhtheznj68Aicbvd2qZAck6SPpSs5veaLG
crCDtPV/tdk99hG4axFrxwbuh1lgc0DiMv3gKFU806zNwLOtuHEnMB2hRTYDj7fO
i1kr0J8Q3KMdBLV/DYTFBbOe3fuRNoKJRRGzg6WVlvQYaZIjjHb5dzZGhHhwITIY
oGncGDWbMI7gdGKPosHIFGjPTnfj5VgMZm0qO+H/akoNwolBfZHoVPOuZqcVptsa
+0nLPq950Yeb/Pf7b1zVdHg6dHli62UHTE7lYO3fZQuJqjBj5nsV/Wv3s4LoWstm
BhmYSbPMPC/9arevDELZgmFdjX0gK02bv6cMWmQirtNjTih9Xlq6hKqEU2hJlIdM
QdlPOMjWpTekYBI8u6ZEZ0Wz5e7SZI5J3rjPR4IRDZG3qcRnip02XgT2YrNPf75f
K7t/ftgFkTqTDPKxSFJ1/iEOphuibEkcvPawJW7CLydWPd39FERmGoFf2SlbMaUu
W6gN87VZpVr1wy9yzLQxdCoF9779z4j0HO03ovk2AbLr85u5rCva9Z+M1WuYywlg
B1C/mmqkXk7C68EC539vJQ1QPQxgrqBhDjgKN8L7jwtyc9xqjv/rCjURoyjG5WSU
vLJwqyBIxYJTFd9bzxx4cXJ0vZm9ZCy52Iilor+RFzHXmk4Im4IJJv3r7ccvLUCq
OVoe7xHVcs7k6+CXDoWhEb31rxmGtIv4bRG0XdAYztQk5NcCItuLcPiBCe7sWGiw
CygDD/n+lAjQ6+B+7THcRZyOC/wkcZH5DgdBl146sp1KSAUBKPd72J1hc/Qz61z3
fV3sZm62hf9WlV7Sw0blF8NCjGF48vt5GMzweZNgZ98u8FLybOK87w0idm2P5c46
+G6ZGGr7n/W3xGT8Y+PnvWMAxNoTurWk19XeskQyVzqF2Vg2aHv1Y2Prf0AuCEXt
hxqAAwNerxqjVx0uASMCXxJHKjdTSWIt6Hjckr+ltd9giNfHXAMmUzmd2BPOOADG
XB/RGcbkdU0IYVcStZvLzLMPSBHur+RjgNs2drCSHPVqrXgKq5s65e3Yr4vzOKHg
1O/MLfDHRWiuiUZl0yjHYGwxyuGAnFdwUYowLpx2ZqtkieW10hJzkcchov9vAF/X
FEVMMWPpGWGjY3D8ANOzCNkhk9r7lTspPumhpAkv/xQ1uSCBFNbeED/SzoqZE+is
nNH9/oQK9qPqN5d/o+2arrMWW+sftjJUUh0r1a7OdrQUs4YqUt3ju4fPhCuWQEGp
6zn1jsWQ2NZdmdJgRgjJn5g7v7IbIM9VNA1XY2SIpjlXjGb8UEuUo3UfnpfKSopp
Gow3Px9dNsUwP607LK5eiYtq3FFVdLO0f4R9bOCN3z8eEm0q6ps8sI1UxPyyakHi
rovAQHJ+jUCTkVQqqXiM0poRvdtdsZUtE25zPzoKUdQR2TIGP57/w+V9nbueRrzB
nw6v79ZUrPYaNMDOxDqmmUnvyP1MXvMn7iZBehy6vxqYgfkFH0f76IAGxnLbx8VD
w7JtgtZlP9QLzFAikhSOJ4DeOF0dSIMyAU4nmmfcspCx4m6Gh5kmqrrmHsR8sfGS
LvBuALpR37jlUS8bR2WCbWZKzmnB3HFGyc88OnXZI9CfqYZhsFLC7pjeHFisIDhN
fX79dXv6Xq8XrqE0bfuHlKf2GV/uBUBG9MQweMGBnaIJ9xh+l/eClHO9zJx8i6N3
TKk76tpr8NimVVbYYOR8DRyiKP+lbbilwBqzfX43CGA8E9zikM5D/bvjD/1uzPsX
kxPtNJ6Pxs5214IGlA21knhfzKe4dOuEZJW6q9ebu22R3FlNbOMwNvH23Lw5uKAf
Wpfqs+RJe3qOvLjYWHYby1rtvjQnaQZagPTom3Q7GecpZfydtBYY7yMDflrNxsoY
FmiWSWffEwUIs8Y9wERquvdHozov730n6rI3KH3JDL9KvV9tPqxHoB4187gbTffI
zg5uNv+kN1WyJ5NrXdqaNUHAIt/2gHsW/9bFWwrQ4Tdxu+hTNQHOvmNYJXx5OrDu
2L8/c8TJCjoEcNzxxZ2pgdKSR1nOXr8dHRgwrB3HfHf2+4z6/pirELE4aW6s1+h9
kbpLP03LIwQsdj8YV3BZOalis3n7R6RXFUovPIs4Gy5Es1sxyefl7+bkzQh266o7
VB/kvd3JZpiYoril5pNuH6S0mI/DpPxLrBCWyGTp45BTj5BKD0VtnhTNVSm2oNCT
Dh//mX2opWFHrqI4pLWs1KCxnyyEIRCY7L9OlgkDCCEZ7eGrYSubfrMHkPonGS+9
K83dBDwrx4UNetJF9DY1TMNnsgjY5g4c0sKcEJNAsVOJzrI4CAXH7uaTAY/nJhjD
hAgs2k2EKOCuIk/RwES+Q2PpyisxVgJY4G2xu3dUTWXz8ho97RC1Isbole5Ma0vv
1na/eO49Jv+f1FTXYb2vTBU8mI3NZClypiZZOj0HQvgFMKkhcH0hULuYfaF1Hvm7
8A5bwLv1UmBsFE98KKJJUzjCzjY/lRdTE+HbXJdZdVT/j2ywN97IxWHYlfrpal8O
RlKB+GMGO7xhjwkLawFjRaG9m65Ip//p+vaN5CCB+Xu+c+jYeXjw4tfu3Pv5Zh8d
tf0klZSWqMueDelRHL9mCAp/+RKMuHN/AZnJaKd6nAbwnjzdBl04Zv9NPff+Cyoq
jJ1rhnKtZI5d9vELGCtiNqRVXoeYWGujOqBWSZvEM0pTkuCoiNGEJyUZmckYTAVq
j+zfBZWVNVLUaRi3qb2mcHAEp2kA3RQG/3VcnHoOeeYpP6O3+L/+FFJHkXz5OAqL
B1hjCexqGAH1bRa7v0ZNsMDeMTE1GW24GXYI+q6VhfKvTb6eB6hzSaQzAS36T3+R
8ZLFnDLCf1UIILevDTP2P39vGYbsCHooNYo08F4fG0pQcJuuKfRlfqRs/CFgE6+I
sVjNW6T+xwBO7sF4A9DjlDLhl390jfdVuXbiva2lXfsGYdkmegS8XEJH0/+Ptuih
gHONtynA411G/Ju9cHIW8/LqFiR4McrcaO0Mc9mL9Six0aEnkYcOrfS7Q4BmM+DW
sjsIpqXH+RD/UemjvGeuyJ7ETTxeooj4Sj1dPjYHrmlhDOboXfmvmuKL6C86841k
z/e0coXM6ics43IT/1UoYmY+4VlIydWEscQYx2EafkYudaDJuGmWcZFuFem2lPXd
6D5A41qMey/UFrM6jmmjnQYyhvvmtNu9NdXmHfI56NdlxyTgQfW4UltB6IHml54f
bti41PQt5U4Y34MNgE7p9KgwDjW1atjxHfu6MlIArkqExAMcEqPFPibvXK9LeWJd
ULLw3Oig/PTf+3EXRSFRQcI+bvh3O+mLkJTKTvEvGMuyKh0jUzs9TkIBdVQnYNyp
z60Ame0W2WABWnew07LcEYiXKb3iuWsQhGzSj9i+IPsKEezWJUasXe8VzhRM2mve
IcsJ6B7UCGuOrTRnVoBZoWlf89mQwviBHamh3bH6ltNHt7QLNGbj6lju5gbeMHdK
XLrkL7ZUFJ+2pewYj/4cFNhohfRiqLZAksBekCFAiRo3d4jQaDZNde06Oaz9tjpZ
lsR/BV77/c2lynVokPRt/H2vmXwPTYGUIyoJjIReNSP+KnQnp76G6blsPeHxSk/q
lhLLt+wMEIYMgtuRy4+8UyqnyAoahD9t+gnpvsD2w4Mt7lU2at11prsvVEwvIwqe
lXhSqHjs9er302K/td0fU0o20dVnb/ypQEb+hYCHAnrJ3V+Xzn/HciliYeHEvw2N
0i7CZJWYmY/rJgRNvLeSKNUQ3ot2PIPSxBOjFxvxBrEHPiWSsyd6rtGMidLZkkZp
LgPYk1lP8qYZS7KCOGW3oJQJQkmp1uwdUMdOonobpvdt8jcCKK4f/MDYf67i2AtM
EnvxOIemKcZsjXcas5PiJCIElfk5ueWLeRj7hESi1ohRi1qgAPH2yLK2JRB3iJXT
wzeOD0LNh1HZ3YQVvuk/iwWUf/wLv0dzf6+iC85ULYLaxft7z4vuJ8yCZeGNCfWo
vjijdl5xllgQLCfHqJV23fa3lVV8e+78FKFTb+BpJBlfw5yrEFbRNaog2lhZcz4B
mAlirdPCF+gc+Cdoh74GusMnno9qdq0sWd/XhFymR83dLLerLMHOeG/9oBFL4u6A
5L/AqDe+qtK2SeJ/pxtC0+fKT31k0eNnzqI+HBE9T7GlIT5FRE43jFISn58Fq76/
fx+Q3pgaOK8kr2XfSUpls3A05LZLmXpe8tEG2bIuL/MWQCxHplTrdTEuzkMNCkgt
XSr71/0fh2t0ZoIkSqN6yvRxIt6ZcOGc3MsZfRHyTdLUovYZxayYBoqHrTRpnPWq
ErEk0lXNGTnV562U/U3jsjpDeJjXdl++Yydf2CIL/mY+wep3JczjqiGDhI619IOC
cRByDPhysMsi2AftiIq2+HwLi7van5fthogOZ9F3VaNnOwXG2fYRImHsWFKsFxIa
7q2utlrZvCxnk9L9+Kfq2VzfpcTiIBMxNCMa40Mp1p5zFDFJa1hos1OQT/tz39ZR
O9lOaiR0YV1wxu8wbt4DciKgON4ASWBiQOt6EIFzGoY1aeWXtiBT3r7AGdFv9wzv
BNfasUw1HpfyAMBAWzHOkGnURHYPITGB4n4TI6o+Ro/W/RyCu8rr6t4WlV5562gO
HN8vVm6zbZhMoapetejWJvTByBaohG8w94OyC4jO3UFCPZtIPGEIFY62FlABiNU8
RlSDli859M9CltlnxqK0GY6OtjWpYwcH3lPvqkD0BTp4wYWN67ru4qpjOTfcWtX7
+kI73TSLvvyMSz6l/Z/zfvr2SuG6hncKOw1tn43c3O9IvaW4k/GqEoKY2Ey3bZt+
uomMWpi8+MiIa+28L7jYtq6NS7iofn/uvBBoyiVwY+73ocBEgmHGpsJYb2sLdZYX
RU5xQCjrYIVFeBMxvYBdzn96R7Gib6SvIJCdx2CFZLWvU8Qd09sSRxpw+npPoH0Q
lowtg4nn786WWlcjNy5+IWxD2RVGH74gSXtMSfUH8yyKYAp3JFI5PEWulso37eKu
P7aRsUeHHARlDWuebfIMBFgBgbYvgjFxDdCnMk2MRXD9JW5IK611aSijjLAz+MyM
FYxoy+13VdEYEGOVHUguBB2JaMWk6aZCnhErTUHA6DKhhhKa26rWss0l9pY/1X2D
GkACjY6gg2FLqbO6Qaz3J0Q63gXXB+VwvnANX84oUNDqtgtHt7FkWIAYM9NA/M6h
YvuevMVjo2THXkoysPi+Lj5dp343A//EyRL5QDFw3lW6Zfedy5s72xO7EH8LYPRS
vnd3G6l12+i/K+ph/ZeKYarh3kmPazTP5T5t0Tvu7pePLJb/AjW7DDJYj436fekj
m1YDMJlcc7nOr/u9fVOzSRIzEF9C7D6wZw42QKrc0xzXZMHXqGSiOpUc3iG7JomR
cuFjTjZ2nv2op82lNkXBJBYqErLLdXFzPy5SIdgfDgNch9uYSnT+71fXi7pfqohZ
R0vJXqJgL2lPYCCsShzA/OCzNKuMydaGzlb1P/PLkqtTTnw67UJtSkDJLOwPgi92
u9hOaHBCBoUgbQCSkMmrPvefB23johHxlMVt/BoFSlZuewA6wYipy6lSFctX5QI2
/OpS609fuqmT1BKptscnCq0DhmRmAnVUn7t/VmULdLVLwb5g7r54h/IQiiGBtwDo
3cT6H0fcLo+1k3sXlGXXuHE7LNXrjWIQgxVB1YGdvA/vqtcyMCHgsNUojyeiuJJJ
G+bjSSGTsvf704gKqrcZy0tWu63WTnr8L4wWMsUfnlTcnPNKRJ8ZQMTqn2Gbq0d9
fu3XdSsSShVkO8XXZs9sAQyn6u1ztDOWNV6QnHI9HuSxCV7978lfQxb+CXulBcs0
pMUiI/45mTR4zGpKDwqGXp0f119wqK0ml8SRXxJuy4LwdbR1V6tDtRZgTm1j6TRf
pIZKgLPA3sEIQMZo/uTTuG3TuNLnSrPrit2kymE36HNSO/LqcmKAbqqnrh+PW+W4
UjUU3p64Ki2LhPvB1IZD8AJRGg0wqL25hujge35wExwB9n8FAA6jP8cegqYsxPxK
A//C9+n5EM16f8EG0AqU1sBuMi9MHOw8Bj0Ug02BlsBs0Uu9fdpeCX71yJ+eRDUv
8Wue0wdWbK2HVDJtEQHtOjXv8hmyLxJkojHiMqFJBtsroR3ANz88/oAyiw6KLWvK
2bjGcflI6nJb59zQeazLcWDrjVv7bonwDGULgQQRnBd7Xq9XO1DOWMJ1Cum9wUbZ
InICV+ro+OiP2pBSh6dfiLn6szQOYQzgjyBqyLm1Lrh3+IYpSZapxGOb+QQWdqof
3cITpKjBKkiWYdUTuyUKoeGtdTqbY02TDRYT/CQEuD1EGNXhMTwRcEwczlBWLrY3
BBykr3iNN8tUOt5fTicbOWLvZhMlhrKVY1V7iKtUNlvIjg8iCu1WTq06rDAd/ZMq
hwxHveGEvRRML3ZmeKbJXXDCYQjwzQOpd0Dhh7/6QAvr7xUX7UN/uNc4XUYaiAB1
82gyu4Cv/BpXCp3WvqKkkmfD/sS3RaLPrTUtjJ6Xsodi6mF2TMaCwGB4Y9ZZuzIN
y7usjv+s54r8DRcfbq7Dl35CLJ0mpfAkDeSWWnM10XIKfvSI0uRvEhKq8OX87WBq
+jd8OFR9YLTKHO4TA+Phlhcnh/E5LGOWvAh5dII5GYf0oSRa47mSNqeNubORnZkB
uypvmK6Se1zKngPZSwp79RyyOSBG1hlxi5FSXadVECck6dlm1kgvNR+ede/TfZt7
rJYdJQOcKp3MogNRTUY2XtPWqSTj2nvLw4xgQDbuikYjjUi1DC2lbJtMd8L8CV3t
OvByMFB4RP+GqTEjK66u+Kb6XNAT2Caa5V1CBm2VwrP7WzVp20TBIvA5wyJX8kUm
7b2XgCXrHw/fx7Q5sRsPmnvuEM09lycFxuI94dLmaeyX9pn5jhFifs6hB8UMBlLH
QRDv/z3NKMxbqCXTvU0wEZB9RUUBE/xlS3N44vWLP3Vhub+nx5JIxqq0Qk02YGa2
aqdUd+n4jTsl8jR3+iKOJyK1Bfj8TCuWai1byMfhS5v94NaKQ5p58hfImC8VQ/II
NAFaf4F8fy7zqiDWJLt2bZQ3E3RZxpNFICPhxpsT83xFVFNWQYmt+5gSn/PPmOf1
YBTP9Wq27r52rPMc9zYJw4/+iAp/3kwx0CKXcKVif7iFNQWImQEoa9WXkaLYoWRk
6z3iZEM2YIRFvk/tvWOfrvwKoZGaJPE1SLYaMSCXGlF1s94m51/aYRfKa15fCe0n
LzeaFGYgxtzPu0ZfFrmBxoasqT0eJApk2ZcsqMiaLGn3RisjiZxjBnSJn618uzzK
DRVElTLEDuU69SnTBHEEZSBbhDhiHfJUYBqtLZmItEbYOZVF4HBMQKVzZ0Xvao1X
+IMfAAZ0UJsV5YawdH175h5ThuiU3jWegJIDUy2dY3j41ZpmZf8XSRoKpNhEGWb9
M3Ch4CmWiPY0yPsKg1ImD403RLqGprosYcBMlEl96UMz6yfWejgo+XB45jPbsmES
ox5PBmO45kcmhkaJIHU+qvTz/SrjLtcLSVFuK7753iDcp96qbsm5JYV9mtEDkx6I
IJLfDqRd29qj+SvmIv3VI9O9dDdCV8ib7QhIth3oLsjhplI1unkXlZ0RPHTr22nH
JMFLL2pgim2qNZkzYI25HKzlQh214YcqKzjLptYMWIsbEXJZDdM4RYatl8sI9cyK
dQ95FLFltQLklopgpQjmyj9AruLv4r4QjxAzmJh7adMx0itkfRLZTwHnpda0EqcQ
pl1Xa29Rc43LYtGx/4ZVs3FCcycfzW8dps5GrjpQw2NOB7Og1pKVitrOdkTEPQ0+
wzefBIfR3Ik4jRHB4H+X5wJFoAxS+JZKHDn9o4gWr1E1InSNn1S59QVmGQ0/91y+
eWZwgAIOUE6gWxntOndh8HjmgmiD1bMHoepan0IWrMO+BjSoYzDXkxNlC246kTb/
mC+UiEl3NeTReGhwBUpEf6OELuCNq9Ymed1QsEQQt3LDc+yhXUsOTgYW7CaCkFMY
zyprqvHq8UZqCVHrE6Vz/HFDBwJtvo5uveK02umXbqKWvt0Mn00uh3TnbmxEsQoH
0r9k96ZpmUyED6wDIwbPvWxudStSjhg+bUrM4Aa6Qs+mF6BEOw5aodmy4XwQHYWY
ATBVfuuMh1XhDpdsIewB69wk/6H0vq7QM77KXzCZ1J2/faWtplKTf57i1D4EO3h1
MsSLizB8G9EyMYa1CzOS+k+9rfKYDUvgoN73eSMXwgKqc1HP5OlHavDh2/lbq5qP
j64nUKYu1T205KD3sK2tYfHj6WFJvtwHAuVs9rzLgv61qPyfD7L5VE4UNYmHoGvS
Sp/HUA/B7lonj/aRJX2Hhi2OswHDXQfimzZkFtoMoxyrQrHozGYBTgmWTAVgA71+
z6GbUVfrpM/gu29dFCxCyvctTocjjLyQrb5YJ1yVI6bVgiICf4YbXIs7p0vh6zE8
aQodulgRECxN2YcqoTezxkzbvF0kBiCSHp8LD26qoiKFAgmL7a5BxgUV+kCGSnSJ
AW2TawQvGw5iIaAuKDDz9ip2qqZdXqXrhlpfbtdYDMLOytM8FLbKfCciy/tiwmh5
zyBetGHzUReGxLAXjf0ilBGdAq73L67nKHDqZCC/SCwuHNJlgIBOAyk/HtlDxhX5
ORGe4g3guD1FYRo4TZ8CNFPvwC/FxeFD2bIBxv3tbVP3LpFwaCDQd1zVjwOySG/d
ikosYJxPuzDQuyv9j+6/dB1WC1hnK96Bx0geU6ye2TgHwf92pD1RxBa7uQc2cRWK
AB/YN32cFpDCDulaP/6qGawXn/o9FcBlz+8zgRrQ8NH1SMIQXHjcEc4CoZ4bffgS
tINr2yI1mmr2c/VgFk2/YOOMFgfzjwKBa3PcyiHXqmGSMVUg5yqwx/5A4n0+JIfe
W744hfqdXzIuxoZlAVuHIYk9dvZ1dezOFgx4JcpRg+pdO4ujC+0mS21ub0zBjNQH
GJH/6jw8wgrZxevk51A7qsBJbDRCYdcX13Ahytn0e2EFqhwDT3Rz1D6sETQicepN
kocVfPRp0KermmPx72zdMBZCOUGIDTYcY52NrCRqlYynQoxcqun2WK0p/qOApmXf
iOWvxs+qjh429sIlf9JrlCNsrq1sLtRHJGdbmyq9DUIv23DgSbaAvyilXU/EuNmZ
u1XrHv+zKj8WrlIsgkDxwF1lDds24WyZVD4bIWo2Eojj3VeW7BX7QEc8lbugA5Ga
yfbY4uE8vHn4dtl8AOCgwPxJ/JqENfAjL5Mebx+HQe4xN0oLW3a38yCBSXLel94x
ZUcESOyJ1UbkVLNPHRjr9Ij8D9bH+0JTLbIzgiCQQud5U6HI0FR1iVfa9pFid5as
OsJ5GPdCtBF7L784n24e+JKTG4kkyvCam1jUviF9buEdfOdmIfngJYf9eOcxeVWI
tCNXMVnNDPMiSSEWC5BToD8lEZbCtq/FZ7p5ZhfrVWkmF3gH7xj5SsIZKti7rASR
9xMvYQ7vkQ4fH/PWtbCVCjxW73nWQW3OJXc8oY57MoxOv2JACTph0GaTKL7PJ9wX
YaN2HlvyUP2ySkHqfeTPos4AvrBNSrcfhYSqwQBASqdhHESeqgz13TiiNhecXu+o
dkPJLIGB22m4iUVMTlxMnh//wQF2kZK8ZceJBDmZm6iVsBbPhtwDmh4WSlnZN1Ma
uDFR0Vk1kK+7awClArlOo87snOVH5D961MBnH0Nuc9t1fr+nwqvIyEZ66InOWsTx
N8WJZwCr4r+PIRW5t0VcpkIrVoweOc/SqeYN7YPQhAG3tDWuHhceN5hekYje/cDj
komqJVrxakjTUUb7rEluPSGrSf8+1ruJXZiwn+Ahv4DH+3jwBGhkeBdlOX1HUWa3
MKlMhhvGirUCNHEjOOfUfnuipEQ8LIHpsZXbmcbNxQyvXnMTDdLOG4+Uo6UJS9l3
HvcRaPfyfUVYBLKAdbcpd6tqq0KJXoucwfA+9DA6GM0Ks0XHfElvkyySjodRLih4
zoNG8vyHYWi95JTur2Q4ixG3gQ6HHGCGet+/AB48qf2NNjp3d61lyvIhGq7nShmh
U4jlN5zZra9QylDZuE0UOv3LGLlH9GfiKopLqLm+3QsKjQYqow7v81SYSuamqVpz
FvaBuqp7QSPicbEnADsy9BXBvERhD/JwQcHlHk+l7KWJ4g8Nx3ll2mm9dtnlxgJC
4ArZ75hKSt+qsIB8PTm/jbWTHNIQ5/q4gTYnl65WIkId5M8eu6gbp4E7KZYu+yba
i6lUg3wyUIoy31wi1wEaISjIWdCigPkSGRhbRYwCdyJwNVavc3d1qldCatbEDbTm
di1+R/562/1y2isCON16oV4TeKuqil+MIHqBW1HP26P9WkLvd33kCaEnlGEkB01b
pz2B9pHoiw0t7aZ9BW4hQBYu9LkfK4XENmhhRlYSR2Va8EOJGYVcKPyYSOr4MPGG
slu91/xouLDhxmUxZX2UyysYY2id3gMskkxc1Q4gkCB2P26A9C9vx+t+I+QTwRH4
IYV6EU/5PAiu/8vWGlOrmecWTc1w5EzKoG3l1fAhWYWEEtZq0cnvxTp/BDbXdKov
0Kc1/oaNnWGDfbdTRJir9zAWIhi604jRv+fyCwxXErizlqVfIh2HyVjck79dmhiR
uvPuZpVKa5fBr9Mo9QSL65HYh9ANKg/3fLe9qZJkUVZzQMK47lyK/Ig3J4BviWQT
qtpPH7ihOXMeD7+bLF41fg+1G7+ORHgtZTGUaaOCJ67hcsFE6d5ODF0swi7/OGV0
nGGUFtutOFtQNiMJpxaHIli+UUUyFSasoBCMI+8p0T3VjSkuLTvGUYTfUlg9iVz3
yTkcy0y7TIyNRQJgAXxPVzrT4oe3q+a7X2aJ8nOLq7CkMa1wIbs9XbnQh0atzs+0
Pdmd1D3L+WwuPVIJLZsS2qfLMFHi7JMybazZeecUh2F22qG++SH/U7TCUYvOQjGX
DucH1BuXK5bp3cT2XjuVMudFNCn+/CgIF+UtRs9xADUHbPR6vtCbTNt5BszwdhVu
om2++FjMyd8DVmFtZ4mNHWh8jZbZm38Qibeg+NDJErNbN/kNmN/92/Xc/1WMhp2v
NnsjvhGCKDvJBi4R8PSd8Mtf3Xu3QVrl3uSUUSAIWUF730W6WJ28WmmSNEIBJpEM
66IDs3rwD7Nz1FeNvjtYePwnC8dv5uwJxPkHrqFzeCov0QBfWEE+OQlb6s3Bh0Lo
Hq6wJeNUlczBZRlcOHi4FPtsJQeAdh8S0t0ALxbuLH9QPJNDVxa4mL3/q8c/odl+
sxVXbYBrHMm2w2iAVorYli5ksuDMu1H65OfeiZlarQ7Ruo1Tyy24mOEH4RjcjLM2
78UB3EWY5HUHwHSoitGPgzn3p6ln5KVBk0nlveZmXrqp1gR4q0F9BVPrkSgIJNsR
8BOX09xjeq4ctYyydXjFGX0OJRST9nis4wp6RyAxMNWa6zMmZYaadLRb73PjfFRL
YONiYmMHHVqpYcVBdK7V25G8YgOqRPJHzVnB/VRqCAT+SupkLwphh9aexeMnDegF
wMmumDYwDeiQ6hHVrejp97YcmVXolH0TNpjlsYkGO+YCLw3Q/AkZWBzs4hyCImLA
x/xoMAFbNpVqmd8MwKgFIyruNYGf57Dg2mXyLQXN9Aw2VQcqu4sNYmm4FH4TaS9R
bSZSK3oLenrQbb+YylfKw9LM0Ee8EfIbnU7y8+EHQ0Eh6FhlYSeePTu145p0+dkv
L7AEDBQFvHoY7thedsnEZkiFTcanTwat85Qnz2mnVh7I2G52SzNixWcSd9pWxGWh
ItvVxG7iZjMP6E+N3YQHjp8RMN4rl4UZdKyRuT01Lp9fNgDnh0O7Vb8wzJjKKduU
+8/VBh1mBLEE1osx+X+L4kP45yGO6FYlBEpxsio3VHNeMlFXa4K9WNOOui7jbPv7
guFNOWDvPIPsMPDUiNFt3GPYl7eF7L+wUMOSel11LwJGf14gQKoQnuYY1Um8uLG9
kF3Vlshe3ddxgctO+EDqG4rxB2K1iFg+rq6+n+URAxW0Ha94yl90mGS2lfvHT8AF
gGe07axVFqlcbD1DmsQjDzH3cjDfvVNmML4sUSaBmLuK+wfhj21CTlmLaW7IxK5I
Vz4eR8b1pc3RDhu9USo9HS75DY7Wan7+aLao5xLuvbHbShhWX9klC3O3YmXzsF5K
jelMiFDoY9Xv/OsWck9fQoYEd3CrP759cM0GTUipcGj6IgOKlMTFWnwKOoCbf97o
U57LqPe5BNhXLj9b70O4xRE2hqdUFD2HzhWOrt4VyxtFbyVvIzlHtnSNKttSNmfH
R4DOkn8Me7uYPKhVMcRXrYsxb6Fyei+GG1Bde+tFdgRtIupQsPJaHRsvacyP7iyX
I2jDLxtwORKnH+XXpJywxHRIuKGOzOoS6nYigKIWhAqxzzgpiJYLGk8kj6c51yUt
pC/SST0hHynPqh4DtYp9+i0lwLNspdEaeoZ/pl2NP54Fo/6+ts9E7OCdq7gSvQdC
Frk9sDLTCgD0AcRGoAhKLozmPM0UcJpWKxWGMstVYDT8xTEZadaA9IDNTYCJQl3Z
qAzsC7y072uzHnhlhj/JPRQ0lcDCxljzWunGFZji0rgyz2fcof0vlQugzYx2HYv+
nyZnlfr49Hk5wAzK9i5SxMWmCpX+20HmCscW1xZSrZTLLYPrYLxchZAPaOGVLxek
X6vjIvRTCJNAyWyrFRAS0IBUaqa/12h6B8noxkOSZULt/A2fn8P0mxQaigjcPhjO
8CHT9Vu2NPB+VD2GeyV7VSzRO+eOo9u6VPQpuy9iIb7rUPaYg7KX/yj+PhE/qYri
qChHqcjMFZDxFxqR6J5dR2A+l+wisgaY3hju51UV3ImL4RgCwkfXWC+8YZKZXOPh
PZ4QelbJ7u99PSwbxPNAZSSdI2XHMJEdgxvUSxHkNnKhmJkz7xgATt+P32YIxmR1
h+UA+oVDJffBfl0Oqgv2SV1dlOB03mp0KVZYSIqi5g1XY/GsqQYAKvZ25IL7MnFr
yMB9LXLoqCy7xYSIhb/4Wdoa20jJSxENX1uaLy94iYGP1VHrom9BMihq+X9edkLO
84tQNgTYDXnxe5fcYoLe9PzzYSAt7mHBJxILgE0t6ow5eGsA2y0jJ46m+RBrhdN5
S5yvzSR4ucsDnnoufEPSfI10eP8tBgC19fmd+RGNa1GnG0+tPB2/pzNT16lJJ+Hj
gnmsnQHWpHC5eWKpQ8fkqmpAabegP5UeY/G1cOpMOrSAs/rxfEKQEe+9oAFo+fKW
4ocy/jff6dnQs811i+zOvOUJULG9fGaAf7KFVe6Ym4mwKyTScWPZvXoYYRzqNK/D
NvTG5gN60eaFZBtvNGCi0VK7GqyNyWIxncBShtkFeg5cIh8QOjECMGbV5hjQl/4G
yefwT/DjMrC0bdgKyQhgwv7/9hOmzzUacnEg7oUXtnIBsOsyUvHy8+RK2/gPxNKZ
Aiore+hRviliKNAm4gY0odt7s/JFcx2hofIKJyNFsomWe5+JSM1fUyaPhxSrQPVH
4pFPLINzuJ5GgwibqrwotABeKJztp84SLg3BrpG4XU83XcwHnCI/JmZu+rcovRFZ
t2ogF81O1ldmQEWCn+TBTdZNhQQhrYCWKfaKIdSscj9koTyhJilAys4c9AsYLUpY
M3z8QEze6XTK5CRzq4G2pyLOQo3z80IBQhIQ5xf2zLxnVhL/zLAEbvqsF2qiO4Ou
V4Ien5hbQDhIsEgRH6fcF9hjM3nLMM9E18VdION0uWmlRv0T6DwXpcNG8oxY2xme
JE4vZth3QT1snlK4J1BeFhjDNaCj4adY+paHozH880dC8WmIRCAV+PgmNmfZVEyz
nQVTmkOoZ1Pm07gXJiNrSjKSs6uNWcskLY7BN19kc+Iollu1MBXphR7JsAX0MYe/
duI1LGL9OS+DEgXj/UvcNbDIefW27WqYG5QvK/aLTzuseCXvXQPpYXYt0N8SW0xA
meCXZvMqTIrpy6xhP+j3kPQ+8UmGTTKSVrx9oeafHsh0dtQa0rw0OvZM60L2jI+u
oBsPxg3RhNfXHyN9BEPcTiJrt4IJg0Jw+YjbNFKzTVbqoDlTV/ZxyP8vFGUxS8di
M75t1p49J1RoTs34H1IABopaB2jMLGx0Bef1cgae9g0Kz4DYGTC1VUD5Lg45DCnG
6nhUrXtndmWlTdkrZvLv20V50GAQlWWWWJdaP7eCaTr33HFG1Tyb8ZFW/uc223hI
a9rA687a6a6SyJKpuZgXOXWz+O6pyreuOoIO90F/teK9TO1TGAGpm5WTBHBlPrrY
XvLoLva0MlKm3Gyvv4lqWdZrjz7Ll3U92Qr5bBuLwiZL0Z2V13vGZxlx3WkIzSml
NE0tmv6IyiJ4Kts5XbMRjVwzl1XfBu65uPD1KrdO3MAx4mA+e4H6n8S+Hy1EiElo
xAUkBqOze54zRdBq5a+S5ZFJRyeHXq3wCKEzErSOMhVz4XPtm2Dt4CgUsnpYr+7I
4kV5mYTCqpJhEMcJwUIAqXdrerFgItOUHfsbyDQg2ZaF8VwEAw7pFMR+Rv7N9H5m
pBv+eg36AOtbMiKydmLZfMS5oyYMD1jduAo5OkiTWLIrmCXcCTUj8RypQOlX5l7v
48uM/4g9tpm74qTohvCvkBcF6igwi6SmJLumgjPc0z2bdrqAQKRZnqRqvPuwP472
pSMM0BhmM0GNvYB8LgggVmCLDrkU+9FqMU0neh+bEs79nCkw97lfoQWFXPN0jajz
7PgQo2P2hWlcYFtXSGpiar3VDI5GEZWXgK466XDgR4rYH6pWN96rUnMA6vRD+lUw
TbZnpJQY58swhvgNkzuKGh4M2Mb0CDFptXg8OLBGivt9wFPm2Xre+sChIMO9srNM
LhGUvn2uQCWSdPFMPkBjWabi2S7pACXheM+AMsovg404/LHiwg50IUTdcQiPN0Vz
yz+QwFfY15PYSVK3qZqYfZLfPo7bcYncFJJBZ3nUzVOnLgjReH64zCKL4GcG9OKX
uJGwb/H+zDBPZHUjiwALC/pMXfb3/BRKxjO14oo6NiL50X9MIiRg4P38Ox3b5FI5
ALdJHPAoUNHrRsUZ6hTyZJfsxTwyKwP59AU8oQn8necwJfx+SC8zfSiVv4AFj6Db
8ZX9bnh/F2S4csHPAEV+37h7Lmp64oW/04x65jPy+YhlAK1/tlLl4+0/xFfiyN8H
KmhCvOcbd/4lQwtLwMb00oDcp6SShoRSATYk35pC4Ucn5DmwjmHCzGVl6qzz3tWp
k+2QDKxy/izz6v4kXm3mgVyRmM9pflVlOq55VgdlSTt+z1+L7hj6IJsCwxrUsSTT
tSjcqfAuYkp9Kk1NkX+SazSdpqjSJdkZhwC6SnExpANlr17QG2/PaRLrzVb4iE5P
WnsBBL+wI4uesDehX92J1wSBqz71sJ52qmYeh18TgVikFKo/lfIXcexRfXxFGqVp
EkHf7hGKywzLhxkCTULyQHMMWH3D3yHoS8D2r9uhMD6Cw4S/juWs5nH7pc/ee0Q9
Jiaj4Ogz9r462q6qnfR5xu4Brecx6gwFP4lg2YTGR8uNsKb/WeW/37/DUIUuSgYd
hNNNb1LOl5romcd8FV8n9WZkXgM2QW+fpucjefhUj3PY+UOGbe7SNhQf/q/mfkkF
mfMfcXjhWGTKu0B7BNfHQhcal8DndVhh7Y8dpASqp3mFRe2/cVZ7w2Dt59cs+Rwe
7WhcHq4Ywiz+uqeUAjG7EFbP0M8zPZDVorsOUA8y8D0cu6K2rMfpigKnK6cIcYOg
UDH/EcNVXh4s8imUxMRWtIbUh3fKUejHj2q7WInu5k8OSyFkQm6wDknQwM9QNYkh
NC7crV3njug3StbFiv/GHauBAJfL5IQC9VNYIRfdKmmph1KMbuIo5Q4+U3lyXKQk
QqGdJP6SqsDol/6NyYQKv4E2LJSWTbuQ3SJidbJhN/3OCFET2jRKNjPm3ukinyqe
kdEYIo1NH2ubrFLhktl8A1d+Oeu/T2l0rhx7W3r1WQqk4pToHk3lZejvfTGab1UX
jzUlWXYlFfk0mZEHyT6ziwbau7EWH8S3+pG/uolQpisIXOp183MuR0eHhgvcXwpD
iQwl5eexhbr9kspMTqkFd+N3IwYC/vFhudA/tCgZJlCjeGO7yBuAIX8oYWwHEetF
ZFpJegzKFIdtjRLZ24aMO/vqF9peYIWHVLITMOs4OJTW1+OJCvCKTNhsTHStO/j4
Umq43nET2TMeWVJ7agORfnfJ4RPBSQneb+T9zgQvYxme5a3yXWL6BdjGDnMNrsm2
mf9PVNElwO5w/sQxH1pXLWUMCi6tRPaVkcf4s15/0H63zUsOeHiaew8vByVwzP0G
Y1hIZDt8x8vpIGjXeqU+KoX4pwjrJwiPQYUQ8TSdBbCLVhQowkp68hQ2rqbZrDAv
wB7tx47STUS+moWwEWpjaeT/G2vPpsZaYsydAy6CNsFNBStnRU9hU78nzS+I0TDV
iT/T3O9L8GWV1Fv4h7KVA5uc07JGLZjwi7g8672/UUlPfnsD5yD3tSGeD35eh9NK
jI9q+GCEiL5x5JXjHdcUHuPhJddbNUZHpAEFH1NlaHfqNSZSJ8BicO0/BQeZPPIV
a7bq1kWgdLxftCszOGP+adVZUbi0ShKBNCfbkWIkmEsPjO/p1AUQtObOl6N8WZ/f
7kNQjnmxbvUYL/msLJOVfiVqiPEMX+tqmXIovhdJRHjmTUZSYB+7tvYZHr4NAbhZ
omUnbccrJMe8BDCb3xxvu/IhIUQKjh/CebFFZwc3ag2A0I8fOc9B+ZEyWrr45OD8
KqDDWMzsKzj9RmxZBFAAvRDQlpgeF4BHwFlHX/YrNKSRe5pRiuLA+33xyzboMsSH
rB6Kt2DfGQgH6ITZtZPpdOAM8Z6YcPOEvFb5YGaFs8Z4dVamV8JxOendt5SaAtJd
lURs/7UUu90YJt9eHNKNBOl7nzrTwpq2JqK/dOEQ5yPkJo/sYZhUJhgjTIPEUw3h
/gWXVNth6HOLE5kwsIhtNhEgJ5pSg6xKCUZDYYPn4ic3Ddfvx/Bg+P3S1gD8uArg
ju5qsY8vrA6/p+MDPgpAAeWcMK8yLebjEIYo95oLmeULRfxavzQvWkQA117WTEEH
Qkm2Zxe5H+2brJy0A7ZMbzlrAMEkHRvdm39Gc/KB33vuakYVvdEK+cfWGhauUxPD
cjccwGxkgb9vNo2ARoi7dID+8Zf8H4xZt3keYYPCtOUSa5ePV+eidNzDCbvsn4Sb
RYi8boSxhbP46T61cJpp6VeGChhm7tBOvjnYjucfdX+AMwVX4PA6rFtdRTllxdbH
yxj5XKr2whEgOF1b2o2ee3dc43x0x+FJOGussXNqVKE16GdJrnqdye01vfdpGAtw
c08ggbR8wJuVspHEioncC1p29K/TnnulTg6AK5ZHoWml9ZHM+xrtJ3zxWeVcTO+G
jYsqSEi768UBW/shSQBvx2rw9dguW7nrRA/j1u6px6o+TIpXzxS2TIevJZUDrjXW
Sx0oOSC2miArBhCb0c9Zo3n25usgdjWWef11H71yz04uJgSsJizbrKlKU2qvyFZK
F73M9QQnmXbTQnvWFD62rSxXDC1hW6dgv3Cc3/ekBAHoBDeEWxL8MRJ7gf5ocS9A
MXSQlrq/Ms13E7ddPJYtQbxtDCzSlDCI9MhHsNKqcsR1SG5D76lAHRu7ta487uRX
JXUD2ETb7FlcW4lfuldqA7AHdcMeZBMnxuBg4+ox7i7W5c6GTwieMTdwPlhKMgLF
Ilgdb+ee45HoNENLBBmsQrpHqcRzQ2CiYidrE7+HHxkI/cAZ9+vNM4JUpooTW32T
foZRiPHGST2SBiyk3NX3hedP9Hu8gJdK0ocWjhQvYE5FnM+kihPDuiJwwHJDHO/T
6HsWHaAtCce3+sJbBXlXRmMH0IZIXx1YUXTp93Li+d9kGJVM0dypt275jSaZYGW5
XvRL0JdiCF7yDXqH1Byz76sbLg7rNZ39L2lb4LNSFeAS+TxY/7PJJVu5UX/9qtjt
IsGyadZRlFyDVaizocoeBeEoYV61/pL1kXIYdGacveSFlhJx2gxLYWdrbYLRa2xz
gm2NdRDRa7RuMe/XhE6Y4lL5/I/L707WA5fjkDq0dYMOSZ3CyJOdZp5ws8a8kC9T
Ll9y9RhlVaNpJJka9dsSJXrGs9QLfhagdK4Q49HPvksl3G3z3oordcmGF54wwC8W
ZxkrppGKIXiBR1RCywsukL8gEyWznrV4S3rgnfh3raOi0KrWsp8j+i/SaYltPXdv
bsp4k0hFYCBWjOX03FZ2BWVDH+9aAF/JC5XZ0JZm/TEZr3it3NiUWJa3Pf6i8OLl
swKQtLq+WsSLxZkvTLxc24vvC6Xpyc3kPoF53C6wAPaNdkDoQ5bEWXS3s4WokCrA
5H6o7wCk9sGIIizLWvXBgWtAbQMNZgyIjb5TbKeUVi4VL1D6vZws1ncBkIdxu4Sk
tN/YooXWWx25yxfmNJcemcUQvIeLcB1jQhG7eRbtXVoFPbIGbfK0IXLhI1/3AaGk
8RXspEL9vmm5TYLmJ8YP96mduon0HcTC4MihEXu7yJ8B8yhCK2ltvJd4ubRtVRwe
rBsiAZv0jzQnA0d1XyyhSWWNlFBHEhpSregiA/Vnbf019SquEYDu0Pg7jNGBQcw8
nIoCIRg6ulKkfu6YbOg3SHLHtLOdnKoI9gBn3rikyEFRfOi7ZWQJN266S2gbHdne
eor39AEVfKzfgyOmKnbeJd1V6FbfePiFu8Mli0ZH6RbIhlerZDBxtLE2qAz81iSh
leqHwuZevc+ZYxRYYQBjQtxsHUrvazeFlrPlBwlJVGP07oIGdPBVBjS8Wr0ZZLvp
7Vtl8BUhngKcMDd2XcIEKb9bZ9P59ZMF16w/bF6L4PQh9fG2+eosjghgFQVAlJhj
ihm/qxIR9G3AX9Zv1iKJDFigtJLDnsraGBHncBVflJuUVHWMI/QKGU/b8FmUuO28
a3kzO9TFhKBx5sKVhCKgEz9frqPpYSET/5S97T6r7egYA18ncmAgJCUixF9bNS2O
/lHO2v8UTLY8YPptopwb8bp1+LJ0y0zpmKjjTGLHEmmr5Z3/ZTtFkCjoNRStfhcN
A88/c+1FlVxmxD1cQSAQ3HH7y5TkHGLSwlhcO1PRFkYZ61e8owtFomV7h4wYY7L7
CqtnzOW0NuCHJh0QDfTxjCh3zfEswRutOO2OnSbnCbcI3ODDkgNUQ8wal9r9+y+d
Kc6ZAzeUW7lu/4NfSTIFoAqL0pbPfl8hgJfyTSjaUyJVivTC0Otn1jkyI2625RqA
zErx+jHOm7Is3Ll2j9UuA3TiH4O9j4M5jNi9hNfyatVBkc2SNCrX79Ycsyvrkl1Q
ajBpl6DCqAQoX7XkHs4Wg/iEkt3oNDKi1g8pZbUFJBqc1Dn6KF7k5iU+6NTq+o0x
BtPf/QMohYR2mDjUfS//7e6m8Fx5uWyo3RRstQK1TPTsctVRW43MqaMJr0TnAqcW
ssSDCsI79PNM4m0WbtkfvrEYsQqeOES1j6cqi0DG9wg3DvceTEYHCyn2Nss4tudO
ZXfrXX+5ELUbQoY1830fcxhf69YskjrOO9QrpbSQoQmVgTY6/MnwHznxgCYBvXCD
Nnu7JwJjxkJ25H8O9yikWzsKwHSy6DJm0tqjK/aLWAvqYhO2m2aZA+dDw2h0pVP0
ypyLYlRvPoJO1QykxRliswLrSH/jmpZcL5S7CpZXGUeuQdJPtoFZa+UvJrxp5QSA
JROt1rhhoH4/DZQ/ouBzqH/Xe0mLdI4oOEuKg6Grw2i4o25Xs0uxy38CUg3f6SN+
nhSeEXblVnpKAc8SoITYFoeycEMl8Pxk1q2GantSe09kKrEExUDUoUpu+1hy7a3H
1qd0xJjASPWVF0nMLmNQvatBe4sLlho+ad39gBOZku9LrPm46P1OqmB1EuSkxD5p
Qvh9BHCz04kXu3mV34yo/m9luBIENs5ae+M/P9COka0+O83zXuYAgyb+Ry2b6kTR
j63hZaeM50IeUB8SJKL9QKOTotcZ1ugeMTTr7VgoXRlhfUGDZbpB5yxhdjfb+nrw
flayVTlja9kghIRiBTVdquCxDA7HK6aQA94+e43V7AUkPBzqUy4WGWvx+w1BG0n6
e5KvCd1c9554DurT8pEHYDCWfE2zGDYd1tf0roj+DFt2UghIUtuq2v2RkkjMIefq
UiYOwdmCJp9keEkTDNFZEz4SGF2P7hC6ZPiHgd2cFV0mc6sGcvOKbrXJQEH/Zbsl
yUzJElqe0znyNavg0t3BJD5FreG6kClDVIXpYjDKM3Dnw4pe3TcLeK3XdjrImq1f
k++prJdvGvhtJu9SmCC8CXIprCUhDwyiazOFCs3NbrNoDkX6IamTqrqI5KEDelBP
BXXu1j5ID1v3i+O2ak/6NpU6OKEfS185zzqBJeEuy88VrMejptLUvrMTAEFdZJ4E
VWHXg2SeUMGc4Uwdj+HcKy3KWlI0jBjssJcovOfX1jwY7SW++rH/h2h3JgOqJqlj
fkDQCjvzP6gzo3FTczwr+3Jo+e09HjYYyq+ToqSAE8xFYw9YIPagOITFyRGNdkYh
MLDW16R1cYx2aisS6WET9f8xe5zCgGX8SAErSGj9RDXqvpX6x3Gm0VhhhWzn0CMR
Y1s12In6qyPpZcEhI4PlDpG2G3TOR5sIAhlDzQf2DA2oGd7OLx9jFXhm7WmmM2EW
ZLp748DOU4L9GfJB0fO+RkYzEHXbqL9RUv4/4ZGlJ6/9KdEeJOx3GbUU0ZnLHZ4H
GQYXyPeaQ02+7ngcfgjhm8Bc+i2I6XQg8m85x44ugAY9+oU/ckNtGp5Y+ucNX6Oy
6BGQvs++E4iQBRSSmqGWE3YDWomJNpJv9jOsht7lfSy9ydATRL7vipyg70ikIgYT
o9LnkuCGK28/eW3rt2CZabhYpU0JC/q0YaD3uV9Mu2yYlvZUbWqBQImGEzflosLR
Mfeyu8K1n1OGmPWTxGKLkGuf9sYt+fEIxFidSUrDSGfjzjhMGzqjQYjwRYt+ma6t
CtvlTJir3cXJtBhLBc0D/rUck3hz1UrYydrGgoBEaxJbN44VhC++QN4j5+ckkeoT
NKmOqYPaaDS4Qht0cHAg3J44jcNCXVczMpZWSFtTl6LKf9j86DTkA0PXBC1zkeGs
EIhJ/Yp19pojbibQdRqrxvk58kYat3oDiA3oQHd3G/NJ8YwY5PNntBmKz0Fqp96H
G9Gi5PGjsrLIUOlS1LC86IUdljkPFe6mOOAR/qNigX3hxCiJbsETmD8P0Gx4hp+7
LKqBtZBMAXhuGstVOjOzqDboi858qhmCJKMK09QmJII9sSgEZYMXiQGG5gCXy3Nq
dOPu1wY3scZgfiwR9qH3KJAmkIXUjtKl0ahA5aXKd5Ms8E5FI8XRAiUo1sDY/C12
IKjcsUgPRYzWG1iw3+bU1OcVBjfXA1LVYjHTEQ/Y9KJ8FUO1/bhmAUK1pLRkebm7
iqOHwH3gRLG/C8lK9bMq2LS6CcBFY5NPHzxepAAGCCpl/Wcwt1ltEr5KUcpAbJmN
LwIHeRhY8g8mq1gqF5bhSpnUUUZPBWbVG90HvV7AhaKz5NYqbEuniAw20yfPb2sJ
czMwaZCjtYyFLEHyWn+dggS3lf/CWoDRA0U8mFO8EOH3S6X3175p5LLzx4SHlmOY
mHxX3Ct2W4MctcCjR1HM5/okHNkhsRIXkWwpdgy1Bv5QUJy2lbhltPK+V07Dp8Me
5HNXRf0yrP8aciXdfFWI/ZlVQ/FPQkqVNLNTC2xNnSU6++2EfJ9xLVs0FWPvQXzm
RypTeR5thKMuZQ3eOblLusnwwfon3Adue0BYj+te2ibLhM0RLgnNlIoacjNYPHip
s6qXczeIijYDsoKsaJC+JiyPzPQTfszoQIGxJHyX43b9f1WhIDNE0J3MToApYj3E
VCR21NiDNAEhpzCooyF1NOJ6BII9zsgD85XY29FOeuyDHzrK787nWoh5LYbNedCJ
CpJMyZog3GUyAY4f7eFh8p0pXF8ZWejf1Z4yG5asyoskaPVivUt6bqUkXKhk4o0Q
mRbOjYJX+NIsgXfh7rlX7rBD0Oro9sTgbKEUTSDPq/Pq4xLK+jUB0LbupjhG++Lu
mN+v4P22hGIDwjoxHOu/JpAUkdomilNtNIdNHTOWaJWGQqEfYCXeO7EYaL5lhXFG
3LPsAG8sbw/iqV/tWpsT/UAvCcnSTCfqL7udlInWFTCKpA3oVMEMJfeIEoG5JcEX
VYozch3+jTllWgmmFKn//5eZw51lbLKdx0w6QehwMdjbJgSN9dw52Hn8paz+/Q++
bRZNtVPyIUEdZJXEpMpeDIyIdmFD5Q3BPs1q1j2KF47sQ9JbnFoJxOwJZqzgnGAm
RLi1AUQbfKX5PipFpGExxYW24oPrXkdhFBooVW5MxWVrMAdGmc+NYpS0RWilYPrZ
3o+SAcfhVdnSsNyavvubBg74a5ygWWZFFC1eWn92mdA7RzsQTNEKDA46GEGdwVKT
nH+hAswtYVY8yMUBeXScy88C3e3Mgya4fUklY2yVviqXbjgPqT6815VdBL6ehcvO
VBtR0u/fyhvwKgVq1wl5Bz6crj8HQ6L7Vm/fBspFZD84gK/stDxwE2DFL73KBf+N
IVFD8GNXZ0h+tkCi/AmSijaOTZnZLQjjfGF+RPpLO+0Raa2fgQB9fXa8CvZVqaTL
jI8nYEmuL8vwocKFHCLi1po1DXSq2XejG5Fvh2iQYpAMQy0/Bk8NvGFU3+AtVwlm
0DEmtvtvDrh8c4Skcm7N2MFM4P9BDrmxDsNYTC5gQIV6kRBpH387bmGvDgCrCxy/
Z4/1SdDHBhlyzFH6RDAhEp/PbOTdW4+fHWvC5FP8jptJ2+uPRnI5IJsd18fBzio6
7ZYQ73dA6Q2nfRWBe0RCy/9pAa1Jfisynutf5bD26VO+K+dLt2rTTGeUP4//ebQx
HzOpNhzay4F7sd1Jm427PxiJsqCg7XyVpuubX/AvuX5U13OJ9o3Y7N/69pb9r4VS
+mmhRrDdEztuL3gL9ZyzaL5XA6hzVCSHajDN8fwhvH8xN1L6ODvJpnE0uNA+0ymi
8/baYgXn7y1jQXWXkK9j+x7y/nqJoxQ3NVXUAG7x08vP0U4ZyMXtpT39p7vsLnA6
LeJQ7xI88cGPUvWJH0L7tHXah7xzpAwueojOKr0YGACXh2xWcevDUnPc0VkeF09B
0M1/SZ0xVjP+l4jwXDYL3+Rdh39Eax8RW9TQBbXN1GZ+FCdltGOPC7M03DduShgD
a5756XKDo007bKlp+TQ7cFOqB4xnfxqH0y+PDBz4+I30F3trW1J0JLG7QwOKEO/k
/iWSQvrDIImfWb1Rdi/1eHaHljPzZPHq9KqMl7KZO2CqDNzbXNFCJJet8gBqqBS8
344aJx/PcBkFzRXjaJAdBLMNfL9iNNm2lwlagDV22dzR1zaCq/diH/20wN6cZAyD
s/keXHVZ79ROVTDvUSO2OzSUjbTSiEocHVL22pMuVmD5yZ66WN9Gl7/oAvyfrDR8
kO/fAHm2e/OXcV577TABlV+geWDoKcx3GWC/I3rk2vMNQv42JUx94KkKV8vzIagn
fAYmjuzaOCZr77wKowVqA9wnitWFgdj7fSQYZr8qrSg+j6fcrQpPyc0XNVhfV5PU
EEWAPfF0g7y/qgP9TObvIDJdXtj875R9YxKFcMvDaZECZSsL05wqdxKW7tRBMw0J
b3KmGOPUE0o7psVMRzq5HJcb9Uo32v/m1/BAj8Zvorsdm65IKIp74VCSCU0r8BOJ
Vyg2aiWJye7uoQpy3DvFIPXq+3EYy1nWJOFr0Hj5GKIv/UeC+PAcY/TNlv/DHbqy
HdADfTCDhX4V+uoR+OV9ouI7pBXKU4Y9Vui6fLiLwdhFuOXDLvwohPfYOctD5PRa
UsXybPoNmqGqKGPpeOjDCRW4ikQ1P6hzHZJbfTcg0PSZ7qV94LvF7YAgaBaZ48st
j/ZDtSJEn6t3Q23lA72IKaGkkodinu3Uz1NVvbkVQCWuPuo5VFhvVzxyYySlYmij
Zr+IATCW13qOhMNEMtuo9GKEWhx1Oe9UDwtRcz5fyn28bU8vAnZuLKjqqeNb8Xhv
WMe+r8k/LjOk1EgSkPb+hKnvyh66dtIgVT0UVVFq9CedlNREXL0/PindfdCbimY6
lYqQ8NqLyqOU14pk7ivYyYMi74/pgODepEZ1QUOFHsTyemTMP+mbMs3lMrTUyEet
LsF4eRDlotG2EfxFqVTF11gecz9W5JfrehyALyyWgEl3bCPXyR/BNlNDO+/H7rDd
knDpRiXnizCEHN/+F7UY0yu9hilCax6uLEjSedWypvn6/git0pcQa/N/kpwi3rb6
1yAxIOQEYxSjgu5LvBx4xGJTnV4XIFZAfFAZubgu/WBXEupKg2Jz1nITrbPj0H27
gno13OUWj6POhMIG1Q1r1mKozwID9LWK9ibOHcq4iRdK5jFG2ea0UuTgQ4CA6wmd
UGM5z7zPDS0JhqHOjvBR0aytkCML4e8LBMuRfUXu5JbIi7jL3mpJlXXaZ0Z1FnZA

//pragma protect end_data_block
//pragma protect digest_block
E5G8sfAdQQN9lfOt93/dH1vBi+U=
//pragma protect end_digest_block
//pragma protect end_protected
