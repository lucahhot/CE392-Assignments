��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�:����R����	���^|o���6��}�Ap�����`�^�m,��"��d[Vr9��r'#v{1ە�^!����d"A�ҏ�B��֯"���O{E�I��qi�[�����\fr�
Ss��V콶�c�Y�B�d�)���+���F &����mi�p<�/�('a_���βԋ+J��8��Vo0"`iӧڃZ}~vtH�6�s�+����,]9I���u�I�<��$�^�v�+�RL�?0�v��	�q�ɺ����[&R��^�\��<Bs�������͎�!���&�a��F��q-���$'<9�I+4�	h����b�=���c9��6�u�-'��s��;��;Š����z���r%���n�ʙykz��(9�ᳱ��v��_��\^�dQ����R�L�yI{�}���������tY=>��@,�g�l VKB�V��%�\0~s�I��.ƨ�?S0��|��۞ב��I�/���(��`?���<����Mau�m�����J�`Uh�>N���2o�p�9UQ����ʷe��,����ն��G�=��0
˥۶J)�;��X��,�E$}�q�p�� ���,����;#��v�=���f�`�{C�c�6�%����C�p�H0�;�ڃ5;*�-"�<@U�v&8#\�e��'oT�����8A��9p�8�>�zT@�6��=���� *���9��n�k��it!�S2k��ž5�s(����o��uP���/�\��ϒ��P�����X���1�b�Kۓ���6U=��&��$0=�^�hN۝+Z�8w�}�τ���J�.���W^f���4d��nO�E	�U<�0�A��-�o�ЕB�꧇|F~#QOp{M�_�Z|f�kd_mt��U���j������uY2�^uf5?!��L�?0*��5�sX�$��5B�����Y�L���2��E�hN��]��'i>�Cf��q�V�GhK� �t�!�~ �]'OE�eN0X�b�V�W�D�����~���y���\*�^���=��k7������	�ȷ��
��J����wj �Ù�@=�'=n�_��e�b�$`Ԭ�@ 5]���M�A�%�۬�q������Jj(���Bj?
6��,�X��-�K���b뚝�涴�%�.^���=�-��%���x#,[IP��Ԫ��_Z��u�y�|�e!�G�k`%Y�L(���Tz�G��~�s7���
����]|�5/����lK.G�����d!� _�~��\(p�EI�~�?��2y�����W?Ev���أJ�8;ء��դ33�=�6�y׼���|/�i��I#c翧����Ά�ɠV\<�p���Q��J*.9���\hhݤW�]K�g�ռ�^����SP��#�;�ȏ�HE�H�o�@�ͧ�D�I��G�jd����%�Y6�,��k�_2�&)Б"Ϗ�p�!ǯr��d��Ҷ6��:��[[Pv#�b��np��[0��U88�l���0��x~��6wH
>�]�u�������s�E����������h{�+�b��aIΎy7_�����A�ۙ}���Z�u���}ϵ�M��(T���,�{ُ��E���CQO�v���v�T���Tt�kw�G�sTaj���v�E��h���{� �)b���̔��=;UP�g�4W�>M��RzGF������$��\�ш�el�q�P"
�j���E[c��^7Hx�P%Cs��8Vp�̭?����s%���޶΁�J4��y�2�]n���Pq1Oڐ�Y����W���w���f��aWc�dk�B�o"����q���>р3�P�f�z�Y����m�� �̴�沋)ѽE}L�b��(rJ�`cz���oy,p�_p�j��0H �x"�;Rw:.W~"W��T�td(�_�,w ��yʮa<N��#P~���vt%��l���!f�,����l��?�(b���@�Ɔ��8��e�)�Y�qQ��Jhޑ���!��G5˶dYT�F5��3K*��9�I/�������C�Mk��G��o$���P����H�0#�y�8�H�x�c�h�L���[M���B�����E��ޱ��&�6c��Z��%���s�vK��x�T������x$���TL?;Ԗ�/$�P�ew�	��B��1�p����3���w5/��a絰��7w����Ik��{��Ʌ��mYiȶ��o�J�E�]����˴p�u:�x�48I�zo����?��b���|���]�KF0��FG�.�.�(i����d���	�(c��72\υ4Y狀�N��ΧM+�z�7�)�X�(�n3�?��A���$��蘥�cbPėz��XҒ�Ŝ&^�C b�?S5ҜG�}h�W���e ��|�\N&S�i�È_������/�~�pʩ���Ū�,IR7�[�o2"�M��R�A;�;��(9�Eִzu�5BR6�pR4Y;��b�ϸh)����<�O\�ڂ=T-u��%Ƞ�T�e�]9����4�ԑ�.?0�[��/7�̧��f�q�Gsj�*/�ͯ2��H�a�\��j���n��Jv���4_���
�̺���;(j� a�[l��V��m�|w-^����x�s��n�f�_���c_�HJ��ۋ�M��&��3�d2n�TX?"��@���	�4��eJ&Sݽ�&j�h�vN*[ժ웤�1I?s
�7��v�A����%���ƅ!���I>�We΋C�a:)�D *�fT����$�z�f�(��t.!Ȯg7�c6y�w;�O�B!5RL�z=�bk�)��M�~Y�\:� K�~��k�փ,�k�����Nʂ�Wq�B�s�`��Vy��6�3�{�A
��Ia�|xZ��G��-?�O2�NN(U���Œv����P�C��^��	���x}�̬��qy�6[�wI�a�{�I��t��ðD�6������7DONP��RL�N����W�����1M�Hk��/{,,CtE$q�K��#��NJPҗ:핶j)��Go7�.l�a�~�}Sєͩ�I<,7�]�/4�,�r����������+��Ѡ�˻��.nMA!��O�
_B�%��?�_6!=�o2 e6�m�k��G�^l@��F��N�8z��WV��d|p�?d��1��O�V�
��㫍����H����Q/��0�~ċ��`�7	�C�Un~y��6�x
C�=���H!�,�LT��Q�vN%�Ӕ^����bD�:���Cv��d�w<J���J�ZN�`�A�[������*we��6�	�
fΖ�Z��K��*Zr'V��c��7�ꛘC� ��!����6��	�/~ߋ�K��h|����fg^�0z��˸�(��1+&����i�\�}��kRd��˛�&�st$K[f!�=<�Z��{xq;�xd:\@HKD6i0d	��Q�N��ɋS��K�k��	�ϥ��gmZ.��T^��>�D{mo��ZK�"�k�j���ǜ��J�ذ�T8=�!�X^�n���E����ЃI���2g~�O���J�7�ߝ�
ԐWifQ��}�!∶��rY���n7aj��NK�g�ϲ�۾�Z�ϼgHuU�b(,W<j[���Hi�����{���S�Ow6X&����Z(R���#k��f�3`%����L� �4f�Y�+����.�w��pn�AcEK:�^o�_VV�te��$�)9�+���u���pC6���9��s���"Ez�q0�ER��h-��n��}Lgv}rå�`mE����CR�_�G�ޓc1�/M
׀ zL[\N� 2c������M7l���ZE����삧��iW̓o�X"�/����|B��ұ�n�D&wY��D��Sg�?kR���$�S����̀�u��Lש� e?�B2�"��#����-I�`���_�/G���J�{�7f�#����	y�&���z��nИ
�v�T6�O	�8�*�O۽g���c�>�$�=x��3����E,���o�Z/�O��:��i�ٱ�L�@,�[�{������c��D��-%��*l�:�}�c��Z�l�������
���|I��ŧ	m��u7I���9sw	<��^+��~�-��K�:������[�j�Tƒ�P�N;�����*�2���|�ɧ-"A@���צ�z>6dO���W�TW̞��c����, ���������*���?q8�D}�@�bnW��$����H��Ol�"Q�C̬�H�:T"w���9���鞴sCCn�ˠ�6��nGmF,dN{��ȴS%�I9�Kc��$V�̔�ު��F D;*��t݃,� �"K��0n<ӣ,�?|�����25�qp9.̟L���&���eeR"ף���`��>�Y{4S��S�֚�_��L2�.=��]j�v��1��9*Zd'*��v�����+L��2�k�#���[�l���,���_$>`�Y�^�8� ��-D�?cL�̥ ]Ni���n�Q�/���x�� F���H=,�YQ�V,@u�>�����šL�K�ONw� ���𚢩�O�XW�&��q_i؃,��@�1 �S�|u��j��ה���2�Q�3�E/���qH t4���}t��l����I�$w�#�9J��k��Iݒ{}q2&v*����a�`eƻw�fNǭ�4�+��ҷ#q9&P��N�x6huV���"]H-�,�n��s�q��"���5���iT��c��3�1�=���L���� '#��ж`��I/��o��QA$_�3�H	`�?@�S�9\g4x�[�@�K%�.~1n�/���5}��94$��X&�o�h�Z�E!���.���' �v��R�l֋_�̟�n�資e�ӏ�ڿG������L�YO��F�G ��sS�o�n@�K%_s�"m)���A�vcf���.��9�ߛ���g�@_彯/��RB�� �s�G2c?�XU��3h�R�w���Ǚ��J��IǨ���B�Q��%��d�����A+܅ts�� ��ڭ���L���=;���	�J�(��Qn��^�k�C�I���G$v��no���>�p�= �>�F����!3��#���A�R�f���@Yp)%mA�F��*;Y��T�{3.@���ǎ=CgS�r�1^t|KǴ�p��X-ӌ��S!d��g%��!&;5�������0�q� �ߤ4���L��vO�	�x@�U�vYտI���֠�~�䐢D�������'���٥�Mk� �J1����.�xp�t�ݿ���ó��"��Y�jZ&���(Y���j�;vA�_+z���rx��4�	��ԇ0��y,q,.��S�?U��7��n{e��^����Y~�����Zz;���i!6TE�R�s[�B|<�h�he���q����כy��4ln���B�kT��t<�ɑ��iv��tIq��ݏ2j�7��+�}��3�q1L�ٖ�W	��v�2���4�i�tx��l ��5z�� zIW��*�,@s����`��C� x�ࡑ�&�䲶%��yL��y���B<;c��4�*�������5�8���
C��B��,�4�L��V��S����S�u�
w�s��rSW��m;����O'�����n��*����20�c��Y�ʺ�ꃭ*ZG1���a��c���j�����jm�$h.DI�]��tci��Z��DI��
�����WD��9��<�C��t�*p�IX���Z��}�?�8t���3�.�4J�H�Wlp��j��o)���Q������0q6��6"��)����f��{��.��e��6�Y�f���IN9t �@)����%@n�ɿ�Y�Ӄ�|/&�&m�MCWuxgn�"���g��>�Er��=VЅt:kF���S�9g����(����M�� ��NSIQ8�+ae*��_���G����E�B�	��rmf����Z<*0�g��	�G�q@���[��I�s>��g��EM�_T�٘**�m���4'���{��K���k�TUjU!V�����f9��R��
�H�7�7;��H��f����}�KFfz��r}�Q�m5��(��Qp��FUJ���aW��D	��*��TVBdj����A�tX	䵾�� �~.pʯ�0Ss�FL�� ��!xs�\�LH!��D���6����Y_��%�+���hu�x6e�~�b�ŲG`�,.ٌ#������H\/C�x�l�Z�:!�ƒ#�U���A�,|�fG���O.c�������?���v#���nxN�6���0��J�'l�	|��L	W�/��tۢ���.s��Ǿj�X��eլ]�?7n�=#2۵͂ ~�zԂ�f� uH�vg�3��*�d���d�ٖtGq���'�]�@y�#����ء�x$�������{�0��&�WJ�V�𖥱��AI�(Z6�q��1�埾@>\�� ��__�ХI<����- >>���pyU�ó+8K?�T��h��|�̋uZ���^��|w}��TU1�|�T�JNHmʲ��|�s�A����1$�ܼ|m���j��	�Ow�v�BLi�J`�
��٦��^#���lo�D2���nZTV��0�b��PM���&��5�'�rP�L���m���2�~SCyHd��wW_j�ڞ>}e�f*%^тB����g������?���_t�9�Ǹ�2 ;�~C�n#�"����i ���+���q�K2������Rݬ��yF��`��׵{w6�gO�i%I���
���_��l���i!j�<�)� �*N��O<�LH6C�Ӧ+;L�h���,�2�!�N�\����&��p��A'-O��S 0�	����"9��ڻ�����4'��j%���ed�M�k@h)R o���:żԪ��0������H\���ÿ�@�D�����[���z��Q���_� �\�=�/���H�3�:7{�)Uc_og硄��(�n����׌��A�彞�
#?{w/p�e(�'�}�x�6�%�&��b���W����r��ހz��\��[����U��ծ~����oPn>�H�����js���,xR͋V算������0����x4J>��
7�abꨞp�e5�E9 G;}^�vbB&%�44����+⢢��(c]M-&y&L�o�{ ���0�	��/�:��;}�i?G��w!~���֎m��0L�5�WԜ�fh�{IY0���M�ϡe*'�:\l��xX�LrD�I��!�	�L�x8���
G��	�M���$>D�y�`$��R8�X���e�v��b��Um�Ξ�G�KĒL�Q�i���	���#_An�w�� [�\
�Va�ν�vNmm�����{Ah���0�`�S��⭊���WϲѲ��n������{��.u�C� w��I�yK��'0��5�Q�eD��w��diC�\O�'�����!������a���n��\�S��3��p���� g�
�E�Zި\,�K#���d5��L�dn���*Ydi���,F�g1Z�;*v��L�1Q7��K��j;�i+�՝'�hd�	I�d�1�c�"����b ���o4�	E/۴�Z���� ����3�0R�.w�VLNC��r9`ߚ�(vvIUOJ�rʖ#��Bڣ�*5A������Nl���~>�	#ε�S���a��������$&eй�*�T�H��S6��5�F�;+8�/et���{.j�� S<pyѡ�~���c��f�x5����Y���!��Qe�J���LPX�2�M�b�9|�7�l��BV�D
�G����Uइ�Z�܀��� �]��`!N����[��MhQ7�Yc�&�'�$�ދ�<֞X�>�����K�3���>�b���P�2��8��q�r�M��׵#����+�[Fh�3�,	U�jO���>��y�?%�~��.诫7$Pk*6��w]�����P2��I �0E�D%��Z�)���z�s��^�@���ad
'%a�Q�)�ҏA��Eڍ�#�����)���Ր��3�*�
�HǍ-[ �k �\5�&�g1�3�%��m!#��ߺ����/P���Ô���j���
UknH��Io����ɏ(�\E�?j�_�����X���4�`�l�-�����4�&2M��|�`�Xۘ�"��i}��0$�>�
�����y�b���!�i�̀ip����)�U5Kd�67R@@vؾ>~����G���q'�����g;��w��ԝ\7�l��z�ui\���i|4������;���u��Iւ&�����Pj�6'e6�`4�u3>�*��*�,��n�8�t�����G�����1g۩6���,A�)P��`�h佮󮤵�Q��Vh��bd7���jR���T<�U	��QXx�� �6E[�Jз�깉��s	x�V.�E]p�X$H��(�ZM_��S��A��+ȵS�LN� }��A��|c%�nUz[M��������?���N��u胿�"M����\"�{��Y6+�^F��3�ο���4/?+�v��»%���V�ڠ�v�z��9g?�ɿ��� ��Ai�?�j���u��	<@��PP\S��++!���J!��t�������%��k �uAy��rq�n��s���'�7�w�Qy���k�&�q�h[�VeB&q�7�AQWeǷ�I��	���<\����	��\T���h/�U�vJ��u���v��3�"u�gʚַ��j��~m��x ��� ��t�����5���( ��B��e9#��~?#;(ұ�;'��#x��?4	0��$��8���������a�i���.c���򧮪�x���16^�
]I�����AOMdZr�k�F3y�}�/�/�����tf��=��Л�gAs%;{+�N�Ff/*aO��r��"9��=->��&7��i�=
������|�P�o�Y6���%�O��y�n�rV���8�9�4�����h���R���sR�����IT��bA0*@5���F)`+-5@��A��"��+���3'���K��.������%���X�3��Uj¡�,"��Q��H��,\̒a�-x�0�U�pz6��]\}{�y0�Mr3v�S�fB�k�`뉅^�;�:w3�-{S�	�D��g�w�M�w�R����Ҳ���-���O�db��G̾�_۸ʆl>��no��(���v�@_R(9)8�yE���{-�����RI�XLҴ�W����yQ��(,������L�-{4��[�w������"\�ŗCtq\���'��>ę��\�zp���N�,�ϕ��*s�C�%Uk� �>~�o�oO4=S)���b�ͤ��]�Pig��̠)���z>z*~�q�Ĳ���Vg���+d'�ʜD�yPR����p5�$��n��/V��5^��A`�.L8�e�����-(�rB�D�%�����A�2�@�xaȔ�$8��m	�|;�4L�Ѿ���h�D~Xq�R�����|�f��t�O[J����+`�~�>�D(3�,���	��o�(�3P�0�t�ƭ���|tx%�*uo��H��S�8hD�fp�)�k&o�@�ꗬ�L�t~+K*��=��>��Nt��;t)/ПE��Ѫ����`8�q[蕋�<�KwC7J�BG��4õ�P�s�����Œ�ރ��b˒�DC� rc7��l�4�~>�r�N�;�"�ͯ�\-,��@87i"�2Y N��0��W���������!v�v��=�ͱ�PIN߸�5(���`�oa�ٸ]�&W�H�1Ϊa�Q��f��D#!�!�O�ڻ�1��+��/ɗ��@�٭�#��<����'����bt�RJ���ʏ��U���^��-y*V��R���ERha�)��UV���Egp�5V������1D����/���_�M�&�O$I�|�!�"�S�7#D����Y��A��N��y#,�3���e7��T��������i�ה�xZ/��G��*Ŷ������^�MH�xf�l�����Y��ST�������i���[��>H��rY�,=~�ן��Ѳ[�
&k:0)~Qo@n���BWp�e���Q��/�m'�7ggtp|����O��P4�?l�,�[�?�����F:B����E� �=�5��Gl��]��Mqc�Ke�:QD�u�Ɂ�yx��F|�~���C