// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
P7Gk+6sC+ephLQs7r96zcQrqwhMzfTDZ1TNeQwQGZL20XP4rCmtdjQI9hdQi7tds
APMmUNrji1MmhWfY8nEJz3Hl/Kbx9qVLVEkxZqqE6COobR0PcaFbFSzeiOmmsnmj
jBSzO4PDaHhju1aT1hwKSshjvjLWJOxGcsZKD8DmTFA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2112 )
`pragma protect data_block
aooWXfjgKRTEFSgei6sU7HmW2K2gTBBnXmxnDOKrDIdoWqYfCNl9xp43XJvDLRDO
fMwOQhJ9Td42IggVAU7MqZdbWsJzMRag/m+asc9TZAXIpRp1IMgwGx8M9Z0rxcz/
F5bpV5r8x8YoPy99xWmY6vspIzGb4B7I7KwCeHM7/nil8D/jGljcqXh5KzfCAIt9
ZRSpDNxbNYdLQOGa4oFu///KPIveg5Q0fKftRhteH5APXp8Mn4JLhs6U2kY1zlQv
lIIA/nKp5b6EqzEZGDl0gj7MAdlAt//kzm/V+ueXlohB3+BAt0kXqylAB12YFL0J
+R6yW3HhBnn60VpWaJ7usaMuh1YG56FcjKTIEFSNT7E4/NU5pEzzf2Ic/D5nwpHf
cASv3l6a2h4+6UyHLeY5A3EyzQ213QgaogggUAPOfou8zh0JZfhYgkZxQ3g2CAcX
GqSezSMIakoYTsV3yMtQmL36sdSwuYcUryzxKI8O8P2oJf4doFtJveIpV8uw4S28
4vI2O6q90gCIU0FpYHhQ/nkb+poYILvkH55aCHyQ2qZaKbj/yn9LTjxQJptVo9ua
7YuAU2y2qUj+lN0GyjMGcVD5a8/3O+qy8pHcbXTmtz+DSncD2cLH27P/9KCe9Wtn
gnVq+sjFqPVdhHg5dMd8Jo/bEaQdkpYYUu5L2O2hyaWSWJ4pKb0tyDs1L90QzLdP
B2KdFJ7rFadXxiet0v3+NQzxDwNLW164ubB247QfHkDeyXRO70NsRYmxnKzThY3i
YmdOag/cyvNmZSx69rXKZ4fdQ0964HyUuR5sX1UhKcEVLJIvMg49MC1v02POCdEf
y8hs4j3AJZhF0ELsVary5J4kVJFuzYrgbpuygdV7mhbNPRcTt2NyKGjr7WLkFIBA
q30Z5YjzckZ3CvlUEMLOEUMK3BWD3SL+Dp2PQZK9Oz2b88a0xK9Z5j6AlYFxTdiM
fSsnv+PI9MDDnkVo8WXnRIdCfjNbYSt1DsT9joPt8wZA9LD1UA3HOVCQE+T+KRnm
QNWYNsLDh+qgUJX9GGluAwHo1OBgRRjknarxWd7AfJeNbTRI9+JqE11V5WdW5GNC
nTEi1hfiCCyjmtXmSWcjz7f+IE2Q8z53ViziFU10bCLmQDPPtqmlUNhjwqUZTH4C
tzhRh6QcyR82E2DDwl1QPZAPG+adGBYvPsO2KFZ/gbQL7KYpOsqG92KGbOnybw2Q
tKqxM003MqLBqABXybQlkHQbWUdyGa57zskQYyaRjd61OpT1d64V5ujihAU8i9ig
m/3+DrSKyL46jqJeDBsdHQk/pb5TDTAAORhGhoNcXV4rpKxPYsahk6Uhqbh62Gq3
CQzgv9JnnZyL8jFiwdFK8n1A5CB8oJlsM3XyAmERK8rhGXbcOX3gJ1Xyb5guD/PF
xxUOWKjWeGDbD+oBtwmig63k8IFLqaFeM1anKsHX503jFFJAPP71Ggq9EnHqhAFt
x5Wd2F0A8e1INhrZo4GUrSG6Tpn+w2c7lNBMNlFQ2Mjwa0MpVShIyxyfFLI4x4FT
EeFuHm6PyP5n3m+jwD1H04zO2++uU5Tez1snIYT6WxeMja7nxQVIgK9f/TXotDcj
ZuEokw8Mr6IYxhfI69Rmy5BkPttqSIfy5ygUCTGFwmaCeKcmJXR/MhTLkhuv8R5G
3V64jVfIwgc5MeNXW7FjmTcKNTfUBWbRDP58eOT2jIZUUerVnp7s7VI+7iyMg256
+iW86bFhei/QSi4SbdLx1DLhkWFwqnzq8jjK0XlUpiWqsDMc+kruTlp2w5IjGCnA
BGwUmFr0258jcqohrNX/Fc29fNc9yq1en7cplxN8a3nGVDDwM0moCrQWvyiptOFE
RKO9CCemLe2EFuMa0+RGp3PaAMuBH1JDrcqM19mT6Mmi25jnqZc9mFJU032mUMzy
ukv9l9X/0csg15+ErociPiHijh5t+R/HAHTp7PZ0bjBGZHfeDJb4RJowZp6xws8a
296HErYZsgQSAUxxEskBEXbXwv5nvV2nyArdV2FaPLklkKFFClXroKTtBbf35EGp
ifqwd1wmeer9j+Xb/LCzhgPsZ6OnaQgyNiij42z4g/U6U/yJEbOfBUeS67e0G6ZB
ARxxDKUltnhMLS6upiyb6VAOrjib8LXiYBIVj5zAvG8tzvEwhbzalCd6jLlfSRK5
8czVMrBlM0NGtJyg7Wsw433HSO4AWtvbaG3smQ95HkDLK7OFMHaiOLTaxUEVjBCo
skWZO6MW9zc3Ql7tHlb/BO8d8NqI1BAwEjliRkpc3RFtTl8h/66gKx0J0A6e8BRS
Pq9qi1F75ubzV1jUE+tRdTz/5jeD81TinyWCs37QmsKVRbMVghme0iH/gDKtDSec
CKngvlsqoy8YK9XF0QtnCqYMVRQhNa7CpF187m0ZbyFsC98k8sGAQXF6H1CiONR7
9IIFUDn93MBJ8rLub+nxfReKRw6qC+3qj3HXKDqLZ41AJdsG50wnVE7YQ41kuf+0
Xma8JMp/GP2jIyRa6CW/JB6HIcuds5RNJ5cdkGOH0AJQARJsK2uCGL3nPufB6ZNt
7Mrmhx/2MkXoSN1d3mT6Wgwn6CkafdTABwaFwtK9HHGqsK3vy0e3XUYJJLsGxUDV
r4gL2TyGMMe5ksu1BHGuwzDmq6GG0fI2LrWqcuaF9J3G3ZWREsPRzYAkpaj801Hf
FzjkbVgROgpLN2gIa9k4pvdwJwj7/DaAJzkB9aLELU93zZF7qBDfPa7qreOQFYbI
P5H4Jabhh+XCuj4p1hWaG+ghALjRpIcV/SbI4c9vOQ6cQsyLf+8XePU8TdjjO1/4

`pragma protect end_protected
