// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
bU9Y1j6I4KzrP584zq4fmlBJcarmrmOHW5b5wWs7dZFdGE4XlLcDyKCeP+SK7GGF
au+cYJJIRomU4kQkVVxylCBcnIj2WdhN0VaxYW5RkEwgl8V2kkisJm+bN4vm4jPF
/Ej80B8kBgWPscQVi/fUECKG7RGBEjWScpqrI825RzhRI8iYrFm8nw==
//pragma protect end_key_block
//pragma protect digest_block
9U3GoKk/1SdLjk4YXcBjjjRr5OI=
//pragma protect end_digest_block
//pragma protect data_block
KOkN2tG5KXsEWliL8ukBodbF51Dmx2otEX3f0v16HzxQ8QUR340EUtp5rDeGBQ3G
dptpdQkdnhaCPWh9Piz8cvacqBc08/PysPO5zz2VHnho1IjYBeb+96Okj0fya/be
j3m05TiXgSDIjGovq/3Q3ASE9u3aIa1RS2np05qwdPuC1MSZPmpA33jKQN5ghJ0h
7bMvT0Ne0ZEPFoUxQa0lFXuA7XCsqCLDHLGqCFkKeOXZoVlDaHOaqxBdUJhmD4e6
r0BrHxowT90sUkfkAjWHUu7CIpv/tJL1My2Quw/xpkm8MGioeqFVRoAjRdJwtZp8
UCovw9wmph3t6W0rH8Gjcx9/lkf1MCR6X9QPDZ3TJS2MjrWwTd5ZngVlSBU87IPa
pMbho88LyDpKT60C0OzHwC3izkP0/yPDeGtMQWrhEkIasFd6ZyKzHq9ShCql2biH
w7xRahpV+kz/SN4Pe431rwq2Ydgf8bS5WW8YfDSX46SyDxHkVd5CMTt7Can30chE
/+QN6fHGDAruGiCUatzftVESi7iNwK75hzgeNZxWZwHJrA60gnS6W+TzBB8JDesc
/FTHYyX1otJtXrJoHUdrebrztGsXIrqgAF9Vz+cv94zF2qRkWuMTwzaEATyso+cI
a4I9CBWKZb0kY14gGX1zbC0h3miG5o/tHQ2bwjGD5UIVICCf1y/haEVl+CZOUrc0
vcOI4H+p5wtPWRQL7Di7T02WR02HP8N/P3okgV63xqt+MN+dfYq8b/nfoxKBIraC
Q7B1wHkYXthZHuqIWOf2scZuBOdH7OXL01ZmKy7p4At18GkEmtwQpguwMmULvxdc
CeFyAnAc9cP+7WuH7JCSsxfLdU4K5PjP/jGp1fvvARhM8HH/6hYohGMgUAYTUdgY
uNVHtrko8FoAd0atQLx3A8YXhHxfQFyaafY2cQX+OtZgyqrWBLCcioy2KiWvCPsD
TlWGmPyiGKSYJN/r/d8Pdh22umIovLo9XsHja7Ha4D6YRnn5E1MRyWKf2MZsRIF7
RnNYZ9MhNTsBMBvCruUoc8rIdbqS21zQjo+430iyng2m/Y5WadWRNL/aGnB/lUPc
FYPb3I6GDoNYGT8E1fT9nd5NsClTeVUmsM8bXkpULIDwAXtqEbijWtDXJLos6VjU
SgZqjojU0r3STLO/wZ2VTOpmLVf5XGPb3p4WKow1Oc96KidWzODqU/ZvaMlW5Dw3
YQEmi+Yk1cOPKIMtJnm57m2+8CQ+Bve5NwwpFEXOohdL7kjfo8ogVFXrkPy9lmoN
llAjxYwmDiieSudbBQF25Fg0lRNnoigLgOXv7B8jWZR/9lLTT8q78WUnoeVz6e6a
vXC7Q7QQt4mXyK4YxxDtfNaQxVo4i/MlvfljPIjRdR1imGGkFuxLAu/qCXB6NKt/
A7u5rI9Fq/gRsqydjdsK+zoePikpr1o27AohYRCsubhbrOCEAcGvyRsQBKE392ay
6oHpMu+GdGaDhHESbyHQOSQSQ9rHxsFL5tTjIz63IfMHbDeXbq2zGFN6ML0DvO5H
h5UI09Ul9Q1Hezm4v5YbDzQ+3+mFHHLKpVBvy5r1k4N/1EDe1juUfnskUiA366LP
f7Wd0aJzT8qm4LtxAvGPpPq1CQ89HLAWu0gr/jmzVcvb8YUd4VDXQmQBq/Hj1u9k
xhPdQbo4D7bu62fwuBDuDLYANBiyBV2Zv4KhGZwl2rH0LuNl8fNzFo9ncXgGPXkZ
yueRUOi7p9zvLvqSMpieqGvVpvgua6qSuK9RtgavqUafXxtO88kiRkqpoeYS5Wie
Mm0KdXWGPUx8UOUrwbkl6O3hopCUx7VIBgb+kNWBQhqikr1oLRHA48P7sTAQ+1/y
Tdv5cvUmxFiY1ZurhHOdaQi3OTzDEc2q33oJdc9UgMFGvI+weCTo/rTIneTriCnt
939ORgRTDVhYBUTrgYokbfewq82E7ZK45pBXlsr9TIQc+cRp0QXX05Ag6OpK1Aqf
FSE0kJQbGapeOjX3c40oTLa4ZRj0lp2ZkmLHhQtH4Tl/pq1gfDKP7qfaTsCTOQ6T
mCGGTcq9gjMz45BrqLLEiqncbFO1WinqkckobvlXoHUOF0C5nFv/quTD149i3aEX
8wDa2+b9tve3fr4xnR23v0gOFUrW0PTf5MakaHlblGEhg0tRnCekkl/AlfkJPBDR
IU0dpsEel+YfHTmAy+XUzygPbVnG8wXXaJ+A+Oc2uRxfbO0z/L2c7EkKbiyvCIrx
kDnkkIUlLMgXja3PG3MgjKhyseyM++QxzQeaMTP76ZOhk4NU0yB8kfoaUKW03Cit
Fm5q30az2KPhlPY/bnTamyE0mlahjjE5PoNboZHu6o92SG+hXgUZT5l92vNdfxgl
UY6yR8qNoL6UujZjZ7lGJtFm6hu4ssb3jaKP1XbyWP/pVGb9qSd20wU8RyIooLhy
yeTTi4izEBd2ZbKe+VWWAcLOzo2HAczHD2p4FhRr0oAFNoMHGmo5oDoAtYN8TDfx
dcvALDwm7xQq5VkVIsVTXdxFHaWmANdoiag4yKBfjHfkiVKLNB7ImuC2ZxpvAyBP
f+qNPrwHY//VFDE7FJvntJ10LrVb91HIwVIUrnYb6Fe7OlZY2JQ9VvWD4MOiNgbg
YsX5Dknc/xJkx4fESMpnrsCZNBBW12vCzST6R4KJdMUPpwLWjELX6+RpnIGivs7Q
JzFNgvCTXuzIWv/HdWUTE8wqJo/qzYzy9ZdS0jW9lxRsPSAmZv91tcxtvtdJ8fNA
knrC/xxYVapqw/Yrh02HeIiJPUKGUg5d/af4REZBhxW6UxsP/nVQG0vKgiekED5b
gChXSwGe6GQH0hdibpEfSQQifV4Gf6+PKBQPSI6P1/eiUHlaOx3MJ1F/NJ+XSw5Y
JsgaOxjCX0f/63E/xhIx+HCxxYer4phRoPEJlXPksu0sH7kaFftyY1zwb9iZVbg8
qmZUCGbPJFF1l9DMriJwfwd/E0hiIoIxrLpMs0+nzev3RILWm+jodDppS1pG/WVX
JUZFlzInZODWzgK2NreuPxVLI2CibM55TZTYRFXFTN+chkV0H0zzUZW54xuQawno
kYqohuSmXl/zjCB6dXHBV78qZiqJQuBNv2F0fNTfZ3DOX0LKJrKFybJ8N46mrqrT
ueD59qk5yYNw76HZN7ZkTzSl06BjUVeDeEu87PJGYVSKoWv+ZdeSZyqgAe3lB+pf
+7gEW+kUuIDKqq002YevjdLAsMONl8b9+GvYTxukg7mt2koxZ5fTwAKmYbaqPGNm
SdmgzrBCOTL2aopuV72GpYmwV4tMEUyDIzC7/D37/s65CE6GOaFn5j/w6qvMzlg7
GElCu2FMncA6IPPxmsSDyjEqgGrJfRamKafxCHMIES/Dz4JnH0N6J86+fU+FAeNQ
kHG5Fhen3qvlgCD3dPl+igzKHXt1ISUswaKcvvyNS99RbWUcudtvPOHoMh3StJmt
r0RXmsqKQcuEESeJwvK8cd5ePoqNKIfAnKWe7grLSFk5ogYAeKK9VVZGzNzawUoC
+e5FWMuA8RrQ9ARZJvetPJg0ggIBumhov7+k/ash05e3RvnrTLqczYBV9jMjO+hP
SbJdLLaxLFnsKsq8dTRnWRameEw1v+CmIaV+FFzxBU+RLMyFGnhtpXfuE2QQ/dGL
Zn3S/A1otSVXoreHOkqxMqfoypg1P9Ao6oL0r8gvbVDO2xORj0UK6jFMFy3avSlV
FRmVhXXOUtznHYovD6L0xBmhKRRXwdaujNmiojrY5XRBzGrn6+dB4drzy5zO5WH+
5Okle/APLsKDCRL1bCovZVZQU76+hG5/KcSVR5Yg/sXgZJPISHDkAK8XV4LLcYoU
eogMwbRT5cpzt+GQGd7vmQlSzOt0k5/DKAwuvl1oLSYJhbMB2GWlXjF/TLAqcb4X
jxvGk/ozpCh20XI3pN0vU1NmZdaPu6ilh74KVavPNsIHG1Crl+74TVpbEI2zidp7
CBPA2msZmGh20qs8j9r7oGa9NWSbQHvXcy8rei4YVVlISdizY8P64JI/pWptUJqv
6Cq83RsJsSN9VZXJhbcAOAEaxDnEz5WnKTNlPt1cTTqXJC/PO6/VjJKOdE+Boin9
n0d7TaZuzEM94WzfqB5GSsfBX57xWl1hBitsXVRXa7HasG3/N+3QTkxg3IFyqtEB
7fdcxG51miRdV4eXEMjK0C49dtx2QcsN2iDkvwuhqW5Pg0vfEm+Fymz7STefD8AN
8nJhX+RIHBMUhIZ/fSI4hXmG6tj+97y4yj0H24e9s5EPjil5FrFIvhcUsn4FvHvm
LKeBqLKLfsD/15K/2aqzVnQGYQAkmDa0c82aShd5CtrlUtBnxPsfc4e22GCbRPjW
uE6aWXPF197J88I/lSoytLT+qZruL3efUeQuTkw3apHrCePqoRBip21+5t8c7/5o
QpaFgfikrWldcuId0PACWX6JEkhDdIw+pgxGqHFMmEM0aR9bpO677KVE0kBvwL70
tSv0JNgI5V4hv8hzK5qlrlf9qLZL4e9hX86OHXvRjjf52uDPjdMsLCkbsPNtRXZm
J29CPDuq+zvUgL3VQqPMswjTtL7YK3bVT4PZ6rqfoa2N8PPuYg+cWgTOoCiYy5i7
5GEBcm1gvRk73GVW1a2WgagIX/jjI/uJD4Cvl6A0yXkhejxO21TxqLsyV1L1UV6S
tX9aRp/3ZEIq9NrSwUL/DfQ7r4ocfULqperrZ65Y+v8gReiqJor3+1xBDESTM8tW
V7enAFgo2GxUeJUMk8ggpYSf36PZPD99ayx8K4mpFQFCM9GK+1MiWPkRx+AejHY/
Z55oCN4yT1VCiDDoHrrFkPdI2nf0CjEN1tcZX/kq2vMxWXXQIsNYwPSrnSUCzhd8
J65X1LqaEO1PqnavpGnbKZVZE+K/ESROwhxZ8nd5D71/NzE/dPqNoFyJQ15FW+o/
3sDjNQmTyH0tF6YJz1zInMFDfvdtk414vUvtWV7ZCpdx1KEYpnFB6Q+tJTVJABmc
ooQ7Y7VASR0xKnExZ+Wz9QS9J0aayQzqjuNhl5dZzHvBZ8z6cGqMQSh1G0N8IkdJ
DE6uXIgfw23EvSw/m0xQClWKvcRnpZ1EwPKHbCKGXSuHfP7iUmdtp78zb8+gj+QF
QWyPWeD78ldPbQFJ/905cxqE1OZnLVuMBrDKD0KUwhfy06ePB/FMrsm7TfxFFYaQ
lke0xdvefveb0MbgOIc2lf7x6DU+iInGPNv3eV+EIhXV/ow4gM0W27jfYoGvzvae
gYTD5rlPPiRuhuN6Tkqc+YVhuQl60Ybr4Fh70UcRpIOYU/778bA2B4Ekpqtj8EFl
icGJrba1NEBZsv3WFDy0r6G0e2KtdjM4F7+by1j2pTU744K2MR4N0lavPbWr2TsJ
6hoy0EqhrZB+mbe6F6wE4kZrK98SEUtx1YaTM37+UL3VSsdcvLNR20U2gF309C58
h38TbdAPhUGAZWlbfIhqSr5ATCbesnfl8Wzi73xdzs+/SZ2yzYg0MeJu4FJzXyR2
Q+f30b8HCG74RVfq4AXPgUEUcILEwknnzRRPcm122Dqr4eyh9hvrIZNa9TU3ZH4b
a72M3yeG+WXjlqeyOkWjm85YRPbRJOad1+JFdYWi24KWW4lS2KyB0VOE7liwgPtu
VWKi9Amdpz/zjk8oqIourNrkgJYwILJHLP8dhFue+0sfBENjjZoxm/rVEx/72jG3
YDh1uMZH1tQVG2GFF5ulJVpJH6P7swj6A/nYbG6miNsdB6g2FS0R20S2tIC5d1eR
/M5qtJpVGnnUKRx6Pa4pNfhTMht+6TmTdX5xSmTcxxlC2UW48g8wVC5hxxXBU9dI
OUW9kbjLwD3C9iZFcIBXa06CTUGIhq2O7YCSL6dFDR7awQRKZSRj50oe6HxeTQVW
fly9ELQj69CtLotJJSZsTtN2dh1AEkwKZ13vpt98UdLX1is8DWed68EH0qeAjQ8E
xtsDATrUfrYmnheXGcksuvUMSeqniZ2OCBmm6UM92OgjdwywQTmIgOYywssjXYTG
MxjfEbjKABfdj1utigJec3rgNGQsZr7ui7Jfj/U+auedcdizet9oG8wTtB+/sXHq
9YZ7rQoEf00b2/O+KB4WJXnSspDBz2qCtLcOnUMlMP0Pg9iToiEaJVs9sZfl6Uw9
8MieynspKT7+oxpMJOVpkFRjXmKUmnOx3EKRhEgeQJNfvK5sZl47QK1yREv/53DS
rRP8XT7YFSdsktKRdcXXQKtSMCdSJ7vn5ul18im2Xs6aVGrIOX/dk5im//0LLRak
Muyfd5ddBhX7H2/9Lh1oBw759wann4iHIoCuwJRqk5o3w4VhM/8ytjDs9UpfCfsu
3DMSHJkVhaoOIkPdULoJ9D1mzZFq2NtI0thI+Fv2hnj9KXIpQF4FQHGjKcFdBsEN
khQvsXARe/woun0e7eaKDlClVuK4sACGRGxktKGHqETmXzBGn7ZVAjUFJNUfSCfL
VCvnvF5HiTZobPXzovo2ttvt063mgIvc/VQ+/SeVDarxQ+Nb1ngDbTNlBkwyLOu7
mOwQ8ablIYRHE8ggi0sfDjNN9EQYbkjuiS6Z8ruwsDGo6yG3lFrFLkjiKgu8oB3x
kth6iRsS2mGs17+dYAyusQO4MT7IfBr7qzYmmCVLBpwVopyYFlMbZkV4bwQfJovD
EJjJdbNMFiWhEwSfQpkBjLLT0t9u9NATmaV2MRQ/Br/HeeWlVgvDYBl5yIWFpL0C
92VV6RPSaryUG8KQOC1u7O9tMMrGdLGTHFRmBAKwEisXITcQZN/PYfgI18TXN4VU
RUQI1jbTt2qL7tW8yCgDV6TKdQ1I+OspJYbNAlPtZQMut5cGC/Sb1HH7S08gX9Lp
ItduWpRpIhDDAw0iWa0jCVWJNajrk0sMCm9UehoiOzVxq1nC3nh67AytRaSWNB5f
NN3dqNz386BJV8UXje0fqoyb274HoR9KM9vhc6LjlbBxM3UzQTvjbS4XLNY4ZsKb
w7Jvtow+t9zXJWR0hkruuNN2ymU/cqXZ7sMNwRfLmmyUvt+ePD0/yfkKO/I7XiLO
7jXw2cu7ScG9W2mHITKQUStILpCJv+ZnmHrxAyQUsAYWJGv4wDJL0sR1MXQLO5PQ
0jStejt8xVwiP11EfgGn/zdb3sTIit9Y+hvRG7rF8fH7jW6KbbaqSUgizlWNRzdg
5MTFfK50wXkD0xnq5zuCIQejZZ5SoC+StFGZ2yil7kdtCCUaQLLZ/bvtbA2Xa5+K
uZPyVHbJ1vEZC5JrFJkY7ULXLy/RB47f6csCmYWc1KjwGvGWmKUm0OOlidqAHypB
QuQvL3TpCd1ADZV9ka5HmMfPvCNXz3a/y06Kf09CgYjx4rTOS5/NVjyGBBRKrV26
EwRF0rXJ4M8TR2EpwSavL1PkvEh+vM7bQGzSQdxR5P/ka3B9Ie0TkWClbRSx2+17
y+oYHNilQ2sxWGhu49iz0inm0jv+Q4vHAEHtm77Ia4qYDXYLg2q+sgdq3j5uH2cm
u3Z0bo1MZarizQgM7p9hjvZX1f2nB5cgdmV+yIOksczHliAmnvnElDNqAF+RDGtZ
uDoptq82kwHQdgUGl0JGzaadJ/AW0HfDXf1AZfjzS8yiTLjSzG+R7lHGFKC2H5Vg
xjMiCAF5c09Q8WG35SOhsuViyZpqywxEc+upniPqwrMjAfHlUr9GDpi225y5no18
/SFUmaQ+caTGxl5pY7x/MdEufA7Kbr6Bh/6zT/IaObd6j3liABjys0iZBPr5gb6+
kTG9q5HsykVhgCnuzh3cLSLdoswhtzRNPc3CZFp4/dQ6zqpikKbo1atieWYtXZEI
MHLCp57XnW8kkGMfGRjafAf5S0I/QPcv4eNM6cd7j4FN62azssfyHIsQlPNqbT+U
KBH8630TTF2cACItDd9b38TPNjSgaOjbQYXTNqyqe/uZXIc216EbQEw8H3fIvsCu
0MPeJtx5bXYqpyUBKwf0AiFM/p2TeH8HJQMnwmi7+sXa+Luj2+R9e1vco69uJiFE
6dAszCYs+SN2f1YkAVoORsGlcg3IdRrGKbi+Voc1K7ldcbiiL8aZig01ss1QYYJD
JpPNKVvwHxq1T7u/1noefeJxVNqLMIpRHuOsN8EiXEnwe2o2LgI4Eg+Q7NSSGkNF
9N06ieZnqNkDT3xPFXgJ3zwFbdpC8vL0LnznhrR625Qi1Zmnk2iWUvk2NEIVbw82
fkro7+BGs5ILLkos6GGHQkDc4iFCalx9igZPe6DH1AvAofI8zPSjVT2vvMMVcfoM
waeDlsRIMyMKMqfuakpwh31NtuOSgjX28fqgqphpqNbL9B8dazXZdnV/ezktQyTr
OS9z1ZYVikQze0oj76zg6nMOUkJMkoRDUYHhdjyEKUwKxzVrBEHua5rZKAN5YyB7
1AYoPsWoaP6geUiGO7mfr4Jxm9433gV2WaKXrD0zLAi4RxoYn/rqgmDV2bZtk9RW
/anXShaI/2T5uoOcZ5MdjVMOLXjsLmZlkoK9j986CYPFAlwQisJw9Yp4F4W4s+ka
ekW38INP84PIovTf4LNJklMRGRqQEq8dUlOaFe+m4HtnGrlwlKMM5CUXQks18gg/
KKGZdyHmSavJiWNSOUq6+y6zqLW4VPoTHhy2GTMZD1U8NlDxTUMJSqjGBQ4FQd43
s3J5V78grFu+/qU7LDqZRrCRyPjymYtQwDe/fapGUPH9/+zj50aYXdWgfWcTxfIK
JmE5DhFd1bmgwD4LM2CZ3UjqXKdPBFQGet3QHjWnzLO6lyj+kTWjdovbw0LhLSN8
zsVcIwo1LSgB6AdhEwrfHxJGsESCkrNw1UcbQaU45eJRpE79qS8HKpKJ0PxtEpHr
xyqqeWcgHuStAeYNWu899LzAibyiw8HxUAewVgKivFMWYZaM8xw0awczgY04I/UU
b4plgL+TU984ltprVn34t54y16IEg0UJC2qIVOwV4B06s2PobpYcdFAS+gMcU4Tg
U1kY0kVmQnqzU/VZiEy8gUhyB5yl6DhNWOrDkEaQibt24H72jmymSDBlMhrv6wQJ
PAyXW9X8nlvVku3pZmzLI1zZF6xQFFNvttqpiDw13bTGSBYK35MeNUUTodFV4S/+
Dvo5bGlq7cbNPinTN90FBh49vp/Fl1n5D2/gzwvIHfJhRIY4Hk9QMu6ztwhZX71h
TGx3fAu5vztPqb+V8IfjX4bvlZHgtmfIsb+QqO89G1BogufcbYJenQBzqZG+9frf
b8nUP5G2xdzQanwyj+4y3HaClz75gWWDgPJZG/IjNzwg5vg18olEV/HQfnF40Jde
hGeAymmbVr+6/XaHDdbWbZUI0Jg+0Vd0xMMjkgktHkfE5V7Kaw0EzsTshn3/iPtn
gQBqDTRj2fzv91qAqzVo0Y4T/88F2SU7nRF9kgbCEUpo/pUxGZPy6bezPBklCZfV
nmtLoOrq8dVshRoHurwjso6BAqNCQBeYOXvRI2wu4ZLg0SZHJ8DyGJh1d3VIAqwc
CN7mpkQNHCFpfZwZzeSsmDfgv72V1KKXvfQzzySbL0P2ymhgGjorQCTWgdoPR5gk
a2yVyUULSzQO/IoSci/jVP8j8uFhYMWSZ7HiUkcGLNE44xEtq79GxjAYPFJhsXrF
CubTP35IY4/xfCx5C7NEsBzGxtxmXPBq9Xss3iDixK30P51E84CBVM4aSyF54qFv
fCz1pcnStsuu9/iX4lIajPkbA/7PjbADeTu3B2BUvsJkPw+IdZztrfsbsyQoM/jr
cEKxrQQxb9R64HNmOWCP7/2jH6+rubrnptyyDoa8pbXHUNDpeuEgHufUQNIIYVU0
+sLPdMCm5ApTFjrtvU3J8L2j5AdE7Iqvkt0/xvPu6eZ1FoCHyaQbwOVttSJQR0fh
4n9B9GrfR5S0CdY4oDgmeOt72xtw2dfLduPn98HF8AHVDWZJuFgZbc9axUscsCmE
1fX2SbfPwhLHpoJdOsGE6jO6GeST10AgHJrD48CfBGTendZHmlux5JGE+bxkOXpM
Km7v4gcauB0D+ENmbcCMFl0oBBxkT/mSYNWYyJyZ1w6E/O3A3H0IuHFqcvDxFyvZ
p2JFR8apxpyOF01ky1/NbIfxc4Yy/fMkD5qP+B3qOozwLuRCyCoHlhgK/3OIBXi8
b5IzlJxkGNIEyQOPscRYCWKQlTX32BdrX4gw3zPV7LtE/ZaUwHFx850+gIU6Rrpd
EXwRDYWcRha7qr9LannfjMdcIVump81mZqLOtWKZhkvVPNeLOE4+b6WAAd31O6Av
3QYVd55dDQVUXq/Y8ciX0YeoWu1QfZcCUHehKWcM8yaf/9uuluhuhPxoadQTNhU5
Hrp74wBTjJLkakjrd15qMoUHCqW4nj/whZYkHFoaG7LDB/a+4hp12yHGkAZFQTXz
XQwB5yIbqULorKfAhk1P3czabuunOt5IGMaTTxn3lV//0HblzG57eYl3rAlEkyjM
jW7fBTBse0QC13M8/EmsOVPC4VwCkCjhzBah4Asf1fWCHo+bBkNnxBNVAUarPbcr
Z1/ihiZu2/VGMwZue0bWjfmq5jFZOt63EjupmJeiY75wQMjVTscx4ruH4VspF5wD
HIynGXaEk6d2lvWIaWhA/IMCYqYIr/dKlnSYeN4IcGYJjOep42tCr97XGir+lUYV
oBM7dqucihXHpacLprMZTlAR76f8Ud8Gn8cIUgnG7yixyCdm4ANSQeLp4WdQjeT4
b+BmjbKFBhQDklF7OjSvxwGUmeJBALRv72kwWCeeRkZxhZ4J3hR/PsOwNPXOnDQ+
HyhP91SG2x6+pbS5qT8MD8xIbbUD5QI/Thy3PxcxkOHaR2TCp4hDpTSrsWcr/jL3
2xoS/4B/a8ct4KEb7iD9505x+LMxK2k5N/EU3hqjnIxxvMtyAYHnQfCB+rQ1hJtV
7Kfu6cHPkGKZUjdW5jMU5WC+Q6CQ+uslUk9ne+MXoThWpXJ63mB7cQMUz81FMAp+
eN5I76B7BkNQhNdInt3WGudr6CQA1j1kIBUrp33LtU7fwclYHE2thju24H6QS+A3
zVf3OuGs3H8XEKwT0viEluf/2RC3NoIMI9reSWQ/mxEMY4vBAm5nWdmaNfMM3p/5
Y3TOcQ2sABWPntzNmUpxvX3VFySFLKMxP1IVyrdBnPyaC2OW6mJHpSYcX0Ey1q2h
N7AmqLsuKp7bw9c0yjkl3slcQz2X/ZsHPIrlkj1m1SzQAzt8fGc1Z1Lx8kPchzxh
CilP2GqO2fe4OzHxy7GkeBBzkOdPHH3o3zsXIR0X+U7JJQuzebATmGZKunmJET9a
OElqS7EXgFRQfesql8PNMbjoaHuUiX9jGD+BIo5AvyPsUwKc6D5WXQRjmM2RrCj8
Gz4DT3sLVNKmsQSLhxgKlKDUlugNragUrrq+bL/oT/bj4I3G+3NLLXqq8p8n3Dtk
hNOJf64uvvgbV3UthkSr/vNe5akEe4fO1N5Xdh0VGOq32MIsC40S+CdqyjC5jNXc
OKsHgX44jJjpL1i5vUScJv1XnCP/wOIJ2S0oitbWKrOSb4kBvDm94rxD++bSrKGB
ce9AgweclWmRxCLgMt1dUD1X7Qd6VUdJQfh9YrRNlc54LbC8KzQajmR/vyjKBMD6
ApyEghUB5/4ZUlV7lPBKdokU1v0Lv5xdAt+TtsAGGi23i2xjZATEfw8Yix6W0m1U
tFmzQ78G8r6ZxPRL8nWnPnl1yzeQOpSt+0EE8te3z5jvwobVmTOJvek88G0Hyj/k
bqf99vuiItkgxW/p/o2SC8jvpwKI4GRgu5QQMOabKbiu4jbN4VzjBkSrL1U6WUNp
FS9pGktz3uzjkGR2P9y3LBYFZ0hrEeQIGH2BkQriXQpxW9kgRPBVyrMXCfzsz+0W
X79bHsvz8PswYI77cd/vfDZWHo3bqba0p1BHTUckJkYD0Re0zYhKgxNq2XnHh3Wb
mzGZmQlUX+vjqA3iZFQ1lo1ofqxBmq9WlLMRlSfpJ5xtcIhxbas1egmoKgO2mpTv
TqQTA0jOvDd64baAXj4TJltB1GXp2YxT0US6NKVdV6iaqUAHoLsmBbC2RY2PwQiM
gVRxs6el2ITrg29RE+mW1XLnUtqiur1q7JxXX49qdYTrexXvQnhKhfPLP6EUI9ow
O3vmWwvIDYyOWLgRssDM+0kZMVnRN9eO+3ftLiJHiwabCXdpsmhpxw98XPlzaGBW
2XFzJ+tCcnRsWZ0/F46vjmE/ZieyXj5BtUJHkg+DUpef4mR5HwgSpRAMMigq6npp
wDyqppnyw1v5YfUlxebaIKVh4aTThy3U84OQ4q0qvv9lrTfB9DJIH9souDGpZB7M
hDWGVns13LzesdIrIXNmD7cMn//56wjFsVhcPimJd0pLhDARTct7oEIYsNq6Hw/V
X0XYfQXJ7mEXwNzDCKKTIDcpowFhUEPKo7Oik1tt7hSLuUcB4WLIO9MZK8AYj+lI
ds6KtEeQONb+gwEM2c2rl+amqojZNDuy7SCxMWr6g/Dcd9qU0noRM+cljCD9M0Ky
QRcqAlcjCbqlNj+cdQR9JRhy6T0ZLieEumiF4DubFVdwWysvMBHNz0ZD2dhI2k6k
oYSk20cZwaw/RgfeQCD+ONYoCPrEUvU9PEEwSwRVN8sOfr3F0hWKbGVu8XJa58m4
34X8pFwSs4aTliG8TCq22rmeJWc+MgFXoowbLjzrHu0yy5HlID3wzLa63qQCY8Sl
SsfFQEgVZScQfT/gmXwFIz01LoTBvBOihVxnYVhFL6NuF6WZJH0dRpH9QKUKGfPm
VRv0EQRaPflEvmEk2mScr7+8SHMkWuGkm6Iy87jyr6ZSimUG4PXGISI8FXTaqW38
21TBOJHHFoT9i6NzPbj3fMgw1CvYEE1v1ur3L67OFMxyVECWxaBztGjD8Nvfu0TC
sQjXRL2FMOdAPg1GsvLpNs4SdHTW1XbihNmyexs22S0JSV/We+ooWs/8DtHVNI7M
97MvrhZGfqinqEmJhd4SpRChLE5Wpob27hVYIXeQvuPjf2WepzA+JOQWlJoTgtSc
ULbVVce3qT3NzP0T0Xn06ev0G0WNw0Clhr5GlobteBgrKdyH1qWIOmww9rx3SoCg
haPpRwYTHxsgD/SYbzDaJGhKHmFFji0W+7FpTagw/UhIBDuR9fQPhkSpv++fyFTC
GSFhmD5Lf8xzdrfRafrxAkVe4+baKEq8RlOBHwIWiUqo+uOoMfPsgRwsgg69jcc9
O5HLImO1ogU0hxD/aCyg2+JpH+vpscqMZZeCjRz2ihhB9mlMtk0Web4hc6K3vYGa
lqn2qsFs0OijfMSeZ1EigBBmGcbno1R9GAp4pURdBm2AlO34DwU2rElBKA/Gz2Kv
/JyfWsY3oRFYxwf5p3bBty8G/O8ZRrQ4eq9LW5T3juQA7yzP698Io9gBXnFx8WEK
PJ2VEneERRjpJGuv2AXeMHlqxdOBcDSR79eO8Zpm4qejM/CEJlwCGflvdCEH3isT
yWJLWzG0qKl5NrThTJAcBu7GoErNQIGcfhsPdje7mxSFFtPKf92ClWa26nOMF5mw
zYIaIQGayYTsMJwUX3SDbmzfCmb+WTuhCdWfws5I2dBHKWnTX/5GrpugH/vx2JAA
Zniq1X7mhdh7lMxRcNtnj8f4zCQ9j0yRkY4wvfi4FToxfJst0WVGR38ojHr3SpUB
fdoWWdzg2IIi3ZsRe0tbnLcXqWMIbY9utO2QU9JrhKmGJDUCUV7luUaIVpUmRYn7
PvnL2mKbC7QloRfsKNjEKy2/J16Y4DQkpQOiIADVm32w+8L8A9hTaqcxhw8g6Hjs
0aH/RqnUBagf/G64zIpHIYG5X/IUcb97kuBplqyNeWWe+0jX6x+P9qj68+Z0YP+j
u8h6h4ESjjIcQFvHCrc8Q7zbnRkjK4FbmildfcoArP7pKy7MWnKI7QkFqm2LcZ6C
ds0S4uHKntlTRcA41lvjCuJwmkIdZfmDSjLocJh/XxnSBeZIQALni1+LuggfnaLN
+80SjUpJGXoxTO+kZHVMe89+CEgkS18IjMi87qsaanCOt+dEuqsJvKMQfBJS1Iea
2tDUKjPgRfpD3siv08ShA2zBzd/35HccGhxwGVWqTZh8DQ0Qd6a1XVJgq6MHxVlC
2aX+wQmcbFQocqgVQuBbNx21c2clskhNZqIVFdyYBbpDljaKbEXUv2EtpsMVK2RW
+djVQCmuXLC0ThaoFAOc7itZKtdJBRJA+T7Rd2btNZLlCnz6A+PSuCuxBbBUFIzE
HkmrDFKehcQLSKMmi/OmJazZfd/vhIvLiutedu6LdVRWO2VbyAnM8CGVsZ0PC0bZ
1jhbNBQoHrFQLRlJdDKWwLkTVO/cBOzETXAF8Mv4fvLCKHfuQRPpWOjnS7ssTJ36
cIW2U/Aiwc9iOibwVooZTnHvKOq/QgY4tVvJs2/oODpdg9RGxvKAYDACq1a9VErh
h22WEKgGi3w2M73yc8lFEufeXAnI2r+orpRXMonR0Pejio8nDWP6QkMaGFLLPVfG
Oxfzzf8LucVVAcz3J38CbcjNTD3IvoBzH8hemjBQDxa7ZRCOfU9Ie5SoYjTrqq/u
HE4evkEesm7A/7f5qonlj+nRvLT3xxZmlhY6KTQKfOfloC1EL2VPALlq+Zzgc87+
5pd8C9XfRbNGNeH9YexcAkYeYEv22FbQ3FKFDPPGqeqUhjWQENZMIcS1IeI1vawJ
8hHbVjKM69qIdbixQ3mrJsutpWCHA+8E7RUbHflldi37itSlNuC4ZgBPRNNF38WA
8Ell60Y+3GSIKRJ2T1+w6Z9Faqgr3zCtc8jYJGBykYHkmRIk75KauSwPxkYPGby1
rPQgxd7C5KfxV8WSAwMEQAhjfFIAVgB//o9jHOy8xnhNg7UkbJ/JUQLFW15W8AgB
3lrIlhYz0SOcNP+jlhbXAANusGvNwGZ3WytzyvZteV9jvBzwcwWy4E8JXdxR2mH3
wAiKVGCAoOyDOEYkb0zWaKr+/DrTHJSVNHoEUHxDMOtH0RpyAKCoCxH/QnL+X5RP
hn1aFcjz4qu5/hV3vfCOfkeIZk3FRTTl8snq3K5mP+ALePCtzIBE/JPuI7s4qGiy
du+UD6usgDcX5t62orLtMfYaV3FUYDVCwgZVcHxFkXhLLZhRjVjO6G/fLB5Fyo63
l3ivqZsByOq7gHwyY7MJ+AQN3GZoPIFgcTXPcL/3I2H9gz5m8gx4S2j9E7OBQbR2
w6sU0HxQ7rEa57n0Q+/g4kceGS/AuL0R0QPD9xch3JfMYefFhi99ffBkSUdiRITt
68+xHQz1tCPTCpf0A5vtD8nmuGRk+c7Ot1aQJV7ChyDpIhvmwdNQxlhoneLziyNF
VKn6DGKKmIL0FJuik4fC1fj+tcllN0rYS0a0PCwiCkPcOVR3mZDdL8iqSi7+ykGS
9Q4u9MNmwAONcVctOz4G35rcuF2BQLnSSLHKf6WuKnYYxmkHNUrQBycyN5L+Zwv8
9YqULyLkdhae5CfpeggJa451+BXopHtb2H5oYP0tl5hcOsKX2497movljECnGfC2
tGIg4pFDrjyEY4KA8n21CWoMFUIGMVVh21hZ//LHheKan/0WC+TY8p6KJZlvBR7a
zkGo0dWhTF0aMRhCCFy7ubCzZ03McvcOxTNMW86ObUt+3rZ+VWuJEytuIHfg2efQ
XqwbmQm9C8bGjPyn4GraZ9ESMbzUrJw6AYMLakYuno5g4WD6DdqNv+p+lxP8XnoE
gngCuZoSqAtS8ep6TrxDFXfszVcx5gBvKZQRmc9Ieema1kZQt9y8cu/yR/N6tv0n
ND0FIAw13q7VuGPbbNM1qYgVLGvmqMrNTinQO0EURSKbjQsn9zGxwtJutE66pMo+
irZZmLXepYHtTKsu36PyFvIBa3VaLA5dX4Vgk11lK4rw8d1NhGpMHccDDkLrJvCv
/lbBnVKHJM974LDuoe/eKSg4l+g7rJaHKrVmxH2Sh7kZUSSUTIu5ZMIrQfWYbZSG
jtpIDVEHncqkHhhOzNozKgcSETif6g9QURBe4zrXcAXVTNJy4UU2UyIbJyP1BTK/
SyVMWWZdANm4s71Pm5YihZZ9F0cG153vcaWwb1zeF9056kAKJ58PuJcBlvmUUhiO
vbV/JOSnlx9AlXpShVX6PA5X02TOpbQ7uzXqTu66U6Gmq2JVfSuLaExu3yasT3pq
fpq69j/IydsgU9HK2O7zicwsAGLufttei0Mln3BjRMQY36iHYyuGfdBv2TyVEvam
GWlDB4naWLwr+nBv+rL/w+NoOFAdbgTuZT6Lw2os5FoLScgbgA6Rk8hmWqG0FtHW
EMp3HDaW4Mr12AxyOKHWjnQQgqLx2Y9iDyn3KzaTEtPQ+HP/uSRaDJNAtQWWtBR3
WrxXVNkgkUJ8SHgBZNn9JTgNsgBltjDQFxAAgp4e6zp/0rwZ5xKANBwjf8v12CtR
4HjKQzm0PUzy+smAvOai9tiSwaiD06DXgmKBf2IDlnDXTpZW1nkLX7JxJgJaE35M
OEAOdE+lBEZMUunnd0Bgp2eUpNfzpRfjUsE0ltAZjx0ZqBxz15ZhszbCj95c9c4D
Jx9GEb1eWT5r8rYAlfMQnQQzdkJuawaBqWkeRpNMaheT1maM5Y97P2d0JNbhuTfP
LeW4sP7OOmNO6DCxdHpLug5QAS0Y8yvN9Fpp464+jH6d0EYWTMX/AT1f49J9xRhF
SPBikGtgeRwi22yNeGVUGcOq8mwi0lufxwjshoYry655d7hSJTXEeSjYOhboue3T
fRxwNgalrF0ZRifUXFV6Dvo4WWmb0Kj56jVoUid00ynIfKjm1TXwzwuu9ogzv5B6
oAHop2NisTn7RtmnDHazDoxQtxauQOou34HkTF/0p1P0YSDyDHrxI4uIF81+PEFM
+wpFPOmgoT4Y1dIabrO2B1vgkKuqIpbg3i9fp/3eUHBtUVU/saPBWkDl3HPPjNMR
5wdjICZfLKJ6she1zyJIJmt37Dir+REMGLER9/MW2sHCXXIutdc2pLyKymci9wsU
l7PpuZxDJWpGMTqi+ecpDJmULnHOIuM+k7ootUmR0A1bjIr+bw59nVLcLlHtekkC
XNz0sXQAO8G+TJvOrkyyChJDL+AdQmJ4E2e6bXjG8f3YHpDaYknrS+0vbor/l1Uz
jnb/YHbHZbuhNpJGRCihS6ZToW9+MiLqkSXGMg/voB/NYkxTPuZ+EtgB1xRlM4Hd
5nZhzcfy0tUpE9lh0q5sYcIhnzx8N5vfLh0EOrG7Mb6XhyQvn6qjbrWNRm1drY9T
5IZVfMjn9Y8sTdm810XwqItdfsexhpHH9JdvLuriZiSZPuP1ZU/HcDjT/aBFzXO2
ANDoGa5JFPi25Cxy2T3NLMnWR2LVkybDe+sEKPNL89AOQ3kv+JzcaEEHIZIsmCEr
tp2vykPXMWHE2jdYhHmp57Oyfjc3U89yFA6x4J2SKSfqVIal17+1I3K9c/CBABDh
ayHBXmY/3x+Vq3yzqww31oxW8qT7u798e2EQX4kI77DTLo1IOyDOu5izRRw0D0Nl
1hhQbeBOiAqthSLv0mHc9MymqJ3j7DLz5yNcyMx/n+3HrRJjnDNJrrwt2dw8pPzW
nUCXiMRUvtwWhXCENWJE/ByPDVBT/fTF0b4BGLEMmsdWTbEm9NThEgwyQTnH/Bg4
r7Z1gUscuiRtUnk/jU061Y4MuE7HS0i/8Sh2icaNS4T7kN3d3gC82TXwXfYp5JNf
sJVOdlceAv67r61dilaNVd4bakqfUSB8DQo3iT0Vl/oDqg3AeHNVXAnQRAEZWXa/
3GZqAG6eWzbeBSpmAvku2z7Iv0uw/KOjEYv+99JpBQbQz+QhrMYOrY8P717pTTjs
K6UisNv4njQi5OJHqt2Aj+6O7Agsyku/hrntIhMJBwZD//3pIB2ywzVXIEoepQKA
uzSB+Kg280ohxEfnhm5olqisve4LH0YyyfeilC77RKOqOqEGfk1R7c2b32/CIP/P
zpfLgsWoVbQu+GwyVCJQApCYa7B3Wdc5dfWEl1/jzEPxdCZC4ynBNmoaY/pXD39l
uvNYubmQJVY3qtZT8wJ7MxzMOssPh85BXjzOLRdW2tYI+Mh7H4b9xeNGSXEQZpNQ
mLHtMC0VW/W9ZBrV5uTazdGAiN6gAEtMDQLQDNKOYksNSyUryJRmzSMbgZkQmzxt
7sOmZBIgLIsEWdgM+5AvYtVNoWlZ0XkoB6aRVoh09qwWdF0+if8xdv/p9gmcd5Mz
YhIUMCt1lvZi2mgySBT0RTmlTfk6hgBgSmAZWHYm6wUdjzJkT/XSY8LYI3RMRudH
Pql1y0vb8hXYcN+IF1XEcSxYPITvsPnKFR5WcAazEeqVlWSrBFLJYqTngynacgFz
Rvq5w/2Pp+UjLUTS3gCeWd2LHk7E0zhp1JJReBX+2AMaw+7zKag/MPzCyot+fa4z
gjjyMp6K4obzH2JweH12dT6G1MCFFGWosgUMkjhZcsG6qLbMnSWoTDCcbgyHXpRr
eFZ1lvpWk/FQgDoyJIVTWcwRXWpJ3LId0R0iNfVgcJNJsUuCB1LCeeqqveEAdteo
oUebVN7Kk/IH+1zA9fGz2+B06YusC60vhUkkL9Jiq67uEGYSxcc+xhPQgZwg6RkR
PvHdP/HpKWn5DO0oNSBTPAc7cLKqVIACyBo9H9nCwol/+xbHHQ6cZZhReBN71HQx
9wFPr69mJLQYjfo6+WVe2YswUn9B4NIUm+TFTT8GimStDA4sjXlbv7g7J+ffVLSP
ECIWf40bgzD0sDuROo6PJhqzghFEjSRbtznOchN7xOLedJsk4k808KTsZJE5CBQE
vTWFiHNeqgjMe8jdl+3sbMhPZFQLhdvemDX81wq9xHtrxXUpuzCKifI6uawWaDxq
sl3hNiCTxlNT9tOpJpjoycK60sVy6FbN/MZq2at9VuJagiDbAxTQEujUgpduxX4t
YeErxQlD+URvV3+c1EY8Rma6OGROkNr16uyNBZPp0tk4/M1thRbqaCT9Rghmgl5N
JISmL4RcHTv1azdygMi3Fx5W85nW41SgOVCqb253E0Qr77wepm16x+gfrVsV6QLg
N8xtxP3SRbNnfIiWhPLRLfAQERrinPbuwKLofup+G1l6CxsN47tcCORTVkaBgzSX
DujvogkRMsgZTlrNg5v01DP+HmnqapYWQFhQwesRAAWLKiVwHVpR2liUsCYE2RBe
EpEV0TEXAI/kSZspnGeeuAhM3CWXh+BSCyN1e9ACaOKWHj71m7u0Bbh61cYTazY9
+hSKAegCoVOXwBrgdUmPU6i+zo9SgwcPg7RLXM6RDKwnzOG4xrn32Bfk1li7VBUz
8LKSImH7JMycHCXzhL6FQS7/oCZk5y6vrGO1pa/QbrTBdeJYXof9JkU70FQVROh8
/fGxvVTEzczUX7dS8AiPeFuJYdtR1+Ka0oDwYcbn/ov0W/Xsj2hRm+CHx7XEGBmg
FaKJqWEV76f+X++Q/W1h8MSM2KCblE9+K+Pb8JLTKfmgj/rnLW3t/Boh03CY3mr/
McLR2J7A75+OOUlmSEsul4UiLgO+VKZnrkOCG5qGdZruwaPH+Th2Am7yc2mxJ49c
akJsIN73LrXPYcNJq6pai8+WZBwt3eH4Z4Ekob0Egz7Qb1y1PupNEcyzjOqZJaUz
FsmEs0eBUC+nhRFeQDCLv9ppdFu1QoWyUY4CIJg6iMnuL5bvaxr/caWcTomV9Rbh
ndN69v3iMHAnxzXYNlT7tWaSgcDDu9XgFlbtpsdKBI8iHPgbHSqVrKrgcboLsFKt
p0qCtomUSIa1kc3kAXggrZmh4k99pGqtD7U1VYrjr38QhjgEi3UvJznKhwUBfAjB
ljbiu08RL3/ya9W1AJubC3CQqQOiLxyqii+x0QgCHSJ/ELyBrxy+YReZSUI1hlP6
e/gnNzwPfHLWI1XUsU6wF+AhrZSOIAcK4OicUi2Bx4pEwZNJbd/1BOENvkpOgyLf
FprSegkWf/j6l8pU7Rc/YocqxC+6/JgdBsKgJ7sjK8fwtNeHXLZoEzn8rawvgbCS
c4RBy9Ry5UX35v5bePaxZkty/9V9wGbzEeHaBbRmjsLzY51nrzSleSq/8VE1lq1l
109j+BOdCChSc1TEIhs36zLSKOHCtC6aj/CDHD+5UH0TvyjM889IPaSBuVbbnPHl
EOqWZTaMt4KYbz6ouEb2/hVNRlU7Hv3B4NC7d+uZINC/uAruw58nQzTYl62TKTYN
4yzv09OwqDF3EtYp6VaFP5MAFrTRwShPdWcMOYIHzRIiCeH9nyFGT2KQew7zQor8
4W0DJiLlbGw/UbEwWVD4wIQLN9Ee3GDMqjL6Ue6g3F0iZJXQWFv/cEnGDkkDdSze
k/1gYFOusB959llZ76U1t0E0uZ4sFLYOAFtN8DNokOQZvi50bqvM+cC3fUTrsac6
n4F5B6jXO8lInKTJopOU/pRGGcn3C1kKJsl1kMgZdXXXCF1T1Gfel15oFi/5dHtF
+yTdKbD323M49BzTaOE4krUijy1XsOHU522mKu+Bl+CAMuKDFuIR2jy8lCWWRpVL
rt17p0mQ85V+EOrSYKbhBMAxdf8uxfM0jR9ijoOZFY/4qYrMp92DIOXev9jYp4X3
/0cwIZP6vaHZ0EzaKJ19ojsBzVuM4cvU2bK+maIlKxTMEmzAnC5S02WnaGrEyAOO
BkmwiEsJGzGmW4+c8sVOKffeqUH0hZHhBn5wEly3/It8rjbiCapUdIsAnk0GvYFq
CfpgfhS9ZwPBtxUjmKMUhHeSHmEfesl6eiaa97/ORr0bNN8P0Do3TE5bzizZP9Ed
fyC0iIkpl56p0b3edfVik6t4dZp8bvFcESYLP3hkX8Ib/plYHAkqamLmSdV0fph0
q0AT20XeKF/Us1psH7O9N+MfIkA/9Y4M7xhsbQ9xFN8X38Y2Rfs4QBFGRBBlcdlm
g3K8kCpNYfnrq6LO0fjqgMvsdpYFxUtUuORn4PXm6E+4ivwtYlC+1aIB+UQKDkl0
Xc7usgxX4xDxPqU1clAtRvrljzIvi1AuDkPXa3aFGkZoRN0BubLyxWY11kRf+e3i
fLm0uY14eJh4k+z5/pXeY3bcLt4vjNhIb/0TUVv5pUtP0zAVpns1vddjgMlLv63X
ym19vA4GugNe3NgmdKjuo79FX5jtXqExqVrD4ordI7AZhI6OGfCwLcR4LZBGMepA
1g6/IHj4cuHUZ2LedISnqtt0OnPTFGk6s021Z6BCIEYIITESFNa9m7PwddFRP7+X
UVXw99nNURSK19B1wKa4dXK6M3TkrqPypac5v/40bo9PdAvE+Whzaxz4FKqn7tCK
rqLGBQaKhBGM1gZtKIV0A89qyaOmUe2avysG8UHwrVUJqtLzl4Pa7hq4h42WxpZy
/7qgMG6bGnZS4ZSdMe8eSJYFwOXoon0tvwcF/lME8DwlvipPjYdIP50ehGhARvjo
FolmI8MPAW6Kh8jRpvwsjXpQtfYuH3qy7Hb1a7w45sb3LqpagYV/MA9OSFxTA79I
BgNQuB+FjUTbfHWlzecT2TxP1NE/BA190MQ5GTq2tJEdYm2rW9fqZV0v5dz2fWSZ
MEiOWsvnoBaAar1cSJ4ubTX9DoCDh7mcH3/MMOdaeJU9wOGIrr0QPVWFUXqgG2O3
SI3tDf90Tf/xH/rXZrG2Ye0a+btujCRsi+h+ywx9w/jzxz+XhHlDo6+34S1tbKEM
1dcCv0cXqqte5Ahr9/nMw2TtH+ggE4OIjRpvolqEcBUr5rv0Md9eV6su3Ywrt0E4
1NwZJnIVDDvRyh8KwAr9F58tfut3EmshHcytt1YSecagtuXw/fRQCRHTrv9chnM8
dg9r2IBZkMhjQRpG59SftWMpo5FNTNaWXfKC0RsCJaSprkzjyUrSyw1oty8VugmS
bxaTcVm/wuw5F2UVPtOCdse5S+oDhM+EZhgL6efazRy7NOJYMstVwcJuYOS5bts3
dacw1YZvC30p+O0zuggvRyJJ5F2jm1skD5PJ+1ejOipfiB7XP1AWc6uEkQm7M0ib
8f1L8e85KtfwZup93f9zJedvTbcQFTr2ism7Rs60PTtfaqWZlC1aUsA9qGw3dw+n
0NWU//fCAQp5Jp1lwBI7PZUFj5KwcFSj3ZtcWMEVc3sVxuoCvB2mVmW3+AKJQoam
/rIzlEvF/r1AL5+BN86BlAv1D75ONI6mMEDuxAAqLeFeDZGDXvMdyuJ+UIJHbzrB
cuF8PeHc8iHfpmMJthLqV3+csyHvzRP5/Obozw5rJjls0oSgEnnOuPV0ZjeQ57aS
bZsr2lHgBWDJ3mQvS10JRZJeKNlfR2HxcJevh5hg9Mt4zFMshWOJfLkr1ODS3nQJ
M7F6Z0V2bZQyiijvCvtpFYuDwGtr+SMMBVhxFkE+dcFTTmmezxcPYHPBDv46B9L0
yIy49XINNAVPIz1yhjzZoX95Aurxnz80kUHOJUShmubtJL9tdwC1jaDqBnYPVoxp
E2UdK2wIjdvTMpuTTAKkLyXTMCFQh36Mf9NWskBdeoap6Vj6tNhJgv1iOLOPfHhc
VktvEUwsnaEeukORs2egLJ6rphP4GqHAxeoHMEzzEE0SEdtC0TYqRb8Hmo32O2o8
qrUEMSChANSpiA5bb/gjnkfG3q4vmsIagAscpBs7YeLpd6IRxTUvlyYCtGXSe6DC
2BnRjvnzXcghB5y7mBB/+EjHpuvVFIkuKGXr+rZfiN9KRWF83q0ioW+/UXyhsSjJ
tte3YDS7OLYmrScm4AmV5fvuQK6TGPz/CLixr93eX1adGDvmcbBbzYIstCZ3MNwp
FZQphquo9TY1gqK16l4yKYYSUUPZtITi+ANZfBUL+SIYGQNntB9Czyby8Rc/CYZm
0pX6Ud2I1iesZZ/86BWzIu5a4lduTlDqaDEAJPMQ8CT5XkExjkLxb/n0NQ7771WP
rH3UXjRUJQl9QyMD9MHClVrXDfgiZmMUlxpMy2OrB03Dn3TDRjtXX0g59LtsHBu7
zCv+qzYNpT0G89EuTlRVdyWHp0IJ5Iihd0PQ5VR7bSKqKAAj6UZvGh3sMnZj3jqO
MmnivaR02ZrkVZ7jbRE9W0MpsV2mqegWPER+BmRoZ1BcYbtIohF/E6dPtc0GZFi5
qUSLrnOxEP6tu6cl27zy9rb0dT5KNaPcLtN2PPgxPV+0JHQsiPDzKRuMG9lqejiU
rYnHaENdR1dQ2psobB5oV+s9WPBucBLQmOTzZ+WJNrFqapweqhuBI+eRoBvpRSnm
lGhP0Qcw/BSCy9LqvIdwMHQbiA8i3r3bJ9EPmPJEi2PPXOtlp+2hU4DjWNqraGL8
kS1XVReNHFatydeC1VB6p/3mjqDUrQWdgkdo17etfSPJokEPviwte5Jm6ze5cZTO
eJ6Sc05bIt4CfWz/C2QZBP6jLgRDNk6lPeGrR3azmC5ldzt1BZ7eIJv+UpBCHCTP
RKRk+QbZSMqeQ6Zyi26BOVxEpyNzE/UICSpMcQR/SpbKVWVDAqdr6VOTl3nIe9q+
gV86sEBNV0WQItGSFWj36XwJkNdtxFVJPhXCudfh/VsiMNLeDC7+DLwatk0ef853
ibyhlgoJzOc+q+CVRqlGQ7HUH2FeVCUY+bXzvDXZA8JHa4AE1aHHKyqwpk/z4xEb
112tbejdDIjfz9PGRPg1uE6UP+lgiI4RP6eXWdCWzGo39qer1+Y8PYh0eweKUaFH
/rQkHdtmKHFRWJJyoP15njt5QJbmEjUk0EVXLoxd0rLwAAuWIyxVoeNH+3yQ2YeK
WG+KZxeY+hsv4xvFIk5FqxPQ6ZlQI2HW/UUW+Ldm29rh9JkiTMMUFZKXhFrD4oHZ
O+38HWXV2Lz6E2LHFDXsx7b8i3Y6K8msFEPdmTQ1PMu9XUyDZbif/mD3Qd2AcWGu
MQAyEQ9r8Ca8ZoP7Ll8dgPQtNQKBYBfrBMj4Og8+wMr3t22bMidi901Mk21Z3hlV
HQho2yVkfQZKZCrnWDDjfPicV2Ewg2aiFsSfYSn/TzqEplpXLXNgzO7qHk6KxHMz
zMe1h5ZOTs+8HEgFbGZiKPQP8hMB0nx7PwUBdONxvac+Ktixuv9Q7tRDK08VTbHy
oboZSROoOkjVm5U6YWVdTsrvArb2II2tuMN5hvt+XAYMUll9pndFpNN1MHv/vPeL
4gXWOKNnA0EYd7miXruS1a5gfGWanck+M/o5bUCaERSMNSCLQ2IIkaug3FQ7nhRE
NJ56U5d2K+3j/+y1173qmm/p8PdLYa9FG85thMU+Md+YbiNEFwQnlpRSC78x1DVg
UyyGzS8VHjXi15BiNn+1ZvBjTpYhhr7TouL4moQmoqtuXcNim93N1DRNvEbj9NZN
C4Niyz8EnEuM/5QB42FRqxTGsAHkhw9Uvyu+ohE7vhQLlpG5LV9D44m4hp/LpUre
Kp9CpuIvnsKRldqixF/5EQ8QhdhXpgWF4+49ER1S6mQaiVmu7rbo+U59WiocUKuG
LZnmT4GkSIOE3vTHyP+DbK1YIDbWbtT1e87blMttJ+kieJH4kNZD2mK8fwZRcvV+
kVEkQYqqoTUDv39IWKdzLKLMEgwe0sQVGThxv5qKT25pGckHEZcEvl65FZI7HMan
v7834okgbQlCwCmVjkRfMst/Ose2S+Bdxdmu7dYD7LDRAJMuxSuKt+uVjF3iI8GP
88uX4im6J1Ot/zXuexa+h4j6bH9EXPqVX/3IJSPJJ/ZVmTIhRDktB3CwUsYs1SEu
IjGbkRCy7jW34/qo+DVy5PwAl/KnUOsO7FxzNQTzJGgajkcrWEarvdlIIH1q8TT2
WGwuKMZ74VHGhV/vp0v1BDw0m7/I4XjHis9YFc36PV7G2CX3W1uBFrhHEorvCQvq
O7ryC3Y1HLFqQRGIhPlCb65p4pqU8al7zsguhI9yc6pEM5kEXrcgolvfPQS5n+1M
c7OZdl82wUjhp+e0FWe18j7c+tszJ1TgvhPtn+EvR//ApdjrAJkT+cvqNgvuTrTb
OzoEKQUybivsGvpPS+WDJQgSCzXlk8IsndOIxByL3ijuNQ0uws8C9KH6MLqPyw9X
T0D+sXjTTx6sMubf1eA/9I+wyTgqobtSReu6iB4lEOfM7MQOxY7pOmFXeklt/FQg
8PVeSU2RbE0rkVDxBm5yYOFuyclZ19dJPYx2ZeQ4r/31yyXQz47uWX+mIdPWlFoA
KinX09JU5QcVbcJoa/WCU2j7FoNGn75AHLQUtzqiAWWOxJGwvIJ1UE2jN2WElQVa
LcZ85nqVHW0JL61bEMeNseBvKBAfrkVglkiS1aOhVg09PP4dySeqHXtt0jdRsJRD
axvEQA1DKguqq/g0QlUbbf4CGxXnHHdfqm8XbZqFSqtRl8hMs73mWDOpnrpFER+x
dTizNNSRqmrESeWAXzl46rtXXbg6hS1rt2pX9KN98NkAMMWKRgsiI5nN5p5ntWu+
7We3CtQj6KSWYyjVwnVx64Rq2aPKkGZ3i+ubxIAhWJn1YyIoUmgvYO0l3kq/PDju
fHqA6JUBmi/bdv+SO3JphkdAKuDO8810f1T3FTg2LGIUJzjiFpweswLHuWtSYAOW
cCHnt2il2c9o7nKGgPAwqb9g05YPvRL327RBiNEwZXsPBJGGghEbC0//Yu2HZ24o
B4+4pRJNjOFtn8hGUrcVswlLElG6O1/jX45P2smXYhzh37zpqSH8DA/IJxxuaMYV
hPNORaj5HGeE01smRT8UhmUeRECvTKPaJ66qlIH2MHELw5Q4ysMKD1cERioK7120
0q9eC5URxvHrj0mhSGmqg3e17UOpNxuS9xqrfBctI2l3ti25Ph69knBu+4lwckKN
7SOMBXYqEnjGbr2+PvOlRJduPHf+edzfGKtu5x6Mv8HZVk7BLlwkayk3WbYL8F8t
ODcOVaKDK4BcAP9z+ZLHuu6dTRGs9nSBU82Vwktf+W5QTn6WqODuYlpvtDQJPGF8
HcZckxoUGgelFf9wNNk2QIRoU+SdufysYoVjAnmzALF/jCMV2TE0mLh3bn8rq0jp
dcsnxRZeajCP7vcj8NvuOwSUAe/eA/p0JWLvAm5MCfMhY5+0+RTDxM1DJm2kQwjn
CdM5fGph0hq0sNOA73yKOWdhYF40bPH/IvTOy/oEUn4oEOukygXlav83Stu6u0qe
7+bY9L0boMYgjzp/WPludBtp6ByZQJjALRmL3SEmYXLH5gkhqxM0K6uXsF83HGZJ
MdinQXUweYAPqIIegLPcSt0zwetzi3XMwKbQKPjh2h6CzMzyieLGIhVLUQluFKWP
aSGzuQndFdZvsV+R6b5gYysH7gl5dJbiGI/eQ2b2sjQ4N3Q5iui2tuM1x2QcubUW
K0OKEBozVo0I4CqK6j2ONJXI64HkgEN9PsL6fo7v2C0b6W7ok1kZ8O5l0I83n/At
HUlwMvo82oH10y9fYycu4+0XsC56vw9p7xCvH5XpGa6YaM8IA3J41s+JB4hHr0bZ
s0FbSSOtS+ZagAAC8tEZaJLsAE2pqf7KV5RUdiokfm0xAdUiIeqo1WqQ6tvKFUPa
EavVmM0yXeqz078hsHwr6XZFBWeO6/Jh5NvJeXyoKNueSYTFpGZw+392QWwRWJwf
O8snWxX1rqXFrCwA++etrZO+N40scMByc1HGx21rnUBYR8r1HJCLmM32V9FLuBlh
0+b882f0xkS0LuiiWmLnpR6N4JbElYimXUs5ulKyx0j3VQmWnwtSQoP+4WuI+PyS
UjedASRscq647UP+ngeOuySwgAMEfjGGkXal+1jPhg7nNZS2aYZvqJ9N+UTRWShs
QJ42CFwYKEkkyvC0zld2O3GBjHj3qU2LzyvSDWCOncMfoaEKcXnxjk51uysVmNeH
SpqfA5QJ3V8CC1t/ib/5Dvpjls9f2mHptq6zS2esGyYLC0Q5nxEqOB7TK24XBBRx
+n5pTfSgNj+mOQtJgauYnBSow9NtLbC99Mse0kTiQvG2KkpR9W+E0KMi1sfgN005
77QT4mQaJcW7x4rKimhnjUwyly0YKUktRyA8P/t+RaDXMnjJnAig32G0yvfp2Unl
u3wj6D6WwofZjXQFu/h+JAam+JsduecHUXrva17r3Pf6G64WaxAvxjasNBqMboVo
XnvMeb8kuA/XAFN4Lof0CTL2S6yFlqDRXR1zEZtX2ViQFpv3iVA0o+dtEv7PtWmn
DblXSz5aN1YbBATehCFgA+o7SoHXFAMNLtlRMgYXhSDeUYOnuxLlHwmCsI4LMuLL
fJOeuf0u36i9rcqCVD7MykgC7CEQU4FS1nknmj1MD56nhTu72Hg6+k8n3D44wSmO
E1YhouU/Z4kZHogv41UeBBXdS8q9VEBuUbrIY7RB/xdieqJEv5cUi7qUSMj3z9RY
oJ5lnenrbaIO8idzoyvwUBX1AxNtex+V3aBAP9fLjlLzZ8Gr6VBpHE/8hknJGqG6
ObzraeQAKWzb8qoNpmPW16LT/RrqRb+8EZEERPDux0xUx96Ku1Up5fgYMoIdKm8V
qqxv6kjDhfQ5Vfr7ZG+R/GNoRJIFrXKpjydz8/ESwm7sFGa6Srz55HOzWbHqruAB
FDjrP1YAAlYkxMWuNnKpzj6eKZ0OgIUGxytUmPaNWRDGK3AuosUTKN/MPYgy46R+
ccjansxRZYhaeuHvYQQSyU4R6cquImpcpwtzTwtsu450L89VeqcM8OlcU6kGAetd
bqd0rrLvt2KKfQhKUiV2mJVdj1FlZFl4+/JYRvEuWBdQ0sbIizKQgzI0yJ70M6UC
C1PddcOttPlnJb0KJDiBi/V8cUUmQya7F/EJ9O2blFY+dPyv/hFgfCxz+YYFmQUK
0gs2nBkLFYjkIH1skSTgNoOoN1Jf/H5BkR3TgXw7dpsD2yECQZvvGY5scHyPSixV
N8G7ywztvBH+AEHV3yT8np6Zo4jcy4T+Qyucj1yt/bbKW1sD/dyfR0n5Zw9MfEaP
UrP3hVwqmRjPgqUV/iCuXRz8grRXQM8oEDDszYs0Nn0N8zeKwgS3s961s1NVW7vu
4qj1E3AEmFjzMtQlm+o/oLLUVW6H7zZUiLaZa5E+luQ6ZCQRoBxC9BqpXXNAAO34
mM3AMnp0i42U/ByoWHFh5XlIYJMebk3dgzidFu55Rj+q/jjdHRxY3+7Ava5W+DEN
TzP8wQYD6U2/axkY4ml78SC80TxFGGX2ZvJ7n0By48V5oaYj3ZvW4Ax5umLrba5E
Jc0+GMY1iFIgvrborFELfSvvoAi+/UVCL+sfOe47M0v6ThGenKQEyLtezI+3uiPe
24NYrVH+A9/7wBMxL6Wss7sk2lcKqdcir/zd5H+kGZYa1H+i1d4hKkIhadywkjFI
rWQfOdCH92tmN5vtxZht4jeGtizodiVbrmBW5KrnZ7nF9Zu25k+ZdCyUkdcnrMCK
fy83FSDIzD3gL/rtgjj2Q9e1fINrjSLqPTXBcRBx0jWEUCX/7CUIgG+eGgR0xN1P
zt907c4fgvnMK6uuGLna+Horn8jxaui8k0xoMZxYQ+QlPKm10ogjKd445VyEi+OJ
QPEtYy6vCNxDSbLcLs7kN36fMHV6uGnq28Ygpb16ans1bWwJFIQ3LAJPjb22NcNZ
jZ5byy5AnTMpmu7qnA1xRX4YhnU3HrCJcqkSe1aYVtJpApZNO3dCQPKgmTqwSLGO
WZUAL9I2XsjtyvcbKzxsKomKLtPhjzYJ1LLsw8fCv3v1H6FOJbtaGDbz4u0mo5yh
hRAF7JQJ2YbeNDFRYzUEE7WLlBKS3IWK3vgCy/i7CGntoPQmK2angn+D/D+rShUu
UM9oqkYN7v8C2wqAO3CyS27MafNYCxI8PcgTpyPxqBYL8nb5RzkfRVjkB3YnYdPx
sb9VjD9hCaeQ+VTwcHawokOQUCvMbLT93qDlzgDeneFKuIbG/i6FR8Aehwwq1W1l
qX8PH9ssLjKsOk6GifQpfVQiC594y5JPQQL9kzztSzUKkfGP7K+BPNk9zt8fmWZB
rdxcNoX+mzifSgiAvQkRemh9e1HHvVNCSaXFzShA589OZZZHtHUH6XFE00ds0Ioy
Nkdz3znL6x3p0qQbVsqPW5AVu6cLXdM0JBA3CvKMapaiKiedxYoCdFo+r4JmZKap
qcYdBSONs7nlZu/19po5MtOwbOzpcw0qZb0/DlaFDeVc+HfXnpsF6Lsj3MHb53hA
pPzNbezTEikbEoruZS9GSs6ElN6/EPm+X0pss8KeUXlk933uRCWG/jqNAQCXrTou
7bfpqQ0bnS37aMMZbrIBzjCSWICD3W38uzpCiWwWhqhW7SQkKwM+PIB7nKsdFRjf
4okSK0omYBYzkTvyu5RzuYJ6h8Pt+nXvvxoTqUr/swlPBe6UshzJJCls+nHG9fMW
/h/HnHppKc1k++b0A5PmaB+MVl6XXWpz1L87NWITrzhR0eijO2PIGPXOyc/L72yU
q/Ve2lNYQx4W0eJP74+/9hOorm1GxKSoqGhc0L8cespaeAj8XPnUxvM2xZLgWbHO
JN1blZw2KpSA0zMOW4aK5qhkha2KYv0HoGSZR7JOreacDs9RZRqIAD/XT4MiDvc7
MtEF3sH94qXW7a8QmBm1F/v+q0MrZv/F5UW9KXoHEsAr0QZrr5DotzwLv6l0IDdu
L22Mzt80y/0p/ipfD+Pk6Nf2r918RhFHq2b1eEhLbijmPn5PRVGpnC5CwmKJKc03
yijYLYB5Wv1Umi515PEqi291pjObRvGyZiygP33tyRumK0HbtUFpaxjtwHA+mDVp
VMn6gCgamIcchEaoLj18PJjLrCtG6EcTb6ulqGvpAe2H/ChAca/fXrTe8IEb/VJ2
gQw8qB8CTZHe8C3lBCEvLNvLHICtCPPnHK8kug6BoUT3owOgAonMqzvAAu+jBRzB
KE2Hfk6AyiIkHnMqIIQNFRBBqmHBHbiPmEAwwcYRsEnYJmD0UEzBcq9oka1ULYs+
2FJuZ7P0ienAkQRA1MT+JmNKLYW7CeCBuQyqNOLgSQD9u3V/26rZ3Z7PW/qdf3xi
X9H4apfg57A+02j8qOcp0YoGtugtSfGd2buTxCpq1E3Wzmqy7S7PQBxlTwu9JuJP
oN515NUlWci4V0ewpnZPjRrgkCcT7VH1+FS37Y8Bk2c7XByBnpjF4g/NGhIfWHTE
lXgfqPG85CqvrRCn2FYX3YQnTTV3gAkxH4qHPsk1Gjhhm9qOgzFqCtNKMjRL+9/E
9nFTR4IfhFr0ZKppxz9M3p5CFTOdoap2+F3BZA3W3IQEabm5nALfwyCCXob5LZ58
HpXwADPpFJjj8HxQCdArJCX8YgvGdRdIhgK0CD5mU2E644CJsoTfU8AWp9zpre8A
JgOvqi7gfYq+6uD6aHsKPrPQSDSt87ne6PVMxJomo5D+88SR8NKwMr7Lqsbisye0
s0TqmVS5YSx75rMs87SW4E/rQzMYYzko7gwHQ8MbxzwQn2j1aqIvm1qyxzIR09dm
WRYVac0QDaIQX7wlMzHwBM13H6vmsEggDm9BcMRJkAes0XjBp18uzksMI7SLg2Jy
egcRq3uvlENnokYoLjbeZZO7t3M7cgfRtZ6k2dbnVH3xrBTb0SNsCUpBjgi0zMSJ
sQjJjgb3A8RdLhsiTtp+oLCVmXMYrDzJIxKiqe6MxHhEMbLH2fVwGa1LBzrgCMlz
VCWbX7wUS7lYxfX1bEFpqnmXfyxMZ9xN+oSeUXMvt8YoZwRWl7roJqezgBdLnIKg
Lc0SvQfxP2Le/HLoORtbcTD2Ly6QE7bim9KigEzguK9nBC7SH48zQ7hnsJA5RDn9
hAstClEduVQIt33QTXJk5PhucrPlTYaaMezGEw8oWZGScdA7IJZ/dRxMhdS2Fhq8
9+Wt3jIbktNwd1SpmlexO5VLUPcqq3j8upVGZLorDF6MRJTukOKGKwOadNpdlLZF
K0OOdOLbyDjc4XSdKtb/bKvoHOvp+ainpySD0vNKC04TfN2XGqMeATs3Dri3/9Sy
cbLHW1DjP5IHYXjAkmA9jc87OqfzIiIeBUnBwsQlEHTpLX6RyyAaQHGhXkr3VHt1
sBEJBOSZhlq1iOT4wRr867shkDVOf97021h1/K5MQBGq2AwtHR/BlMB0A7xcPfcX
0k+QxlWw6xBTybPEo249JwtcV3AxKmNYbEqpNbJt2a/TdnbENmEs0k//xjQbg4G3
10JYVrfyGTFu66R4mL8HBK7FGxPopOFNcLRHGFQFPkyqnxXpc2QzaXe3MwVPx/OE
Tvoc0GR0pjt61JBSPh0/kpchWXHINwQQlIotmcU2ziI32Ul0ADWG+ZSQTL8QNgVv
70XF7UyX9lJvWdZxQbdpkV6EvRrsqyPwrVUQCzGUfXus/DccZ82IfDF8Jm6aCLc0
oi6s+I5nja5Lfj2DcdkZDcyh7lNaYzaHDDqiA0d3cw9KMhEFrYv3jYOr1N/Ds8N9
Y5ttfyFTI5secfBOfyS0YlHiBP1pfB8sApu+nV3pTIJNArCJRZ+Jb43d1ZeguLvY
oLxQpHYJj8NPo8t+LW4Vmfhm2OjeVWA3dtHmo7cCAW0hXqzna07doiYJdQZR+ax5
X3X0CPjpkHNjTJ96qUMC5FPdIFny33Ic0wOBnOhayuc0TbGYjPSVEDMRZGdmPyKU
V9nYbEps5QbITXVCKBJ4PU2byefKY9cCED5LeEhxAjBlFyP2bCgaiRz5U4/lJnc2
VxUipIFY7+IySwy34iCxvN6I9wIxlmUTJQMCDoW4gmabjTpkFmlUUzEZWGkOpTxN
bROf0FCFsBSZT82fRAJGuoL7Ik8SXXxu8agWctlJQBm9MuVJHA+iXjOImwGm8D5T
Nf1/azO3qfzRIfrcSN/+3+4Pxs48zpADLw5vQxd27arkbjPDYA0H9qDeMMDWaV9v
R2Dkza0yHZyx/5QyI+B+YksUu5niJbpnQZl5p3h9W0wzbilS6drk64EsxIw3RZbf
tPIOrM/Cp1q8MWARX+MS9zlldEKBJj6gxBxuehiWqaJad3XrMHaSUXrVSlWfaZS7
P3LxV4j8HnqM79n/GCyYHpoSScK0lR6M/eJUdCqMxEmc9QqxAYKHmI0sk+jGrwas
rBJZPKfEcc/YwSnHmEW2uVlLVtRt1lt7yAKXAKHjx0I66B1F0529Ur75Qagvf9qp
tHytjJVBPVt/1D0drCwwQ42U9p90WnLroJ8C8L44vv7HCcpWAdJSqgnSU51wwYjI
0jkisHm9J+jKMylM/0IqvCiZ6fsvkzZGI/19XwFe7RSPBV1E8pCzS9Q83TT0W0Jq
QVyF4bn0P/wPqzYAyCjoPBPFwJkfCBt85KVtURwPGVizaU3GMIy0+HpR2ZTB4jNn
yaZWEJhZHvGXMfIz/7qmqjOAGRhCnVdbGrfN7Ot3VfYwCVppSi72djlZ7gZSmWvg
Fu4gaW+04aAzWTSVPe1x1owbuTqhG6QNkcpOaMKOmvov43sED29Ao23cZ6+50YyL
ymnoi57ygNu0iwbufXW1iyEUKwdJj95q/huXygBikvPn3tiufVaqqNWLtUN5DOdG
3h31h4ScyyEoupQ9r7jXcSwEmcT61zBnK3232Iusu9NMK5s05X/I/rVPMtyb7Qgq
V9x0pRKoLu7Iu4hSVabXUI1UDJV/PFroMQ0cdD9O9vkWgFhkKAq44+Uqvl+gHcOR
ohYrchjLGnOCUQ3YkzouYzU+XWwLdIj21OEbmCnxNr6MnZ1wK7U+qzgNwyVlmWuZ
uVMQx0I3LykZj+z1Qa7eiWDlJwB9oWeB1cd2WOTGcNTri2Oew9m+67SBd1TFJa+0
3GPuzJYut3vW0eWdkS7iH+VsYiVscaQg/ai2mYbft/6m3T6CFsMBWQfytbv5TkwA
q8rnAv+tyRwhvdbl97t4R9N7Iu6cgd7A9Gwwye5QiffYbKPVgRSZvZje594kn6JL
tyDWEroOzPSShViwgJX52/N2rDfcfyiTghz+qreg16HOTJKrV8rAS3QUAwv4M22h
E2wHpPI8liHXGki6NGWCqG/OnD7AqPjAiQ1+M90RxG/l6RRrMUOL0QERXVsyMm02
Lkl3RRYmVrsSegIZGrYZNVRXqwIQtQ044g79Uk1aIopfz3eevIMpGrByXGlJpgwd
KWOapnVNU5G6NsU53tqbUvJl25Au2eYJlmfqWBhdfnONIRD2RKGUNHxSvhcoy23r
0n4Q0KXN2C6yEduWVz1gd/6OaZj5PfAaLMKpoOiMFrrbZpKj62D6iiglWMdAbZob
G/eucwn6nmn86Tb2K8hI65QaH1rhkymoKAydTQFTXPQ/bbNYeSFGsHxj1fadSyuw
aw7Z5220BA98iFe3Gq/ztY6FFyUxS49U5bAoDdKXKcsA8vmVWCovVH1FBECquEDi
cSyJwqDLIb1vyyPaHuMeAyBbZ7i8GJk3Kd7i0Kvu3dXldSwOVH1YAcWcQqG+qlBq
kVJMR+EO7iBNEwWOwld+H0S6EjTJGfOffFUfKyXrVFX+4sGQNoDSI6ut+ExL4jTP
goJciX1+WlXXrHdzU+Gm9R64kyBzzbCX9MFrYWg1J19G0Fuho1YJTjbSkDPWg16l
vKivBqtK9B4GWw1QXzncLF+rvYAxlyno0BDkL/LRYAUX7h7Py0Scjb61QK+aXo8N
5aEzm1y3hb/kk8Ib1zzbMZgVIYLGWJBl38wh6fHM/RytHU3M3dOc9CGzs6Ymp4Px
jdRH37nukdjCXGMYZ7qM1BfZoulTBJcQGXm+s9Nf5r7a0gZt9xV6Pv8fE5ZiChKv
WEv618hMQrnBaPFaWtOZmpETryDxA8/aMMHXuSJ+gcfaqGu0kkLvEOcEJf8EDBDy
yfaWJbt0nFauqPS7rtvxYmLvs3sV4uRm9jhO02cMLseSw6GJRh+ld/bGlddefawi
yhHRXiFa6r44LNXUnfZW3KEG/wKWX6sUGgnKcz2PXuRXfJygBlR8Sjkc4BO+2Nej
5u13JysUfHAMvcR3sw4qB/fLF7mcPlvwqcclZAMqjs8UeVTsN3BnO6NuTTZmh1ID
ka7/AtDE3OkWW4HFCOIqJzqCAUrBI9y4MfrO98b6dnZuku6B6Ao4nyt12Hp3sQqO
klB9HdctPWQ/w8xiyBVjeondpSJkQ7Yf1g3Rs+X5RBxoOhVdMz45lhwvH+UynnPf
c68ln7F6tII0Ll+lxVstIQCq7Xh2M/POfB5vnQi62pXZVzj5HZfz+F8FTXLreoam
MGH3fBrfL4Apysy8wVGNvODa6II9r2oFyhyj4VuEVx25ytrh7SCrOvV9qzk2SJrb
fP0q+hnMthbbpeBjlq/wNBXQ//nTRmb/3QnvDlsc4PT/coxKm4obOk5My6wQTInK
iP79eoSGWcruSO+89a4fQn1XeV8FvAtukzTmt4Pq8Rm3gGv//O35euGWUCz8NmGG
hkvKZaElqXApUi+0aqiWulMdQyc6IwOAuyROqPfrT0nV1yBe0JHoRyyd8zTSuPZU
klNWFTJnuh5XrR+yZhpDL1WfTxmDYlXCwpRDr2YUeorUo5ZXf/CkEPaV4kB03Eqn
a3pUQMRmbP/ZnQqWEN9eNSuJz6NXVhym05+zRZ5ZfZPReEw0VKjypMu4491dgyKp
1ZE95DUWf6ppj3OKcOfb+CPuh1ot5FEv5zPWbEQMpLUiXleH8vLmrkI4TRNpxcYD
vD83yKKpz/eJqiGyb+rzTkbiNl3dTpMa6IXrss2v5PcZC6dgdh5m7B3en81ob934
d+xjMECJ6EA2Yu41i9fD4FstuVRqEi4XxpUtyLeplY3hzyztgfQhFqLGRbJyxnw5
X3h32qjUb4aJsNupkbM/ux41DxOJRRNYOD2qRwbE2YU0q3I7s3N0u8pjyTgeIbpP
NZySz7YIJsYTRpfkOuBCRm1xmT24nXIpPtIwJnGsZKXGVfvPPS3sLYJ5n8XV4OLR
o3NzUq4ihAjaHD079cqQIbRgEl4FbfiB81D3+n6pW5OokdXcLRfbh1jy5N/Q0HLU
gMxdq19YqIv62233Nx9KQb5Huu3VLg02pmo7c7xympn3BTG0tPbtWJQCx2KdqdWD
TcK8Ie8kpEgRxZVDvdCHk2DTZp/YkENrAVS/1vBbqQUjEYddnUAYeV/CdqVKJlJ4
THqg/WhBIkmCNXSIe/PZSk3ipTDaDtCLCtV4qNUydghRB35lvX5ZqbfKVkdDkk8V
Scb7olEEigIisIjVu3PDRpff7D55OhrSoJMRDvfuQfIMToc2mAkZuIYCZ8XsL+mj
JooyWNvwsFePQcFkGgOca0l2LMyKuac57dbukuETJLWp1Dg1EnRko9r2bH25HyxB
k8qf6iMZ+ZyYkno76Dk0r9W3MSMBwquFgaQ53V9c6SYywdiRPiDN747RO+BQgwbl
cpfyDOqJ8TDOx/Kdfwcy5mc1b7mmsWWBgu5MtpgoyRkrtusXmRgB/ILy9RRV/fCm
rQPceMy+iJM/D5L7CAWF6wMWEkpSJEf2rIC2LcGicQ7OCYPo8JIKOOp0uWTlZspu
9AYpeh75aqOKuhXTDZMQmFqUxQV7++zlMQHO8tAYibrMZp2Tb5KL6Q6i+KFxmTuA
Dl4NnP3wZzA1rq8Cd5xv4iuXUQ6vRv4N0qjr+ZyrPPUyTCt3d3B6hlOQSv/nbJha
pUzcvv+2pydEC/7NuJ1oTuXwSkbQr9nYyyv96h0hcLs9cEON+H5cD6rFwN1/oG6G
Rer+opB7SqPJ77aD3vnCDxvJnQFOf0j6Lzln9Y12mNfXqXmKE83lsN6ol236yfOT
Wg3CxCMUgEnY4HCJa3wnGNPjmHq3tOXRVhGTj7rULWISSwjHAO1Au5bF58OIssE8
zhAZWptl0TcVsvPRDJ8WadWpqR2sqc6PIqwTmAApofVUaMUWe+HafxUTZrd42H2Z
0BI4F5TMchTLcm7rSUFrvjBk7WOU5buBloEGyPcEauVTeksYrDDCoUDcfk5i0Sul
waRTxaroOgCMbLTqvxJeH8BYy401k/pIg/3XDv567x3ECwfkpizgTisUg2MpQLEm
rSI/QTaidNNRWCDXvq3RQSpkZ6zLYbQnBRkmuX5vfVgxb9I2OI+KMYVyluBT06ID
DDF/r+nGpSkLpusW8fa7i2SYsx2OGZvoAoihTPKGuMow4GzGnj2UAqClQ9Mgz9gj
K+dg1Gd5IsPSaRn8EbCH/idYk5rDdzQmpztVID+SmlzvfAySn0JN+5e3GOQk+kE8
tMRVrfVyKXkz5sTLgVPC1WeMWZLvmc12PBYMERP+pyshH/iW9sH7lp5Mh8zOk2dO
1lHNAykgT61xkuPLhtEpQ6Lk1Tnz6eMcrQ6YKZnSVltmTDsbDCNmrW/YKg2Ooetm
xOLuNgCiSOj9XvipqkDt/INrOqoiUS1znVoN91a/AwtarpYrMvYq51uXP14IeCoT
XM834UoefLoL4lxPL6sQhaBPqAe8vvLaxVOVDmPF8kqhscm98gPc01Uc7P/X5O4j
GpHKHPJ50UQfi1z8hOORVHEmuilmJX9d5adCYUqPTefHvXAgbbWryOyIaSB9WA+W
7y8kXa1JIx6TG5OUgE3ajY/2mPH1/J4TGsYCKt7Yr3lQ7L9OEl/DUIrOHTsy9iva
OFmcm3rWF54Rd6k1wW4nQ3SJWdyx4H1QeP+DMVEsLjx1NslDQ0J3T7wRUFdF4JEJ
sNqvZZP7eToCcXdCBB/4dNIR0GalWItoAOVvcZSMxboEzdvYshcJ23foSNIRoey4
211HdY9lsgkJrzC+f9hDzLrmz2c3612XKZyRHkpl+8uwS2N5e0rRcr7bpCtHBkx/
LKp4s6gp2/AJm/01hYwxeGVag99PfnKBUlvrEQSJDaXSrIrDDtTuFttUK3apI8hN
nIFRIBSoZF32Jn36FaldEWECiySkSO5774OivTWwf6FzVAXPJtbx5M3w7rLyRXw4
Ulrdmv+ut8k/Jdttf99B0EDswC1pjId9NtTNgcUKxi6wBjGRblsrs13ChqaXCOhC
CvioEdKOgACLjf8NuCgsp4HVj8jUM4V1CFKP+a1v9TyyFOmx08oVJjF0HGd47oxp
33s7dv2XKdmfq7P2qXoTG4fhODEeThC/clS2kkiU6bxgxsFqi4gvV8uEgXbTahMj
cMZ25gY1toFHsiDsaSGnA8q6wQulESEHr71T+4EBq5TVuPQipU8XUwzIPu4qvPv9
MA/i5YtJls1aW5y9QFnMjP9cfl57GEFy6J0D/MsKoS2DDXHLcmYO1ZyeGT+YNL8/
6erCALVd/BAh/HX6604yBfqHQD/GhWkpolPakHdBJ/foj7EaYUfPQBqPPQ93OZF+
8ehDChZmb99Q3TOMJqYYry/G3W3aE8Gg3ToudkvrCXiKEApPum14iLwz03w9uz1C
J3MWjpcN+TgxQ48JhaO//qx/lLN+ZqcmvsX4n8qOYdhuKt4Gt5nTLkevbigof96q
G5MhSlTeRsx6uiT915r4gIfBIlBnbYMQLoJcnblmgj6IP3CiwgIcOpxVlWbc3EkM
7794/we2RenY1ehJjvs8dNZtpPVh8qtkHK+brApybxwiXJT4drenllgVqUAueed0
iygpdW1p8urUzEnCAlzdm/qtB+gWw7AZt28qgBMrCyeSS5s37hMGAqNu44z2uAIV
ESNMPYNsQ5m4aL076djaFwyUcm8AKciTfaCIesCjnJzCdkSI4Bh6JS0fC+2pjXih

//pragma protect end_data_block
//pragma protect digest_block
sxhBRm9alZx7cwacGNorz2lXEzY=
//pragma protect end_digest_block
//pragma protect end_protected
