`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JB9XRmdjXyZcLBRMdMxImsGB3aN44KDjvU1qxMXunnPAWrdXtO9pLBHnkQM44uhR
CP81u0M/l2nzF9KaTSKg17k1gSTljTsrsRhbg1wZG0VBod9orCUERl8ahLbY+Gfo
W+K01DI2MZ0bsa2iqE6WYDPHPVKwub0KQ7LmlNoRzQI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27984)
Hh391SgBirNPoYB5yt18zYetwMuf+doiGfVsOpk3O8p6VG9V6H5hiCQwd0PaOfQL
xdT0H3jBVb+f7qVHgWWLuEUBhrYuB9X08rn9ONiP9ilhyKgRWAE5upkHOGdecDYn
sgEcUogxBkjTEVkdts9JcByl796e/Dnch2my7T4GbjXQtka7LHG65n0CqcUmLPlH
a7I0IUI9O9Zy1FNdRJzZl0Djd6mNzqKXFMTy04N1Df3HDRIBjg20UpwJOkIfkY42
Ij6IgUqzFtOcohFoS38WvcarQ6fZTkka7xPMJEGlXEm2/i8fAmyLGUQGsCql8fUq
LT81VQSgNsaE+x8UoctPviHN8nAOqHFjffu5sbsjHGkM+ppFbR9oIXbnp0x8jN1g
eUad3s1V8+LPCrovMHwMxiWKNWEr/7hWdP4pZFXkPYk/gJ4hrFyMNaD+Znvo8U6i
SM5OyhojrKvU1J88Eq7g8VzaSgVfZL8rQFpijf16r+KGA4Sm7JSRDF4UXsc7vlR2
yUWAqQx2u7qL+UpIFFISD913kgCs7yDw+SCLC0xiy9fQE1XHiTlxtAB8TEaymSBY
4+XQbMouIZzj1TLYdCVQZWo/FKqCQ5+w7aY6+6eZgS2/qfeS2RD7Vn+7ws2gThHa
hmpqgxThQCDbsRJxqP1UvnJPsSTipugchZQXUGXFxQ4ADPU29YksvRkbM95mUvIA
2JrIZ/effOwrlXAytzl1Z6PooayKErpPdUE8Uk909fuGo1UIZi08ztfKb/n2rjEJ
xNXZZHxbMabJuRcvmPeXi6OenyFiUqaQpDRdAk3X7APch9ayeBCuCHVFk5/xurWt
mfjdSnpLJUElKT9irXRDXU76YSG4xL3LFrbe4gm15b90AAVg1+mH8NL1FwSZZ5NB
mT4xoYi7bAiGI7rVNsWGLNR9X4rjaonK+UeuqYS8fKbPy918wz9bPgNB2mpi8oRT
2bJocFJZo5lKfO+6VRuHG4273yj4Ej0pTUxiZ91t9O77ASd2KMpogBTTB9RdiHZ1
DO3qdMAO4cAr52XHzr/D0Wf0eV49qcaax/76noplrRY/vADhgOPhurhv8LJ6pxp/
xF7Lr4/6GoO28UEvs01CjdoXE/0NvSL3C2hTV3/UIRtYuKLKWVaxijsKUEWv/h0l
ZyMVCUDijTzvK63sO9xsy1KOiDbCZ9C+ob8yKwa81Kd7QWI1NaIP8ZO9ujWCEOWv
EX0X+lTbzDVgiPZ6B4RgCvIx8LSpUYmOAg6l6qrfO0fMN0f/J2kl2eNLXxXGMLrX
ucrhkRwHjwpy7w93wn0x8PhJ2+P/P1Q/IDJYfY+N7DgmYzEtBrEtDIJmJusRz7+h
o+SR4emS/Ym2WFG5mQwC/0Y5w4n+pG1RTPreRDaq9qsRTWN2uzXGoJi2s1EeySby
qzOOKz14s4VjUea9ETdkdRzl1JzX1MvFVcegv1OLweFhw/CarRSbgMYWg3OMyBPy
4R3hg21wnbIkvndfhWeUGJIsrq+cO6Nj9obRopzEyTrMFu1Kbh/SBfqyHoJ2gbFA
nz5vPoVw7RicA5Kr17NeI0+le2MyIbXnzxcwhX45e49s/7/mbo5fyihIAu/Y4Uxv
uEqQcOj2NQ23cbmQRqa3m9CBRgcKkCnT6pszn+6oWXb/oqdv7V3BC3IVFgYnwQ7S
ZpyXM8l2u7UlIZhp9Rs6NiAzmTUPqR+ANzJ33rP9PEdq6VvMh+TPHru/tMYXLJq7
iIEAGo5ubY+f3tzme0JKvy1CeYj39dSTD0anFGwfth8gV8504bMDxeHlMAjOdoqq
43C+DThDd4jbX7wHOhB41XGIauuzvQwLYGQubiknTR82LBY+qptd2OrPFL7Oo3TF
PnxS0ZKEk1iQ9n8qrogqDMipW7Re1eskK5cvzpn3mWovT6qtY6yCnCRblV6FgABq
MUWW8Zn1gQ8wyuGYvzVPKP6CCde9KnsZbCpCHNYVrwltRzC+UbOwTf5uCnbhk89c
h+TJwAQ3dY8qiv/2+gskBhmZRQIvzsVpE311cGjSwLckQM8iZNoVVi0CJf9DT5O6
Mt3gDGzpOMroTZuT82BzwD9Iq5bNWaUWxbTd0ICtYp3zHuDmz537VsSmSwvavyVh
x1vCWkpoBxO5UoLBXkmNbXrLob4g+BsoU9BSxazNMxxE0ljMLVi+NnJuR0Dqbv8S
8e7u/oGMzSUU0g5KY7+baISaNJyGSfitE9vyLdcS58HnPTCHEryGj1FGdIsPayIH
/xtbktwwYf09zcyuaVFNWANOMo9qx9i5LhOF3cABmXAYvo/tvlE+gFTVQ65ucsCz
AOSCGKtegFWV7quEc4sJQ+r3vE0zWrnywcOqlvU2UEyXvvixmJ46aTsVdPAHVQEe
SB+KdsWKrEa0fMLDKfSd+nYnl/4TIVeVoq1jd00hktOe/knh09wljClToUuWy+JH
6K6xrY7O7SwuZEukah1axtnS9irepMQzWkQf4thHr47et/X4iynoLlyggEyhbDDU
+QS63Wl9LuPmPhEDkwRgFUDPY1fBhp3iI1mYJ5Ey1B6pgesDc5ZdM/Sj8FgNNBGE
t2ztvRXq3CECGbV9V+ZhQpydHQU/tbQ0ApxW/aLjXE3DW0aZxckHmqxrCqUSZCjo
GvrEzjTUy+Vjj9S+NvX08BwJPkzPEPwBgS+PZvag1/9TdbuEc5tWEtQ0FpborNrT
rxyAKIO8QCCmG98hUS4beFn7NFzn1AIZ/a34+WxMMPy64e1VwUe6uEZpBGQV3vDz
7oET3k8N2UhwGKHGT1QXt1tYpWDCp4rUnHKE9ki/dQl997CQQAulLd4XFgaUa5wI
Lji9dvyfni70nlRjX7MzNoi1PwUGD17ugHEe3SwgkvOUu/QOSq/IduM7ptECkA7R
lOf6oxRqnbpl4YrEh3+Hqx2QPM1uSUTcZBfInYZYe0/QbgsBDX+ZLCmakkvhG7cT
VmG5g2efDuvoA+/mN/H7Vx5LwFQ8iULK1F3CF4TiYZOtb3suVX0OTJffJyjMz7nq
nn0WXUoZ9wnRusHgL+PyFQRWFYu5jrSK9SI9PVrLmaifKcyCSN7eWdluDLMOmtnp
/Oh7weBJk9NnV6IeLuIJ9k0UQIChHma41NVqswEhVgxgGMhkiPGBV/S3rrjlZ3Qf
z1vETucGNtx/J4etAwrldhz87F3+94nGnG9JdkTphGVFPTvxB5HnOAafXsFUX0qo
Nech4WtHo+i81L36OaiDQLDzGejCxQO+Nr0Aewil73otg/+jt1hKt/qnHQgk8+wa
2YTh8e9MM8UzZrqaXVbXM3PxoXgLHjVma57VSssuPP+6dbhA7G7PHzSnjGEjy5+o
aWC1p1YKReaOsaoU+EqFEMIk+K7RPNLRVUTrPoiHaiGS2BlZB3vKgDoK660RXl8o
6Glub95fMl92x1sII1T77igKeCvVyUve7zbtGzNFlWr+Gii8s1BYaEjQqOlB93SX
dJ/5HcFY+fAib2nzkf5fR3h4hrHQT8NjvUbmyy2DpcE40DiZVKLsQb0xpR/Xnq4Y
i13v10w9CuVsuW+y7BlTN2bZ1EL8OnUG3LHqFMWKzqvQopbVYapAMQtAJLU3JgQx
Es+qPy6cuSaskiqxzNhzShvsdokrpeFsP5vA/kXbTqA4BBgBH3VvSL1mE5xQ6ZEV
76smxjhQDMW4QMHP4rRekbL9iqMWJ5VxodDr9ySYyypVnSwSM2yxm4EodxPhELZy
JJls0D6baJN4IWuYZGcdd7CXZl2d7SvsJZUAnMn25cWdWmgx9S1/DOqlHdW5C98U
yrm0LVJ5pKNMxH27l2v97gTHRdV3C3IjaMcz77IdG3PtfcloBdYjgV/cpeXGcgYS
Xi1O3gSgwmOhJZZ/GIBtNEjgSAkPDTimSu3417FW5CzciYIexSmndsVe/vryT5jN
klp6lH6K7HpIHzRCjSdJISAUNqd5tr1Z9Qkj+Ig+lD6wmuNEEe2/J1c21Tq+msny
LrRIIKFmPlHe1/YIF3NO/FD73O8gXCMjs7Rg0qQANPLBv+0u/27DbGTD9rgKM5Cm
MPyKxIfC42a4wyivRdhoDbB1aAbqo8UBxQMxu/GnFm6g7iiCfca3EVb8Qy/BrXu8
okjaKrZyAWTZ9kGpR+w94vveMrg2bvbsWsVBGAeHXYdHYzoT0PlPvsI5JCzmjaZj
jtDasQKSu6UZHDwzrRO4slMyQX0B6aSgJKzZgEkmJZd5eM125kaWjgAH9g6ydXxf
P92kGAeM9KyHaB8bTi5F7VOwhKQRlW+f1YRWSlkSeirlmmYDr2lBxagHjjVkcBSp
jVmaZ8eW+6D4LRS8dd04+Lx0ch7myVTortw5ctRIAzG5wpHh4FIssme232Ct8DgW
8dJpyVdbgxgS2P0qig33UkH3jm/PwSuA04M3eThN3E4sF5pH2IoZYzg+ZIdP0bVv
vkA8MAMp3mK707wyckvrWYdZcq5eJkv9oYgGWmh+7gdJ5mZULKMbDA9XVNTjM15m
FRsMM++fXs7aYdxGuyzLkzyaXlYV3tCFf55ehf7KqeHs567fCkcDOBXGyTjGNvZ+
fN0GZVE58nrUd8QiJE0525d5YtD+4/kkbghGVZD79NVrGhmLQwB90Kvo8d+D+fBw
ov3Kt1kxVrPYxFWd4J1IMeNbdRshN1E8xtx+8KlXYOKh40ReVR/dZhwqXoCab5M0
R8O/cwCxjZotLxLvmhhh/PjqtfsLSlOM3VgWot6Dsv0JRzT7FiXvreQQoxww1bnn
dXDuhqC84WnCsfYNzlgeQ5BBGsQXhBQ/KOCb97eZuAOC27tIpjOTNkQ/57s9+clS
7H7p3bv9tL4iLGyQ6czmxgd0nKzPPvKhUX8BINcrHOFvOpiA2Im3k/a2ANWlB83H
epUzjU41NZOAVBMEBllfBe+tQWLiLyOTjSQWYfMhvX136KyXekL73/15oAZgi+Y6
VxMAea05ixqGMq3nTZXFvyqYaU+nsqzl3XekCR6uapFwTCdEPYEugWdqyz/uwrUS
TXcTLsoNowey7nglU9+KGxFN8aQtjZRMOD0hpEBA3fFZTiVFYTxZnEbbuez8/MKg
wMjUGnXPzCBVMmz/AXkb/n8CIqKqzp/vxg1KAg0xOopZNl7GGVwzEY+zhGaonGny
VFkCHYT/MC1WsfSr5yjtWOZQUKBij4wTMWABNELMc0xrTUrlGx4g4v1w5cfQbFNQ
p+vyhghtxvWhzFJ96IYuqkHFYy+PuaS/XF1gomkTmZ8FxHhtw2v8McQvzy7dhybU
flhoKShXgRUaHFJqlMSac6MBdti1M0AkpGAuSzMQ9piKSqtDL6lT/HJckH34O4Cl
nFFtYeKL/3cGQQAnQ7Q6d6rrl+15GxJ4z/MACvwGpdXHBhPMlH+g4Yh2GHnRcBVB
O7OgyBSQ66XPV4VYuLk+2ZtGVNUFP2GWJJ1MN+ReWKxHTwSuU5LPHlJPkXm/uep2
UcF4O14wpSCTPs/1JxW9PgIA6gpMx2twVmsSMXBsDJyTkwdUQ6rXP1c5ZcXm0pZi
La39RcM4nHMhpBFvOxQa30vXO/tgsJZhvVGzFNpf9mDqPRZhFxTQvdZnsS5+dmfS
QXet9SODHkPmIW/K+HTpD5ymsXx8lEzultUFL8SQz+1fnbb0USdTQpKJL5hA495K
AeqSsAmkWCs344sn43FQbtpCVJsbMYWkH7VhDorEXpaWCBCyr9BKuq2+yVDHVTT1
Vl4EVMx7KU/QOFe3ko3Ze1/MQ6h08kFj/KwtBOTuX5C8yS16vK4fKguRzUN99ZtZ
51FMcYyCweuS3hypwwhwmpZC5T3Wg3UralMNMr6+/sK+tWK7PgRIYZQ4HVLykIti
ZMD6ecMUxtpMR02nkURVcUC/Cq9J5fEhqKnw5eB6ulLf+OQdPJEFkVr5yI7lNumm
2cTCfmP0RDAZyhQNVIqMc8OurlkpJEZa/N8Z5X7RC0Df7iZPoeCIy6IssEPUBm/4
sDVIjMgFdeonQCjBlkIO/Nj1pi1DlNOXbFCCp5CiclZkFhUWxSN3xxcV43gqUVfq
KUHOuwlMjPksxZyviAwqlxWO0fJ5F1WugGjb+oVL2kAzWLQ1RNfmW6UawdnUAHgp
vrfelenXNYwMyMLcnPUC6LygFlAvMBoKdk1KQhIxyRQUcdR8hZ2TpZVYDoLlZfg2
ST9mJWiQM1MALtudm8mY10y6xK7/l6XpKpw6X/1R5M0Ys4vUqAUKsLkJlqyNlMsf
Cb3/1jdsgUsTyst9EmHIZmSYUyh/hTAYRftz9ivP1PSzyWJCX5Bm8WzZY0xZRi7o
h8LoQ4+7ySa0u5x3S+qufnsBTvtOLXAL+4I4g9++z54Zmhj0/SEzIIvh9MQiHlr1
gFdpgDccyY1yaIvv+wueNRBqc8joWmY27BEMQoyIUge/rI/RLgKBE7o5I8Vcg+mo
YHSGR2gQ/YpM9Ze2R4yUw5RHbsv2PbBceTHjapUKM8Am/JNwLwDBAILkHNkKR9HU
YTFFYC4IIXkYHRmF4B1WCo8vMmnyT+Oh24odvYFY/6P7VyE8Eurt7IZVcBA1fjuG
/iMB5En/fo3SiqNk2K80Bwcmczqi5xFshOiBpLkjsN3sJDPjCV3NpwHLqT8gFPTt
aO7X3tU2gEoCiYw2TVufvsReHDB//4ozH9F5yieU8kbPfsfCgOp33S1RXPsmXmVZ
vx9B5kcmdlUibidMuaeo4TnkkeY5GJD3KuH0i+7Vp4Ric9UXRzNwX0bRkgx8fHbu
giYBpmjSLEKsZsnCYpqJNo6nOtkZqIRY+pWeMVIGH9GURy48VqFhQbnta75IKjIU
87IK/LvgVmINpAqdPGOb05y64xFigQab4/vSOnKQYWZsAeXKI7hZSsuxKhDUtwXm
qGwU8YO6IrAOZ8FeGDX0yTQboNadWkt7tEa/7Mm3x7rVYlro0eV2b+FhYiSeu2al
c/Mw8XXw7Hefljv98uuoAQp5Z34pzfMxnTzQBXQ/YNyG2INbhi+bGm7Bmy9sn827
JptYw6ZitHDeD7D3qAv/FRlsy0aChPcNgvddDjDUOqnhM7O2NflQEmVUPwD53e1e
yacXLlv5P4ahmMkbmgDw6dVyqwMTAXaSvW1zOZoF9NS5ZJCv1RIjpSp00RIldDsy
2fymN9NpNyZyimBrDMWVJctveXC1RhFz2ISseSS0WpImrftHBZgA3VLBYTLAjC6R
crHjvZ+9QBmsPoJQXtHIQh3PRBc29+kr0mnjQaC5GnAJ6VcYLCikmdcXq0KufN2X
UC0qE0796SebL9y5TrYsWbsyixxCd4J0J9V+aKjed0gqeci2ck/UwJyUtu2xvQb3
hxCpzIJdNOROxcySQZALp4dJUmlK/EtnhmnHjCRDu+ndnbg6Tq1VnmpRHbiU+nfN
gVuy7sdC37MyAqFyaaL37PkI/Hd2YmSkGPwyyecdpSV9o+WGrzkOjl4+18j1ZcU3
0KQKHHJ0GCjPoIAk7c6N3CdF7IkUf6wZ+DIvIBMUloMAl60Brde7Iip3AnEXWu23
E5Vl01NDqbBIRA0EEViP63FNXl8DlTfWVQYPM6aXmf0vT6C8PxF2dtLcExFx1/+m
AQrYIHZG0J2wAcKeMesvB0j13VlrZbU0UaklTqYXf+agC3sPtffwyy/NURR8Iwu1
U0fYKo3zmM22RRVyejiSDVc0DI2JhfkyMV4SCiKe6fvIsPsK4r9aDTS+Q5erEQ06
h98YXTjgGEsgHZkKY0JdcCQrDlbx3urrUo3fkNuEYi+PZXynCx5Y5N9mWkwLd/Ly
/zjBICApK/+9PvnEHdij7Hd12eZSEqhbK/vnaAlRX/NJRRikkWydJW2VahXDH6Lh
nBPtnoo4+CQieNYTf4CB8XezAaLUlFsLd9WerC/cggHloshCKpTBJVGXr0xvv+QO
TSZXCJN7UD60iKxJdYjBeJi2MYAJOYC5yVluWJTCOM7HviNsgoB6X7GVnpVLOBo/
kc7S8bhnLrpEtO4SRbOQAPCgJyyl90q4U/zZRx8WrgWSY8W9103mRf4jVzpFjPBg
WcdtgdXD1zz8Xov78K5TNmqfjgoJ6XFnNe5wKObyBCIgz5cc3be0AYfL4/VFSv5w
/MQsUL3Ubg7qdp120LOfjx4hUQQgATbgIIozDjxeNpXSTzTmE3VGDRNQf3MkunKG
eDoewF8ytYzTlV3r/3Yzwm7PtJ7WROrTVPbCm8532L1PWlfXOPHs6n2m1wBpXe9P
K4cQOEVYMnSu+6mww76Y9buten0b262voGwg4yH/WM2noqzS4PFpQixy8mwcVa1M
XR5a4pDKrfAO80tiGT0S724dF0zCS9y6xIvyzmwTwdm2VYV5Btv/qqbBKrkL4KHd
MJ79SguZIsKGQT/KXHiIZqfes+oveMBCDpYIHF8SWPYjwdWLMF6cj6gmavNU/zMS
bqrq7KU0sxQkvw1CtrvEKakzppxhsJD2IVVHMfJijIZkvimuQyLc1PkqOZEfnlyJ
Gv7Xr1D4d7RyZKDLa0lBsvs/YO5X0XHyj1E2i1SEP7pUmF1NrNoGSz4USWE1zeok
CgWOmXEfn202WaeAKDaZIUJPMhYh+4Ij1ZBP3h0L/PMOPb9yYnso7ztZeTt5q5lY
NHNTX1gNWt8ezCw6UJ31cmTBRZmS/WEc5KlYsxElTQB+Vx5Fm4cKgLnqlL9mlyo5
OXVB1M6Tt7fRndNqIC6hUMwoojqI4PMIxNwD5Cn4ph7uI9Ib0x4h4hJX6xrM9NX6
gIQVDk4hiO/7yyCx/dRxfs/dXcmy5BCw0S6pA66dnmfx3OyCffR211UABpSBHKag
2Vxkb+WYsNIobfUXh39ZQbMc0vjCzlYWn43oYjakdtNO0+wKvXOKNmuOe4QMyyhH
EEZgVurQoQAgVCdZ5X+l/vnKXnxTtkaUneRkkkYHxLxqiY27agIL4J6g959C745D
d6L8UXu37CUPTo1drfD+fRFamoyM9WaIy/cVgcASn4/CvKlpUPFeOApgqBChPllT
CdEuNtOt66i0qwvHD4Qe2/TX4N7yty/3yNeVqo9CR4F9HMiYdsoNX1g8IfByi/zv
+r7YYvmzKYgVyQSBN5VEej6rec5PI6mmTYKg0HLOB74xwLLEiN2y4n/SxrVCxzU/
a055uU1W5M+JfyNDkWF3ykv2C0x5JprFnzqnuRKTeWM55F302vDKFemb4LayD+r+
pEYFJ/NEogCwBZZZ1rCFnxij4lw/Ac2qXaA491ZqlgB9gxCX30INcH00Z+NdeEd1
s5OQufppWC2KggmgJYDv/CntPZzeH25eUQVrJr8gx8/H1LW1v/FjWqJMKcA8Icmx
qVutLuX3xPsoKDnOu8dxCZ6jGpzZl8YmuBwcBQO/QRdYm06LhhRAFmkgLlg9ANYt
YBufN80DRf8UWI4m8p68O14hVWE+BykJJOuL9WDFHtN7mViqErKd9lJpg/TiIoGZ
VJbFskXDJK9hZGJIOoaj0lwkuV5Fa53PD6Nv+MJk8depY9DzE6fxciShfFiXku+P
bpf9zpASVCGB5Ua4yVjCRG1Ok+eYFB+CgsmnLaSYAmzu9dxeq7wtbatOfySqwy8O
Zmz90NJ+v2+FS0TcTdX9GjvyjCB2sGjcIHVUpOunu8tRNiuWOWoSlbOprsUMUtvN
VZGPEmvbUg9N7IqTCVY/5xoHTtLhDnd+V3AykSBc7U1budmO6eD7NTTzEL5s1CBN
IOkRH/jsaYSKHEGOoEmNgn+RUZE81hpN4feRs8jKQamqxKuKcQIKg0LASEe+AJbu
04gACpOAkxI6bZcWmaq76Iz3HW+NF5Y1Nov3aDx+0uyFCeIB/Aum5G3tSkPGJlLt
7rzxIqfqWdjc6MtNtG8dz1wNs+zfEyP410B3YadogDwNTTi4axNfQMrebG+znhLP
PwNek9kuK70WndYdCMYuMYtNE+Z/XyIDy3ahOWePxrKm95WxtPGZECDx1DTV8ZGG
sbz9XYQGNTvVqeBhkiLulvim3pqG1lABcte9IDYpkDVVXqBW3o6la2fYtjESqYQq
fGgyIAzQcfX8+KcO1Z371N9oXRa00XGBGgzoDvghx+HDT7zTvRCDZ6eDpFUUwP2v
1YD9DE+e0g11lPwonkylxBMdJ2nfVbuMm/fWdkQxvXKICzvdy7NOCc+zDDBA3vbk
XzttIa4Lxnh8JyFBpQtLGKJFyVEgdc5Y61jp/Na1YWbjt53iKBuGOZIn5k6ww501
2ePQ72fELLklEMqvGUvTbPHVxXQnBKmLi03hfBC7oVV9sK/inEaxTqZaQ5ptIDLp
idap0IrR+HQig8GROQj9rkBmKiOPVCw1VdO5DtJUn8x8SKBGXSTDc0sjn2c8/Sqc
+8sI2WVNWTJ+c4N5TSPumFJMm0LQwa2EKMF4U653pn8EMjoKfYQp845osfRuaW/a
oQW9m7YKxi4U/RJR/BDook5TsfzlBGs3yVi7nYuofn6TadlmHH52UuX5AxUnGVrK
OXuAtBIBIjDKiYbgItMBh742LR7cCfpeSszceHd42WU4X0RtNgGSLAZkbAijCnVm
C1p2NHpCPMeScQCXgsv13m8IIughfm2mhBIiARd+I0DuATnmssYHsecxRfXFWJGH
oP2xNVAAxs7eiJk9yKYGnJ2q+Mh/sAMeh24e8OeZpJwf8nEHsJkoh3hZdwttkQpz
QP2VwyRM/l7fBYH712oZNKUt/Ibe16RrXCLFIHLjM6gjjiPW27AeK26GaU0GPj8L
HLvCCA3heR/tbCfA8ucf9n7uq0jNWXL4L96JQr9Mndpb4nUWOuhbvOg7GPCUbrwm
JFmJfPeH7f8EbXW3b2O2Rpei/Q69Tg83LDDL8OlqE3cvPr6w2IN71kMSMD8dSzl1
d5PSngQPtItG2fOwpT0cP3a3EjrQ2zg0FnXyTpUEVev1LkEHxWRgPPTw/lA4/Pws
tIDa+rhk1Wzu9jea64BR0DpRvxwG5e8EvnITTvzBFGPQO5tu7D4auj7iasRmawuD
bEr9Uky8OGL6709MjG8k1XOWm4FXsyUoQkyU49d6uaGTOYGYHsnRtUTi34I6Ox5R
b/M1gpyTXTJJvJmsNbiyQLIE4B7c2l9fFW9KfcRU2cRizX9J0zmy7bbLZfFfa1RJ
nep1dTYMMXPnMFN2btIhcJg5UCWDFxtC0q7Ba6cMRn8IIpgvjrbo9/ABd4aRwtfK
8VuPr0Ffl18YRMp/p6bBHmWkmmUCA/OPHz9TaqRLCmNufxGiTcFhKh71g0vPU+SS
Nc2qoUdZRBOWuTWixmyLjoQbLLUtnsPY6dbwbLw01YbBPTBnsGPLi/7ZH78Pdoo8
imOg4ND1k/L4YZpgyIr71GQ7ZpRMECQGXH0ApY3HsG6YrvX72tYLcJ+FvNQ+EijO
5dD2yp8YylvBpDPS1F64MwGP6pZvA7ODiA04L9Qv6JlcXUZYiLsIzYzvtRm5J/BA
0GY5KicF5bVEfuDavb3qmLRpfTqifdb3yGkIdo5ecFa1aLNH0XH92DlP3BbPwIb8
ixktM5jS8Cs4b+kD7Ar0APp+rL1H5EBZbfKAjj6Ena8td1RvmHGk1COdCtBQNhWR
VU3ULpTup9SmVkEiTCSL5EUoga8UjyExF1HYZ5gZP+HXTBr5anajMZIG6zjIJUTB
sIVpgVMCCO/Z+JNtY8VucWN/J7JoO0VxqV9AtWTA+sEkBS4FoHwmaRYUhTvrUO37
r4660pIv5DP4A7jj7NV0UOAwyGoJGPVCdrq8DIr876jkrwEeUJripD/+PIOrFSdh
qK6m2RpkK0IqTAPTRTpbKHc50N4og9sIytWNq4BG+v/x/iluF1yshV0FOSgf6+jn
eUVVSeqSeAkQmpYV0NdqMaCeCoa2VJMpIIhEJuKr4ru5fxjXId/Zy7uMrLYM5rls
e3reRSc/DoBj7K08zwmWpjoBlU6Pli8ui/eAE0jpT8CBILlpbMl5PcZUk71Rjw1V
apx+hGuB2cx8ProEa15Ud/fhrAduOqDgmEPV6RC8SDPraGgz3jli9rYOj2fLAnZN
HbJthZ/ExwtbIwdJMkNE0VNqx8UbE0aPyGdYtGX1tGcujRc7S2ND3/hfUmiICsow
d3YVay5/Pt79c8Cwh59nWSivEjgKljz3xHJIQ7uhwi9bPyGFgVRSR5PQCTwNQAwg
MS4rny+Uxpd1bZRNjrcN8QUZKhl/Ofc0iVm3cDNlAVj6q4raG+VZeKfN5XOxox2z
iXfp+qdLI9p4W0tjxmtL8jUDbZwZVcfLPyYX+GcvIR0wuXfOQxfUwiAwaBotEBXA
yAZvYJD2GpGBpuN8/q5Ikh6nc53XBJz2G2OOxkaWdiznnBiR5/kXGvFS1OEkb3LC
9fJ9u3lH8W/B+s0x9hY89bl7EOt89XjzQ+5hptNYtGmiLj/nKlIMY2OFN0L77QTr
wT5qRmrTbxXJ52DgDQQq2fec1brI9BXJsdhfLrSF5PX7qhj/+MoZM/KbvOVd9TVZ
VclNWGBtUdXEijLrg6GhK5LuhaNRuO3XVeyMXjeRK8aq5QJ8DZfITTMlKzs1IXPC
iY4/k6kUsTjs1vSgPf6svTHq546oGrhYLvU1+lsxyCLp47yE8wti5QItssTw/8At
rAO4mVavZ23bFQxgWkiUjw3HGEwfHpzjsjiJ+CFGptLCFnk7APGmDu34dWP0gQ3u
3a6F2hVtL1xoZKFNzO2kKE2+WbgdLApiI3hE3rr4vq6ztCUkBcKaKKLX6lKE/PXH
hgRFby6nHQzgEppEOb9Na0iokEpywvYffF8/s9Hmmr1jrCSxHfFFgX65r9153aaq
UK93ML+HDKKceID7r0YRU9AMOGb4aBDeElCZGvp0vehCIjap6UUfP7VkuOeO9fPa
OdIMaZ/OGfJhSbDZg/ozapmULKObostXw57J7cHk+lXB48fohK/BB0mSBtr/0aTR
kDNSF6+SVtvYr+E12oEc3xMIQ4wMI4+jbLzHO4U10nDX5QVePe//yd6ZjmW9BNuR
u9RvaHarCVOyZFR9m0MLfechCQVaM3rBUyZc5H7afwp/rvZCCERf/dtbAPKpCyEu
B+6MJz9JWOUir9xgeuKWYDXrk00bLWjQtAQX8wOXQnlTpWYTj+nSPUQ6j+h3bzZM
2oTwabr9guo0ggHMijlE9atZVuX5G3gUp+ppxIHYnKURA8JzaavJAf1AYwq5DOjo
d7+fJlFuByam3xDu2PWVrs0q/QCDNuejUxKsYc8aLVWP/xc3YfMYg2beJwqFtpYK
bPPeWwZb3n10MBQMwUvadP9x7+uulewphzqlUwtTpKAuZ26kNShK/jKwhu5heckI
5B3O2KN8k/U///jrsrK7huMGBHOm88w/9FCWtFvYYOarH0YZh4uzbFZ4C4WVGGIA
Bo0FNrdmiWY/8CQ5OtrUBkYINbmatjFYbZKMhK3ytVSoyyz1pbblyXD2mn4DFBZ0
+pwEB+Gjy3l0wqn3BC1oEW2ZakUdik0okN8T/XnqdjkBNS2vjVNmay/uzhxdnkO7
dBov2Zf/fZz1tSt4E5nSfJXMEn2hiokCKaBnp3JO+KQY2VYc7Ch28X/lRWf4XxIR
fpt2Gfdmxp2Fziv6UE+5zok61vadeDhm3aAMQuIM3prSafWlKCkGUpU8ZzcQtKWO
O1Vgw0Upc+75hajtDiaV2RkzDbbiAXY9ALFXHm7YUX7QuXfBIl7lMco+IvXInuiT
hAg205ITbxauIdJlIAk9C8umKa38TbiSvNOI9JTU9Fcppn66cvqF7yyGA8pLPHPB
dHcNImwb22OBKi1Mof6pu9LnSzklE+pMM13IwSUEthpVSXNQJzcbixDLzqRmG3Rc
2ZU6T8ReGyqpV+xiiHoimZJOfCeIxqoB2kHGm3he495fbzZp5ASd8XmPPrBrjb63
sdVT6omUG4E73s1uwlzojEB5o6Aql+VgqvMsxQYOdn3Wku/padG6qmfkDN33ygu8
MkOWyF01SzlG+aTnKI5uu93DkCFwjo//1Sk+x/Ov3QvTCQItViuyD5M3vDvblvBJ
dywKNQJctOzZgvSEpsPDo3TZneyw6yUwhZANDIjtgZCRhO3oRX0MCKjBZ0QoQrFS
5OnRz0hZL28ZmwnQ/k93/NEeY2Cywyzg5uiLS3LITt7sBOyNcT05eMeTD5z/v0PZ
i1uWWvYzf5TmgJhykVX/Z/QJ4foqnvwiaPeb8ypFw1ZCpLIGZwtZDGfPy8w9+mEG
64Ucu6G/hqIqwENzlFRPsBtDus7bUhehYd0zEuIUIjuAlX5JNgHm7EQwMjjKIMIn
fQGWqRX1aqvALb6BgcAwEpt1fHS1PEkYl3JVSZDIBGpNJKWiP+M+i0ecemAnaLto
5kjFb0mcgWPvd7fzq9U7IlY+Y9FniaTC1d01njM6IX3SzV9Jlum6MhEgkwCuWADV
Pc01ARPXF8eCAh7Uz56RM+oFv/mibKz2nii9swqcxbjmqwdgyfdZyk9w9FL+SFUw
5eXlSErz4Qh47yhEkai2bbxuUwCPTK93a7ZPASjvd+SkXcKxPXjHMrurUSWfkHMj
uUoEEoVlsss08hePCPC584KeGw4X1CrRS+2XVmanDDbuZuZ3CDkTNgSX+r/vviEO
iU8B4z+SOhMOk/zXo+f7UU5ZKn8rYjjqb4T68/cky9PPcyQNKeGy4xTOGusp3TCJ
7MBoZdN4Jc3UymDFMOdJUZOvhi7rec7uWat+9glH6PQClM6zQsun/i9gKYVIMbKe
Q4brmR7ndSElaiGEDCd1isCnV4H2M5o8rPQc89Ozj2pJol0AtV5zkI2CtdntIe0x
GTUO6MXphECnlRQ8bOFA3Ywsn1Y+KPjXua7DcdC6M3NNggweSMi3r4NAJhnwJ55P
EHtNmSvY91grKImhTScdDygNNfUQIAK3NAGqukjA+AyAEjcSlA4XUtljn419cYka
sznWMS5vQo+52fKaU3PpgSGI0qX8GUoBp4J6m4g1BLDVw9hjzFhb5YkqUVmz6S3w
yRcavKFHWg+Uvpef30HjgwRAyu38Som+WpFTVDGpJGJ7V9WaUvr/mbW+X2aODpjh
xc4YMb57FO5oHeH6IgjEYs9ME2fEKkRCQ5wEV4Z2FEBVSkKriwVUY3UIEU7UdbJe
PgaBXXErErsKl9VAGlPOWhKxX62bbfPNCiiYY3M0CL00HaeZfupE7Nx3nlbjFsHa
zyXthDLO+aQauc5/MV1CquGizs4PqquT7L816E44a7GcbpfXZelIiFg01PV/lCT3
loMM22DZDnzaxaQzCAxJ1JY5hsXaCW8m7dOVL1Zj/pPykllj4X3YiBag03puNOuu
h9X/W1RzDMlmtI+db7/ZGY8aKTw40h9GJUJbikKaZw5mPIx+qKNjM4dPlprcUend
ecNwlNRiTTECN7DX8Euqz359/1BzbmpPACuCwhCXEDaIkd6N28n6yx8fnR3rXkLi
g6upKS0yGqKiegO7rp8CxBmAEIV1Jc+9Zm27oxBm8oXdkm+/gLikQCrHdkims4rD
vK82Sa+cn955t1pljcecyTPy2Jctfj413O6FCeCzqhvczUoUnR4B+i0uWE2pkHvR
qbxP4plxPNEDmjGhCKUG5wDNJZwd/l7bYGpdM0VfhsFDwCctB7nhrDb0duKaCoyi
ZIR0aMwrL0dOzR/Ti0nThxAaWRJucjbiQfhQ0DNE38AuXp0fAtYBqcyRi+3kuAS+
Wr7Q1qU7yEuhdAWApDiQcBa1KTfiX9wW66D3gDOWGaLHHP4vLNp6P7nQo4l4JGGi
hrv4dvTqYqvCOJ+B6Oo9HU1gzP1eMnWuCFgx99EqZr/cGCX3eojjfokXLM5J+yFK
jkiFx9gzYCcPhPRjC6Te0u8PJd5wVHpClGDEmepBJfnNaRdBgkaz76YFLlI4SBq+
RgRFKqiohjRverPcvTGzGz9vB9VUdj+TqYNwKL4TBNYAscoUxDarEJcemn1NSI41
IeqxHiaa9vMkZxLIf2lZX52kuix8j8IFkquUwQmRkzOxLMYKbXeGRvktuLIyqHcy
ErX7czPiJbWFl7GyPwrHOa9N5oeqvsExUt6RYKZl9rF+o4w67trK07ny8Hcn/pn1
NhWeQhn6E22ERvvDbG5Z4H/cRyPc2p/q8TFtoRIcqzLI52DKW/iVV+rDR8I9bx9u
NHMja5XjdO4H5i1aiuZd+/lowY+fROV0GaWy3Mykbvcmc12094C7mHM56kdtyrPS
quXwTS4n05Rxfs753dyEAobBoMTuRWFfMZ2fKTB/1S0WgaTRT6AVO7ZFlyS5i++r
vXLfCGHnDRQAWeqvKZGzXaAwEEEyvBpogkiIevdRKvWjcgH7qUuHu7hWx6CK8UpG
rnH8jRa+88EtFXWpy9l9BOcKewHYkLsy/4u581frSwk1j/rmGbywsBNSTv9n+9uz
V/4cZIusfeW29jTWOlwJanqGNJCQGsC6nfagfOc0+cx/dPPTRNN3AXnb8tq4QpIk
flT/8LJTHvTjZUOxTD44NB/qn8gPXVXGqpIyYNvk7DjqatFEzzCKmiQozt46tmkj
/PrZ8sT8+GwfkNCEVwc/DJIinZAJvFHpdZ3CuFtEPhGiMH75jujHiHb+isQZDIht
VZzhSMW+YcZU3jMg1tGoBFwY9fR7TjjidgI7Md7qxLG8G3MZzjhrb1+c2JC16CIO
msR3tDH/jGD9jI76ZEzliCiMElbo6yrQISAT+MdbXMXlnzGXPnhYgA7yDLIor8xf
as4pNG3mQoDwJq4nemzzaXAwrSfKRQnDGXOWYgtI2OYzRGt4+UTvtlPJRvdJqy+U
vfVCy7ZOdfo4W/udFw6O21PrpR6OdsT3lbJMj3hIB/5DvI2ZuAPfh0tWsdmc2zSD
otn2178mqSj/YRjxQ9sOIDUmGwSYz9P5NyDHRdZlh31E8dhafla3KEFP9uJc3d+6
czAm/Bd9YVFZZ6blF7akSSpT2J3wouL/Y3eglXdBD7dFr0E+c5iU+ik3+uAIzyb2
oqRGi9SKDC8ehJi9ugLvvHBuMwGxHsk6Q83lXXiUBYGnXJRnVfYufXHPTaAVeg6p
cw3Js2XWPbIJb2UbIvBrWKqbCjwMrkM5D7Bd48nfxZP6Jx+/GtliYWDSCCtXY7Gw
HZifg4A+WQr/YeSvwyN0MvLV9SUhrrVLkUdWTSeKn1XEDAZCuK2H15Ll+z9GYZqq
pximCvXFgWbVhtlvWXQQpteUI4AZBrI4vSMCA8vb+7Vcswct81VrlBgos7+q+jpu
tbn+lRm3RYvBJvDu6Az4ZXr+1riBrkoEsbSpx53fEr1i5GOgChcsBf3OCBlmpcNm
RC5IEjuStLiwtSmhEc4rpZ3ooBLGSxY4EB6vzlfM2r5cXeUCkBWwX/MVuroWBrS0
G1mCJ41CFXl+u7b8jZPKaHpBbLsRyYjA4lf6RoS+m4utGgWADxdNDJWtN1lIEG/R
Pck4fE9IapgwS0/2iu4gneZUfgb19wlNozcaxypnUvDFYt8AhFtd1SyyBSXPmmGM
LGXrknlphKhtijae5tgOtK5oEV5VG2X3jy98Xif5y9vPS9V2v+oYRGvLrpM+Q15j
9VpWBRKqqEsqFfWmlCSMEU9M825PrsxkuIkLGcIJyisgwiLvSLFxgV1hPRpZzFeq
R2UUA6PGwrESNaGxqSgpKXVN8FtMg8GfcRzLd0QqVAjEdiwT1PFcHl1KRFSREPPN
5441LEUGa4R6jWL/9Tbd9fflazluRlspoC4ZKlVEAAEjTCJF9xi9a7u8Shjtm2a2
6Dn9jXOXWEMkHGLgevunucf32WNmKDIpH4OcGhfBEhD4kGX1rNhW4EdqmZRrJamw
9fesSVASDf5fgYPir9HTR+6uV0xoRE6rRJin0wRWE7itfxYKIxVXLDmVd2gSntWQ
SQ+BcheagHhq0BaP6JRIliqZ1KKVWqNsHzvnzKak2FjlD0pKTzoXOPuKZULgrur8
fo4JM+H9E3rqD3J4pYN/puSkY98e0XiRgXFU8Ad6JvlNtijJ9kxpeH3dGinBqa6f
UAJFsMTkJNCC1gxaxAeqCyyU/FcsA0Igo9cFfVr7qrdgkGQwWCaQNBx5Z8TznG4Y
dl4kAFhXcUmGxN5ybA/iQLKXVWCjrILB3on8NZjGvY9yFI2Z+9z3bUmosBUbNjY0
zjWkO8xXrf+coUzjVhY4mqPJrnHChE/SXSS6XBhrljwEFEHcb2wfDsPCMak0VBGy
utXtdduAkiB5chUK1s22NyGIKCqVN0tyqN2m5FTDgEk9iidPi0ESG0+BveqdCppU
DePcIMl0OaaRk3Mj6z1kFZ3OFe/vbO33tGn/HbGNyDdQVnZyULy1FN6ZSoNHeYXq
G9ajXCsK4sgVixOF681Mb5k5MJlTb02Ru0UbyAXBtOoNmpF3TSP/krGQ+R/omc8F
YL4AdT9CbB1pGhNm7+XonKHn5Ta2/RDe7go4uU53qf5nQJ9cAdyGDYH48+g/2g8V
FpOYELi/T9jMivZwpAOxsCcmPOddl/V2wVbifhxWRhtm1Bz7IyqxnIPnbY2vhvyj
aQPs539Sz1EsApZJkPTJ0dSiMZ8VWLVKG1AjP/imS69GR5lv68U17du97YTJD9yS
YJp6D3S5H6Etk2LD7tyStbMZeVLS+I57aqV80rahHBrCVe0hfiKmLw5XBTfP7uCH
UqzFEyc6bJ+s2FmR21C219pYcTtFN1y3594T2tYKKwn/dm3Kev3PEY1X2nBkiCS5
wS0cgjWbFz+h8bZRiCdCGsj765egMbTRLt8CwC6qP2DcICdtFxXXaV2IzgmWg9nB
YTEfxkFfRb7FuHr+ntiwz81GRmqMKhltan3bgOkKMkJbWkEkv95keqfYT7al00hQ
nVSDk9kUM3KA50z2TCHy27uhlF3TvpKq0HaUdUyQ1EJOALL8FpMzP2X03Obkocc/
7JmIePzeEoIOTqf5TVsmQAuwZRG/Ob06iUFyovP+bwf6812yxmXDunXFKPW+oYGN
HBu4Xk4bndV1KwZNw0qpAbVE9WFBnVFhhzIt52H4l44fx7wWXIhnXT4LE6y9Qaze
Dvn4P53WsV35ntPahAyfsG8/N30CT5u6tmhg85887j27wY3ll0kS9CIqfwCpludH
GcaZaCumFq0AErrDTGdOp2lHerCOTkueqcfI8ED+cPYVQ08PJrpn73+HPhNqnuRG
Umh2sSmcO0TKSo/t25ukYL8QHGPu19e6BZi6u9qDIm/myhUTMQTKSuHUsxZS6JhQ
c/e0Ao6Dv1WMFyCRjupfnDlDBlzntB9HvBAUf8La4aGu/uhGMQFERZDBlu2HffIH
I6wgjU0NeDLkWW0vGJjelOVYzHp1NXLiLoDNWrN5HCXUjAl+VD0gmarOxpjteKv8
pyA/BNcPRekRfinO4FQCya9fYeLoU6is7RFkfHkPmTvIn1qKsEkZgRH3OlDkAjEN
20miWEX9E2OLxCMWjth3tsFyKeZ9sXoY+C8F+G45RTpDdzmE+20E3ntbWh5HXdZQ
7axcqzSfy2PzIXCBY1gVfGi7vMNmLdUMchR41pNsDWtpw3Z58SwvWSlsswYRFAaa
UW9D1oU6M0371+xExMACYOngjxakPoy9fwYKBnsyw3OgjTbUCSjr6LWNtqiNmrVb
OxQkBvCjJuEJzPubG2+2Y3M3jx7RfV1Z8wt5Hp5SbFTZAjofHoGqkRGfBXIxT9kQ
xI8YFJkp+PL3qVGOPe/wmDxJ0O9h/qF404BewyPeyk13UZFnHHswkpLTXeKU+jik
d2oE6Bj+/OFkprvTyVVTUqFITTvuD8t6SsVpG6wr/wuUrSxaZPx/sVR0AY7670QF
6a8+I+WBsuGn36a/50aUBMFmNeZa+iTRu8iN461tijWXNovXH6E4hjY1V08y7fG7
yZQzvfV+XDyYV7p36Y/riDdldP4YpnHWpioy3quZjf9EGu39nU4y7DHGoAiWRZVH
eqxDBeFiZzFS2DjRTpXMVGFolL7G50/sTVH7NNxw1g+xLGBmE63LznyCK1cfy+uT
05tALWD0Kx5jb2ZhDyq2ixxGZEtzeWK28VluO8kD6zCIJbAO3OdnNsJ8f3ypNRgQ
F4fWFtTCr4+Lr5oMepMQFX2K3bHPJqrGV25/Kmlia+xryBB/DcWT/Sp0//PyYl0f
vXqkAVU13vHjHLmeghMHWiUKz6B8olyfpPtz1wIdgEBFVTAAUOo2O22Vzn79wKh1
prUcUR9ILzZH27NwevuCiFnU3yobzxoG1IKTAn+IKB83UAm+cW4mEJ2FMxwnUk0n
MtLrIziDx5THMzO6nDk0T0m2M+hl5yq1EEBs2DnxawM92GcGrNgnVWry6wTyJVYm
gg8b+WgsfSrMBbQ9caoN5AGOQJ5hgtFw5Z2ElUvEpPQNe+rbti29GSVQ8xJbx2AS
K/c89zy5exzFcwi8RN0O2JAcd8EZBdhbIaEleNdT4JvcrrBunxLcsxGN7tIYAExU
GNWLqNpdXwmvt1Sg1xfeosxY5AV6sfSxocZxL0H+Pq9FfYlUBWCtiH8zwR/dFNmS
Jrcr6/KUYGL6ker3reKhClTJqMIXeM5rrJOJutKfZFA0N7ce37WT9u8b86gwnWgN
fV34C1bpiu33DrnTuRonI66wpAc6pbj0zejxFccVCJLdP0+vO/fQjpQBLQNYiDbM
hhEK/GoxHCaPZzs39TvNn4grPFRFXLeEM2zrCuqNwntBVVCF5/B4bcdhxqGtEcDf
tJiBl593d9zWd+1fKJ/AteUxrf4p2Y7xQs46M0ghjGce3mVwRsVHc4iMuw9w4H3I
RNp/ORdlo58g4Tc5O8LmRNC0P0mB6VN/VsP4Ph8OzybSk9FHJFeotRHXgRViiRN2
zp1LjAlQtyynRpHw1AB6fo1UTQ6FGIvCe3ZaDclBRoKnjZGHAmywbCpuc7YkTh/d
Lfor771cCgPvL7N9P5HOsgtce33xOGHjIPi/i+JeFvnOPMdbgUVaGT+fO01eA+Jt
Lr7EWQXTYlg55ebn1Uw+tq9aOb7eHqlhz2fb11/nDZ3Yylk09yTfY1l5AMAx8+Z9
amtkW9u/Qg2wMHyVozo5ao2ERQPDI4cyUlb0iSsQxeaOTj0Nn6oIrg0sAoCags0a
nDaFFVU18ivwRgXsJaDmBZVVlqrfBp5aWP1u6T2Cn4Ig1tSS+HYar+e6Q4Q0nv74
EzMyYE9XMEWvbI6vKZoQFRJWSorRurP4AgtVyv1BxLoIfSwdEDqp8kREECQn6Sel
MHZYQhz+GLm+Xyq/cDtaYikxzQzfYZyZukvPRy9gBW6zfzmLDdOQ9LCKcryZERmg
S1BM0duYA8CVYljfHBf3HjkhAjko1H7dDWaQWdezjUcNWBxWLl/71P8QvW4ldeWj
YhdaI2oq3mtYLJvKJUxs3ZOlmbJYNzDSN9x9N7IhFQeRPT9SFhBduBCi2dqhfPs6
v/Y221/u/SJ+WHVvKsT6CbDrFlsgj+INXGTakmYALBw/ZqKsdqkX0xZP4hpbFoDh
fplPmIILP0RXwDYjRWXBGIwI8xQfMo9m1FNxyonvfkeQ2aq6qXmJugsa3vJjvX2B
heOVaFLV/LmxTKWrSYQpPfos7t3ZgH8N/Vej82gZc9kKe8wG8bSkRHw95zL4sEyZ
bEYVLYb+kYnScVzbwOrkslljkTH7GtapdCj4zK/jHYYKgb2QVTMEnB6XKzUjrdI1
vtcdTaggXlwHqdIkDGO3dlWb0nAPAKRD9MN2lOy9DszF4+IVl/HFqZySAdCm+0Ro
UGZULqYmgpwSWIh5Zm8beE4d9Fezv8+mqz731BuxzE3aL2FmVw8P5YsC026ZKBXy
WVvmOH+X9IF0qnZFxQZLY7+CEdNVfWmFnfz6Aykb0RHXf5Yh3R78IJv5GARIXwwJ
h4YEP8GcuL0aPHgOCU7W3R7kRd9MMt96SeDiZP69XxsFVIccGXRSm5ZAtp4t0FiM
B8f8C0UClVWF7obP54aHkVLuD/qLoReQnrAla3YfKurcRmQ1E34XSCxUcpoH4EEp
OQgBShVE5uuQxCnwr4hio74Moc//Ezz/d0sAM3C0PvqpZT6X8RQVi3EOcWn3QcvW
N1O1mvcXbnZ6/E5aTCzOGorRzCt/FxqixrGZs5QsBjBpPWfxcin/x122mBfIg1aH
werS7+nOvBvgzQiE67n8qfhR1oaYRp3bFSuYXm5XTOXvnjdoagG0lVCQJUeQoIEy
1HmRTYcNFJZeen4+PQgubMMpvzD15dShQ2fhp0kRCYI0ACnGcZjNya8yTw0rrpvL
dOGxi/vDVmJ1uYoVPsMv+4VQOt9jXGvYq1AiRu7a7xDYuV5e/rghSvMGo1B/JAks
/eVg7NZLj7CiJAAv8K++3Tv+5176xIHPuGQz8RWSRulLz/br5214zsuh9PKt9Yy8
DTdRDin2C7H08Lvii/sR49ExA4BSiMGhjQ/eHUkNikuFV9aZkXhefIe1SN4TcDvI
7eG4f7pxPXrkZb5sF0uHRHQfvFNa/bQKgYtRnAK6RTaunzpqn2PHFZ+LEUSRtBfb
uI2EzsU3YV1uZEj4qpH5D/8HZt3f/zm6iIz/StzboextG8cCVuvNJVJs1pJQO++5
Tb3YFxwedXoZx3k0L6bzi5BLr3bpTWY74hEbpszu83XEgkUPctczh39fvVd5cTME
oKNbvj3NNp/i8G1NJpPNf72WA3ci+cFJ6bB0DHXNPexVxgGSxKLoMJfg3X81oCpr
b4rgP0JpkertxW+mcpDUxgmqr+b9T1TMzCB/IqQ0B88abG3TvacAEX/mzPHjlL7m
qAixdjx8hr0pPqK0HEO5/Kdlvb95hzYTxepSv9zOmwQnYOqwrjZ2ZwM27hFGiWee
d3M3w5TuitD9Wed4Zv2yhNdppD5SPST8iGBB0c5z/Rq0VH8wraA2e753TijOa9i8
yUpZmaec2oepJYZnTJ3Cw8qb4UpmlV9UO+D6hvDciPuZeKD6yBLSKaBSRLaTAK49
Wri/dbTDx0y3n824fR7vLRoEmk1lGSK1HcCJ1TbHK0+ma8gCM9VlzzoLe+sO5/Pp
Sm6Tb23V2a0JKOMzctSAhdjxIzyyxCD+GNtKIzNCpWY8g7Nd99iKU7v3hdR9y8Z7
KI186SELso6cPVLO4wL84j9Aov/shrQnGldbBf/r9riTlb2LuqSDzl7zOn1fFTTc
eHwUWYBJwmd90cs7MNJmUyTBVydxA6TpLzOOe8vb+9hbuyS4HA6MHs7ccOxrisTo
PSZAFNTk7rcRBPIugzQtKH2DLQjN/LsGs7+YSDr/w+uo7j4Zcs4gHGRTf1EZ0UF3
DTOCUdOaWfYjSZdPxoX/MbL/Q9QhzH0A2um72n0O5a6+sDUI1X2rP5wTcW8NTYWo
P16SvKoioasfJmh6aPscdwTE1BC6POcVrxTKbVVBEX3Yra5u1karpRfxeyhr9QWL
jFo1B3DnEoPlyJTqot21/8DhkZz4MmEHvfE+/ZATjz8uxuD9/lzqU4cblndpjKMG
djhDb3CWVwaJCVfji4rzOc7h5pfLPIDl2wVp/GW9gaGFdHdwiCjoMtT40qgXC8wg
9YPpbyGh/a1td4RPjLLapTK/3jFk046RikiRPaavfT3789YTGnUIWD8ednkO7DO9
my839XhHzc1tgZwowK6HAMAzNnKiWvcTS0vOwBV3zzLINKPIGtAE5+MDOq5k+OaL
2n+UtQBQBxWaU0LwkXyUa2YsFoh1VS5HcqrL1j7XJV1ZQDbkcXinmfBvvUWRX5+3
lxm6dDVmFd7Jy0JM4B+GacJ1br3812yFkXcJADKYbxrpRJMuOYydUfIvtQeiRE+b
IE0ibpciD6gYjaKJRjrElEqh81qa09kmEbckW3uXA3HGDCh8XYvvQs2rpvfwhzwG
q8xOTjX/UshEjHjfaUGQrBxAIDhb532k5kw9clx6IcAYkMYUCKJ7fql4a0l+eO1H
TnsODEvubxYo9Owb1f+ef4tHeTHFfvv1r5qSL9atFucPFR9wDN3+wT94ejJqv4To
1oEq9u82qOtDxUgxNvRRDoRPDAM4nAlBOa7DI20CrQuSB0jryl9cXCN7M27qRJDi
kTL1eiml4PFLTAmRoU1yzMGIS2IRGkdlqnlBomjndrT0XyI6REcY62QavBGxcwct
xZH9QoLtpM00Q6NQvgAifL+Abrgd3IthHoyktSVccRs9mFvXYttNEXZY6MM2SemM
sWpENIUG8zaYv81Bb14R/oUyJBSgGR8E3pCQNUk1hFzn0CjcUTrY6x2avX6cn/9k
ey/mR6Qv0dciFVqt0mR+3g2sSm4cfFsEl/483XCJmSx1Kq3urVPceYK6zKt7L11D
piP0+LmRCSknvjxbeHlWodDCQN+x2EWKnbwtDqqiMYrJRUvXszq8hSt2RqQTWNrQ
/LlY09qlsNk4ouqwZrfe+geoplCC2vEV/bYlf6M0ylunBoWi5tbw0wtPHXPb3c//
/zawdv0ZymA4UMR6N6TPYeUZG/kUKBLwophA+nPz+RcRrHIrcoAhxG+WHZCifzhO
JBLoMg4+DmpP3bYh6zZp5JtqmH8BuCIEdVAdCI0cCozJnNV6I6rbgHfi6TqBRWhT
tf32E8qnlvGwp8OJu9YVWoMDdER+7dUX8tUl93g4JwXBY9OivUf8ArBPMbAq/tXF
+EXJ7W7KNR9kEOk0Z6J8js+75hJHJY+61ztyGSHbYb1ZrBw5XK+GMPIjEB+9wWVB
YRkwj40kQj8l2tqNbBij+enLZ4kBFNI3inWU0ZdotbuBXWyuPimKXa/wgXnWfV8/
eiO3k57rA05D9dPahQUcWuJcLdHim9M0qDpfWktUjNOHvVsmjFFxO8ZOaYs9zJV6
Fwn8o/9RYZLJWLSuT/8Dp63yQKwBqDG+J51Po7WS2vaVe+SXUSo1T6/uf6C3shZF
Yfw7JLd9cqQE2m+GeeT2JtsFbXNOz0JSmuA5Gnb5Tv9/4LWyV7mCFTbtPddVob7u
NT7+HIuyFzmVhci61UcLUcWw2w4k7MKBQqGOq+3SOZF6VIxGZVOjxekoXNmS8hKI
YCDP+EEQpwLSAlVkvq81J5GXmuCjQsN+MlRDVE+POqB6SeCPrjCDE18CcCPR91eA
ACe+LnwjakdNVVm4oy81btD1gPWRJpR+MjhhizExNr7iF4G+IUZ3n3Up+xSOV29P
Rh9ZV9IDY+xGLjEeFoGn9OFjRnTUXXr4epIURfv+aqh6NYC6i/0hPbWCvfEGcpuQ
FzVFTMz4AEn5ulKehQYpD9+XoNlMRArW4rUdvN41FJVxCRUPiRcgZcNDVZ/PlbIv
Z8YVhrECMd8qt8ViJ9T//G3ewDGRtNawAlGMXm74kGf6y61VQzowP3s2CU1pfh8r
uYtGOoM3PSwEYyVvFDrfcOkR6LQcUMkVS5wy9gW4hkt1HR5vVTXK+RBjY6mowQv4
OG05YBdLODIXfke364QFnBd+nGyuuGvHlSLUHATAf0f0tkOkMnKdnRfMYjXrKtnk
Lw97VV0M30gt0+r9CHROIgANDxjz1QP0+2/Q7cI3IWx/+Vy08v4+CkU1/lJsB0d9
4vHfoDtWVDF2Z0Vy+U1VOm3s+Z8Pu+DjpCHHU5DcpYyHb8SgNRk5u4Onj1qdAWpj
NL7wCbtfNllOf1JkpEewpwDLI5m6RkV0goZ88NslIpoM9pl0SBOnE4eY2ZCqKl4z
wXpcxi4po0jFEaJQcy9jrCB5Ye1BFR5iJHNNcFOORDGyLB36q06siubolWs76IYZ
1S0q/d72TwyO/bjyIlhVivpGhRAi0UrCq8vVQT07HrU9ViG2l0RJ8OLW2vqo1OTy
Itx/oa5LP8sd0CMzFNAkcXA5Lz4P57BpGFhb6TtfvskiGxlEQJHLy3A97pkXiND6
3YBJQjzByNANurS1uqhmiDpYDNg8LT9jvShY9ZTDk3RVQhObJ/UKe9PLEGH6KIKO
fW2YkbWJzIgonpokFTmheG5sMzp2FRoIS+sXPdwW4T28bRXuikoub+29DXCVsUdy
c6xu6aBV+P7u58HwSLn8PltJ6MN6c3KySywIKzaJfyuAchykVkrM9Bbp4YNq1kjh
8ISV5B803wW5IYgtJIyAWmphHdWGwaSy7AAbG0jm+W0k5Dq0TLnk6IetFy9KSr2g
UG+BCrTmi6uMnaOW0SeWhKvvHFOX/ckSQdMqxZMAGUBQotwUVwy4eK6gNb00DxSm
c33zHRpk19ghJVBP8477VczulolFt997g2ywI2woZ21MMGA+HcXm6QeqT8IpefBY
rIGA51lgkWAHMETKVm3DX+mQKuPqglRclP6mKoSDDee7bDVBN/gX+9sqo+GUV+hJ
rRlkJnO4z0ypBRiXYV7rqGPyMN8udMWMJgAJ3NpTDxpjB/Ezh5qIBtj/R+3FSS5v
xQ9TGas5+frSFVy0FGoe70/USbsXXGjaNMgGfFC1AFA1EvQtB9cOXlDwIB5e78Ut
MpFU/Bwglh9isByyJIFSqXPGGavDln7ct+nbdl1npjZWhMGm4od6AdWdBJn8ZtDS
NSghgCC86h6IYTkbh7i8Flqp5kpYbQ8SAfzb+y1MNYa6YMcxr07oRfhO4ufbUs38
Ooa+CP1kHq52MZZyabbodkuZhMxidUzH5HCb0FPVLVR4uoTiaj0ew5pk8WHRX+iC
sfwWr9FSHVCMScGynDQoenCXTxqrLXQk8H0FhdpRAY5IvMm6ty9MsDLQaGzjfTVu
pjjTKdndIK00u8Q3Qx0YSUJcV0wX+zso7Q91q3qQV/B6zgaHJCZykQ0sVPlfIjiv
eRx5H1BQh/zHQG6rI5l9zRAPYu7WA4JPkgwtTZH7wOPp7TE38EayKP9EmpuxOB/n
pTrtWFYfMkiqE9Czoo1w2+T63DxjASmzDyO4oIdRWe8f19gkG4jsjAHIGqMMdrXH
CZSDVJz/OpROIoWTTmzkR7vLOR4H+8kPcncsj34DVKYz1V4YZkG1RuqUFLv53VQq
ATWdtTEB80JSFT0QORc9WDjW2p/3OYpKnsYKhZaBEFF1ZaGEYosEpb1TT3LJPZLn
La8yIApAceyS/HqfZ0ai1jSeBiRsKH1Wuqu9sDKoZ3Npq4W8jBRQ93fgfYXWVdpQ
IMt9h5oRgVOfRH6k+CCKmvOAXZRj0XUx2iWVW+owrcqfOz+YSENbEhFty5u06Wpm
Nff8G+GOMo5Sa0Vsct8Hx8VpK89ewVAIuWzybJ03KP6DNLnHX3vcV91w1OT2h89w
RDyaOsH0b55lFWycHXgxXClIkY8vL7OMv2DozxVz+KnA26ZuQp0EwxB89Dr/fRc7
ZzGgFrZoV/lGxNCGMI6j5QOVg+vNE/FtIJOBWTwdh2teW+DY4IFQ8Ib/DpHghPlJ
+EccT1AHnmp5SS3/4av1EeOdsWS161bWvkoZpgQTVq02Pa+jP4nmATX2ETLHgaMQ
nV5pVorD+sVX7dp67N6E72pJc2vYhOPhR/EGgPI9OaJsEOgwY4+vlulCdBN6WGoX
TKEvManJ9it15XlxgVg2NaBc4j5Y3oYaQe8tAcDB2J9jQfPxI4kxt8bkojboXreg
8qw3ri0OCwr6yOGkGxhROWLuG2er3uqwAHsCxNZcjKAVrZVjZ+vqJsX5HjjFRRQF
oWqNUwTIEWqwmOZOksaLtl1S9BrF1+wAGGw36kK3KY23dp3Wwj8ADhcMmvVgKT4j
8eGTygnfW1X9Qrt86+IvVdbdTgpXC3OWz/7ZQdLxBv9F/HLD7alrLdeywXVKwsHR
Ka5PWVrMV7gNTo+6xUViIcjBjc+7kOlFkj1CDHUPQPUadJV66hc5b0c1b8CrchaJ
OvIuSDdAWmdzbhybPh6/Yj8xgIUILulMdP/kMAK9d1JMAMEBPX/bHr4hXqkrhE14
u2iN8s2GXlar93ZaZ3KbqCZYeGXiYI3s+3YxsfgnwLuFbHt5kjG4Yixtaukj3qZl
Cam8sArikaA7fzUeTs5+goI2roEMJng8F1XpW0uKzCsxjzK1j5hp6JqrGjktVoRa
5gfNnTLOWHBvaPxBHsPiW53DaDKQumJsdIQjwoEcQuzQ391jNquLviNbm7QINz6T
CwhBkVM5JTxfs+mVlvYgxrFA1DT6sxT5b0kwAj8JOT5BMLSUq4yveuK5PMREsB+7
Za9hTApy3fQDoC34G7AvCJGltwY6SSOt1mz8gx4RZHvU+BDsrDGX13Hd7yKDzU/E
b49sg+KWlcO29mNN3ZoXgjsH4CTuZ1UlGKiG07GSv8PGgiwwhcC1wtKrI2k3DYmJ
MFTBdhsYD1526Xd6n7pI+r7oCr5cg0Yw2wY5R+j0T5T1lxLQFJ9nYByWz4zuu8Zu
cIjmTsgy+lExxeB3Z95egfWdfB26k2EkrJPrCA14PJ6i39FZoNpmKsE0IBIbYrT+
ZbpPV9bdCBcs4dQ12Zq3Xvau6DboXfNdyg7nALdkA2EEbaNJ8JmkhtozQUS1hH2b
QJTPXXUz91jkM8RfzuLSkkseiaY6QadipPrBlu7pziYMlhIZ/P6Wn3dhsKDB5xdh
AMD/+IeDtIAfHAZfjRjjfSMimL8HvEKVkkIBMG6emdJMNxzbu30rGtcMQiGje/2H
BFU/8uZfa5+LzZnU0g9J2CBtcN9B5jSux+k6NOONLIAuPC7jMu8JywrznnmUh6ru
206n3zFU7cu0L6VQURvRDkYvBE6xWWuNzQibq+rAGMcGbTqXa3GtGPCSFwavMCdO
XmNod63skFqW3BnbW6PzRXXyE3yvKjaqbeSbNxR+abJqYPcXi8nTesDwErVvb3UV
0tfW6anxlC/jlphdaT46t9dKgj5m/2hILm0af3i7BD1jPaPm1+onIIx2uiMDHTRk
23FICRxzDjZBHiiPnjj6U8fpuM+JbaMqPueNIT4O/HXPLll9UuAbqIIIJIhs9jV0
R2fYs0PeYKthmaEHiioj5nN4zBjsgB5z5YCCvlbTSxJIrUeYmAuoqZGhMBYGAAEu
45cuja2gT4SNjPVePPWWaerc2T+JidEeG1cPNXIwB94sztf6RqstVPo/lBGdrRE3
LxUB1VJg4wMxYwOxGGWUMQkmZliopdiM9lMMB8KcTq492B6pD3Y7Pji4ixspyMRI
O1bZnU7YuVJTFX4iqYBfUrhu+tOagT/TJ7VGEg4S9sZrJmfzPSVG+jEVqDRpPSpF
2YDqH12wJdUecIVsJPWicc59qPhGrISQQHZJo/jq5DSTOYuMfdk9quoHddAjEz3I
Z9j2XVRmhlxvkDgpcbW3tPCzZpuNcOogtzCOuojIgOajHM6P2miF7EMhqK77zqCH
/a7p/5O+YEhUrqBSWxe0qpNorsIHyaDlpHyOJHlk8q/vSlVV1QU61bwEsMW+rxV2
pXeEzx53f7Hkhhm4c1RH58ljc971rtmMXvGmXxglrBdLA+trNFXpdahCNSzbf4RB
rGoOP2orlXQv8BGKCQjadjuR3P5QLpDiXP/NzhrBMJ7WNGMVkCPU/qCdrIsUwXlz
Re0QrcqJCauwfhVtIltXsv367YooZ46YWdb4xa5nJBNqwZFiFe/oZlsSrP4d60Q7
d0OPP9FqWdAjDJVj8FdAekKpNsgPvr3zCsDGiEewHSPusWyp20gKytHYnwJbYzN6
Zp0dePvclfU5KH3AKWPDpFE3Y8CIOmtSWIwfK5EgOaM6Ul1XkB+sQKl24vrF0j5E
V2xApvcO6sdjCeGe7abx7CQBp73D8yecRNdKCyVzKRs4jLAMeXFi1mE4p+a2uBLO
NIdbG8wVbIUzKx8qSaeBILkKPFIQMBtmZT31SuZoWZ4VTcwdRBlkBBtdTzEcOcNf
TjRUJTq28cbVjvzfjArdRz1QCVLCEh2f64OeHjXzovVK9cMaTjWHFeE/amgzvbHB
kjC/aj9kYud5tJ5YaZEe7k9hbG74Gn07EBr91hfl/HUnv3j/2MHA6M+CjPxppSnl
Sl/SpWhrazJV0+uk4hI0NhRzO2R0gIQinFk7ULI+mJwdZs9gDn93Tfh46HBkGAKT
dePrb9I04XGKoUxLknkh7S5p/7AlF76YljnKlYxr2+N0aumwWVELLF3KTjQIxerV
/rzESHAONY0Ul8niCDnVTJpPLKWYIANmeOu4E9MEzoDZxDy4CnX5WzaUbJvXeHbo
QSGw00P2Rxb4a5cZCSKSb6YQA2Smu16JDKzC3+EDRXB/2TEK8DSpqJaUD0nyUFHs
K3P8e9AStt/51MsvYENBPj0g9/ewo+5zoMmyk4tSKQdChx4giyUohvxcG1KHqDNf
EbYNN1x3wLX/qZAaBCHRsByHkT4ZMY3rr/UP71KxGG+LdrfwSXf7T+Zzf8M1IkVB
NHwStU4KFnzdy9GRq4NgXoYLKuDPnzi/EH92WcE5dAiaeGkeDjN+cdjnjQ1Uk+I1
cqiubz87lCsxw+Z2IT7BdH+7VE+8O0CGvEf+aqmiJdzeI+Kq/+KkBWCt9Fj3uOoU
mzwcZcnOTueyWwfFmk2rK1jVh+/zJ4CBYUTqv1OV6LTepUSvJjXQuurSGMEayktt
UPu2eYWNEsI4wTxXcLscixCMa4fkw2YcK6zOQF7STK2ysNoCI33M0VPkEE27S4FG
AIBPA/1XAvnF+JZ6M2WWPdPQP7GG2aleIkwpgsmCw5n9lqIrzD1mdut9sA1lTIDC
VAAxEuiiCVvrws8r8j2Kr1CYeWxLimOJIpE3f60MvS0/kHovBv4d5t/+rgcjcllh
4MaB2oquQMG1JRhZHwDqzv4W+4HtmNIS4TUPRms3RcNT6lzA5PLeCS5S5hX1xVSn
JqwbgIRnY9eVGSTGvg8iEt7shq/TpYolS3iAKuKAWT3wZCC+CaBd4ngW02WnkCKD
tqLyUYaHCPoq4a7t4n19LohHKXw8yp0H2lT9qBgKdk/a+iEt7rBoZiFkCiLTB259
JtQdHlDx2Uj3xDOllq4Ux9V4ZMBH0IU+tIHj/sFk8PJHDhB8111Qzbs9GNBHf6fY
PKAuwk0iRWSWo1didHV1Q/ybRJvdcdU8yyQHjbyx6rsAisBDhdOADTK+Z6VEPkr1
0ff45tDagpx+H7tIeKwjBfIk5JzV7D6eiG3FkcVI4pXvkB2yB+fhFV3Ws5EITMcN
UBNsFldU4xLskE2792d2VjBf2if7nJ1p3dEyJ9ZWezi8e4RgGO4zkfI/ghOamS3W
nbVFMhU+a/8fML4u5NUsOPVu8SDpSEZ7aXAGW0Twjr1O3B4DoHYK+a85spoDs7X3
hx+ZxA4F7gBncn8DDi//yw3yNLX17ylCes3L9XRKqD2p13we14lzxDE2iakSxibU
Dk59ZfJVpFWHhHLWCKlSbdW+MF+HoPtsZst0fdJS2R8VxaFfK3ehV/UsB+Wzro/U
HUdbmwXrSYjvzf/C8uoD6/1W9kr+LvZ4K3fj2xUQA5oBAaBQQLWX1+0lfLX8imbc
/k+oeX0TPUWf3L7nXzDU1Q31/SuditubRUc3Kw32aVbKQqbB0HsPjQzONfomkeAv
P38FYoREHDBKRw5zsMXCooub8/Ioavm2iprgHh+zrBziwLtjGjlJeHLLGkPjpTuA
cKUmmBqcXwy++//Ws2hHIVJfMvsyYBfScNT7Ky6r6NXfMk/mp4IHEJyQ2TaycoCj
qAFxT+L4tJd0D3i/2Mv1FlCirF42sdUmStJk3bOIma7Ca3S5yCwtqLXAIIZcyTP1
tLYkLLp72uBuEkvzmdlEHGEwKKbqEqYZcoHf1KAcNFVsEIxvEffoEc6kHBbnpYZQ
DJAnHmw6fdjIydPdR8Prq3Ln1eivbkem3F1EOcthlGE6V5VPnl27h0PKuW3DfRNO
H+7mPUoGlYrtdN2FrVruUancaW0sksEm5pKEVc5mLK03PDV7nxhJGsHpR+smsxJO
0Wq4y+ewD8SC+m46Fj24EwRTwvtAL8pOHy+Ft+nBo5s9D7ORGN/hr1/uJqXqSJ1g
7X/Pq6cUf5sP6opZF+bfWCqdcr43ANj7FoBIfbm5AYqreWpl4BrTMFTAnfvGNDc4
kl7oYZnifiMBoqGummh91n+98e6Sp+cbH9eebrQlIiaKP0PoKZD2lhzHxpE3EEoR
vOi2LRRegVL2WRyP2+DMuwIG07+z+I+QaEg1Bi/7eKfLoggfufPlZwawGgxvFeDD
6oqo1TWHMf7KPSVyFmBHOjxWvQEjDwQXbhNpA7lnMqatuUFH+clIlwD1k449xtQQ
Ovvl06vTwSHIVbg9uzibMa0TL00303NmMcv+0RHbe50RcDLBdzPwu0hoLIm4jXah
+8gQxvvxmfYI4zn3yvzup3J1uTd5CLJGQRjq51YvJcqLTxU1jp2pBMK4JtUQww2Q
9rivQ9xBwFPeLNx1V2OCQSxrgJIaXvJfKy0jpreaONyRHYSo96Mfz499bdXpV3KY
IxOQ+FdwZfoven3FZQTOSztBeHNogoXWVhFG5yLu9s/ywkKClmK3pKXd88lnbCmD
JqIEN4EaL7HdaOmoo/6EMD5qUcn0TFp2PM8BaaaH00GAI48qqIR4cUeSKNDQvAQN
tgP9D90gBmsERB5QB4n3S+98AlEa+8j8taw4zWus2cVxLY8q1QHzUvZDNJbWQVfF
MGBSgFZKPGm/uVY5sh0tLnC4rRKS6ahBGRV3672QOkiedT60zKBzC0C2XbqA55te
AjMF+/dIwdkUX7G9+RGoXiqtjul3t9oeEOFpIF6YdKt+j/Y4ldSPObf5KF5H2ZCh
K2pUzRG1aXZ84ov+2KHZEm75AK9SMO8tEO3NQe7v40vQONgfxJx0g5QRNV/a8CUR
vDforrAhNimjwCqOjxEPO5ePcJ1bx1PM+eN4qc62jOrzLsK88F0X1R8lS24ZPYvz
sBOMb5/NM+YTzqM2Lu63eai4Ophrb6k2Ui323NHYdC269jOdmy0OkUhZYqZ0lg8z
miuq6HjxiqTpwfYFUqX31THt9aElG/WJiE+XYNPRAmvSJS5nIg/2u9A2acS95soN
tIapGu6i+3cZx+nSFqYQatw0sadKxyQkwyrEohYi4Gs/ggDmBxHTr95fkLJG9q6o
dfdRGVoicwxN8umhuhZ2qe8LdcrVyp7Vh3OzB/gr1C7S7i4vVuQQ3YproLNfzr/4
e/VMQNDV9hh0Mo/vw3yTuJMDyc5gtbYtcskMei+H7GFfVb1/bkuvvffuzf+9a1GZ
0vIZOyZVf0PkqQFuMhBf6glVfT5LmLboAyHk33n7b1aMaXAz+OxexeXSsNOhy6xV
qBV+nDNUgj5OwCJMj8Te0nVEd2QIyBQcZ8lZitwiq2wK5oMFfrEtkN5y0jjT/BkB
TPGq1yQelJrYdL7XqCD4xHiodMYE28ciUAq36UbDzUta6GFHZ9UPjiG4cNfkNsJ6
bskPSgZclj7LzS4liCodCsfT/TYtTAM13205fGMOzdv8nh61eAhvY5t+ORJduRx2
y7m8AFLRNfY4Tj28p7KJZKS0vL4zJ6SJ4u0olZp2ziixkkqyLbi9Iku7xt2WjHP2
2ZgG0SWmguAELfED7nAtX64aLsmpbsknS4tTKuRM0musWhjf+khQc8DQdKY7lupM
cqWi4hAgKDzXRT2ON/50jKQjI2hwRSzucdCnKoE6H9UDY2UcLk1KjASl2IkunaD4
gpdyRaWHa4TRNQsQYEkKm6wcxxnNdoY473PNm9Sp3AZqqkJAepsTkjOfvMyQMmn8
QIsA6JkkAz3My/w74nKzOzMLdH8JW888nEqquK8nLnTAnhnzOshRabu8Krq0yg5e
YXLiGCkDj2Ib4WdD4kPrkdWQMNl3obGonMHOec75KZ2juJKRKVfsCjuBTbfnHw75
5GgODnh2Tg8/nxxEVC9tWWLJhDsyBfL58ARji6KOc/tzGfIDo/b1LgnEs3RDvhN/
8blRvwXcYMtM2vc1kA1juEqJW2vQqrLJTCSVebv7GaxWpVTubS3d74aRYpJDRyg2
3zOPJe9NMWYlK3goqJTZS9dG9vztjaGECHHNVFjQyC6Yk5ZkjtgzN110jP97tBXx
trkIKdvPTVcf5Cg9auK65F63T5n11bxD1GHetwEeqY9PL+Ya6w8Vzjz2RpoV5SKX
hySvWXZdu08HBqR5yXTPqTz/kBmYr5ptau1HgQisI/rA3QN45duuO7Lpa4CmYQ65
w9fWu0D9dLwGERGjp1373CwgTyf32yjUm4Zt+a1Yy4sNn92syb73PI2YRByBUbAg
Gv7xez1AjM+MhUgBneIntMO0Sted0EHBfDC1ONheI3HkKEnxvI5CUnYvxLyg7o+I
i7ura89JzwAue3yVv9+d4g6rPsUCDkxJYRISbU4Lstq8rojSOYSr/f/kP2a+PQRl
NOpJ1xvRw2lDmyqBLq1nRQdGvzDDfQMmhAoaO8SFXuUn8W6GwwHfMrldrGxybFZv
zc42P+lVua6vXvImVyi5U/VJ3/7LLJPLt5C0v7eHLlMfbTwziddeuxZ+4nvSx7IE
7ynJ0N6uTzBWV06qAirZWJB7pMiONGt/sa9rSExXbnw2VAylKKpfJI4/iMvx0Jrt
FrhyUXDcvjrvnf8GrJ6EV8oLDz0Xi8jZls5fwnVX49+utljfQwNSCk1enzdapCqr
IHFwdT/S/TY2kk8FAprxLLg1jbgY6E0/XTCgl4rqYXsX2n4LswKPqY+0a5b3KP1L
ir7GZq2VREJaWLIps7KmMZT3GhSt/I8vekJ9Q65BhR2x3dEFB+xny8EXi0Ie7PkP
hUbdSwZbXrSEXKBd6PJ+TavnKcm1vhyoM9N4Nm3LdVP7rycd4gV2vbtzZFtXGcQT
h3lOmMOtUc1jLZFz4W+8J0zRdIrnsHzjrkvKJ3pBiyObQAhUklZyDjuRDSW6GrMl
MmfDwFO2h2g4Ruovru1ZXsfiqMR6SR3WExUJktzNlM+LVeGw2Lx4A0cLvDVUBJkg
YBnwxg2/PDjWp71TzO3zPGLY18b6Mvgn2jmSi3m9ra4R+PDlBopYcLdxgKfS/twG
SClN+ztLnYXZZyzL+WlJOgNfOj7SP1XgqpQc78ge/ZxvjinR0LJp3GoVYyXfzgFk
BDNYxLQsg3ntJmUkfr5R/bvP+XSFUrPEEjj/gmL+FQ67seU9g1x7fjvpv1M7OcNM
U5YImFC3Spg55RRLGLZbBxV3xANUXVlqbrZwVthay03O+YIK0JoNEeqtDUAMt7JZ
8R4G205ZBCDpOP0UP+ySRF8OgGAG8yAS0HEy67CrBERhMnL9Vamhg47xtIA8POoP
13JOFuRYYBB/HSYHRVVeaDwiAxSVKhSb6Her3WEwsn64zDcKabLRZQzJGz507OPG
SgwVvm4k//p1u8lPJyOg3EFnztGlXNKWXbsOxuiJHDjbtZj8rOgqRn1nO17eMRxi
QC4IOUItQb0XOXWlEEq1so+GbVWpqlw5X4C921eHCyTuTu22ZAovb/xyZPXBZNNW
dqNpAMvbvBWX4GAA4mQ0KBp1POgpVOcH+IFc6p/oJEojwdOYI2j1cnKk/DbB+cTP
/Ta25pVTHR6LfdMrU44RGVdbbVqn7T/X6C3Q7tYULUnBHI+kBJH7yc9jPa0eyRPg
6WX9RlBnyoGdx9dgraMD8zpI9vvc5yW3GWZK504QwLbfHl54YL/RnGRobhzhp+js
VN3FxU1Aes8XIa97qDzT+Gp3QzwZv8qO7WPH8EPhUEyx6+B3ZaoZxcfqOsj5/UAC
+8orCJCoAeeYlImWHQioUscxKinmZNDdPjgRRDWhfgNfltF0V/iZfmbfXiQGKrpf
faq1E8RmtjgQIWwpM1GlBevmLEROUHauVCMU9hb9FKUJBAAd+iU4HyzP9XCrSTWK
OiSRqCgEV4uQwmu/bYGX//rhLyJYtZ4relFfaAtiD+S344DJlu4Zrz9DcoD4i1O3
JIarpL8xyrXFrOOqQoZQMZgV/aAZTVLssvBZe4oYYW8KzJaCPp4PCmfR/66io5RZ
JJxUgK4hLAVGSRTHNq8OxnCLXE3/kew6bzqOTT1yVMq5LCdx5mkM+nS9seGNeNW0
/wh/HKzwKvW0Fym8yhb0vANh5zm1cPNu8JxDDHTbdGK5Q4FkeRO6WxiUvwPagqHR
mtc+ztP95S6JE82E8rifXG7zc6DHO4AbHbZxyTc3Y91WyI2KiCGJvLElskH6C/OK
1QSiGWB2oNo3GU7DjWpXhNHpJ8JFV34Sm8+HdvnuW4LvsvWHcfcW5ib97cXmW9Td
isVHbMR6FKUTosz5iPWkes+K66rxjv1lE0zbAtPJZlKWwo0A2nv8a0pXzYI2AK76
SqUk86N+KhfDmQlicUaLz8O5BFwK9XrIJAohuhFOfkE633FBkSblHSL1RBaePJ4v
p1tnzWgiJxh4VN2KpqciEiUDdHAdhCAHqbR3BPbo+cq2pDo3P8czyvTFSQevtsSx
58aTMeLCE6vYsZPltbPtdvSVgpFHYXSk94fYZMskcBOy0MbhUPAUPG5VAE5pXXHa
L/l3BaF4KJ4KsBM8tarw+975PExwN63Jw/2vs9vIWLii5co34FvvU81G5iJI4Bpb
DSQeHkRNf0KfB+2cG1fz+PJjom7B37OG6ONXYDlH2HhnICJGeVszP43Vl5J/pmpZ
cbgWq4odN/MunW5MKqNewFwiZAm40c31UW3veI/LdBpRcwdIqGPmhOupAjQV20uh
Ub7TeGoI6W7rDc9ZtVnkzsOUaN4DoG/zUUTd9MASCUzQ/8S0R1rBIvySe3BzdZd4
BlqSLwDFhYL2NFkQbmvpzP87A01e23+6B2ScjWuDAUavzdjpr+ZQNvV2hmYK9VTM
5kB8PFLzPTaIm9aQqvI3GXe0tLZNT055gzzSt0dSmHdW07NdNsQARA/OF47r+BW6
Y4IPk2Xf0iszvzAyP2DVjBZCU9cjO468mkrNkboPKW2cmEs5ei0sgze2uRDIQdQf
q+/UDKxhyUEkMF9vROZoSwt4mMf9pP7EHbfz3nzDi5iqmigYQiY9Witwyu7uYLRs
8mkzCUNGNX7Kut1EWA+Ie1cZaV0Fsdmavzae4IuywYgSRzy9gnADZwYZ0ebaefhf
DK8vxqW78DMicxQKhitNWr8MMLaR0XkFMD44huQbAlbDKGF0fElfpyRpbLfeUo0t
Dpd+eKoQK1Ou1K2loa01vgnOVF3JdGF4x6Bvu1UVmysH6G8FOv2EIxLu+vG0D+Fp
qc9KPllqIAb9/6INXPV6kORZA48Mwra+W4zxMbM+ycbFBbdJaQaM7VCEcigu526f
nVJCOHeB+UgIE8hjyDFbneEZGB28GU3a8YXoBdPUX9vM/9Dt8ZZR6c/cnF5gF6XC
sXX8YR8PCQm0naRPwUH7tvOY94dvemnEPTJk6T/y9QL7x2hz1r8mWr6xV9kAxmn4
OYqgouxP6OnVRl1eBSfr7Nb/urTW1io8+BQJpqSkTjLDyjhGESwABTXu3t8DLdXK
Jl1zKZ3y4YkZALZZDsUcKdKSaL+hCn+HBTThmPm8qyK9CPjIv6F4L+mCSombKpu+
OoDc/IV3OSjEscGbXC2RtK4/MXA/cUXIIqu7O0Ou+YdOGp9AobSQIcF8qa3rbMVw
`pragma protect end_protected
