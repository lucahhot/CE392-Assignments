// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
p8qm5HmL4WFgazr1dnQOdzNNStEwhh04xS1KIa/mhDBaowGeP/Kf/HuBrdcjFaHcQoPV5tbmmYaX
TJRoAYLxmXd3vcln7HnshZhvRIl6Ty7FmAf0QnOpVoeM4GRhudZ8eI1cpNWxPYU8w42dUapZKpTE
PfY0iI3zcLiq0Go0wtW+5inT8+Fq2vVkRDxZrhz+7ht2FVgM6Eb7YUY5P9dmEDNAD/OsrDp473sz
S+HWl8JpROho1vwP9V36nxg4gSwh+JF0UhMBga/Yf8hK5jucjsK3tsKfnrcxGaC54BQtrIlWmCVV
fCZ614HwhMpnrcRX6oKPztikpb/Z0BOZJzIIWg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17568)
4m7j09slgsaVQwPvfM0/rx2HqQpkp1Jyx38lYpuFk4Ls+5MbMjv+pNxP67GopiQBjswYUHFdqDIq
2lP4bTpjLlBrvkq3MAmsbb7nJZbosdFWyh6jG1Dyk6IvNQLSsuDrtzxwYs5WRTUBFjW2geg2lNWG
m4oZ18PzvtqPPH2bqJCzHpb7+vWI26V/Gxhk4m8Cb4ftn3Efz4GgIbv9KymBj7cGSs3N6bPG1eYq
YzSZoYqlEOdMkaaF7OgdSz9NKlK+bgkyqM15nQpwZqlh3ee3SuUIEu5QLV0CKq5xBQAt9zTydf9w
6SkWo+/yaoRhdKA4JbWyeYM3aCjS17eSXx+NAwi2LZRQXyEFfdvrh6roirgjuUcH7iyiaXKwEXo/
56VvUE2kysDMEZoEGpHegqs1O72nMog3PkCpt3wNYs6K+/uj3nJYeIYHJZJTdkY2OQUUO2CejudW
ErMmeBYVV6cE/odAew4dWAYgt9ATdtuB9OImsMVvMq6cWcWGu53ZmLM1jwAcTvGUitYo0tAqj7hO
NYYxhlNOO/Za1fjj3Z88JzYocNI/JnTZGNCxScniAYH3APLm0rFHnmDMq4EGUjDpH/7TZwN2pgjJ
BL2/865sgkXMfZeBi1mrMDd07DguYvfA6Y/ITGJDzWViE+d4ad1UzsNEGhG7RinTOn1EM21bQICn
wnazxGSbGVO5Bs+2GxnvmldVbu1APjOyaJsYntEwGcWoIgS/G07E9kP6GDRj0/j9LuGPewnNSCSz
0jgZmPFu8FkmvNGVbK9ZAje2qm6g8yJlQwgAnRIOQvM3RiKhmrWPWMlmbxqGM2WMHG6EOs8sdMyZ
Xb1r4oEXfn8pbqNouSVxpk9g9h6F7gFl6USuNWpQ0oGBVrZnvw4cgRngDtE4+n8MKxdHECYU0FXB
GjVS73asWB0rSpTlEyj+qSsFtXGeOl4yoyPJQ14SWBr9Tu/+0GhHBdPwWC57JjUYUKaLycWQ8QcQ
IdK+JLbVl1tm1rI9F7WOOAZ17i5x8RFVaa6+qaVh59tntwBuBQDwX6dznUYLHATUhESyEt+LsRYD
Cv7k6orO3MKRaFnJIbhEKVQ2Rq77kWAT8KVSoiDYTNECKTgMLApFQZpk43VsahSGSYaQ1phfgh46
yNv3c37PNjLhzcZq0i6hxwS/511zX+d1VQCB9YShjtMGcyEiVWiyqdruPqAincAlZZfSakyG5hqg
yZwa97P95FTzl+1J4Z2jAhiNCKHbP2m5t6fBEua5tIEN+uW/peDL2xg8EsI367m2JuZn7eVaIGHL
ifvIPrR+UtQMcX6HoRWePVU6zRMzPIZlGgCJY6Dq0JJnpgqAyCddcX39GGraDJS728gFFD4P/2PL
12iTuV3xr/kGv4xhpalVE00FPAW0YmH/GeeFMMRuF/cLvU4I5dT2zNGk2GNbVF/l7ZLfsEBfx95t
WHdrv4lGSWbTE08KEUMSV2kEiBBGKw5PdwN30rIJt8vg8bP/l+jZiI65P/Bpnh54irbEM1EIq63p
Ido0TYBG50w/W6cDs3umejfK3bLnRyy14odkcODmfXu8oYJ7ksfIPud26O7qqA5MZIKWl0OEz2MX
LMbXVgh/K4jffunaVNirPF0q0DT1VDtA2TwCyTpqDHp/hR31+OWN2KpflUg0WlTLip+yVetRnkdd
kF7S0mEI3ehf02U6VwnvSfVylW+VLWd/4CSuSBjLZtYTSrrFVqmDjCxiKiO61f71djN31o6aVtvv
7ul6YXRNM+3sTAeaVcfzblVOHhkqluf2Ava0n/a+WQEPDhLwyLHzVnHl/uTJTe8i52Kt4e3ti7l4
MfLBWWQU3ymL38ZLh5mm/W/60/Fbcu5HBRxjxLerMNhcllsMFde6b/btyYknH2LeLlPTpzZ12WaJ
9zPthB90l6NVVsqnGSnumQv5EcWgQjbpuxQ7LWL1UZMAmkrdOuhfJr0ao01+t+6hpvkRsGYsEq+U
VzjRlzfgHDNN7EaXY2UGHGaeDSxG/W6S1U+GsTNbKTfnPa0LxQM2bInsMRu1soJL0RTuCOWtkH1y
F03zSxlREP4EQ40eQpq+MTLakYe+0EQE3umeSkloqCQAxyZJJUMVrGYTii5JhgSM3PFCyNP/5dit
roTcsVb7Zq37ottwt/1WftoCyoqNjwlxUVTJf5Gm1gucPQ0niE1KpxWyf2/sBIEhkIW2ScCbmWtj
MQc8DHcZgjveBlYyusPTDByxzZIfwbuu8m+mZcIkMaAEu7tE2sfuq7ZsmQw3xaMkB4HKE1/V3NhX
cVs8jVSUfEVQ6u20zavS0jye05CXj8fH2Qflp4bscwJrETcnzqJDu17DdpIeKodKfoKMmbE9O1cV
qRXPk1H9AL5afnjuueWYChgj03mcGMPbGrY01hwMSNTQ8AlWoA1CvyTZMsCQXougWR15GDcmGmpo
/iQd7oTgHRmjRuw99ioPlJ/r4x9uxCaXqQ6Mh82zGpIqocMy7hDTl1zE+2U27Ojnbtply0xbvPsv
CjEsYZEZwaf5sLFM53RFkt/8MbW+/yb0eClU3FNMbZk2hPdjhuhY1PlyIo0sgnIZq8huLucmmSft
90rsn1jhbr480k340yihEkavOMqEWQBhAt2Edt1ms9eAGe7cQMV77qGdVHeL+vvIxEaFl7ikIZRh
GU62Nk7sW9YidP9h5GdkRgdA2+Y8TAhRHj5RavOtJRmyrn7kPvmggBLd2sfGoIWGMFXZwJ0nzdF+
a8yWAgF2OkJKCmlnG4HTdMEmW47pVsql2q36uwY3sIV0ZC8hM4gPxtRcWhPi2HnnxSphr9ChTTG7
Cex3aZwGt49uvX651YgCzhfEIxJMxS/XU0kcpNZujzOBmnUfba/LJJ/GSfyqS9yGPICnTg6uK9Vh
U3YZC7wUEQtCHXekGtoIoZIE9VL0MRCSSsO1TQcUkjh679Vr/KY7ilvrzh4PTRCJeyV5SJVjgnMr
6XPa13Ggo7w1AiMze/tZYmZQ9sX0jOmNyVDBLZ/m0hkrXQJXdtL671cr1ygI4WADKBeWSofkTLHE
pXEGkQZMBuKZhRlMKqzpKXxq6GgsvexJoEoLQ7NJhs0pbyiguCNM+tMGjBzP0fDi6OrDh4pEUqwQ
5a+oPlS2y0r7KrjQgEVrYaQPwoiJ6EPIknJnJa1I4NOMu5sx8jTIymL1Mu9uSRq3W+N7RkfJuClL
m4skNEvEPam5dhSOzE9kEjoz/0cI6kL2h9tWCHu8lypghn68Jktdpr609UetzI3B9Kzr552SkNbQ
AZgo+ZeN3wcGrTQimGYxx0d0R+YtevsgyyTLd87vOO8NhFljaENQLI6qNKL8SJDp8Dwispn732FN
uIZr9FrNkoKsDXIHmkls/9rx5s/Li8mYeDx31KUn6wHUFiWU0+VXOMgPxrE39cuD1mJc3MLMqttf
GO54x3X/ARQJN4Y6ttTMHTpx+em/lhYJfReHNDb07p/b2RYlOOEnQmjTXFcrKBmMWnRoVWywoCJ4
wLdes89pbeC5hwBdp8D1VdQE/UOmHt0Vy9RRCMpc3fe+AE19uAkdvaYtI2JMD+X6PjVnReJsjBLo
Iz75cxiHyusJWqimkJZopQTzoLOO0hfZfU7r5A4LB0UGN1Umi2hMzgK3IcHbssQ7O13TO02+V5yU
f/rxXjo799aRA+1pg0LAPkpvlU3sANeZRp1XrxL1NkTVM3kcysO6u77dSDg5lVd2IgpYHEhDhNI+
BCbuB+18jmozTsH+yxsAw0aNTQvVEWTVhDSSHZsTRfqEn/yxTbqMN6x7wyJqm4hVWCI9Ixggmg8f
9T799Csunz2I2JP88J0gh3taU//ckw52J1K0m63QqlU2rDYdBNaJZNl1XbDSCwyIqDuSgojR1yix
R3x7iX8TuJI5rupZQIZfScODjpXkbGQSCx7KOf/diAoSjArsLJU/il192z4L13LvSzYgsvKIZG5n
aft0URvCq2V+Onf88s0dj6cwJcH9ZWpD+2HqvvrKYS3wLjt8bFA40qcZEyygVLlPGN0sFEJgNvcO
R6bhXe4ifHdoM9c5EUFicOrvpFBaucVZf69xeWxnMmM4pVNcb+Ce4sPT18kWs8Z4KuDaA10tHRwK
F/uzviymqQxbpNTPWi3Xm92hwGJSJF1s2yXH2hN5XKX4aZwcmXdJ7Kqby1ZOp/3ti1k5P05uFvSq
K2td/fR6BREY+0D7SpQRqq1OyxcS0TuYcGMquTbhvdxcnCNf7fzonLadZoZVxz0GT/AwIkJq6TBH
3CXVWcIAoQYIkIHymJZvn9rl6YOHcaZRPQTYeFmfE3HoeRikDZ3KF5kfwY8YpIlFO2W94FlWkej4
xp3pJSahihxobm2CUsIpNFA6UmM07JhkPMIj94DIKIH9geoUo9OMigD01OGbJzWbr0vg2NqhpK6a
tud6S2izJrQy6psxGBK1UFaWq96nPJOVUI/IzuwR9vko/3yG5qHY4v9cU+slW/S57iGTTBZ4lg9z
G7kG+TXSwWoyimpMaeDdmHGHu4XTgZVBF0F0r0b/we7BVoLZFZoS66/eZpVWJs4p9xq4T63ON931
6eoqlmAWbjrKHcgXnz4669/gYHWMlfjafo8qU0nQwMA8WkpSpGzU41zg2vFLj7JXW1y5YTqzON7M
T8rNn6npkK55u0t56sQh6CtYLem5F7hzF/JZSu8TBvSNGfRk9QUQmL6lJi/osisolP8c0Fnrr346
C1lNSwBH8czvMtogHFRMR5AWPhUscIGUBs+PbXp6vHDmbrgW9fIKS5ZBFL7B3nv3RIW6/m6YISxd
V8+p/iASJRDhmjzbWpSmPBvWFZe9f8ZTYx1ko/j3OT42tUklMNWu5VUPkUlYGACMoG10PgKoeSyU
U6gwnkN69BR8Z0l7p+itK5P3KNxzcWhNNDw5brtfH7ogI7Li856S1XubDxsU5xuXLNQ8zcTyMhpg
D9+LijuY9rnHzgi1Q9sAMnIZX4I0367cQOMEMVtAuQpdbzPTXnz9M6W1uxQ8UslrqrZs3OOodbB+
c2zdibpnnhxPNdFSfBx8Pk/ZsSx37cI5OuzJgceOrwk+Bico1Rs4by3JiFRKrBIPM4d/YBqaO6tO
nyqcyHgOYnwXVKXnAHk6puvCvvttEVCzL5r1N+pWPxOPbbzNLgINbdIQA16xSvFkY8a5iRmA1naR
iX+hLpX/9iwUs1UAgH0WeE39ITjUCqywpZKzRtAp7s5xEjdIkVGWUzIAhkrsAcoqEABPUTWTaVIP
Y5bhb1BykfTrKYxkXJj8OdJLcGOcttPk8dZyglavEw1ynx2JuOf+yY3htyQd6W9COM6zgEuzBRqU
mhw+QBRRAwaG9F24prjMEuaYIWKiUBuG9xdyyvnE3f3WTucuQkuT2si2V5gux5U9bMXWPmXSjz89
i3vK1tvSdzwdxn+U03j1E4Vs5UXpYYWWwBkKDAzRR+n3EK3VT9HhF6UPY+arjKkrV5ZWO/dYhS3V
NcOBqIKEYosfNSTwpgoNDzVaPbnIwkoEEzrU1ta7NeFU2E22Anuj8Mg7boAjLpl/Dvbf/3RU+cHa
I4mHXq6u8E6Kf9JwpD8y4BaDtUgvaXRmB5FxPUW0LFRRvlwbxqMGz1wfsRHCI6zv3gyMaP28I6k3
/5VvuTjRFFGv2YeDp/o6Ifj6IPyCz+vcsO/nyx2C/2V3nqdSUDFrfPvRhjabiJPYOfU4v6/eLlVp
pL6KBg9WgcvqAbW59GKZ5s1mEvGt4zwkxBM6GuKKM4oSqgIQcudnrgqsIP4gOvytjXazA1dyc0Yc
ghCQSmdh0SzlbpvmezW1v6PMRrwdgQKTZW+SuUVnd2u2iJeQ7FBbzsNEE/DSMCslZuCLcQoXS9DS
UUg9xzg6V8a4FkJHisXSNAipFv0l/qXIcbQdDuA0IV91AWFVoQFNbV2yIkrT341+lgwIa39DHWSZ
UegPaGxJIDgxbE3DSXulRU0f3s1Ri5G7nRkZN1elqZHNGP2/byuh5PazrP/th+9B21pLS4etlmwZ
jeVGI9/h2ysTo6C07jgMmC7GBnGsZblgIZQTauGxraukA0ik29um3pjL6VSlx+M7WLaBNQliIXTn
UnwpuF6P6YRDuLlzQ+NkY5BmfYlYY/5kVRLhc2LXJwIm6o+Szg0g+yLpbuDzJScab8q19PXXDRi4
OrWERSfl1FOD3QO5W8ziHJ41B7qjI+hOOex+Im002YmlJ9BwQF+N4mE7+P6ZqPuj0Tb1LJqUBR7r
GuySN+C+TAc1TeebgGCL6Cw0OsjxPdkxUy9r3xrePle6oo0HDBalDAsRd+Hqq/stjxxNOmXVM+jy
W0SdEqhCA+b0wsHKgBy2kRHrDAzx9smW8CdZLP0GIm7Ig9rpXp1wEtMVLKIgkIaV2fdPUY8+jW2B
Sy1ZEtOUiVAW6iXoISfNyyItWEjYJ201L6yVaUCjWghZfKtU/SRznIkKImH5J9Y09fYHpEJyq7Hy
0I7F5j60aA6ziL64ww8BTg9SjcbppGn94TT/1zpg6AnjjaOaGXTkO+bz1E0MkqjQSQz6rYwbg7/U
NEn0kZUbqvb2alailDBB3EoIHYXBwQtxXVv2exkvuwNeAEWJJJnB4F1PyE+I2+wt4hjjxx21lztf
xlhaYYHaAFwQ2m5Et6UAOMMSyr+a/KhVo02m3omT07oPD31bs3uA5tiXV0DKQqK+4j8j8HLbrBaP
jymE9Uwk0YJaV1A8KpVhS2IbzuQnrmlGTaD0md0oxfhAMJfmzXRKHpThruvY9K6eEN4EC5bUTWQx
q183qRiVBhhVv7MtoJ0mg8ahEQMSqQxUbFohTzO8nq1yHZ4u+Y9+qWXDpbqBDjk+k1PoRW4RbwCa
o5Ab88GAG5vYWRrfy6/WegCbXViuF2GPGz843zPDHLZiNIZH4mISJ7u54TjGRaG/xI9xdpiq75Va
bePCOgUjr7Blyplx4HrG99EB2hCvwcAqR9aquuSkLyURQ9PUCj4KAUtRfSwwnc6PNpDiIvw4WS31
BmnTvNp/j5lAaS+UxbnFV27dGjG7nHtD3lYAH8B45fHVDtkZNS0JEdM/f23G2emPmYH2HD/KE9mF
qnEYpA5Nd/yQKhZf5RjstkJTF54jg0Hi7cqE9MBsyfJ811Le0dSWr15A/Idm5LUIvGiWCd8VhI6D
6zRdOxCr6inrnriqZcZpH0QbrFz0rwEwyHZrgXtyxchMf99o5vK8uRolv4B7KUTbbMLosLxLIOEM
5zzZ3iN+B1AKjQt4xVk9qG75seUdVYD2ScabkMVyvqA3VkSZ+c4386xcHeX3UT8Rsu+JOV9Vhobg
urwrswDkLDwInnjqOOL69A8w1xZEXPgMKVxYO55roqK7MLClaxkNlSrmOwATZFpBGGRVNPas6dNF
ri0FegeSwlwRF3pnS+eV93QHDOnu+q2MILOXs/TN+zM3pKgLaawpmY3jPkJQqZkTjC2kGqw+7cRm
DmBNBybQAk2oJa07RCvbgpLoidIz95KlUK5/4bxH5R29+AFmK5p03DFietokGbSAWkuJYg11thK9
6fflFJppEvM/2nDH/nFfqkFo2oWQcaUgnph9yrbukqIB8kndj9r/VzzPXKuuCHr3xqDXVpoYaxFE
ZBnjdSqaawtrWXrZtjQRibD3/mSooOEwA6QMweGh5xVTgb9Jng9yIVB8h3mS7G2i6sIwtqMb3Xnu
bfU75T1pDRdOmZzJzKxWZXac+HI/WbLNzaL0c1w0Jp944dXzTcohraua9eEx5m3YMccnL5llNbbg
XeSKGQOIYUg4855Q2/qyq0x1zm9C4S0uLP9YynPSpMVuX1/S8e13PjB2ZGAdDvC10FFET5NNyYcL
GX0phcDEZ8ngDI1X5O0CNlwpxxex6oVUNm1v3lY5/XD8A4koL/8xbSZLot3lNmDB/0aL18UEKIxw
L/3NKlLfpl143qNTubJyCzGJYbYEL/dGh80voR5a1JutqhDFCXpJguSJ1CsgcvLFvjk/M6Gl6tgt
VPDOsrpQOa3eXEnr2nc9HjYqvFbeRE/TMQc+FXSUAmDEC0+8VSZ4qzIB67G6ayslR6XPu6bvKZu7
OfJBSCRI58F2LuRiZnoPuNx3NfulDa6rdo/om8wyvT+vvO27442xO0Q2Rripk60ZfijPib/whZ/5
MueRQkeoEDVM6eElbmiWxjYgPRxLMTFH1+sYlacIuGq5ekR4AMTq666fHGr4cic4baUwMTFbyq7C
7U5a2dDf+zd7nMf5K5p26qAFdagMw694G3/DvQSryRPSPW7Jb4JxhLR9afLBrGU1Sj/5sqKzLplF
Yd6/adZvR8sBoRxlo2/M+MCdQJp8HskBpjd3HSbCs825dVrcKx+paBdGs/RalzZPDbbndI7jrULk
JL7bzkfWY4ChcE8+DtKaklChas8W1FUBp3n+78buubKohh3JVPbMjDe/5WV0Z/9CRaYVw/HXkCjk
wl3562Aui7M+8Oir4tjgAbCf+rXhvTecckwFVoalglEwBOujsJ7fikD6HRNG8+hsx7o+37DTjWdp
UBpzVuBcfeKU5q9sTjDY0tSGOe9EZtP+2Mz4Wb4veYS8VUv6hoQ4gRICKziyEZSvg2jI7nv+zSAs
R8Bc2JXUCWj1j6YZAYwxW22wJduOhh+74DsyHNd/WabXMPRZYACDXz0OTDOLQmZ5lYTMd178Hb/T
OSERyrlUaPjzJeizgUPO+UUxc416mGUDfc2AiT1ZdBaXP2vYuPv6XZ/A37h9tr1VJnr6CX0p5tR1
zSLWWXsmef8Euf6duAVAvMCXj5v+4jeZXAiVvFxLQOo8YZj8npkmP1hNSVxLRNxR5E+0gYp/IuYj
A+Mz2Ha7XD/hiJdrbVbAWqp7pWDyIUK+DfNIwdwhUh/aC/jzY2evZV6WCbERDotspEJCQFzRi2aR
oJft4rQ8E5r9Aa99+KhSwtWeSfH/U2Iy7bSh8Zb1yPly+hNkbQulOCMSHG2AMh7um9damU1fBlLh
OthvjqOpWHqOaCEPdzdZWX5O1YbQtLr91bcGtdiL3CuhsSwYbkBXpFxNBpgyZN2gKu/Ckssij7uX
MHtecZYMVe4ly0g2CvDHErt+wxZpiIsDvLCa7f4LO8uLcyHYRCVV/eVYXzU7/WbjoRt0gL/YUw8G
8mquinzDFFiR85TN/9WhIAUXB3j5zLI07p+IwxhF7JnlHi1kK5vnZpeuGQWoMOJ5M0pxVPhfHguG
+k8JGDyhcrMzpYpY07rMo2sA+5b4NVVdn03QV0gtVrH5+QR7inLDb1inPJNk40PDJzuFOc2ZiWbK
AZfrOaRvhS3As3G98StbeeF74lnG797yLXnSb7RZNtjXSyeczjd3arqILo2a35ELIOcb8c4qau8I
LsJ37GDeINgS2EI2bg6D1f0DNB8+u0lgonnN9LakpExLdquhVfK932COaAY9a0pgkBcTH+r45T+C
kXhEvqlaRazs+UYOitXvH4m+6ZnN4akFs6icWKWrPWxaEszt1DY7g9ue9tpgFKiO+pJj3tjbaGzB
mzJBU7Uufp3oowiJa+q1Kk3OKft1nnX8Kd1Aho//lmPhwLqlszTbQW5Z4j5h7xxkv8ot3Itc8cSw
jc6oIPod+6HYVdtnP9rszOrjVBcsOwLPL3Vnu5PqeHMRi6Unl7jrVULJkQaSVLoai11jESkSNuIC
oPJMVHvOdxhb3NGm9bEKE1aRlAqNArAG1zg9D2M904rVuXJ7y73aZ2dIc+LXbFOLcApyqqOtmFJ5
61YNRjMiOT/Q0l0kBuxtfbwdYYjd1RP9z/M4OXn5h6FyxBHMU3kFyWoE9mHva8127PelrhtYPXkq
IKe2YrwbSC6/3APPpYdtxhyD4dWkISvD4ft65oYK3wb0lvNaARA/zyFeyqFBnw6+lgq0Xw82H2AI
VY5NtN5zPFkvz05pMWyUYs9c8gygXFQYXe6RQmdSBIoyCX5nrpH8Nc/q4ZajAVgc1eJcOYOA8btQ
jeAGVscVHWNRIgRMGxUVHlWJ1RvJwy5H07SPkOCq14jOz+N/Uxvesapk0Aw7ChK5fCxVLIEWkGwU
sWs0vYXadjLWIJ+QZziBzlofBO/eLzXsE3O5YLGCGXrjWjIhGH/zHRp+AXMFJLvFrWOFr03evIe/
ptKJSda1IQsd+WOOxs629FxjtiMRRDeXxE8XEVGTXVbEvYRiMITCbFRXpwtXv9x2F/Ur1jyCWQbW
pZ7CktahzF5rBukN8OE6dJWOTog9U67w0AikXR2x3oipNYcerYj8hoRVKYiFrl/VK0V8XcePzEth
MNbxTgTSUJZByRODS6ybYlsJY4wdsbkr0sBHyJ/kvLPIhMsVfI9mqusLP1spJ7uqt+aSSEH5bQk0
yRughuySS26qbvGc8FvHA+jUX2/KNk+VTWEQtJenWp7YWa+wDlZo2PyZGUYyEo0qlQyABI6baIa8
6JWDImDIBQJHAGMub6PHhuxm5kclazHdz3jRSF2K8/D8fnc5OrJvp7k1oN4E2vgSvwdfQGrNfF1U
479C+WfreAhdUCQSwYS/h97ZT84uZvsC6iFwTPe+mlFTA4DLb+hdgWF1C2eRymHJzbnnXdMcDriS
rac/dQZP3EX2iuKxH6yOz0toW96WSUwNzGCFfI6CYk65i8SBZEdyNqCs6Nyer/lBRkf3tj/vSVc0
k0W6WTBiUwQJM8wfU7IULqwK7KrNJNs+QKpxuzDZrGFz+o9nMbkURCVDTLPDUae/2cI70z+0uwyc
4twQS8Piqpi1BWUOVFLN/qG9i7dZjsyPl6I/o9OY0bUErmr+gIaAO645ECvB+x9pv51S7knTTnuV
CBqbUcHV6fcp+ioea0fhTYxB3brMGLVY4Q9GPPpFO28EMsEoycKcb87RbsqRTikMg4NkRBTyxH9G
ZvfUX37EAsnNxLZFu5CHNNZsKVRxoliy+vN6hbpy47JVg4UZsjCO39eZbD2hKXSI+Wcx83BNoSPx
IzqZN51b+yYWK3C0rGXfptvDn868y7piYFC2OmXWCfN4hxy5rlmYOgym8o+GwniyOQE7S4Gsz3Zo
CY1aSPqIxcODsxw4rBm2rTF9Jn+c0E9NjalVgWLQBrbNWFKsdAnW2Yst4VGQrXcWp+vfE8XrdA1C
ckF6pAYf6+npjbkBxz/WJEn+xxmUiZPPEgYESKdXk+RTTP6HnFp+evxN6LWWXOVJXf5wFWG09aff
XmMwYFQH338ehWbpD34/UXozM52gDawyp9tYCXjxAJLDurDmz5US6xls3G1xjs80N+8pAe928Ubw
VCIRt3xOis/F6OXy7RMVBhhHF723pChXLiyEhyqCuSFwM6VL5+jS7i6hpID4EyRsZ5Kyb6ToQgii
ScsYzvB44KMrWydfSGK7PESiXu4zpHD8bBTYAljdOEbnY+81KEbkUC5Vb1AHeU8BosceWC0r3Mjh
yUTPoYP0lywka4mkOZ3stof7otOvSX4VfbpVbixEwUjloTpKDcOUgboM1m/PmdhWtk/+Kij7G2YX
QY5E0b2MabxdjUISEpkKuZC8V/8PmvmsatGckWaDmrpWI1CsKVbxEbiKCkCHkblKWxc8c9LoUrxR
qfybPB14lytYTdxuxdrwXzfmBRNRf1fQNhwoz+r58KwSGCSEILr8MleQA0A+DhsJCRT1/g4BJj2B
6zDYFGXGnLxzl7P/gRthqbpJdSZYptIzLzcumcIk94RDC7FXG/KwcqN7Wwbt9INhDfwe9+/Ua657
rZpGwCYY5ERR+R22Vl4FVTz2+fIsLeERxoGIEgxQb4MLVagK6pTeJx1CfKXxXvzjQa+ML1DWNJlg
oWTTBbUP2MeletdCIFrDMVLHCzH1AB4WoI0U142q4HE+fxFNIaucdih3tT7opkw53pLJTL0G2JI6
+RK0mJgmf7MnMX4p0aEii0yRNoOJSi+N6Tl2agI90EacbLaP1Ums0VojuhQr2VAVg2cFfuVFsLUD
06BwsSZ3vqysvG6kfRIv48JGPcYLuilM1X7ARWrQqEDAiI+q2DvG269CbHnMcF5yj0nkB2Qx9lbf
sn6guQnQWqk6p2RCm4kcr4ztByeDp6oYuJnFE2Z8mx9xYyPMiD6y4yBv9pWwIpL0ZOZoNh/fvR7V
kFit9jf6dONS9zu1nfsiN1kzf7pVjoisxE0c322pPTJmMOc+4A2itqCK9AZyDlt1hfc5+Qaunx5j
nyCToW2PFXntcPjT1NRJ7GHXYz9k9lNGjp7/E6u1ufdCDQaxD6lujzB/B8dIHBX6wbjaDLKa5Nla
6K1sgjIU1dtyMWnMyLOZDROOZVW2XsYgVvulLTi8H3FrNqKNTWtf4s4o8obq5rkbVuQNx6QsbuMD
1RHG/tDuVNinReM6i7BDAsoYQgjeoilDI8r/RfUT2mYZNkan8VPokhJ2/d6O+ZIMpV+FAdW4a1R7
fZKvGocQAWMN887QihoMmhf6+Afgb98S4yCLF8CD4GPwDmq78hmtFe5k3RwTopfEuCWxz0uR9wut
AT1tlzfnZyKEurGMLnDj065KsNFJ8DzalQRAUfvNQyCzDQDCw6GXNsEAyHlNS9k2+yY9LuluBJ/9
TMqscYrKCVPrEuoupy6XcLoiXkae4irFIfFeUley2FBN+vcpQ7qn1ZiT9Cdi+b7tjY+hTDUkybp2
YlAxqg0c+ogrUA1zWndHFktDKwJvpajLWizAMSEliUctOVqjfZhvUvC8Lh77Wq0fQyklEzth7AnH
XyizNskxVY1b+TVmI9Eg0H2Ki0pjLNBjLJQmevVnHYxQYWzmo7MIh8Ndvwpt1ZSZt6A8tu8QGPT0
am+nn3GZwgfy7E+abUMZGVosZHqlf9y6sBQLmqHFamOJjvU0HcD0M9PBQqT3EuXCLIdy6Xpi87L5
sNWelLWXCsuJLiip8+mBNAOC3HW9WV12sEvpY/WgmDCC4ada+8xZmEcW3yCNJD2/udD8W8GVFS1C
Y0bkw/5A/ILnh+Ya12DCR0JiP9euBdui/KPGTqx6XdoXHqCwBVH6CnBQcZsryhcQaqLEkVxzKhz1
TwL9fnsrf8NMITKz1USlQuSew+D+LknPhFdQnzhD3DbYA0P6xJoMZPx+TFB0as9clQsvRwiPN/Oq
9OKA9U2bJerxRBxJCg937PVt0tgSzlr+haLwj6N/bUBGGyhqS4uGPCJx+nNxWxtsnLmWxJZVQD2u
vFV05B3sJjdzRZcmQB67Sa5cm/qptzd3vmtrGv06xC5SydEyU9bKeX77JklO1NBPuT4J1Q+4cKs2
scoYncJamlQUstx3YkwkkCkiyOx6dCZi7+AKWboy3JV/6UA9r9N5Aj+WkZAlFUADi4+IsY63OLjz
T2urSGTZV2jVLs8I7il5M4GRYxUg0bblAn+j+q5Tal8DagCR9t44OqEZ7qhhjjB3L6jen2qGB1OE
EaEL1RVhDC9VoX14B+Th/phm/nuWgpbsVZqGcjjuzYbkZalGCUX7eTBK66LAPGDoo+4T1S4Es56C
J78P8r/glQLYg4IeAXyf+ubs1p6sWKWhXwYF69w7v5u8ZvH50+3Lx7Y1DiWzSUYr2iJ+HZjJybHS
uF67TSH1iNZ8RwBWATlRHbyTrQkzJRSkPtZkpMnzvD8yXsV695XSpiqp6Vu5hnHyFaNW36oQzTj9
XIC2r4wnH1xgvJYLysueSLu1ghm8+MrkPcFrusMOGt72GvSSjA5xYxvTundzXN7hkuly17Y4a3PC
M5vxMofyPPmGAgAmD2stYUSlbD/XAKQZo3YyI8p9S6bjxj10HmPUlicZGSfyKqX0yhczMWJq0P+v
p8BqTHePe0/6KXBL6zUbOQ071l/CZKtMgQ+1u9Tum7DQGPp/6oCsPrLyZCkbdMNIyfjq7LP4jOZN
DnjjaWeSAlnNc9s/gCXoTB49sIfZBhRVidLI3JSvR8aMCUyiaLmBdo93P/Pcr0peeQwe855vHKsf
3LfQzv0GQYAbG+114cqE6XCFZFzOE8MsKNN8jbNuQ3uKu9PJcRB/cXEjnlHjGHeLPS9zEsLtTQ9P
qTVrckiNKIvlPnOG3SJ2WFk31jlKe52WGgKMU4jZKwwmn85apFMj+yAol9nrsthT5CVyRL3ffcRm
RnTalzJMRq2/2CsauPi+f9LbQ8LVaHoV2EYk4VJzYXm4ij3pJVnAe5Z7oshUA91q/jEU7f0u5MAV
X5mKN1DaHU3u6RjkskmLcPbsDSGx0m+jVEvh+JLKFsDI8oqQS3HNCGJuSIlIkgnA1sa831uSLTcS
QTiinbEwBj9ONRnauZ0l/dP+nBXXhsNBD17hb9KSKf04uPgsPVmF1fi03EeKz+N3McD+9kr2PTXS
P/zORu6sxLpRG4kKBCP8ijtzgAM0Q9PjlT6piEXg3vwsV5iWyKDg9Gydn0bTAfZ2xg9sQk6O5Cwg
WeSRLbL2yR2ReaRryI16i1Q1VTRXe1FDn2wEVZUoWJfbcYE0IO0W5PPkHdOJbv2gVZiRHDuzExlA
uFQQpbFRXNfpUezHiOSVzi3AZEstKw/ev88WuaBVw/SJV0PXZCY6CVBma3Z7TAtxER8ct+Iylkx3
m0f3jqu+8WGOT705Lujv2yBHCq5VRBcU31zGoAb3NfydiUzBAUrgTRNUT0FTJ7WmSdDowMmhapJe
b06UY9Tb9aBMrKZw1lAAUUXa62Ki9MgnAbj0+VGhQPgflO9HhDqV9pMiTiS+hoGPAxvOgG9hqckP
4MUHVldSNpPjsdf79NjDguZuYiq7JYVYWXNE3DbERyFPTvkNG1ZCuK/PsAnUyhdIwOHqR9/iAqND
Ks6+QBehOYiN2vDCR0EpI3jq59V8bOHivIelCOV582lIpJfAuzJvS9WMkCvPj93JamGOc/j42LQk
RcJ9oERIBgOnQl6u6ft09xs2lDA/liAFdbWc1AoE86MaKR8palvTh0ijux9RqHwfVpIS+h82C+t9
rNsYqrtfZl0mTVTKYDEff7eosOVwXN9IaYkxV01Ey3SfPYzWgUMAKdeUQseTewRmoCyJoAB1+jcf
JTfWbLD/1Eq9LTOwcVTNcQSzRIQ2/jnuhuQxU6O4n4FPgUnXqTGjFWCj+NkBwz953c+wXAKwgP9U
pQAFscXg2ZG6Ve7B+vmhCkl+EN9aZ4CCq08d5H8jmWq2Q3wGzcEBLN+i+59lBZ8eTydCSVHqaJk7
KTBYQdN1DxucI1VuqjK38nQELIAsOq43XxfZOwGIJ8nYj6RJJ9WEo9fXg53SIcvUPlrVxQxqedNs
CsH2RI4+snEO0wABu8dgD6HieJI2ZPwfgjQknmd/rB3rFbpsktxR45YmIuf1x839wWszN6CEXtE+
7bxM7OCfhdZq0nPm8H5Sf43wIAqvtfhC4T5FKkBST5g8zRPvdvvfJH0tFE1EjVuHFayLc9HnIxsh
24gP/w3vDY5yIdnGlzoLoTm3jYB04YXOWQKJf6h0OomSwHCj+3LbSPwImM8EW92FZiVa4exnAF49
QYmeETtJROtomUlHjKhPGh6JN3YULX8C4vz4p6BjGpnUbbt31Ito5zknhtUngwmGOhY7quBMCXvh
AMMyRG/m56L5rglakE1trODVK11jQ8aF+XCDCiYT+rjHAFr6teUc/kS+gagNRBl2K7F8TuDdeFgH
PmpYpQkYFJJ4tdz3we80lKlNG0y3XJCUZDNh0VX0UHe5p8IP/a9dmkPXORLjb8WyvnNxR9/8B0EY
O+0GHujQ6jcqk1UzItTtbF24uFCdozbpOfbMtonVrtCbLMFpZZpt4U7JG4yjOD3JL6Izx0vhc2jS
17B0MrHTCpRSem9yBw0t31yshEOW4J82C8C/waPQMlWCxGBUN/lDjrFDS7lYzvZ/lg6hWaZU3ehp
IebxFSWYVU10qjEpmFtz0rsrOUIgsnhHFFBcblPzNiftGQh1wTPaNrGqTTHmkFPDTP/dQKDGD9et
joppHJ83raQM1QN/bKKA2OQJ16eww+V3+wTkhpr+Z5wMDF2K5PuoqJpJfJFHyW9K7F4XRTx4rlEB
MzLgT7qNJ6K3IdptbSiJO6UYxz9eqOO1Bsyf2RxOjVSOWk//J0Nd31MIlRkSoecHPq6Mrwt1o0x2
lDpKCxlWun8zeTSXpgGLdJBLv1jCLmrsQZ0HqaU2KXtedIA8qtF99UIYAaHIz8B5I/vSVHmGW/Ae
GZeH2ajeNDMIdUGEiMr+rbP6LY9a47uaf/LiIZh/eHjRjIbsbqIYtrb29MwcYDD6ur+wOyuwFjFS
h/qnWwvwfxTmtoU2e5tBA6o/JejUkKClI9kzoRqwL0jWpQVVhvV4uN1ZCC9+H+7xcXdlx0he0JeT
COqz1Cs0GGboSXjtixv8L0FL99RR0guvj2v919nM7xJGxBZPLdizaWhqnzu2XNd3TnmKaQPvAtdb
UXlVMqJ5CaMwmQYcvoSUaC8sXaCGwBJI9TwXqVGyY+QLZbeHzxw/mgKwasFxtzwSfv4/EaylIi2b
NuMLLx8H2hXkzmRzZr9LEbuJN/LXxO7rSMob9Tvd5Kikqup2O0GPjKosVx9LQT5prpCh7GhZ+rmv
lu7x9ipMpHe34hCW9I005VmK0Uft6t8gHBTH8dLHUactEmn8x02thXNysExCkCTXDPlZ/TSSEHeQ
80Tl4Ht4JvLAjizLF9dY0WkOqayMKV2aC3/oGjT8xsk1OXWhJbcV/8e2/FOBinbTPs5vl9HG/BjX
ddif5OkrHNm7UiI/asaUKj06IRs4+3IEX97ExV/3DJTeSDAHV9pRZ4ToT94hTg8PavOV954TwvGR
qTGJQIElS5hgysHnHf+Gm6Ovs3ZmXbI+pqWPc0no3AQXUDvOmX/6B9nZgrl3PMpdPcMeFVX2u+rS
F0eFkPq5V6Euay071u+hxkxZYFf8OdkuEsAFXPMF+TF7e8UjOFwqSSC+3t5Ke5j2dpy6frS9GplG
suk8hczKy668Re55rw2kDt8JOUdSeG87P8Er/VgSW3TjYFeBtUK27mwAEmFd05RwAjTB/UGt1rcP
JR2VPpHijDfgzrrBN1ehDSNQxrp4+zUQtCo558Q/XkSq1RdRzLYgMEzWnoO2DVxB2oBPcb7prLzo
rFoIRulv5udZdr6o8NphhUi28fTVc3cZ/0G1Pdc76JP1Df72fJfak9gC1uM1I27S7KG/iAA679mw
MkMCYQORuDTfhbRFEQkf13r1M81fnXrkK6JKFq8sXWsM+dzCo3obed8HwZStyfrufL8RkzxoYMa5
yGc7FQmOm8BHt8TdfwcxsveuerUK5iQ7Zt4b1K0aNElQcCNF5Q3tfLThcyqm/HcNW4F/cxvksPcK
y65IVvGmHTSfNFX7PDmJrDpyKkUXG/v76PHo5gQRBqOvv/x+7dvuUf5SVzfsv/+ijuxORGZmLZLj
ld8W67g9XFet9gXMfiWUqze6KMo1cajlgn1mtVULxiprJ9R3nQWbr/8Yh8LrTDEHZdJeAVT+3Vk9
ZZOXM18xCTcIHrSVy0eZ+MnZoFx+GPxAfoCyYK53rJpWO7UtjQjh4E2k9uAlBmRtKCqB4PsydUZN
IdI0tDmd4T907bf8gNhzJcO3Ooub+MYe55zSc0ObnhSjqkbxS+2Lt1qniKTuVioHtn/MgS3gCvYV
vEKxAwcQ31B0CFk+4rjJpUGuGK6AxpeJt6NPwELaOkJ9T5/R5WNVtDtZan8nKEXo0B8IV2uUWfUC
nU6vG/2EBZ+uPvYFHRgutwNvAESFhuu4kUXnp5u+gCm1KIz9DBkoxwWsr+RLyfTqDw614Uo7UYGC
BubdOEHNvWXxjLndS89weZfLQgoqyWGAd6Jixp0Xsjm6F6NIvQyhRH+Oqz3ZcnXWjFawf56bsDRD
ORhhhYMGdhPIjdQgUexcEzZg7+xAe4iYbXBD+jmpe1oVY2xYxAw46/nj0YThBiFftL9ny2TAEcf2
fi4OAKgDHI8cZavfxSfkphGAjRTHL9HTRPzGOTDs5qFAHhEh3V+pLRBNkJ7xNskgY18+EGCjObaE
Hg7G2A9jKztslw7XvSV/7NtpzbfAFD7ZI2qXHunOlvEx2Kesx/ZWjGVTGK73UDjEvubAc0qys+/Y
zi5u+38F1Rbeanzbo634A2vWlQSXAq01b26F8TlWU8JkzXoCGjiRYrrGeTHLbCbhUS8KIreF1MNc
zCl4Egn4TVoPhACsgFdax1scbR0oZE2wzf/3bkolqKFGvll6QaUuWxDLyc9Au8l1XYWnCg4Kq39I
OqjATdxPhH3wi1abW66woddlPVyfk1d3PIOvOMQGyFJA9zNlcV3j9eaCeMU/JOGAp5Xne/7dgvUm
bg7hSlLFZ8rTwj4UpZxdR/z4XsCTbYUQR1P4ERZxb66cgLNzZPxD7ZZwQGWiV8bQ6F+ELAARfLVI
/W/p0IVt602kgEpj9gB6+niEJf/2n0J4lBMR5uppN0OpTZaqE3UFjHa+Z4DQQQG0f61yXVW1HTY3
0k7wFsHGcRFCYJScDcEButNPZo7RRzFwim84YOWScP5Udzmkoc2eIod0gpV69eoBGv9C4P6RPn9z
Ows8+B9mrdW3LPqCF9fuCWyxcMb8eFa2a+uvYBGSCodZouHHVssNKysVpLRycw3k8mWGtbrjzl5k
bcYBCTWh/mrqMWgfWRUdTtv5hpR49lGIKqyN4ZBBBOEKD6EP2dIh5sYQoMmtI+9xHD1pjTwLY5mT
J63okgd38bUxGXnZtP59mtj4QkmyIUjMGr90kroURnsgu4l1iCotFqufxsfswE5vu2eqZi30Ny4y
zM57yzeJhK3vET9IBi0moFb1XAzVKL9ar+dSKhU18id5+uqDKTYHQjuj+fI1x7t9/ll3u+V/Pg/n
MTlhdcjmVO4mYDf7bfrpyXfDqVp72Y/IKwsmPiAE/gcvl45ZfhYoWfh79GiwhbvTXzmB5d4AV3Us
o6HB4huFclJJ6x30Q0LC3T4P2dPZiR2Ur9nbJo3/TTyxStahZr8q8fl6Ecw53GqgrcsEOE+pvBID
pxkniOiDoBD439sEsQnT2Le4n1PpYFdiAX99Nw38Hx8syQTQKaAqRnUKZbsfe0GVp28I7JG1v56z
W6RAkKeituphITOiKzXfsrgbHdZBh6ed/rWoqW2vM/SJ4tXRJUWo3aUVcTRfwYxwZt2ni3+QM53v
cHJI13aJpG1IQ4Li6FfUp6SNLiNAQCv1nJ/u47bLWRsvNffHsnAYxAxFO2+rCTOuNKUxZi5zDQmS
R0KVWgACJ01E69xe4EwxfL27t2rfFeVQ6hbtoezKePEiRSH2pT3WCnbmUXP7lJLXvToPuV9ChaXi
mHEVL7sCyAvd4AliRdf7JCSaNuovEredzjJM89/iU26aYWJ1L0Z01KydRYecpmGX39eWxUe4C2AG
q3D9Vr0MQiDZaWRzy8CfUEeUPcRUxXXLVxbzhxpA/qCYcqcpAbcpkPo26D1CbbRD2Icikf+SI2qX
tJa47ebxCSLn7bLnYcMvMO90Tv47uCfrXVFaCZZVLjKvjMPdwyTg0ybFikMBa6Z29CdxLm1l+Dnj
EJ1wbHsBSkQZsQZtfZiYHaCDA1xG/lwJ1kucmr1vVpi6hwnVkG7BvCfvCRKZYjTI6esXqzMHwwnA
PCk7MJ/5FT7bLz6Bs4wXVmlcx7sbrqVDlGQwiEZuGynhRjQ6ihCHxfkmoBBpPo4sUUFJif3xz4hS
Tg7AbUtJCZIHxTEzfmAQ2q+yDqKRVU465P+dsiknJroWGFJgMXFUimfSd87LTmGgwHIZtCVPU/GD
Q1zsOQOEAiWartOLySaylFoQ30iGpIJWHbHbITlHHqpHaSdcmqQHC3gWCJ7tv+DQBVD6Qq6TD71e
JWi5H+XKst2aJu6djYcwhWTIZvHZZjjMBP41vcIXD9W0WAAyTvG3tMzh4hpJmGgNdsRe7AKlRgD0
JQwOoyoK+648ts6MKD5gfC9DLttTBzCVXnKsxqBLfN0kAzgXZYNE5yO9bay0yW7dbmKfSTSffCEq
xoK1ce3bIChKB2MqvWjhC9vUyHTtRCWjnf8Ul7/lhVfWqoSN73aOjFgg+rYLKA0pFnZ19xkRxaQN
iryDONudhW84oxMrNnKAw1ZK5Dw2LcZTM2i/0frF1WTXY00Sx/J16EVlltR/D2/P7OaAJol0CWSx
bRhFtK7KYfUOCnkYldegn1wMsoFs28SMUg4CX1rPH2ycz/QKnBH3OdWSK/QSzSwLHSun6ZPg6GAp
NijpbYFCSgJKxWnaGsVoYGJe4L7L8rF8/Ww4rmyDrqWYoxQuR9ywYNZhLEb9ooM67m7TqGCbLUw+
CLDfnGY4tJfo6lSJJaycee8pD8KGdhRXwUPoqHCvJd1Ki8NIOv+rBZ4YXjG8mDx1W7iNPBS9lR6c
QGGchkum7A9phmEKOSuVHLfEPIDhsLmXIfT0cBvVBuKN80B1GdI/CENW9UxuSvZwEsQIua1Z2QWy
aa60NMgazecPZy8CYjkYZWxfdvOPQG1vZUuKLrbVULic1klufTmEa32Wlh4LBwI0cW+G/Gj4pCoj
SXyyr0/rAXLEN//4INheDiD9Z7+45BVLjdc24cFOIyEZFxYFu2vTQ9iyO9Ovx7n9ITVKujjedz/k
c1V4FwIha2p/bBJfoqj3cB0EZBDRekVWTdiDP+CGs2PP7X2XvqhayEkkZBYlrgsMf0H916fBtxm+
cZam3HlIOo0rv1L1B+YkNozJFlYkADlUhF5VHgvTjWAYp8KSQwO6gjByqc5lWERWQCVGzXnJ2N+T
5lniyh0ZWSkoCdoXlTeF+3H20taJVClS4J0oupRa3ulaxnCi/YrxjElsGJ8OvbHebwn5Eh7zqBXY
lZde8NDByTA3bKW3MgtkKwGuljnqLoCLE34bG9tvmtHEmETqSOrO08vshOFuinAEoxI7PoXK7DQJ
MC8pWJ9BDghMdwkF0jBsxlgXdT6B8OQaaNzhVRaO1Odsm9wvydId/KHNc70lXXOdYATbbLZzqHFz
Vqu9l4pBvDF0QDs4y5wZ5okfc4LM1SP2BiUWsR48Qzy7hRu9FgL5iudeWJd3HTyrLra2CCxSbhIu
+EPwA2xuTeswnsjCePsKk1aa385TjNQalFTncofXUT7+lIGPVsXymlRhMXQl66hu8JVm9g3vZa6W
O6SZpML0kF3Aerk2bzbEWPYDVfRt7OGedga8Cz8iRwwSXl6OZL/oXz8QAjFilVRi1kjo4AGcbnQQ
0NyiYFH5DyFcZR5ja4YRXq/lMF6PT/EfZFCouJdm8c0H7Ay5ATzXxNIVTsQZBVxYfpAtLCqq+pty
98gqpyDI3m3Oo6g7kMhbzUdm5xyGRAiGov2uO/7FUV2f/i+qcK/aDIQ1PvphSrJKJpQleFXo8JFE
tcVSKueJbBSVxQ6FJntci7N1cGZLeIVED2aspA6uIB4O8/EsXXenlAZ9H/3wmCZ5Odyg52ghXu84
YorJ7snZoA52vXClICoQoDHljj/z3ig1zIWof7SUQin7Ak+EXxaT3+FZ9mA/1tFb7P+VNHgzf8dl
5au+5oMHDgOE8uM31SLPwtOX1B4BPnoPQ0GN7KgAwHRzPvYSPVVpUqpwGyIyznOgTzWTMoRIbGd7
qtR5EIaqYrQV7UWRTvEOui+D3/SRWr32JhVUiVbKz/4tTd09ohzoWAUWILcIs2USu7o45AnFM79R
DhLZUGSdbg7ttioVWiz6L7m7vK2hi6Sh0dL3h3tDrwL0pgJAjB8C5tc9YL0N4DBdp3ITi9ACweBs
3UMu92vy3JdeX5g2/zFlczQzTrGRODO1/VwOn2qfTBK4kCt+5a5cG0Q8teIiE++neLhCM03WlY1h
kgwBt4thQR4p5Gr0SlsqUsnvxoi2yRDDi9HrSpwyes9K70EIUb8ErR/6mChiuVp03QpYGA2+BXnY
mssxS3pYvHg8s0Cz3lUgGMDRIfVrk86T4uSQ5VH6rP/m+m5WmKfQ+eg8ZruBELh8zqYfbjIFDcXz
oWzKyaGm2quC5Xs/m0XbZGBXR7Y9e3dcV0elt/51GRj0iUFayyZcp5yes39dSeo+g4CMwZbqnTUJ
Af04rglawaPngY66nyoqm553gsfdKgEibLIk9KO8xWsKWMVHrFKtAqkCTD9ikG8PZd5FjGZZTg1e
IKKERZEstb3qa1hrQ9jitakA5SsMRvNhS/6mP6lhT6XQvPjO/XzRWAFJ8uY5jcrGw9JgWsh7xJmz
+YNsaWJ7yqi2GAd4+CVpWOPK3P8KBUEqTRUsEbSXth3EE1BfCaI4HtLw9d1lcdxIjVRkAtfmFWnO
DkSXv/RqCc5Zv8VZBWG7FojrVoOsbstnLY4L85FfvMVRA6b6vkd8xcRyUVf9KF5W4G86bTBgNkv8
XZJjYI+w8s1yHK5pCXC6Laqx28/Q8aOVD6Jtxt60m9tbjtnvmW76jxshPybOtM2/0RqYt5e3EddI
BRWoVAjYeOjbZJtmq0m6F1yAD1hv39DCPq1fiJGZANHu3tfjNGpLmifVZLLineugkUHF4+V8rur5
uaaDYrjgY4ow3WfqQOIBi7qq/c4Cc2PkmT+VMBsvCufETebxQ0OMwb5ZwDSHAvAQIrCUETrVMfrj
ycu8PfUvZrwyhQ3xQg8SZp6s5fy8CpnvrlridxxL7tjiXXu8gKFC/QgoiecEI9uiscLaGwcnhry/
MXL1nFGHgH7e6gmnnwst3/cp1oRJ75KWxjmevR1HfcaW8ec+b0JVlt8Cf3jUK9sInWKizcIt21yU
iuxuJoqqqQLBHr3SvtwpUiC+CGf2Mb1aOVvO+x7OR+EEfhWFwuUj5BZ5y+LIzsyAEQly8dMigd+u
bl9VqEyiqBASDQUEeW/CxcEU9Kx0M851FvgOzWrqZIpPJ3AeUcIXsUN7vVH4coE8AoPbRw1+W62j
iFM6KJUp3tmPJpvJeTzRP4Yy9W1aHePLfcTLJhbOlx+dFpo4Sd+DKItf31EbS2xEPGll6TDFQUFw
DS8dTxIazyp2cg8uvzD9kLfF7CV47wGJ44fFj4+qdBkVy4HQVKeU6sFjOC9Tjx3IRVhOcR0g3261
vS0HkS+A3cFJfHJIDJ7OA/WNERFSYB28cL4G2r7aAMKmBf/V2+mNph36qUb9NgWgk+8vliZsvd66
Rvt3DJSKPf7E0yRpVracviWORixG8vN7NQIB485vNdE51xlTRHRTpW3L3jG7LM2YOLQGCNlbmN7F
vaSYWslOhm3gamxkqiLNN+tAzyd1FiBxtFu5AgDA++p6IkaiurQx7J1Om8AvbfRMImhGBwKaAUa/
o3BncQBjkYGuV0/xtxuGYZMIsrVdSMp+vNRkX8CktcotJsN+X+rezRuOsjxHYEEjhmLW0sXI3tW8
kbpYwliku4eC97uxXBhcUGFbLHAg19+MjY6vlWgeF++tziziHlaSl0vug/U/eNLmYEkLC2WDoqaU
6nnr5jO941yhBggq0IG47+FRP3x6AmGW5WfBiiXEkg9efY/p2njb0aSCZZBCOlKYdD0m5jc9DDiu
b6WmqYDJk12Jc0j2
`pragma protect end_protected
