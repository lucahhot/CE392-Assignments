// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
LXilXZKgROHcx2DsfxqEXc8gIbqHiBKBPqxtD5CKlJn5w1Is1R1TeGqJ2ORGTUPhArKkX7RNDbSq
Htznh3nmw3jP/pIJa/+15s6rTl1pOd2nuro8Om3/3IF5Osww0Pwzs1dlL/Y5EJ/JAz6km/yL/Haw
4pfeQE6Cn4nT+TKz6I5Oyv5sNhGKFYi/TCKoyzLhlFEE7+8hH0WiW/FcE3sQVHM7ePacag7YNs6j
wl/o5BXg1UBwRDEKRNkvsKqpidJACqLbsG2g5OWgnoLRTu/7x/aWwVbY9FIk6L6uLsDsgeujA81f
mO5153UHnLRrcumb6oHRv9CNi9hVYeEFm7aYKw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 25232)
UTBWPzWekxGuvNHZCBZlNFrjFnMcdQ57hJdyf8Cs9pkKpXQ0rPX87GWQlZ3cyKUjLusItvnmcX+G
xwBJoD75bM6m756XMHjEuAUXY8Qa1CB1r2Mh7backglihCpJLeN1Uh8F8KVrfHo+tygugbCj52SR
nlI1g5GIXXwqSR/piyJoSG3OWnPW2GtME64cuTE7i8gJ5b1uw2NFVcJp4OYiqqARSTsHGZSewSf/
ROifjVeG1skZDKlCJtNGrjTqmFNqrWWrlePnNYTzp/nGzYYqJTOkcosYXaZle0okMFjcG1XqqtRf
UcmAJ/6wbUoU+sMUKEWY5ftGD6lMgRW487VeSHHfnNunyXO09KJKk1RasGtV74ipr/ynH/qp1kyx
NgchFaiIZXF7eLyyfi17riJLZfaej7O/4BUgPjqgFWYZYDI0n1/Nt4taGHvR/KykzhYSH8+3cBab
MOr0u+K/my193eeGcN/UkPKu5Yjx+GGc3Vd4gqGGdiWGKF84cNAG7Mxw4hHONsYcsuoSQRumU0yg
K81xCi73CGIZV8AkGxEYBwH5WXKkIE5NXVRvGxnRtv87g+GoiARpt4Tn7wSG57OBP0CucFjxxTR6
lHvRciAUDoubhK1tpWOCGU2qOvPGqm+JQp2Yw+mx4mT1om5IxQY3pAILkkB8QDFnd7FeI5+axyIS
rslDd47pF9rbAybqEzW20skUT4zorZ8K9iFCwXfwSPnXRfD5E+5zkUAyQ60mqRjx+88PlqrKAGzG
Ypv51KdkPgc6A/aiXW/lVSFDQk1Ofrb8UI0iy08jiS1M9p2oeklX5m0gXE+XqHFzXheZf8nWwZR/
alm7e36t6JDUXwLPA6p72e8fqY8Wpo1jmX6zAL/g40yjSySPn/ET01g9Nxir8Ji5WvqSV4NenmB7
o5Q1j9sBYEAQHgGuJUkw2AzLf72/BTwISQXgJrQpGI0NUkKYXIohKGV4WzZsq/TWsJ7+2CpyMdux
Kq2uQuI/w3b8wIftovOZt0kzx/Whi1wtOks17cSyeh93MWVboaWzYqpEd5AtfFNnfCKObaHl8xKk
9jfZX94Mek4T/SO+V0JvbJTMJgpvF3mEXNSkcuRrFudPeMvCsk7eOVVosvI7fM2eGhSaruH93YUZ
f9y792yW8zI/v1zy//IRaK9imTG0T5AMotwo/0695/twZQnLuJxV1As4cSzVXZLN6Y7foLj0saHN
eSth7ZX/34/6fhL3TXwkZB1yv+iBRX8jZUQROpt/WGjSEAUj6guQWWXxN50byPPS/wDi93fK15SU
Dy9atIMbqo2ZIJlC/DHRv+08uVVMoC94FF/vqMAsadYWab2MQIwYFTHCoEFlhgMMaCdsBKTrfc+C
vD4Llr34yNrRascx/9BiOrFEg7KLpzat4UTNtM8MTJRikKJmOerxo1Qbq9gc1+dR3pMYYObNIbV0
8BqQGLyouNhK9WhpmF4wOj/CbS1WwU131AJLgyfRi9qxOJY8xktc3V4QHZv2tLwaadHNK4I76/eo
4JoKmzSpDvaX+ekHwvV8qBcDR8q6zSMSAyoPrabVE6JoZ6xuJzo/qXlOQv0wPuLVywg64jXakhP7
24R04lwWalCn5e2BGQiIDMwju+8gFVHfisX4VcfwQVFtIc0uYEkYNQ/lgSUAj2q42+P2txWvy0sd
fvwpqgvjcG1TgCkSyQXLoPTlPzFDVAP4gBrB+mOw6xNDXuhSjWtTrz+ucXSh+mkLkvdfU4I6/YOL
VkWsrHSj26XBBC9d7cpU4bS88qyZ0SvROfqy/KCo3+nmxWEfdH9gY5aHqFwPeexcPMitM7w4R3zg
Md4jGGB/OCXajp6Gglyzpjx7tjliTCglt4ve1GFW0nxs/N5zio87iPd0PvqweoAuBGLC3RN5fd9o
GgMED0du6Hed0C7aSHLCncIvcltaAFI/h368Xhwh+XTtgXIcFfd3fFCHRPivVEkF8rf1eSItgXsY
/W/rDwIHMUZ3JM5V3qCd9PifnEs5e5TDLqzsg0pNcEnK+2ZMJTgfoquWt44JVVJvhUWmGSkOLC/z
ROsNZR1FgesZ6xbnZhh8WGjPYCPubIXsg1ZXgXcpm16sRtdvINVsh8PDt6SuJlKw11BnjAxp172Q
lgkwVemO6YcVhwYcl6AwVOouyVQTcmigFufKIhBmr8KDOElk3YukKYhuO+ha/qP5UsJE7cW6vAKq
F2XVfKoF6x3B1imdc3WqDZ2iHcEA4v152zVuVVyCM/dgftzjq1+Es+njDmBNezo1jzhUtHAtq34f
vSmYcCBDeJJg2qRnXIkMiw5dkS/vlH3BoznHiKOJOGnWquOGF/P3Q2Z8PMxP1IvuVkzkmIzvGbA1
C2Wypwf1jlQicLZLPljjHNVwCI8jvOh2KG/vKyD5N9Vz0FIcHt+IPopYKPOW+Dqs+GRmlRu6Z0ut
f7TPuI+/lakEPFVj21KtXHMF92VuJy8CozdpMMS2KcFTmkUuw0VR6IB/Lpnnv1CiXD85hKzSu5Tj
PFvOUvBrkuJ6FM3g5qdWjwFY1QBszNH8Nk54s3E7R8fvcRCWdc439+WGiPgw3qKFuVrHK+bF1fZq
4Dp2blP4N70rw5Ytde0XAsQ6AOiqfRWtizzq8z5sbktREAFdEeRUIQP3nFwrVqcxfBPJQI3E5uts
j8hpRlAjXLT2vPTh9EHh+4U6Ys/QTzCAMn3lkTAUl3dqGLSLj4INxx0N92jiGZXikRX34flyVS3t
kj5qKrFHhyq3+CpXEiGJiNmfZjTkT+T2Zu9GXxEuNBFVh4Lko6OCsYyBO3eNO3A/DoaYg2BMUKcI
8X8kyZMKFXJXYIi8jidS+gk84rIdqIVaY2V2lQmkQUmWrxZK6KtKzk+B/6pu5/hvGFIS5HYZmKJ8
2IHM3Aq7dFPc5p7Y3dgGHnGmimKeWeuSlQ8mPHOoUciz8IZ7WcHr7FOvlTAP0XZ3CuxWEwVMt+qx
Spt3lLIk5jhXbEsHepD/2DQ5QAY0gLhXR/Fr0AMPM+JgKecbQ9L7lHkelIvLNmDkq8l9HqbpQlhy
U1qAynbWAg0KAtamF3Gt5YsvbQ+PPzU81QQYUO/ZcsHtGjJfPNQvCUD/7MRaWl/JTLxjq8BhTvGW
2MoPwlTnq3uSIqk0X5K0LvMstU65aFW04vL8EyCZnF3TgbKCx0JNTHbkaHKNLowO2976w6YyxBHD
N5v9jWvj3xhR0big1xemxDcV97kbB8RnyVNjikaUmEsOkCj7Ldy9SNNKjwDRqkSynkpimS+k8h+V
KgZ9Dj8j6SFI9EL0KDTbDrKQUj2VO49JpmI5YOCdW4v41SbluWIO9U5loS8SUEXAD33S4HT1OnRE
REYXrjU2lP1MmGSdNUSjmMoXXOzQND4R+SlIeXaQtS3HLG8nSFSUqJBSGa04VDp6tibpRNCkfYMv
wF1cYaV22fdWpUZxfodI5Dzs3pwr+1HU500qP8lPYcmgID+EAJA2Gz4k5oQU+61co3Hpp80Z5T9k
b4AxcB/U9Gh9H8en7QxbUdgBinUNebpo2H4G/+IenxrEpZS8bT/Dcc1E+KDhJsZxI2RqIt0yTEkZ
fgI62vJfulbbOiXa5qhIi0i53VmnbXXyUnWnqN9bj2pAkU093P2UPkDZJGwKsPMOrMS/6Yb7U4S1
amXPFW7OMZzLh/yCM0DHBLKUKuCxTkRcD2zCLntp8mkyAsvrrH4JnrVywsHP4Km2sq8b3D9JStB5
mQzKc8GW68ihMtXbk3tTNoVMqfy8ysb/m7qt9OU330Tuc5APEGtzczidrnH/yQ9rHwKC+LQZvTzy
oBJU9C/mz0vB+Wa4LIXtnB0I7bc30SPeAWmbHGIQOD3LD7aOgFOoDO8VVJf4QhK8RhmXn067gkv1
/ZyLrTGHgcO2eTbW6CIBa92RSw6WmfMfUANIIPolECKUkOgljfyQ0fFjOHUO2j5n8GsiZ9wrjGvr
Jh62BZ1vSXKk8F1hK0PnG77Kuj+IlUTkX2o5WsOZ4awpZWa8CkXsUS/EE0aB3KdlPzvPUm9ivxDe
c76Bi1cofVvuacLk58XigxwnL28sRZlzBWsD5lJ2gQMvVLOpLP/bweFztjS/nbOBhoxixmJVXeoC
QWHCfj+7CU5cUQAVptoqpaOtNu6cskATZUXUj28q6DXZa0gbXb76BCGkvRv2xnspeIPQpU/bCqul
urC2SkzWJiVcUqrcVx3R0yWTXx6VTHUJMfHH8woSkyV2qNj4sA+JK91lshvT5fQQIgYsh41wIdcy
k5GeqE8nu7Pohz14zffOkpia51X0dwgOg/gRGhg9M0NnQ0No/RdXiCcQxCXH3Ims6yH5v5soolym
KXsf3KtCxwFMF54xvLMW85rRb+wrRy0ROocTJLibgtLJ11WK4oGGUpQieR+PjUJU9f6RxmDOwMeb
ne6ovkOJsIVXJwJCmuUQhWMm9HkUPKHukDyD5IMBQB3MD+Pf6enFKCds6dX3h/ckZE1a97SzzDwQ
yDmX0zn9WyyR+OUfL6qLXm3ZIvs60iO+Gmz3xBYUr3Sqh+Bq3RwrEY+9j7z3Wfi+cNgmUyM+Isxh
xlMO1VeLhv1167g18ettNmLcaBxXp2uyVMfADqDmj8KfppYkhGriiuJRGeWVER2GoS9PDOK0kKb/
XaLv5G5K01Ra9VXY9lFTVdpFhXWPYrZO75H+Vo6lJe77AV9XtyfHlZwDpd2DpxwxISqf8lKui0eV
OmHB17lMAiV0ayY+eROSgC1Vd6T1sQeQHKy6DHivuvYMWTr61GwRaNurbfQ5rK8IGMOb0gNGefwD
UmTMAekDAzFaSjTMiaEHoL7exTi3WCNtYZa+2tAph8UW7oL69K62Z8+X39+GpJ3uz8Rw5N79GrOD
qkY2CWeLyQrMUe5wR0u+Wxg2JtFX+COBdkedebgU+7tu0iay5Jt9v/G+o9C3c9zgPlslevpcU8PW
UnMfppc4zTVWQZ7YNS8jdsz8jVtisxDRFDB8qMlkIcLPuYBH7pj4ia77DA1Qa27nAFrEVqyEc4UV
SoEvJcL7SA1yEFZACE2n7CMS3yuj0l7irFVpb7tVuWqyL5Dfur7XUC/dBF7ss1CGNc/MG4vf3V0K
9kTWTqJsUrCjE7tPd5x+ivCL2Ave7pUdmOhOQS0N734KbjKYG6hq6OGHtw239ROyP3bWSdq5yf1r
Tr0vUnRYEUgpVElf5FUQNhwrBO7cC+UQU5ngJ+wEsV2VCy26/JtvEVl2Nk8oVKuJyE+VnTqKUb6b
g/MkQNNY2TKE+DL35OMxdVMrP6u78N0vRGzM6k3WaZ1qynz9m3c2jqD2wKxF4cAVIr2r5yPLSKSU
Z1W6xed73hGQAgois1I/dyWdv6mJ7e+Twxcs9StHuilTAK+xWKZezxen5WdxemTtQ5WjUjX8BTuo
w0uKoe53Kdx+3FtyAx9G6APEfbp0sUaPMDKhsqSVkDdefCJKaVfYWlrf2Iza2/sYEHsAy6/ogSxt
4gvT22LkMkRr5plj/SYInZlItAdZYpqfaBamP4rxCpljn7zSQikvYzArwUqT5YR3DFJJ9co1e+79
ZOxZQ1h8AiFvI1NrCcPd6VgeCLSpOJYLwaZSOzsoUD1SNpmVBII1VDK/yHDTBfGgXdC6w6UqqJN5
PPX1vhhZl/11wwugyRDHKqB5DK/35nXBAtD5hIWAWMYqlHxsse61P+19YXqjKDL7I40pE5kH87BB
AIbPbtloucN/pz7rpr7dwhKHLH7LHJdJU/n3EsnWV1KBAXKQYA8TcRzneKTNtSIf8GxWDZcg3gRJ
l1mgc8qu8scoJd9/yNbyvbbb2NtxGGoLDlILQGZNSH28WI2ACPcRngr93heTdIJ9wyWFUBSPYrSc
2Dq6Bo7r2G7wEf3qiniA0gn4HO1IYxWg7gIKT1OvI6mAjl16M5LXVY2m6m+01RU+7UoKyWA88AkA
DaEjTodl7A4BvoRjlsS7hRGgQix+p51Fvd7abMOTNtyvTWpowKDr2bApYQjcx5b//+8dChmotl3z
ET62r3HkHTPOsbvSLGXLacIinZxt0Yr7cJWuX0O1Ikosm07ioSfDkF6yfPXPaSvjW9tOmE6bb9Bo
TqTEIS63u+MJYr+pzmQlk54n6eaNv4JC4XulrK4CJeSoub93uY+El3LHlTtfL8TcrhELQ8KxpVxd
gMkU/CjDCkhvhfVl1el8F/tvY4n+ixB0xYxhxpHQYREqHiJMcj+XBOwqbnhnmR6VSj7wqIy3uXrK
jA3qDyhhTKAhIhkTKkc8b+9xJXzbvrwhsCh+pIWLkbUi+pZ7lgLK4JFfGegKtejtV3j+2wIHHdDq
0xdCuOPU8bVJj9U4Skxu5Uyf52t3+2BIRk+ccaFbUxbcM+x4B68vI5s+RKtN2fDR4kr8gCAwlXfK
Ai4UiiJswgzGXvMnj6JyvrRNnElz3T8iKzYdq/rhnQlaC/+I8Nz595UDqYEG1juvFyOme1ExwM8y
7V/wwgEKe165EVnkn8KiR2g9pKtHqueB2NuWtx5/cMoxcv8BWuDvKRaFwBUBvAF86L9MaVjIQjbe
f32Z8vwiMDX4vAvnR7fK2Di6G2cXVUxrRslfMlMsd/EZ2Yq7ojh11tXrKIYslEZHY2+bQNFNDDdf
xWU2lStt/a8RKcDozo20gzOmEQOzwW1kpsbfk+/pfjZNwsgshBk1s8JBvIxpTyZC70wE2+g0o1wx
l6UvnERoZABLfmyVDX4iKUfzBIcLHX4HJgLHmXI43F2E0DyTYpc7+2LLezGqNuhQQUh50w7b2was
R/6SsjzG3JyzL6eKZ7XLIKLHShpSQw+sSn+EOQTP4EFDe/8rh/Byd2E4FEpIZX/PKAcdZ1le9IH4
rUiEJw+t9smO/TX+HLbgyR3uE8yJVIIm3RpFxabHCEyVL7yyUvXNr0UjZJh4ytbkCbuTLchgOMJB
clXH8y4hkubzv3R93ShKHhcHA3Pda+LaLVgCKVaoYRQqO0vbsUYdyPgAffgw1XTlURHk1pw7J+Lw
HHcIgRdysfdPXCvUPFfAoL4UX4mI6KkwNAZv/jqAz1sGoAaTru+pWBmUYFcOE9NlEvZ+e+alG6e4
BzSkgqW3zQZmwob6FzZxPdhj34dT5pZbrCC7oC1u9djzuliVffa5vinsNtHnKzGXCDSDiKqE8FdM
r4iUV+3AgUuqun4PItLo6OglPlIpLdD9cOFVtAhlgX+3kPKFb9NeWZgfYrkYhMxcY97/jbTTM7+m
tBsivObB2xVq1OR680x13Nmc30DOfqhKxsl9ajsREA0mo2lZZbMuhgx28tK3czJTJt+MbnoZiJKz
qXeNWLU9bCJMny1T/nBMLX42PcohEWTb0qi4rvPNeMOwyEr+JxhH8FweKh8iY9m566lV2+K8hQWo
Q4WbVc+P7oaji/8KGQXavg/gLP1S79NJU/eomIolD6W0fYBbU1DCAQL8YZpsOwmMwBFtak1Gw33/
nbac27yVRavwiq4BipCNpIctZAoMm2BewOGtB++l2Hd8iYYcUNrfRk1brteq5ISs1KZA7qWbhjt9
pVCPL6cG15HzfvywAVD0pAMJdKLs3eE4Up1obgSgyBoV7HuTHvbTT8g5izMjLZZYO4lPkw6F4V3m
CXJ1IPlQEUZ4v7SI87w9mPHSDod2B2YbMs0phk4kGegAoY22rZnif6RNYgdf7j5rd7iVw2YIAVAZ
cxMhSUfGds4SHyiTooV3WXHfqRstFdVngfGHRla2htxFozcLaepYYElIyYrqxKX34qMG/TvUOavY
HNSU8u9ZFvvnBvHqC3NHaQiUZWbpMcHOmURafSPhebeqR/3Sby9uFTiAQlgS4UAkf031evBKfczV
3HJCzmFiDffbSSfLD1raDPGUpzWL6RbEfnt56xPT21iSPWR6fso3yz6Ll/KMcjNGX8tQo3nz78mP
6eElgIN8zm0tAX6T98ItmdsP9xJNxEyHgSSdSot2onXIYOJJ6IEKG/POLNWbhetm7P+gnYuVtsx8
RksHTJ7Gs1w5PTLw+PvpZO+vENt5ekA/NTPWnxczLz+rWQGI75V+UuNJkbWAEdwmdmMP8EBIAOsm
/nokQXDyEnlFVtU0hTCLrm8qeazVkSAynMPhaVs0dpq8y8H/bPGtKu347zKt4RHrlbgWLST6hxVj
XgDpYuyKBFc6vnjNbG30nFfB7hnw/hsObinxNwpJmmgO/oyP2vO0RRn9fVMyf37tQkvmaloDZVIP
L350qJR8v8VbsMhEHOPpE094xmVhAo5JgVfJmM5PwJNmGpDz2uqOtGGBKXuwdDetzbDo1IhfahEU
HXwvd8VCIlHMxE6YDgeD+6Akpy1fEnkfTvWtEL0dYLuOVgRuU4mytWIjA0mihSc3/MQ6FujChNR6
05sxSKwIwiYaIlEbub1cZPKqHCgYNkEiGrazof4U9YeD6BKB2LMeEPT89sMa0f4m6I3TDQpdUymJ
paS+MTbdHE0jufjnEu3k5+yjIrR9rCSS6aF2IukRQRz2gwJRw8SI2BbTIMV7Tjz+XX0V8DvaVzie
j3y1qjsABOAITZeFsHjC9teqzZBg7rB6o5+1m0i+vzgVvHGzlEva+RC3RElQ01vlzA+6SZKGpZ/Q
CujpXGm8EvnSVjNLGbq8M6L4Mx8Ow/IuyXDyyh9v9tjasPpHP9rGrfin4vxl5Pv3mru6W5p3BoJK
mTzEEr2pSjPysmkX0bdbZc4KSMH5TiTqmTyKDjAFXjKDF7Jm2OjKRb9+1VusEH0Ew3hMJll6nHiD
bNTMcH3wiKLmjPKHDKECXBGRg8zprZxy1XjfpbL9bcquKDZKMFDIGVMsOZ3b1KP9zK5HTA4v2faJ
v7AHD9bb6L/4A6XPic/Vj75H1bofN10W6R017U8IoWeRG+H0Ny3dSrYh5F4eO6GHpUEsB+oakt6o
Zzy1OaftvzBFEsnP6v7LlMXGj9wDKeeW2bSOqUkpsOGtMVlxHzsI0HlDEnY9UDQUdNA87HjBqikQ
6QS7UaAFsyT5G/EKOOwMbyIXVPWqexbXlo/trcXVY1+kHfQ2aLPS/YMB1C2iUKj3phJtsyzwJ5bW
3GY6fYtQwe2mTA7oL4+fpjED0t9451gXuAb/omtwrGrEUykyCT2aPE6cQFsgm04F5WXed1XDQAGt
7WFxBBczXRCXBWGdH7ZDWw09jIwLLL/gs7xVvu53Td6DIXa3bR5IqBNNPHOYvn/iFjg3VbdQ7aKW
6xIFQY8zz/zqyxQlpywYYNORC3jgLRFYGjfllOfxijDJRq399095+fC/b0jld1fulpTSG7aH+qfn
dqcXmG6OqTyUJ4/AxirDCiZNpXCThE+q5f0M0SOPcWO/4v3m08cZu19GAh6rmkPOkRF5GRCxj9z/
DzeszZxO4jb1IxB1y9vmj/V6x/rC3zgcUR6Z15sNZ9PjOm68Xtp85INHtDr/gcwBoFRDTR8F4CAi
ebjmauDSEz3Jz/pTOpvOuxgMKGyB4s5Qj9yMgOiW1wLROunhSot9ndAVhbSZjckFNNDRSZ9NPuQA
gSJR8WgiLpNAijK6sMJZr+7t4p3gvxccibPUu8NeFtMsX9SjKUpbbMmvqGdbeh0hoJ9+0mq6GZci
YIugbDQoMbD+ohbpmVf5ShysrqpMH+uBar+odBF1MZJhhQ7MXSrZ8CuXI2i6K2H+5l8vIIU2kS8i
yiBQpZNfmRkzaL+kDZT6NXyCjZLyntuL731FdKhpDjrEETpgrPTetMJcH3UCCDYUEV6FGaE5jK3r
5PuCGaoLFoK+W85Ia70PVJoGsqLh2cljUF6MOMN7ipM/A75ov2eEkLSys/302M2+tluNZgqPKJbj
pdk+mIbQBPPuoZKFtcA6YXpTryNSD/wI9jIIVXGNMJ5bro/0uEdt8nCDDxilAPYF16RP5O09NcJ/
t95nc399c5oKtlkiaqFQhOCKOGBqIY76twbCV4TkWxqYhTlNMHJStm1OMV8XFVyk8fTQEErqx1gB
Z7GGolvK+0T0g6WMrgC0RA+sJxavA5ev0Nt83TdA5L8MmOXX/U4nGvdfX3ETyg0cH9GXRGKaLT24
4uERnNIt6NDcREu8Nk8LPVwVLuxx5M3uw/zCismLSjf3ye7F5n4W/5EC01U3iE72MoaXPY5GHss0
Lg7ih7eGmNAYIgppLLN5de/oZ94IZQF6GzpA29Gaq7waRLtq4A8GMS8kGXLQImoegwQL/zqlFiWl
8l/IomzxzDDUbI/rcLNbavHOeg27aH8u/co4xvBPVlcojZvx7UWYR8TAoA5enZWpeY61FVgJz4Sa
3nofinW1fYFJk97t7bm8RHMMDFpchdOXxVAMTU+wQE0WJVeZcA/lQ+XVACn/vO5scqwXqDwBcgVu
4Z8eTkCgohcgoS+rziXaxeDtjE1PSvlRF8EiLQEQAs2UyiTs9e9+yHSLQ6InmGWAhgFQHexsffGa
T7G4M05H2bdjfLyTWXkjoHITqhVzU0sVkv+Lbpx8TnxX5fekhDmzLnCZ/hFrxsHocE4agrIHqS89
NyRhxQODT/JLQDv1BJ97puLT0FeT8Sl6ML9u4mhnPzMLrnqbflIoz4QWmR/Wb858YeT/H9nuCUo6
DiS8OR5w7h2SN303/slZb7O/wnXWAHyHGUPyNxxphNi/fS+REcoHyyaFaniZBzAp0on+L18Tr92N
6+erDvi4KILzKtlWR7LNgIXdTFbYW7jS1ecf9XuTHlNj/cSV/f1tYrfXISjEHSxcokWc6CqNRtwY
bTOQC9cunCrBW4CvMmZIzAiGIdV22UNMIiefoaXlPmMvuQGQSfPcplYQTNBm3Sm+hwFpomIIw21z
S/nHgqEgyMKukWD+7tl5ObLiIN1eLoZw5J8JW4nhRePqmEx2mMNHSZM3GpgElQCqpl6Thy7keMW3
YTMZ+Qjl4xKSso7tpDqJrBgE/TcC+RS+xg7CZkZiQUqYoxzNKy1X5ntIQLXq/x+qUTneuYOhO6Lu
l4Fq6jw282S2m/J4BXpopSJtt6i4EbdaIHN/Zp3phZTxZJqEjd51uZYAEq4sLDkLwt9aVvvb+JeU
LM4w0ZL7jnSPPvy3XiCBl6/B1uRyKtvHqo/YtcupMG6nZQgPv5c5DD/GgmsAjWplcSjmRCX/Z7nu
9EFMclwodNnp7gdaLppvytJHdZ4hgkarDM1Go/kzopJU5AJSjlfg19Yr/U5ERHngDuYYTBuf+YIs
h3wrRgxqBwwQ6vrBfWsFoTfl5AKqCLMIZObOobLyGLvNaKrAI7YErmy3ASkCxIsMJGUboI42rjVB
fl6uM1IkTTbUmsctpjptptAZ5VHm9zR5HmR1XmOO4skpoJ+3H0Ew7mTuE/HCWRhHGAj5bAwoIyPV
6j7PhmMOcIKlnhH2QvQTR27Ca39ix6979NoegI2Ca9qz2Ue2LZfNjoPLcoHRkgxhK1mH5FGBFQT8
G5BdTCk35IWyzmp98Lh8bR1P2AgMuCUaodYMJbKCKRK0Mh22KESD+7pnkGv/EUFfNQbPYic54o5h
fqqS7bMHhIPXjT01/5xdz9x8/2Rf07bTEgs16WdCLimXwoXxHuGMT0a5QxBtzjXuyrDPHYI4u+4i
WIFstXdr9SypjDTF8niLZIzXON15bZ4svX+rfq5dMMxNDVwJhI/2h00r5TJ2yx+9aQv1lLtcrATj
daf0VnZMz7xWVm9rIe6AjjXHtAzj9VdSx6LBY20utalnPm4QS2oSHLwFDLXEptVM2Uce1IOVmav7
rjsLxMoLT7GpQ85Xh8xhYoZcKdlHM9Kx0uUAQ1NCtFGw5Yl5zECskOwOlRZp4PlJL2eJ1yNjZfr/
Afz7wlDmYvBH9YG6zxQDLCSJ6gH4kWZ/1XNwgB6r/QyQHN0XKtam6BCZA9BcNzC0DxtHIxTJGHFT
I60Q95DUBcmgPjlf2D6u0CQ/qTJMUR59eP5qXK4Nu1GTie9BB2D4AcYHMuoBzPI+hKhNOKyjUhYy
B2B618KdmWVS2jxxSaxTsFRCa831tPCPQSEu4MG+Yka6xeQHugwV9/g5oHEScd/X0jrdEo+WuPuK
wIKj8j+wBdQwADswcoQSWW/fsX2/wT+fTm75qNz5Y6Vx4iNdMVllar6y9nfyuBNI+TSiKMRxgfqO
xpy8SQHCmaXIBOGJWuLO0FkeFmFqwHjuR+s9BBSP2gBWEbQUCUK7zPDKtcVnns46a0uyyq5F/tPm
7YS2VLA6t8vwa52z58Zqmy0jLCH82WykL+aHEbib7N1jIXzmPau56+nja2ZhSMjbDgX5Z2SiSqUJ
rjHMr8Q+8Esz6SBWHSh0yTAi0crCYkAlI05vA6euNPwqP4CGzU0jX/kXurOopzi4YPuR8YBBdoqL
jWFLsCxtqmYesgLZG80ZmsFL56Y17P22E1i9hcGSmKJ9eFgKUFJLVhuxQwAst9OHW4ZjnPwRR7cP
QuAAFHdddMAQ6SaaBjl3HbaJ625MzCR9dVYpT50UHG0EREEF2hFM4wyrLylmC84tmx5ET3EhtC6S
oU9VpB/1lolcIIRZT7E2V/ed1MrjaPOs91P+cWFA/japudi8gLTFU2c1cBXiooI+oD16e9mtYALu
NU8WC5cQh5Xp/HIp6f9QL2SrEsViOeoIarAh8MwGy5vEMaBhkYCiAPLrseCCnaef0RQe6E6ap21D
aUxBTwt2+IMHQFsLCl1e6KMee1AcJAdfdVhStyS1cE2AtUdDm7kJuvjwG06xfdRrSzmGbkAAV6FZ
8c5EFoA7BeNY8/ut0bvXxXkTEEAjFUe6nfmRq2bPHOe5hVwp/t6WSeHGpE4FPixGyF361WY7l/7O
pc7MrMMQZz35KPolpwllIVPFIpyhagC2g5/YGKOhueIn9iXZwjOs6mknNy262uMYXvrDZZeUv/WG
DLW2T4/dHIP2e6y9NN+xVhmCUl7b3stGIqB7oui/OmJ8e6AngYqOaw8pqswIDywznYRSt01KsVOl
Ikddca8N9wPwEZXHZKlS5rBRI8Dfl2zoTPCaJLsZotTl8hZDsZ5rKiuTbY+CC3YE/b2szVViFung
iLc7AqbTheW0GwjLLjs1QLd9/xAm1cXt39b2pf9sb2gsWgdLBJ/Bn/TnYrG29Kehi/sxuR+7NMJg
QrhbMi46+19+lYRctpDkoxMRg16YT4LDmsydhdX5cPH6xvg95EXKEam1c3NhprxXVn50o2hHXX9E
Pd2umr3Q75dfTlRrW3sGAfTuR85W/mcC9V+9rq36OQbsfFs9hz6hSh7G7uOvrw5pTE9m34UBxs3w
BXjm8svTg8J0uo0F8ynSvdKy0DD53QQr8yOnLOPPeOQSdCQF8ndSGFZPE+LX8LK37iA5ad95qZ4M
WCnK/UK3UjiedilvqB24C34ngrsa/0ZmlcmU4lw0vwgdW4zS9GCRDClE7TJFdbHivafpvdj3MZ7V
e9PlF8fVBi5A7QB30b6vfrCeRqdYZc+8ARTMitfYi6yu4CmnokNolwteNXwnzO1+/g1ktf84h4UK
vdHwEbhslPQiryQAeNShomN8uMvknvRu9oQYBGCa69hUijRuXFatGUw5KsuJzqXubYor5GyMaG/U
542w8SlhHYIcE+Nq7n14zfHxsu+svVQ1I0JB3tNKxeSQ4t/2HbpEwGohg9x2h0VymO5eDiVMmhnh
1RrrDAsRTXHXynr7WpNHpo1GfhuduwxUoA2LADsdTQCSRq35grk0mbGcfIuIug/qJmsefDiJHb7e
O8rsxJvpuvHgWC2QizbW8C2UXZITrA8Y2XSG3KdEyPoYnehtr4zWlx1hvnfYptTCHQtSGLe9h7N2
V3SwnnADKVdSgHKK1sparwg9CAKwCigo4tNMssLZez2JYWH56i8QD+9bCcb808mYPKaE9+p7ujF9
aOXD+4U4B2vcMsjPhG/UXwbjcgdd0LXsc2vGjrHbQYJEi8SbY3hgS034cEyXGvwz9N+hBPWPEidm
wrRbKdrmAjfeGgtZYBFFdRniW1Iq4yd/fLiKqix0TYMuCll+hXgXh2rFR3GXrySPnkIOjvclLfAx
NOKkpue52kWeXzaTQfqufvfltjuSbxUI/Co5lOvRmTjNiP/gjiIyAkeWmBCaNBTrct1IgS4891DR
TdONuQtwK86braSADMfOZNsQN9HkTzkAPwh3XhKS6rpcvoxKnnYRW3T88XfXadbUjyj8Gmh6kobi
XK0D3IMmntiLJ5iWz1qi9EEkL+2tC1S1MGNYxIWSzcjVHeJJ0O5PES5poB0e4NBu0BzfRxtWNh0D
KP9aC82J21HVp+yngHIoDq/jVN4nMtN0X54oVcd/89GgnnplHPYin/8WSZUu80VvDy9mNMHWV7Pu
uK9atWs53MaG1elq9ETIWcMKYs9Xf4ccvCQdgkJhnrKEI+eg/tlIBKagK7W3Bx/KY/65WJWtPByo
ZOZLeN0ACQtjDo6FV5Xn8Jh15Q5lNBZWTAEuaBeUhX83fg5yZx8aZzQo89e9tSpFQRTG2Wh/sEvt
crUJCqIIufR18nI11Qxy2JebEn3Mi/+VN4Yn9EzwAGw+d+63w1fC1AZDTEkRJvhufuoVq5kZMY+K
uwC55iNouTzwS6WkviTN5Bf2JRb4PU3n6whzNU/ZgP9EClAE8h0JK2jbRCu/ufp4pL37/K4WeU7r
0uo11OMOMSe/zInptOlJfoXFlX2BKQchbzH0by2ed3R6c36YN1/rcnRRDJWxfvvV0Tyjcm0nfuEc
Rv/fhJXBX4WbjStKTay/OmtYdVDKBnerJogY/Pu3CXdXAqIyGif34rYti/Z02fFIFIDrd7w2MnW2
C8lsUkcMuGwJkpHCfX1Y55C+0p2cid4ijBeVOLh1cvD8n310cwD35IGCsfhsCGDM91AiUjIFk0XC
Un9V1PReTXVcgcJkMPdM8kjaCeRzRm2kQKDmsUAW3fslhGexqTIodbsYOPSIhRFHO+aeDTamt3p3
QC2EjtNMwKAIIpHlrAybAuwwQ9JI4dsXFWzHQUQ7RcracMVTESV6YStwdxyhlgYr3pDdYBI3J1rC
vUienH2fXI4vH50VBQfJjc9Duy+pWT7zSbGT4JtAqdnyggV6ixzqSLh3RrlOuajTVz22CgjKbTCv
SlTvgJM5D2LHH5DCCGVUgJSiMKIPJu53xRZKu18WEWtCgafKAxAJHT32JqPpkQTImA6KHeJQLop+
m0FS0PVhxRrX6rq6KomKOekRyiMb5Vs4t7bA8bxIEheVs8JteYAHf+QGNJhY1NxHzTfwV15ojx7w
itFIkA+80ZaG7Z8T/gBQNnG2HrCc77jlqf0XN5/WaYtONEVF7tGAO2tn0GDd/M9s1f1Z4ZiZrbax
1bVN/CUhUeYuLk5e6hC0r+rVyKxWuy1ZQywjJ2crTilzCQB3C3ZLXJPb4Q1a5qNktRIRQolJu0Kf
7HfYcRK5m8houvXbO6yJD0VYWnIf02c0inVrc/UfYRpEprZVCiq/jwiSHMnEoyM+sQFMWPnNcKVc
O/otnQ/74Rgtq4JBJDbuqPZjQ1/vMyJC+VMA/QgMnvSyJ7PuW8nqbPkxXT9CXpsUInYsCqiIS9na
hQvUeFUsc8XJAjBszZYmpHaana7iM+vcpSWaRrIhSU7eFmsUZDJGQAWbLPavex3OjmFJV8HCZIGF
eCWv3TliNmfo6wabC25pmmVxmfTq7QH85TU7C1fQZ6LBjg0AnfeoOal5enVERYize0goP3PFsoQK
JDs5fxmxkK3T6SBTt1IyNSqlWcaZGEwnaXEMzBzFDvrjzO/NNYObkZSao4w03gT8ooiph9X/YbXA
h1JgxEY0aXx6s1R1oJJET8hSGnPXdjUcqhIOqOOsIuAj98JSkjXkAjuMkuT7MtP5znHxwi0DaGT9
Gi8wO776lj0mBTWIa7N32volWmMADb0eYN1pHSP4Gl3vo5OeMV3sB1MTb0+GZaEFfrV42FJTvKcg
VsC86POdb1UdeHFPX+418iCCPS3kMHf64tRqVJ1QjJ6oAPFld5cfXumlH6qo9FBKmP45ZJ1IesPK
uh+BTayCB8j/uxDbXMOX/lSOK7QfBVb8rrhbxvrbKkKGNte0nDIlltnB03FbWu+1VQsiMVr0hD5D
JpwFRChUaqYudHiIkbOaAn5W6lfNB7MdteBmNnbpo3I17qiuOPP1xOkspHfNZGRSni+6GrUxdjeT
urUq7FAcGN07z9qvK04SbjF3Knge0npVvQMZHGoekNZ/Uj6TH/ypBXF0RgQ4xh6GCADF6YhF92wW
0XRH/qNMhrhpuqmz2NztRywhxS2qg4uhXWySBbcRVYgGTX9hjHN82Y7UehfsCC8guf7PMuHTKW1c
rG9c7jVS5O0Ar6+G47hx9rKu9lcf1TX9wgsSiObhZZ9rQyu8zWRMwT1jC6LkMob6Aaw61e9ramT+
B3N4pnehJh6YvOCeIelKi1wpbwTluZx8R6k86X3YtUPARN4HxzhUtYfBnunw/hamvPhIe3nWPfby
xVsuAyLIN0HEl+NfdXJU97xHJBHJyFu3JrR1ITNLUXPOl4pHS246Y7mes2ClOP68jnfmsNfUDt/O
p6JQPELUfX1QdAvlogmalg6x7RC9n+r0B5VKSbYAm+f8CyD+O5hNUQEvW9yb4Yg0PCQIrHFWUFoj
bPOSaq8lnY02BE4foMfeGM9M/oO43yYn+Izq5rXD3BZaSFvnDBHHq/zI7inLvgxN85dZbBVjUN/h
jFvQReZKHztLleB1PE4gBks1UVRgL1E6iQVQhEdehHLLawglIjMFNvKwn/30UdjViyAcnwijPfz6
pMPf5l7opeNE75kXwcSa1u31KQl6xKq+N9urf2SIDAZmt2RTToaROtI/5XK5o28H5up8EslOUo5F
8ePF47KE1ehjQQVcwXxo4yMrFuAnnsV9P6zvS4nFyPvqAh6Tib3l25oPgL/vaZXfJbAc/bGRWl/w
oSyVPu6wXbbXhBhiGnK8/gmh/iyNDjDI1ku83r+wjU2XXQBE9MB2P99kdNxFzY3qvi9F1ITzuFtP
gSNJOXbW7TqEvDOW6UCzNrOGkonIBMxukKEkoZ8BWYDeAwOrf/JkYqY6gQCicOjbCE9Y1sSDKQno
kIX5KaT7mt1oMN7/FZTd3L4zdOM8s5lB4fYRFJYPYf4sOH+6htTOK6tw1c2bGhXlOX44GlOkFX3y
WUn1e+tQ5J0aJsQCu2Pvl2mqvdraL6B8mcycgtR2l2gr5+zPzD66GzyMAOanXvnAysTMCrKJIx7y
p3gR8pbbQ7iEpeTpfa57L7mh9o02aSqkau2y+yfs/xK90hjH78IAYe1zKAtuwDWHIAAJhe9R2a6w
hbO5OutyFGiK5vl1PiEPTn7Ob6b345Wfxic019DKlfWYf0pC3bxJ0J+pz49qfoYPuD1are6qPYUG
8OE1dngoAefL2pHcCxuWSR7wTpedf98inusuSXX6IF+lc4hg1lgPT6bMWDm471eTCNL36ctaNbfO
AMh792DLQEQdpRw4rxA8UALeg7XTnuXCpgp4NFYccYDr3lgJLAhQ5nkf6scYaaZ20UzNW1vVTfGw
NmeUghcfa4SIz3Ai/70W/KpKFMKf6Z9upSimVyZ0kEHSKNpW94ZyAwyo/fYalRXvfKGYsEzZFFK1
8CufVvg7x7Wg0fVTcbXIYHjX3MBODEVLsz7FyGFnQjsrDih7pltlEyhK/aUuEYivll37FkcsnWq+
gfMV0lOKVrZCxdgoQBFffN3YsVAmVnbl4sW51uPQ7C/gmATztPzsOiJiL4vj56PeWMsC0Lzszbs6
SXZ6PuBK4+5d1lrJ7zXrwf3VyiKdsS+zgQbqdGRGfj50B/aYv1IfVcHT1rsyu+2HYHG5qRM14REW
9tbP6LLk2lUbbCWjLhQNrxK7ccqwAKCGtK3zI8uWryDOOinAMXK/W1yXzp/zVXV6INAHLQPTXEWN
xbBrnPCT//hvHOcl2wVUteDdFy+3EtNjHMLDFp4OcRjMeWZlIxUdYoaIhjbMY001q/A6kH5pBoeG
ne5I/DXhv9PNwkwluEZdfVdo0u9vyorLAMpBbpMn1zZNSM8YZujwvNnOtla7gm+AzXWL7CGFaGvl
Wo1cw1FFFXVaGjyvqI93owNsCf1NlgE/toapT60xOnAmRqxGc0NHh1YotOyNl6hRjvS/O8QWA2wS
f8jytWBicWPmyqsZHnjBvh4xtalYKOhlTOsO9OE7Q13129FsvATRx1WL0wn1pKRtWNJiGLsvPTtY
wewR929mQhGIOTzlJNuEIkIz+Xy5Kes4oYa8vBg/kKBt/gd7UZmbr+0Pe1pckumrFz02aaDdukSn
rGHe6jMwUBnAin2ORooYp+nEG2XMDzNO2D6M2C/hMYXrdotYLYjR0LdSzZxA99REnPcK/4YZRwM0
oLJP7IPqJ1pLMhazFI0FP8N7u59iv8Yi13gSJ5gg6r3fi5gyaCFtZwaIdYNp3gRRp6JRCk0VTFLm
IYZUVNVTK8SSlhk0a7YMcGknC0C63yw2DwxzBhROLsDFTzPitfSUcsRN0LC7HImkaTLbcbbMSrcv
D+7PIEvHjGyQ/Zd36X1Crda90dodtXGL9zPJebewdfh9MPnaetZjV6wKXDRlbwxlEoR8P9WGb8n0
aQ8opQDGwA01prLKjv36bmnOWTPshBrG1cp5qZlDXGl/nwe0FQNpuN2qiK0u46GgTaCs/WrVZoYL
GfZthOA+CAv8oQdqyKEYvjF6LDqyzhSqA88t62BeBO7eYYHOMjSsHzoMcHKGP1+UPWfbpdzdfJNO
RdG6qp+QOSRI3y7rFcDs7uE1/zR5TFLSYa6CdIrH8dZ9GTTtOxLJVddg6k2ufiCSqcTlTDNkxJ9s
iGikHVhb4DP0BiYUcTEQ6xC9LGKfxagvqJf+aRHaXeyD0i71lMXBN2CvXTQi+P/vTzYlEyCJ/kXw
BYZShL0jPdfEg+uTI+skZ6kvIsDoOeYUCidZ7UUTLZHfWDsHC4M6H6KxEszW0sXb2ydhxxHfTpCX
su4Nrg3sGr/SGgi35LMUgvovvlCHoMWgQCtZpUyiXGqKJTC2i0b/iRNxMu3Yll2pQUurZQ9Xgy23
Dmu546QNExbK1JqFyoupnkBYubjgGi6dir1IIucIMrA6tACshxaNd1yu3VZlaqroCx2zeA242BCc
qIW4fnViTryocDtmtB2owfI8HV50qgbUAn7VHQiIB5OeEwDS4DyTccrJQGT+eFeB01uu9hguD3Ql
/ggdMdRWswmvE9FHIz1RMuRPQiy4M/UaFf/jvFRc9x5KyeDmF9ia74DEm+9L2SUmjmAClOWHA/Un
To8XGnLZpVF1WUUXGw3iGS8DZk21P0DApU2jEG1kgAqphkA1cuRunISkTk+72Tvba43S7yRFJg5r
uiOCR+3ZeSgT+4v7I28vY+zKbLgxjtE8CuULovw17T+9IRvVjUZXQLDU/aziLfC3Ya6aUE9qCPyi
r8yQRm0j/1N6wCjE92wcC98hIlfp6ZmPCE7tsdt7eeX1b3c2BXZ9S6RzBacDVjYEG0yu/olGNKHj
5uxG15D1cgrqzCtoxRuqsNftwrj+4+77jjPHUmU/5oIbHni1RRXpHVFGZmdHiUs/xB9IIxu0Sd1j
UaBUr5UXxWkTCH9SJhVtgXjNtu3FbwGUvhV/CXgnYSaBWhiqSXD8QfnRr8T2CpM1ffXxUa7cScKW
wnbInG/kZX/1nYiMJHsngC2brkklo2KMjWiA6w6BQNmghoQfE82qFnddjRngGCz/ru2+hYYVpPB0
Ke/ppQJsE50917g4k3kuGTuXKWRbEdyV5spqMyARK2eQobvgxsY6ZhmnnsIIi+CeOUAlud//tQAa
J06GjlJKOEfIUG9MJoekQDGSS0VwxVDUM+EeyNkMytU/BcY9pjeUo9gjMBecRWv2BtlivRdv0MP0
T5/MgMyyN98x9GPeoeIw4hr4yAwoR1BSuML/dwAjUv5WO/vFpYy0T3/GK47Q0cIQkRdfk5y+1R5O
D2fDYdDuWbeMgvooDymb9e8vJznWOWieP3e4xaBz38wG2z7OZVz7z2mYxhPDSiwVtynAwXa58aCc
fspsOLUobIhX+UMRMOSlcr9R2x3XAIFmsoCRJOJso7ZPpfkDIGtkoskiHOhSZytJl2Uxa9a+Wp/E
8Yex9cjzbmyIXE2JieU1UipdYhYdrfS597kjmrvMyPQ3dOMjNLR8IGqIBjWWWbvL/TMgMzY6D8pE
0oxB19r1oWdeN/sqrWWkRdZK3Jv+kVlYwVXD0U9ABtAPBjm9L6u2FtYi4x8Bb2KNloZcgP2zlkcX
PxkGUOfYq85j2wLXp9b0Jic6tB6xFukGAhenCaKxA1saKUvcwU8HRylRESrxJyUFGzEPkss9iyJb
UKP6Wrs2b7y+aORNIEyVJIfkvf1QhwS2o82CAs807kjAqXdPfQsKibRgqlSPiwfQtKivXezws+Aq
rzT1/FdQG5lcvHnGx8cBKCdUL/hUAlGfIjKYY24K2quCsec2JU5SaiLH7thI2Z92S1PN5vThzYOb
DATRJO708XhypuJoRTo+QZjN8njBvVvPprFJGNxTWW7yWw2xh0+KGaMfMZ+52eIykl+cgNhvfYHb
CTsUYIOEIew/CMW+BWxK4ALlpBXI8WFNBr6edEAxFCWnTTi5iz22VjCCn0MHrPRJjxALNMQsecFK
j0IPA8sIWIF6z3USVarlNYmTs5OPii3iqEcnWAII8nYCrv290T+GUTpPvFD+hnRMA6A8+WX/GIEC
4TpRBilPiw0QofzRzEwTCLW1EtlQRTkD4GhgVVw1VdGpEKJTTSA5OQW0Q0cNpR+BuU7QtZR1ISJt
RH9NgKVn269R1j3FC/cK07B1V4Pfq27sRIoGhfoAVp9XwxayUDtdGLk9L8XiHSt9WKkVtmHgQfPa
188LLKs5Zd4WK3rFdZ1thRr7S9XZskIw4KnxK9XJWV5C540EB9e5+xFLOlGAtErG0i28OSJGtTFk
2dc2Hfyxc1jV/kvOjmSnytXNgtxEmlMWdxVKLO5+/OXFmDPO7HPOGuTAHOeFcTYh5zADFLZIlbHD
cSYi6Q2Lztkn1ye/0whQ4hJ6i8VMNAFgvFujuHioxdHbdlng7fNl621vzb0UBDQbd3pjV4EXSmVQ
r4vHH7r4lmJtOE+KH+xombcAkXPT6hurqCK0VDPT8sOK03JFs5VnzXOVT+wqQg64qnVamO6DMi/g
8KPgbbid8xEzlZZYbVbXhOWYjtvsgusBMg5gQkOvJWy0q6rtL7stSscFmeDTkFZFdHnl/oZqnYE6
DBQC/19FTNn2jvAJfQ/y34XLEhzGKI1paOWTAxw+A7UhYRA0eZKnkghB23bjwBGuSu5fEupkDU6H
c5E5N1rzkyRYN/75bo1cM1MB5BpIiSLcSuyGRePGSwzMx4n8WnSzku8DuDsAyepCZ4hbhWHNTrFm
InRVC7Mi4RJ1YI/TXN5i+LkOjqeemW/NVRJIeoH0nr0RDfRKxnQOzUVEKlJTymDpj8WssC9YaR+E
EmfYr5EW/6QqW/h+CC+0FuS6N6fP17NDq965ZIcfTyMmfM9VjLRssztxk87dRN+CdjTVhoplQnZw
rtyANtI+RL9K4KnNQ+4gE9SbPac9icvOmsRaADe5lsrKdDR/K2loYKViKuHZPCxEcUmCIJoEZUoj
M1PGez1RQQOprtDoZaE36AT7TsXDOfJoZ/2VCcSQ9995DDuNb697D30WfD7A96LBMmaGQSZA13g6
b8EjBdXsGnv+HByokgC6AbdLhMW8DZq417H3k7A2g2jeikUiRKa5ZwyLZH3JEczqXuobtAxw2Xzq
gXtV2sc8ACbWMNxrAhoaA/8D+JQAZOpZchGnYrJRLtiZQydmZCesL5/zsoZpFjYPWjwhiXGaQCx9
gzRcWXQPh0eMCc1ui+opDsFTazG3fianPWF0rAGu1kQ55zAipYP7wCvkZ0a6QZCRtg4pN3QXIiYN
X+Bzyvi6xUu9CCXHh0l+jeeJrSwGUShyzs7OMJaKx82ZHOeheBlOJofxlZAsAG9PAhYsWKvjDygz
gDpWygbYYFiqdtOzn+aWHJJCNkRqkqOgFJk8M3p3vr9EKhqQYX6WjVijVxD9bLOLWJ9XBsMVjXuh
BTPva1XUMLS11AXUCBs/SNWMEyX4iolyj7a7DcTHEy6S7jZaO4os9II55RQfrKAr3+Ij6zxpj6hA
tYICIoH+ashADLh+mUtYAb7VopX++quqFhUmBviD7dk8Bn0XI291+vSC2FchTajlf3lH4Oltq9uE
Nz31xQd55q2Y+JHNHcpitK4QvpWaYfH7YfSRxaLwDV85mld+Mc9Z/AVFp2pjaP0CTN5qoYpo+pLL
9fMa+K37CKdLObfn/uYFHqOjboaxfSYMqpOhfqUYiXJ0+xAjk3FAzDpsCb0j0ZDxScVisseHSd3f
7e/gqzWNGtTnz4w5g1Eh+K9oE8a15k6CyuGwTaFbaqw0yqs5aQOvIqxB2eqQb3RTSEeMn5GE0Mp0
gLWd0Uif3b2qRcOyx8QLfdAa7J4y+TFyhj0K/O1OAb9p94RNIvzesHykFSpa7NAVdHSFtoWKTBJV
N8vIZM4Jq8BLJYTGNlSDioO7knvyG2UaO8SBN7YtMY0vfKruOrCOCGcAzlbg0FVDyxGxqLwJqwHS
+td474Wxv34gE7vcbvIaBesFORdQ5ttkWITRLlSrWc4woH3gpAoqLLwowyH15bO2RqBGDJ3i+iwG
oCcb5LFna0k+XDwbLB0+JdzBJ8H/Z/QpPzHRshPTYh47OWsnIZZ9holm2mXoSMV+qMFC+cRPTzyS
X+liWP1n3uL1cEcgeMeUF0C1WamWUxmeo6ekFwC53xxcxXCIYyNdSOl+rRxTwLpXNvu65TqmsOOS
gjVj2NjNUzFdug2ri7BFoI7a9937YT+zvG1kbUoloXvUb1ZjYVl+oeGNlC+XijU+1rtHTpEmCwWE
EAh+SS7RwMDSZVVpsqBMAe/FHaHj71txWbzElqarYHB2svlmDPS24gJ7dgBD+9GJITLgRd2MBcYQ
nW3FNMtZQkFS1rqLfKcJGOJRopyOT+9TyCMnMbtBFwsPPGBSww197aBHCLOLcSEVWF40TgdHAzeA
IW2YqRNgpd4+e0bktItxmH404RhvaKTiYTIaSwPvcN+DHMrjEl0ndTbQypnaKeMWhDiOvWw3pVTo
9i9etlHai7z5JD6xuli1y3uOOgrty2fteKQJg78O0IWNhmFT18YIvuy5+2jxj/wbVZC4az+Z6Agm
yLQfRT/T2BfUXpjCTFVDDBSa0ANxNFxfoopk6tyJyZUqHf2SWV77uIcL7VOlrt09ekkxED4ljuX4
1UIIbQCV2QlMEYoIgBls8Lmjy7DsQ4b4LLjkPU7rdLaJl65itsJtsV8LmhWRHUj2rPfQ739/WJnM
Md/naBl6eU2+BTIsqrS3wgZBv8Rk9JpXBCjNY6D+XzZnC5buum8KKCXBVL5ndxdSTNTUo7AIoXuf
DrihRP/+gYUwexI7qTWLmU60xNoRS3f+kPyZwZcP8LkuThQ6vIHqZSQasJ84oiyousvW8dDQ6iPp
MnGvlZVzocMekiRqvXqo6W0IpsejUd/a9P+nlqGENkuQoexNKcmbxzP1bL1rWQS9AYRHADJQf7/2
otFIV4pSq7xjPfPwnEWMwctbGjXzEyYwXiedpn03xyyDL/jYuRqJqiDGKXhCWyV+dr4D2fP0N1Co
sNZ1XyuthmFDK2gY1L3aEsyNw2K79JidiZse/wYprYhX4bn0IpsuHroGmk6y4MgYtH0dzSJ1Qs/O
nKZO1520nhe4tK0IFpTjZsRGj7Tc8PH8+33MsGyCL8SBtf/7oEMSjqolXKDYXxCxcLsIZfH4Xhcq
bN/1igh4exZOuz8LLubYt1k5T55PsKv9GhqmeYnsjFpwAuGSyOUPuNxgZWOMAT4uYkeQrrtU4AYR
b+NBpuzBA3twyzFmyzNkiYmftiCElhs32JXoHyArP5z3g7tD97gTDUKlaIGYsSjJtG2Kwf1Wb6TK
ZFylcy7x8UNZXPgFJrM9oc4osxNkB8v3QWxiRf8VOrvNyuk3DLe5JI2yf72KVyfylNNUF7TQLTHr
4QYXwzEvuTz8IAYmgc4nti8WOsdOKCO4x8a3sryuVi/YLBkFvM6Do05bBVLgszEm21text/ZAtJv
49lZZoB+0qraT6wPmc2iw/KQIlj6sIF/hjRhsipSvKYvH2yqeDjr1bnOntg8kY1MJ46ADHmnFn9A
bOLjScHPnhpMvCbowEx8ibCOIywvL3qwilHkOuYHziAz9g7ZsoRVtUBL/kkSoWNn1Dg9BeAeFRL1
LdW/hG81/Av3iFSVV/+NY6rx66LWYgyHkQ0NkzF6DFsmfk55KubfWZ8sJZPKhbWvY1kjjAd6D7Gj
y7XaElY/UoZbrLjBkG+x0HKR3SWGQ74CRCP32L53fRSYNuVxL9l1GeD6+CmS8GNs6c8uACVub5Qb
VPPjQN8CjBrTccq8VBsdxOEo9zv/U/DL1NvCEHPOE4rIJ0skAT38M8MN087Yc7tXuw4Jo2jB/czz
TwCu88rhlJy2459DSyjswM8AmQEVV0uc+08pQ/Z/GMXw5z/abeZGOOZJ8vSItNtSbW4f4hVea7nu
VriE0FL1AUyXj7UdCNRQjc0d403w1Q6VE+0EOow3x2hVsYBC7OOohFxx4aPQnXxcGjPeAbKn7iFu
EFWdvJRy2e+HOn4P9UBYde3CidjhojNxAJJAgxo2TnBVk/FTM7pVAO57+sprRyszNkbQ3P25peOS
MHXLRXLxEY+bf5vcAvAZBdgQcMv4fxF8qfLxWT9CK5GwA9yCfEokrc8XM1nciJQ97mTHlHcX9x7h
7tc3tR/WCqysEJaeeOpu+OmFaCH9dGqtHms2uyBTMSsf2A7xNHzyp2qe95dz6KDD9RN4EDXE6nKa
FTZa+siVJ3wQsSPi9FF+2tfB3k/Nce0HLUAjcLS+8wvuC7MfkammP4bQUq1JiNRKRqo9bXiEGWfc
C1RS/DvCmBOFWbfbyd3uRawSR6+9Nr1wTW2lr1jnHTDaI4KUqdDPBTVLQ1dLmsNrvgr2qhMVgaG9
kJnhg+V+GLp+FBW/ZVyCwKZaVqBJmRwaFWgMl6ZQtQgV+CS659EDcl7XigouKD1yIzNfm0yXpI8X
SZLUBNeECxMTAaQeWWSH1OeMpleRPuUlggxvmLp6uJcxknCLKbbg+ROf3ifRROj5D+MoSJtk9KK2
cP0CGcHW8ehQWoeF7kaFIJ1aTXyZJexy9EIN4a6wTJFSIpOhvRaqUszIVyWNjW4Ro3m/m5npF5t5
7cAKAGD0bpbEa/e+mfECwG6pSOVJArWdlb2OimX2Mso8XinOV1PJrnOjRMykmReA5PBzopskYP0B
tUy9/J5BEKR3wtLhKi9r3Lo2U16OH0PZqFgEOySoNOa7VAFKQ8Ni/8FbPouL0kIVb8qVXx6EpnUc
C5GbK7zZxKPM8iu64xDv0RkUq2ah+qoVfnNHr2iqJpkuWZlE0U96vKtmo8O8GpRifnArf8lA59BJ
bhd9hNFpuikNUwv7aTa1KgVUAKVJLbmheqX5rmIKFur1FVNV8r/4dXgR7trrVgGPLw3ZbgvQnDvT
PODrvxoFeZ6HJ/TA1WLmLLJTIXmbJ4TKi6OkykNmjQnbtAkrPUa83LlGkAMdHx97Tynp2YNQkR24
F70cjXxdEx4rJS7A7KjUYT7NRGDvMjpupYToSrztXhNtANF1IttVwp4gfMLhku9vY7ATLL5ztDjy
GYX0G22rCkkqoGPZBx+o88pCd/TAb72RP325aO7M3zyq1rMtThJ2NG1VBtjaFhqpH/MPW+c/l4XW
ML9zQ4/a/u6bO59Yk2EImeQCrE9ooOoVOXzjfbToE2cWfkPCDcozmaLpksQzSnafTFhq6fntPfCP
ofzvzCHBlXzmSFrsS/25rrzbIMsAanYOooSctjkUbSSQH80P2Q5Jq0kSJfM5KzYyhv67mb5CenNT
yRorywyNr5q24ooUvB1zipK3HbJApx3PGYxakaNI58/Z/bKHjDlQ5MBoSs/i97COcSTRuVOSLreF
ovYilS2tyO1CCh8am48Z4Lp+sNDN8Qhyh3U47K5x4L0GxLMFrG5a5iXROuG/tcphO2UYnN+5//DG
Jg0/d6ELefEum4aZI92MrEjNqxggQH5hs3vAv2lMxBWs1IU0vcfLP570RWtw6ehrqWDbYvZUyaZT
DW1Bw9xysUnhV+Cid1Wc94fxuDQsHa6b+2evUkS/TWQB6IzU55fpX5bWlwpoPbL96OqQon6lmGye
R88SuF/cn6msViSTzIxIFSC2d1X19ssSmeeXFJeHpBee3NdUHd5p/fvkWqdhTmPTmXeFtWnEQ0wF
ALaEDLyCHZpOq1WokkXMpWg/8R/8s+9SVU2m7ev2Uz5WGo56s0OlHsmACj7if3qusVHrvUxEhVQR
ypaEWaI00JxaS2/+AXQ57ypncufzJ4YMGLsxhwEv604UVvkYLUtvMmE39/WHtzTAZNxSUidGC0vy
3R91Zp/xk83YH+LmCZqjh/QbVLTkCL9TnVWkCoU9UftkkMDT8YJjpaTeULfb23RrBnkkoP+9K/Tl
gxXYmujBIw532JZrJ8qWdU7ToOrrdavT1mG4UHBPjzShheMuguEPKzkygUYzaHVP5qE85onkrhhY
G70PW72CGoTPEH1ZltyhdkdtiGDZReyZGXzOQwMm1+u1dWDvSBNodBAYECM7Q43ptjTAeZEty/wF
mcV86yqgblH5DZ17N9LbIOiVkVYd6H60xBlKqm3vduPGtwtfOCsMxlnAzV9n9I1lQnB2gGfUtqqS
6x/rawMTsj9Uzjo0/t0If2KZJ7AlEOJozyGqEKqsS5ivNOfgJsUAxXhcmQ7m33zq/eBBVcxAzTpY
38Yf8JLktwx7G/TNRKx5BEphwvBZMSGb7YLpNrMR2mwkTV4uqRIE0hJvByTI/Nq6cMckjHNV/wWr
QghNLGy3fvdI+AicHJWM2nN2o/ce4fiUooI89qHoiKe2bfpUbpI1PHJ1ld8vsI/YJETC62Rm6WnI
ycVsdKA+eElJBpLWX4G7bQBkPFzv0MYhk3GH/FfiC/ngPjcyqUjYfOz8fOHc2r0W5F+TeIngiuyR
XoaZe8YJgQYTC3u1MAE6o1B+tFRXiSoG88vU3Ykfe9+xia9cBO3GQVdTzF93hZYZpXtGscsEwSro
b7JuRZmEEUi9SXcMRUDvqWXUuHFdDruC5ulA+r1Rke0cugHPp3fs/cbmovTbE4a1sOZPzFGKUgKF
0QGp6hTDSEAP5EO+6eM8rzmGnaxJNLLVzCn5GXjZK56yP14VqAwsWPeiENNk2sBY74wbdvxaolVm
LJZmptam9wCJ9FpVJJ2FV2WW8DcWDTqvVDrJaFQ2izUUhhdYX7c+5e3WTnrlI95jpdFHqJKpKFyD
GDzoXe8SXl77V+xAa4pLKvJT6GfdlL1YKkMxY6rbUYzKpNgVRx85UV+taFkumVSnmaiMRYEWkC+6
wabYGB/B6/DYFWnmCIzB69WlNFX0I271Y4j4OI4jU5XRhiyW15XJynfGt3+qkQH4Uhpzx5OUcNv/
CWKyPoGmKXnjY13aFRHcZVrxi+39MkpjgGidiQqDC5TctBpEJhcVO7x11p1JwvZ91yf+h2Fgjau+
Z5tWlPE6RfAE1kK7AyPAABmXyGoQatZjbmRmvS2cjnr8T/xYCqCAcl7Th6IuXGWBgrBKXao96Vff
Qcqho9QxFtPJvqFkJeowzXWDBx/JEiRHmoHtmBsdnuSrml+Pii9Q59MKYpJQfTfSABuKOMygr/mU
TLgrphsd+8iYPY3GchvrvmoO0eX/cAof+9ml0qFsYo8QDDdSeYkf7te/6UTPqqmRBznl6lQd5hXl
FPDR/cH+CKkIa87PVSzgFP7xY5Lij9sj6R9dIaImdo+yfpSkNFO4rWQFjVu+Evpkop/dvqY0mbyg
Qfm5lVbyLgEWaMGXSi9GclAmO06scG0EDpbbghg6toZeE7MUeQst3RQOgrDCmDgSQFFs58MI4FBe
hMkjs6XT6cQqcRK3VA7OCkjl3AyaWhYQM+knwRuEQ3abrhMTIOt4jqsecLhyCQdJHqaKHX2Es7w4
PcRYYHtJL2mgE4mVSDQ8dDH0i5nLRe8D2r/zf6WB7GA0eBCr9HGRwqBpXRV9IHcc4MrM21n5AaWW
bi9UA4NN4SoOZMBrofVqff1AdKqXs7rwzB0yornZb81y72iVQLGOUHPhuNl506KoZ7Sf488Fetae
YL8UIxK5V4WB96uJGgViLbsdc3pzYpym9zOYqxcVVej1u4ousdD6RYgy4R1W+TYBVa1ptanVpKpb
YaaPB5HMW28B5DhlknthNY56eDpZxen0oV+3XKygRNPohzIMl+BAf9/DPI5LGPc1ke2nBClbTU+J
5Z+DHc5D2QwDFa4RtfBZZIkpQcAN7ECJSsJ/dZ/Umj5Ypt5U5kvaAtmApJ5B97GDMLDBNnzrPsph
o55bz7f1Hfh5qwiTqbGdN+o5UgEicyfbIJFcr+whhkz28Klm4xngb3bX0HWn9x+dZrBAa2ncE2C5
tkIAyDHGcbRx/p4tPmSJCyaJqxeE30lKperxmWrYzTq6zN+TRtGtdypc3SFJ2Se40JoKjSzSA9+p
+Pn/2MmnocUW1h0DTVSQwtHvfc/Gd3j2NI35YW7pl2tgPCDkH/19Vvhmu0scYStMX76Tzdo+48H5
6m2IZKx1KA3VT0Bev6XNx2tPSJP2gaLucWD3jGKezj+SnYvBm02kOUebCkUvTTWt53rOT1HMUGhi
3mDas/amDQtSg451tnoEJ+ZafX0pUnbZweTyjdvaHl97ahICUQcniUCXOGQCqrZCxvFAjEJV4l02
sBBtxNUPEHZ+pjRFAT8G6CHRmcXev1soe76ytba3UZIZocZiCsvMx/3Y62oRIR2HjbCucFNTgWLG
tTpL86BKPt/Mr8l/lkkA3U3Oz9ntNdOkDv8dMFpkd/Epcnzfgk9wytS+APrjySxOqGfqubIE3Tud
PfoG304Du7SzcxkyGpTecSB9u0tEYrJnHlikUxB7JyYrbQGLAGEt0eyAzMae64RqRsO/Pnw9z6HO
pnxSIdCQdSV8XEoJqqXObu+mcr3I+J+v+WSalsYbKgxogETk7L8pIrCSeA8++vMOcbb6+X0p3uR8
8OiM+wSqKEw+TG66+c0JZrEmv5PeXozYlWL6QcnqxUcu2dzTMMjAgsY4h9DIYgwyxc/jcnXUzOOE
Jcv7+keJXY8aN3Kb0kq4SD/+Ma6YZ1ZVS6kbkCOZceIoXBvYDR+4uIpd5xTMgpzS2EVTgjDliZ+p
sFcWafc58pmVclr3I/rhDqrym+PwO8UU8WMNRs8NmCJyl7L/JeP3CnHMIYxZIC7I7OZUPjjtvzcJ
yCE46SoDGxL8MjH5BIyyVLj0Ql2G0LFsyJmwMqbxQNhbs7VFuSHFnUAsxEo+oheQFhBdy7Y9X+6v
f4zPUX25AftoZp5x4kR3Jno4/mTs9T00B1fwmNya7FYoOXRGroYNWdsLJ2iq7RXWtjShHtSSbzxT
MKI4wOs5SI7OOFQ+S8jFVXQGxDyv7lFwgVSj1LfIJEPX3+jdYug/QTe2EwllhYJgcy2qlrEZGZB3
lSQO0KpjOx3Mwy9L8AA4iGLxVgA2yJNYMaf/SH4gkCOGUVdayJGujAcRHQbJNfWHaNnpb9XlCSit
9nX5j5w55SwmcVq9ERTqJBMlBaApSZcaM38Vocs3aHg9dZJXHBxqbmhrtkAfAAjaPHpG4iUc0uuk
Fl60YRoSWIgz9ACj1knWZUisrwdoNM0IqkQ8YBUzFCAuugFvlKz4ZKuAVsXJ1xnZt9+aZ8d0SnaI
eTn59GnP90sbrBa0BrCHqGyMDdALQjCf2G1QKdmzA77T7OpNmiPNQmcITFg6D+/H1xm0fZ2zkmVl
jzMJQHekJJxjtpLIdF7RdFFdP5Uwhx3Is+zobFRH0M/4WhroCyuhAhbgidQi+y5b8KcTGJDs/c39
oVMFAUwerqvkKXKcwXiNEJm8eg/FV2RN9YFh5FwMTuj6knPaOh2pwFDNkuKpK0OS8GWwkDVf5Omq
q/Uklodxr6e0Kwy9ZwnoAn3PncIpqoDst23i2YanxB6/+feVUMilA74tFMSzAB/fHe2RGOkpQzRL
Tj6MiqaFpDW2CKLHA9aHJOp0jAWLkce6cokclZdpwEvwJoOIkKR08ACdztDyT3PHk7DVdsqdr7kI
+hzh5EW78BFM53IqBUhhKKIr8RspUd+6x1vEKEWlBizduJaThFlthnSVVPkpJlnR/Aa6KdOYA0Nh
tR+8MjvcnYKm1FSBjxmAsSHduXnSHTayPjLIathhqsZYQHrpj7EHssV5hOMVIG78m4pxBmdW2HXr
aBqxWaPRox8kCqQ4Oy66wu9Qc99qr8UhAnTGkWTxCayBDvK1KNpzEvQLp00g1fpuaBADZsi1ALwX
qwNxJxKujUCl2fJcxaJ8pMfCJWO6X6jSewdig/psJKKNAREmfh4NCS2a5WRa+n6LQEVcIKqyADh0
E28dmsVejvLLv6qoWPrXTPv+/0FGdiY0VMipInVSS+v4zEgeEtIkJO5CsysLd+mfAUtwcHFi8c4S
cTlPE9wRyZhbQGry2ghkGxKrLQO9r3wuT2Y3EFRzRqtvDmD9OimsWv5K32eKCzynq43UHBaPsm5v
uQDQpsE9eYBX/VTorrYm3s0iTh1SlYDFUFdD96F5x2a0HQnqO24VCL56GW8gsSSNtFz6zoNdAtI/
YzVyuWGCTVndBD2o3iXwcubjmNt97z9YSxDV1d+6oaRNB6NVvuJEhg4SQPD7hmHJqZFZQBHMX+Ve
eBXzpeJ56VCsUwoWjJ4VQeeeBuDAmXHzAzHelc5QXD8r2R5lbbvGcPj89ZtzVNY3idt0r5+ZnqOi
gBlbHX5qC57Bg2KTNKgQ7zBo/+XUBK30VWbwfvQmPrpXmTxa2iEOYxEgpp8acPVEbsJllRTYSprm
6VMn57GlrRz7wY+1xAmF87/h7SloATqeAN1C/nTBahjM0qbP6GLOoLKSGOB407KxxWumSkWOTe1Z
Knp2XUxRklED1gaN8/4c9HpRMvOg7UT08eqclp5BNMgZcDSTKOqtkn7VNH1TZzXoA8bUD2PqR8G2
p8zcPUY1KzvDc8v1V2kFdXUlV1IxyhqIQRgY3jJ03B0L9j5eETY9s6A7G4ZRJR+IGaNU1r/D1PXF
uuC/S/dvg5sN7i1NneYG2qr1NNb1abK6ZXCsKDbv2O6NqM5NYCM0dFIAExMHVtm5AUMLySZZlIOo
Zc1gK5MkAj+oUFfDRnEnJqV1lPi3ZsfvGPWBs8IP9ZfwZU9Dm9BW3qrg3O4ELy71uGJaFdriPK0+
0L+n3pEvuLQI0MJdYB5XZPb+aKRqSN7T4d5nylBGgjbhCwoi3uHLZHrHr6//Q8HbjEETxLb+mLDH
QeqGneXNnZ6E0v+zm7Jv8OXKTeNEDgD1LG/KqSK+jGbUEh9fJwlRUM2DoezVziWO1MnxcBAEpQeX
5qOe99x0CeHyDhHo9cYARUa+TgyO7OnxdveuDu8JStsThXNdHecRBP8fGXj/foHh1BRC8WZPMzgV
VABVMD0au3oNTJbGQUpS214CKAhbG6Rf17NbVseMR84+Dv414jxiC2/h5BdoekgA/cJpua1ULzts
FENHpHGEgMr9eraxVI0DcUr+OhIs0ua8iDJI0KfZkDmCMN45E12YcYodcYpDGo1T8w+SozIvcByC
e0wHlb5uJYWGySyoVVaXXG/divi9qSeSAZtMysXM5ddiZWvwKSIkuNxVGqaijdUAJEbeoQMghVRV
htnDdODTt35nbtHtIw1XSwmWBkz4tF1PMDGt9Vefk6KGdQMez4Vlh7fqPTQOnypddpq96ZtD0xH0
nnASZRBauxg8P0GsowSqNotFBSxvd7LjQDV57dAr8L5eLNU/tcxyE3UKTN4lg23RRIvkp/gBbUQK
MXSMF+myjWbpmBhDvSpH6K0hTK65XTBMHuu6hUyKx5x/MMoYI8bUfDP8ATp/MrVFsV41TZnLpbGy
SQpdDwwDlVQGmxm30ZjdMC1urkSSv49Pwd9vzbPMqKl+KgymQr9u4aSJHSEKF0iqKujMCo1oUdlx
RMODDaWmtG5exE2XwVGioA3v1WMvPKjshCYNospCGtu+recMP7CXyaad7vRRAvHgidAiaaW8qEJI
ZGksYZajy43mBCdv2X+5GMsRGHguRMNCQRNEPXtz9dyonr7DPGaGqMESCVun1mITEhznUZTNoh6q
/fqDnGFwDCBzeqrpA2p3BMmWeYoJleDuZp1FOfL2o9Avlnz6j3eAuXR9ja0IhXmmYsPWHS0MsFgY
i8zuT+pWdA2zBywZWKYcpzGcTUHq4b4wGb8RpETDwmJ7rerl4DjRpeEwxj0GfscPz9dyQyY7j4Bl
XFoW3NQBbU56I6jN6KuImK8KKreJVWnB0nqQrwbKaqmwFQqezwnJ/Yzi87Golc9GOkmNk7T1bzX+
pT8WO6eFD2KpY0e6/kZRKPO50Z/vmVfAM6Yfs76QW4BXoAABCCY41mQy2xTULgdjna/ju2EAVQZQ
WiaYoEHwCFnKX3t26rUjk0RKlrvPDaYxWxs7VXo/vvdfAvdcvlNdJXmDdn6Gtd37rru3G2hdbf2V
1Pm04lKi+jzKuNK5MjcL+LTdAMNBCI4PS1YgSIxeQWiloA7iHWdVhSEG5GnyDY3r1V3lzRmArkDy
dLZYH/FypJ8p9IRWdFDqvYYlVmY4BBwzcBxMFgFLnZpa4fT9fKMkodYgjk01sVrA9TVHpydZ3KUA
gw1KKYokNSZx0MXGSRcqqQopdZ0ZRJyP5DashQCvLGJQufBr2I2NYAsXQIhAprDgmxNOUp/iS5ws
TMrlxzXos6va+ZYq1aqC8Kar0r+cxFCwRw0VN5I10mKrVnN2TJgzDIkkbLVke3xEU+G2QKlKjKyx
bdx6Zjw6Lb6EVbPHpDCaN0O8yJOUsuok69L7hVnan1BIchwLRmGzZv3ejYLy4tLqpsjWZZ9vIlpE
ATm7mVGMSuUVd+ry2JU9OZU7qrDyl5FvF7zvP1+zUQDPKU2+pvNzlN+GGyVTRj2dzBaP+Z9lNPoP
CWtBK3QHU5b9TLS+vebasnkh6GrzVPgXDwU3Ka5Ani5+sZYXy+LtiyF3TnqVLHrp94KwhBRESSiA
/E1WqLUjiSO+iF1OklqlV157ZsQegvWiL9WS9gIRd3PM9JrpiWzNAru4sglq+9IlkH4EybOnEW75
2OpFG2SRvcbkw4lG3bWYdVoQyWrzD3g3LvL694L1ROEzUnzFVpQ+TqN5eQtjZB+svziPQyxIkB26
Ni5QunZ7wo2ZDQsbUGnog2PCF65FlVb+2ou4FyIbyF5rwoRwX+B8YbIX1miGIX9XRdlnsllhqHoW
k1rqVNkLtzBry9GbFEpoUgLVz2PER72zSrT01y39/gcOXGlRQnn/SQdx8Y3O6frfCIb4+Qh++d5H
O+2AFn9KfsIqUkoPS2tt4w8W2OAz3NkAcHPP/M1OpZo+f224w4Ws828d8RD7/YFiyRNxCzjG0f/3
ftmr/8W8sWvziECdoQ+VZ4iqt2fY/NSRn5l4oTZlh8ndumLhAItqT0kURVuP3AVK9SH8U/1+ZWRq
gJrhfd6mg4JuKbyELlZ3NdlnnXtqBxLUdTER0FNtwrdnn5VyWNc=
`pragma protect end_protected
