`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SwX/8e/VrS6Q2RZJEo7S02IgVvXbzQleMUnPDkl3hBfRwxgtun0z6fFjr2tNwr5p
W4TQAqga2UbrpELyI5+P0CfBxjqriXg5Y3IjuSMFUHw9jSclto9UiWHqQGRzhT2X
5MFGHDY1NqdSMYS5A4PSMFcapAZhRYwtsNhnIfcfPYk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3056)
Gai0I2wKNOaX73mp6SCM5VC5J0n+VCLi1oQK47nSJoqIkBcTupEpx/Mv+NJjhf+j
YMSREIrXw0d/H4cFaSIyjQFKdGDz+wlP8EKra//iayNQgeCYxlu9yIipugmKtZh7
VWQj6cRuZgOwT5TX789LVIa09ySRNe57h1CiwZxH1Lp6UN6w6P6yxyTtkwz0vQs9
/2nNB8PFv4L9NbgcL/WSP2tdH2Z4g2ibaEbmq0kX0yIBVvC/LgRuTCBJRqb2b6xH
N010tsYNPm/G4DFqynQMhkkU6Cs7DfWLQMjJLk+ITsjlVeCWlVoT5j104ccGArT3
Pj9YZ9Xz3EnYJlT5zI7TaJaZpGX0haYSnGFdSpEQNPiPpDuX4Wpp/EXHgc/t4Fxd
rWQE2EjpxIvY3qI10JQJCuBUzNfH4p9hXmY7do+FJxvUZC3MHX5N0y/EbYEbT69x
vcyl3p6k9LUUszdFugeWMB2cYJXiRB7iUheoWKfFwUl82PK9kUdCLH0a9dimzb3R
BpAMPqjYhcOnYRp6UZvIS86/J9BRgVp69SgaOr81RaZ2R5FX4gG7Ozn3ZT8um+8d
gPmYSnRvAbuOjKCFwDWHKFVYMRVur/v70pLtJ/zdNpeNE6S2/HZHTrZ3hMsdXyyx
UsItxK7a7zkxybv87TulK64ZuhXTVJbG6QsWjVu6K0ttpGwC6Yh1JBToNP0scSm/
3Tc5HOPOhu3n7fxA1QrgOLrZvdAZjF1gLj75w8gS6dOql6X51xNs5WsyXGbsv58z
PrhHsgtNuR5haXnWPfUKPGexlovUJLhWCWXeDhFv9/rD+5ChwIrhjbJK7jn0tjOZ
VsTbK+XtiLy9wiFT75nZIsbluiYjJBSkYJa7/4z9Ut4ZMv1j/mCwqxQkkaJqAJa2
0fs18geKMXm5FQIpTu5sSERt4Byk6ZruZqi3tisPgPYAojZ0DZHNFx+C7GypVLD/
8lMVpiISJhQN7Y2187KFeDgIcgrI+bKbPvsFxkbtse3rdxthOaYM1UuOqGByncvW
jGj5Gg+EN4zbD/i8s3k44tDmKLlZoVQ1FeVXzoHIAuv/xL+BXkDEfuKbi875GT+L
/+lNn5DbavklIb0cP7LTwpYmLmn8D7hUj+H0YQlDfVkA9x/H0yyU1r3upO/qrHyR
67+JGRF8Iicidgpc/8fBrYaxMQDHup7ImmweLjaUbPrkn2q7LFndt8pJ7bzsBX3Y
7xMiTD1SQCtw3OSMFuIFfxDV577uFlFGLdPM35mebA+RM3ilx5VpDUxlmhf2xVf1
c/q/TrKNk0YfKsIPnYw8v5/Wsvki/Aj+kcL1MoN6t6lfXXEy8TY97+KiCImqe76U
EFFiWGZhhQDiqAxFyFFIowN6oCkA28Ov3AWGg8BEOyUOqzTbI6JuXi89WTyvhHIV
4YrCwVIiNwS5uRzGtbcS38ug+p1Ae0K7I5qF0+YdNnidYrRzLiUKfNFjJoldcsr8
sL3fnzcYdiAkNX1hRekUIEK9QcJ5Prr+3sm9JSstpTadnBqUiB7ay4zCf7Mfr4Br
fofOSHr6FDahmuip/c8grgPSe6kFa88sXqc33C3OiCwksFbUnvAdKmyOgGElBYlv
NX4ojqrZUzHQz3t+a4+q9q9PPfONu1ZockatN8GEThRQkoO4+leamXvIE2jSek9k
SjGBEFd9IlFtkayvFSgGXZOVU+HH6nlPPaeDq1YlNu6fwt1oEONEzgH2nZuIiKwc
PWsPtf3PUnJBt6pt7vYXMBpMRBr6ZVO8WpV3xJM6FdtFpS/CJiAoXn+WHYf75BEd
A2/SsmssFHV9EviID13yBRbIW3+JSpEn84qDSH+MxQCWDg6elaugig3OnQ1VxZzi
hg7dBdKGXVtP3Cd3WiYhtmJ1Fe/zpceCTkUFb1iDNmYB8wYQN03fSt5hybfse14q
vAjjyyM1rW//PeDbguXQVxTAA6SNex5DmS7Gh0AvjyNeWqNjEuqIyC7xy64Sc1Hb
sRMYO0JLeRwMIS3DqFtiyR3prb6UAfioGKG5vsGQrzwSAE2yTMrp/xki+R4Nb6dy
zuNYulnvyN0DANWuCN755wgcXYZI6aH31JnLhPnnNFcBxCWQpreJgU3zctrqJBrG
STUDQR8H5dkCMTLDppe2CyMb+x++5Xo4LXsvfvHvbUD0+erVZPzRiESMX0h5/nug
ZwxhlGQFFsdc+j63ASAl/HgXJCujjjTeEfZwHF69YYYR/xVq41oO2lmJwEMslc3n
hw4qSZANsdguRI2WPB00WYSmaxbKo0Z6PteetOfIUaZ9bA5yC1MSPgSDIMziGoEB
FjRCS0gVgSbi6nuwLE9odtGLXoNRzI/5Fg3FLJ6hN05Q0eOUtHm4zJekybg0cemj
LuSgIfws/07Iskuo71AvGoWUHZeyWE86Hk4RqSMt0ISLAlm3W9RRW+p0g6Ok/Xhd
OXuMAv1/SxJvIMW8ktaJfho3qvjNCCHNtKugVpOh73M2wj2fgEfGuAXiMO+a1yFj
x74h0pGB4xeTnz5cNUdrIBCohDGfGGgSwQfa3yGdAcEwKTiN7hW7dAzUJuXu9FQx
F2m44QoqR2dl3iP963qLaPD/ArfvObCtbe6g3ofFeEqsrZYn+StsV1vnIITlwBN+
+5RQwf56MWZ35ewI8yFNs+haks0KYx6SRKqlRE7lIjqZT2AIg56wZyUqQ7Ozbmgm
eX31uQbzMPStAx6qGWKeQqwEWmCnpPLYWPqY3M09VvQHBNedBLvQaO0pdnZKdmNT
n1Btpmx1wod7UQhmI0vRRjpNzKOUryN36Mamybz6ps8q8mk0w4lvrieIo3R3TXoM
9gG0w5n7KhrkypBvn6wLzLG5pCTS/qUN6fvUNUymPSIH2vVW1Ofx0vDQ57oe65Hd
1U67ko91rT/Ymyah15YrhwAarDryAhzLOWM53jaAer/55hJQVUbcxKPOu0lKzenN
RZSHBewHudbuM7BJ6Azcxm7UjbbcWNdR5T7/aOJ9gx1nyNUcubvmxlktDL3F43LL
o/l5arf4s4TBa4V051oCBDmqqZ0ctzZiW9RT/LmCB1pH2aFclSm4XhhcGrafWDfc
g1adKICddHKs3WrGRj4bygG+k1uJv/ZTfw5LLAmHNkUanUFjyxn27MA6ublOW2UE
598zAhwigDE7BoYpt4qeT4ExlYIMEWBDTH7eLTsCphsmgBN6VGHDOTokvSHd0Qcn
9Xg+3e1lY406APMxTMUVUrl6IhH8hPYIN6890tEKorzu/X0yiplDrUo2X7VPWtkl
MQ0OAcRUa1LSneIO/tOWynIqP1CVoVUKvIPbUUbYoyJEZiPNtet3vArLmKigt4lb
yibPM8C6DNcdqpaF90/R0ro3coXiUfcOLZFB2aLcDVpRGdZIiCtV2/llkcGuH1As
w3JCVjx5kvvpqxZphNfnx179N0cMfiiyqhQ/9sVs+W6trAJNoC3SYTdSli5fsnTv
nEdaJVeKKzPuuCStQkYmcrmyZTjxZRF+tZ8gFqtT4EO79s1LxNXBnB6DpedRwV/1
qCo4ZgSEFzsxe+Fq776VaoGAzYTHoFjSBoe3p/ao+vr5rusltCs5/hi+dRsqeBA0
p5Y1HZB3jl8CTNHIxQca+ncIoZhXI40+3ST6REyJv1ty7/egz93+/f+qeytkIUCC
w3QnynriSXv/2pQteQzWfIFBnOMR9JKEd7WMrS6tSh9qvPSF/V87Y0ok8K7e5Z7p
C1YWkXIhIk9c5nHvuCyGL5OwGiRQGYO7MKiYx6NYuEdK+sRKVh7dHMfzKsvKvK5u
VzNF+zzbkNY5c5yfvr5tLKCW7L1kcoJNUwuSXLSMHVu3QnDr0G9UZySbsCDYroh+
L6qL98j90LCZrbkSgE3kau4v+UUQLmWb9md2KUG9MvcRGKQRul8hxgZVH8OeSoBd
k5tOFkh4yIwMU2OfN5v21il3fVLwjwBcdT2N9sRT0U5CClloS4JCIecYBy/OD43C
t+OVrKdyqBqTw3EP6kCawmJMvjUtG9HWZO6/ufcPdYm+iSiZo9pakObDeCFBvsuo
AjDRmRmrabopAw8/5yWeIZzkJp6dasYc6khmgyCQtfI=
`pragma protect end_protected
