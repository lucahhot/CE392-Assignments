// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
0JxEXD13B87hICW/huXPep3ZkzX2WsxEbvesqc9cULET315LdJmqCuhkcxlgWcQOd2WhS/MhdbSa
CS/7JXR8zWBkSoj6+RP/0eE/cuveTjaraCELe3Zuy5c/WGUWR2yoOJR4F1aHfcHAvJbOr9gRnG9s
8rR87TBa1IJ0FsVIYM4SDF5rmaDQjHFBSILzFJ75s60mJgslr4RYRF8U3PEpn9z6l96yoHgHD3+e
CwPDXpcZQowH4cCMMH1/9KxmD+pu5lmohHo2UTiHR4cYovaA+alOudBmzM/tV8KBQtA6LchVzrMi
BKKZ094xWPDQn6U2ubx5x/2dqvmjCJ+LYRh65A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 26656)
uE1C36A4g7q3+FzeNGbVM+peAFwrIQ2uQ5ATMtf4i1lE/uiuaP+SaLOI/l7VKfa+e3XMMZ/N3WRE
f9s5AB0+Tc9x/z3j38JwZjgp7dZES5NfgTlp8u7SZ5ZgKYSVP12JRePpPlnaEfPbNoutOZMgPDJH
O3/VjyrTJBSORV5RHtMNtlW9UXSNs+ZQtFgAWNXQrb4QLFcoD2QqBGvnMUzC3Y8rpvA4iUOyEeD4
KlNqyoLbcNuOSLHUpdAxnymxcWSYxpSpg7aAQjj9cIu7ylXjQnDPjFpU8zV8rqEYhweCSxUIzPst
A3YJ35pIWISpR55AP0ndRCMn/gKpxT4MhV8EPwXINEpro+y4I2b2PM370n5tUrBbhTeryXw0ydh1
CuZ+Qt4h0gtqY2imodQOLwF6yJBgaZZfRW49WmEJ8DDz058YFIh5YnSTghuxBO1miinLNwoZ/w28
Gpb6fv0uuhWXIm0yGgjkYrNjY23jTl+D96gxXQ4LCDVORMMyKH8aSYC0m5+yqiBXaZaXdVamc8/W
jjui6MSjKCs49z65nhbXa4Tb8pir1JDWs7FYeRjZ+HmELiULEHOXIRYxz656WNWC38KsMTHESTeu
nC1m20JnRpRnwFRh905xVqlpPcIvrdPCgpLXwD82DRUTnBDs/XB6mxlPHgIOdoQ2y3V7U8vLoIVG
sG6isxuJc95DHpVHqaK7JJG4B8VGEa2qsWGUyywlHXEzFUkCGBIzCI0WiGFc3Ne1DlErH0nS+H7a
JiCK5aVxrgKn08+dXmKxyEoX1q01BwOy+ffUzBeig2mxzPoj5F2O06SLea98o8KjWTRCMCPSEY1u
+kEBgYxMgwRN+Q/6w293zscvL/QcQ6tPApzCYCA1ML8DagUjfLAkV4c+ERDvd88vR6DEQ+zCwN1l
uIWw77YPCW3PhshWq1HuXjtRxiv6DY9I2tRrpjVf/6+O8fDChUILt7My7O5XvFknaZXNvJ0MAqRE
xcq9p1Wu6uvzRiXJOoCYbIQ8E9Pel1WCW35NQZMxAQypFY/JwWDLz1sV1FhSXHjXyheuIRzfNVYu
kPCOeteWoUae7IwEWBS16ULtFCnBmB2gDuTddcuaUxsF/y/N2EliHDxIOhEWu4EqkV2M8yJQ/rJ9
ZwMkyVrx78lxJntzZLcr52VvGKewE64wFe5wHkKsuqRMt61AhssBvToOw7K9Zb2P8xdas6zZ2cJi
CO2MeRvth3cMbKqXm7B6pDtk+O3lS/arUHQKvXvORkY49AETQM+x5s1jtEon5ZlXYNCrHH/sWlEn
VM0+2VnO9my/5EdcBiBK98cRWWV38nmnLlz9KWm1ONwQh56YUXSdF531XWL13rcGLFaD6AbjQ5ap
VHw/7zuPY4Gx4RuFirPRmPNidfuq+GWIOoopqBv9WoITIKRfX4xbHPsgkwSEDOVb3oZGc0vdqqSE
YoCIYbDWGaavkpVnRA/b/ofi961HHBXjd7dmH9/mAiRdQH5z1AgAjajnhjYYdZeu1qAuaRNNMSNN
5UfDoMVo5CIyfUq6/TYLVuuGu/6tByjjKzTqEBhhLamtFJyW34AwaRUDmSzEB2CqWZiqrf+Objiq
ztIJJ7jnkmc+FDPStK2KjxOAvjavhoM34yrCQ2kZGO2DI3Pz0HXQ8nfQ0VsPUcMXlZa5+uWjwqBv
NGPxFBSUyceJQ1LTpw1ZPa5leG4rcIzR/sVN8SjhAl87w5HSeksUdcKLSuqVVYxFMDFh8MUWOlYP
CgNG1h8Jz61gMbAvAeBClORjF63ByG85a9GfUKO3ats7KHs1PeFty7fuWIVUXSE9DqZGr4VXZ0vX
7uLgF75ANc5gRvMgsuLwvGXKnm1/55USvCJ1PjduRstG2J/5g07r+WfLVKgwSZqs/ZnhcNTm1zz8
ro+7SVOOFFyJQ10EQ6FKCXc8FLxxoQjrFnadC5FK7ASkyDZ84XNS0/DwCqzWlqnM3Up3wMtlgRiJ
R0zSkEZUqO+OiYoLLfHrLXh4sLDmkDMor2WFchh88Pd3qWaQDa+fADtGT5DMX5ZURZtrwJlKobqm
5aMoOXAJz/7faxjDSRXZI8BYeiQAPpJWZ9iHN0KCEaiqeSMeNG6ImTamesSbWqNQ2DAlAFrM1Trs
LnJG31lWs4RnVubXktUGUks3zzTvdhXaQMGv94T79aT2aV6uzKd2RI6vLsxJEvG/Pe0dht/XLc09
foiqZLcyXVXiWAoPoTY90mtBZqsySjzwVL9r09t96qamWWwW1ZT7wyiA5xTQD6KsH57cnGHVaTX4
Y5q9Njn37GxCMv+1TqZAk/Pd6w1UAbkQzJ/6rNrCtwUBZFp38tQ185UAXYzOhBJtHIiDPq9bno1u
PYJmmuA2H+pUnBXIuJ+0HgBctXyXA5cEwEuzKXqUUZp2iv2efP/Qd5Bk/hnJBnPNUUaumPQsuBEx
GuN8wUt6+/0+c7Gtw0mKuv/35T4FA75SkmhxVoyoVBPBqpIKbVpxcfI76pwu24zrgieuFWPuDHCr
TqMZhPn+eBw+uLdLvYL++q7DXyN9pQT3w12lmSbEhmCuIvwyq4CUxrSnBHGMGGuXx45xP9kX+AiQ
AUDDcVLVSziN8v4wNq5z5q+QF6yxHumXiqUuf9mvCdp+mxSTChMnQ0ZciCDaGE2flNEVodHwKhQu
CgkUCqKu1g8bdK3xfo7JxcN6yXJGTKFA35I5uUzvloGvfRv9D4SEtbapjQ5IZ/rSGRYP/7FkL2ik
2801aAxZGXEjFDE/DxJ0lhMIa9i1l5VySHhPHbyw7ybOxbxH9COI9gKnm0SRfJftxxM+DBZ8PD1L
j9xPd7NlFEJ5XUqlqpSqJSlA+Km4JcxCbo0da5n23qKaOA5fsltgbQh6VmFc2dlp47pZR5YSDzXk
J91+XVCExuPdIo8lPIZxEfcA1AM5fm06xNNc/EcFi087701IZ8QCPTa4GvX4yCv7GNa3e6aQYPNf
kkECQQJcMYDzNd+TfEeSS2VSrkxV0ccEsGJ2QpMTFLqCuzOWLu74yoUQvXYdZGnG8/o6x/ZjWbKR
GJYHmQyGcP+gNGzmthbHaLQyuwsaQH6YdlmSaAg5+4QHs6je3nQ/nZBlD56ov6rY97A2kwIR8cYa
88ngBpAMMi9p9aIT+2+9Z4wzAAdoyTsnkgYlnlCeP1uW96WTPzJyPjgFdHci1RzinT3hvQSunlhF
WMKAGFYEE1Z5cpvNfYRwDISeXHXrsjJDc39CMPJ25kP4l4EsZ0nVcvuvlVhxl0MIqpBAQplRGpvn
8+afBat46Gclvq4hitBckD4JjSqhFWiQCwxBxSreUoXi0SoYGVv0yVnLcCZcpdAGHj5lATQFmTre
BoSluPyBwlEZU0CXRVLT7viA+m2Wrod9pNGgWPrCHgiMg7N7J7KckyaIY3o3lCGgaaU8P9xtfwYA
h5zwMl4jyfg7HTUwuXMRrK4/LWq64PHfzbE+om2I3s3g7STQUwTYpEM7JmtvD+AS0Csj11+CQe9K
on8Zv6BHCAK0hYo7H5JdZRDq+uKvohkextpgTPasi56yURZgE0OlQB3f1oFPMmR3sSZ6SgDsjPhm
Swec5BM96B9vR1kDoC/qa04iEpklFPtqMJikgY80lGhVJuqzkBUQjtTk9nHEclK8kgBn5HXGG1lg
NwJ0wAm8DzjUeQJ68y+vZbpJxSFi4+e71CoFSWPew97ARdJCyAzC/8BGwkkZce9C6Xi8Q2H3OoNV
PJLa6m3BSANah2ALqtS1ArDgWhpHF0dZnr6sDbGf0QTZc7kvYWpohzygYehMPnmWSHXaOV4dPruR
wXIlHnfmXJoCATCcND6vdZ+SG14xUgXpVU5O+zeiLkpKroI5aFow42j63Wm1LPGv4oA206bHnnpI
NlJ231KvFS25wO4W4R/s33ukbdqf1s8VfKukG26rq+0URFneLwgqM28lqOGI69xfjBY3hblpMkJs
rwHBT/NwqpZlEgEFtDRvRH+IDw8ciXUFooSxIXJ7NFkSwvHQkV654SbaTgCx8/Wms0Q/9+XrXNiE
/hcaI1UXaYP38PccRCDa7Q07qpUmLU3usyfXVNw6vGw2eEx6if62gcIVVHQ7rFwgSggWxXCUaTYj
dqdf+TCWPc6fu8j//V9A0piKBGwSjpdlPJmZdkwqvG1dPt/2lJU9Gw4x6LvAoRc2Q/ckVBq7CBu8
xjZYME2PFTOLzCCeRQ8O6Mqd+v8EdE1rB111Hki2PdP475tKAluFopE8SbCtTq+b9cAdQQxYyr/r
XzQdRjNLIdFBdT8FiBv7dBqEiN1uw3slKqwZcW40mH3pUPlhtM/y+QlBnV1AMG7efFm3w8KuOhlb
qpVnjwklIwIgSW5dNISLC/0kUusSpFae6IdFZLyely4Eo4Y3DIeJV5yBLbQr4nTAA/IyRdVExark
0tZVsR35Rr9P+w/6o4AFllGG834+EGdjMEv7wtM2SiyWqt3/AtNnII+9DQgukXPpBjBt7xQyCJEV
vDL0dhBnX56XAy29g+aBlXd1xxRiRdKC8/ih54wbawizZuFyzixeT5aPfgkcorJAvTvsA6K2dN/3
A6KQsoHXAKVN/8jL6onwZVYAhLQ/SfMSyOJbjafZwRFZx0QcoieXtquAPuWhgDyH73Es5QpNKapY
sjL0sOdis2YyhtthPd7OP3rOKpwooHPRvGjGMW0FRGxvb8XgB8+OAtqC99OZ2C5jQu3Bmz8bvqO4
6LNnAeWoee3d63Zd4GB2ozM3PKge6pSneGNcOykx0YgrPrI+g3W1UIBOpigg3NxC6HvIx+WUSGea
WgxW6OqABi4vC53cl+1jLqC2RJ5hoDF0XAzATKSupTsERzSRS4ieK0wAE6e6XW2D/T82RyFsDdN5
w4pO2XeFSV41cP+O843puak4qG1e9wzvUBlHwVsN8WI7noxpF7KpJgC19uNT6Bw2czI1pLiu+B5e
TFUtk3aJFiRYlniOmMmkIfSn7xBQa8OoWOiwc8KSiHqV79hjMHQnhqwUhh9lB+cw3rHoNj7aNUct
d5dB1b2T0ddwoly7Bg4O49ZJKhPcS8zVwtRxxX0+4WWwaOlDvEVh3/kPHduAo14NLy+76IzdUmwZ
DFtibWOG7Ft38AHpeMM6ykdekNsrsSVdvpbd5y5oZphg3tLmj9Zvz/T0koOuB87OPpSz4bIbJlXI
bRMoqmL8l1P1tSWOUIqguX09npBME++Aq9xqoLWDOFigrmFAEXY0T6B14cVbi+LUk0VznGrbo1PX
blF4bfBrLeL40A5tQl9xiT8CpqqCgJ5LqTNtIB04rpPxxuL7pcCD7Q/L7MajAjTmBNCQnI+gKtlC
MkQ50sO89Xg+fA4vnfkRWG30Xg2wafV/HRT6cmKdqiE/aLCGAbDRe9i8KneSA2rnHx7vzApGDEWK
Cpq3gVETzAeDdKOUBURoZZXByC68Zke9WicDUtCNDRfKkFiVmCf9JWWvdmkiySt5JKOG7of3Y9+h
QHnquV0WtiVDFU8bv8J4cqtQRI+1nmNBGoK0K3hHZZSa0uMR/IKxHJGX0QGgLW70cUkwTIBjTH5/
xgWwsy5boZoLR6zVMUEuueOI030A3Pk2JNscUefwCTdmU8iNdJPdrzahtQ5wX5a/U+UGcZzcQesl
kY8WFw+iwAnudemOYLNKeum9lBmBtwcVxFZVg7Cs+BAQavrLscmXjlFeEp9vz3yMuN64U7zi6XJd
y00U4UtVjR4BG/PLx2VoGqgqhPybLjeStThLMCJE25khdUhVdZtorw8Ktt49K2VoIvjPNHgzWXf0
IU84t0Npe/8NV+l0+cXBT3KMg82XjmJoKHc/Ve+NVVjfSJVgjCTBehO04ir3Pi7QhbkPmnbpOvN8
MPtqBsyjFfalZgHt9EyBrxojDIwCPDvvn0qMdKbQgcuYsN9busDriELDMfSxwpR7mCSus5qT6DLW
c2Rh581I7/1qWYkk8oKHHw+DNuYri1iA2fTzrl9H0cMbV6nmSL9BBMjFYRaSrDEgMK52r/dGaalt
P7rjftPmCgkAnblgEOZfwQTvxzXcGuTil9gO6Ow6hxXjCtnWEijzeFhxJwGku44R0ukprSVNCrdH
lBM1bOVlZ7c6M3QOUMHPk/3Aet08AwfDiB5XDc7O23Vc1Tm3iSK+59feZkVaKAVwy797Zr5rN6F8
V6HfzZViYFZM72eMUIdhotOUcmE/ac+Oi3x4LsJ2HiC4uqArkXT9zuiYAruxnjePtTTF911PBGWi
YSuwGtZoqZX64qP7ox0NRyOxa68sMYzJYeUL1dfYFoO6X340sjXoyXHOnufnDXVqFcJq0FatepKq
0g7h6GAAw0WiGl2+j2dOhe2y7LoEoeqicH7Hi4mf8Yt1PuvkgYSln+VQ0djupZ4cPLdyCj+Y67jl
00lhm4sQEcxw46cI/GkEgJgAGDEr50ydvpE6rX342boSHJElq0fa8/UdNZO9CflKuvc0kHHHiYZ1
O6JXA1kd+5+cGtqJcSWxPKTSWmnsm3nqZO610DzcFqtW0YCuF9Ic3bT0ZY6JK/HbrqkwIHjk4RQ4
gUFJ8RuaWcZ141ESEA5SiasqB08QWa3/KJVsTwLcHDgitnJ3xZsbtP3uYAFUzy2maFGouqAjn4No
VhE0xzH3EJlnwIjeXUmz7j4P0eGtpi7EuvImQz08deHj8ibIbLe5YmDcIdbxkT8Miq0vAYXpidwC
K90xNC1PIL0OQ9BmWQp7BSWFPNTOUpRKKY852wFotaZgtqAqJgfKJSqwcCTqtJfUYDp66uQny6AP
oTNfYaeT3jtcljT6Slc0vh1UZ4wy1UOnAE5HbIxs2vTUsVlPZAa05F0NIGQM8D6nI6+nW9BbZCMO
MeOiGt/JlvOmoidOuh9N4jN3HSc2XedgB/w9w7619niCleIoxZl0JMPEYYWnMqprUiRoNQsf/0jG
AyHDww+Pax2biVdb1ipsUnbv3KGRozagLZJnrvvs9Kf/PtEiSOj9g3bdVsgG2IYuW1IzzagONmeF
dqM5zlzUEAXqJy+Qo3GqDG8Rjb2A69xele5Fbp6ifx3xjz1PWCwK+KGhnV+7zeM3GGQ90eJHlgNL
hY+6UNz9o9zkT6RortNtt2K66mAJIwEBLabDelR7wA381PTo8HvFsnKCQ3hFTcxNcAETYgPdOlzC
FNcleqnU2iy/IHJmTc0ZFQ8vqXoYH8uMZcIdjl1qKNXCkMEz25eVYz6I7g+mLeLEcJ+dAyhJelxn
qbU1sPkBrvzQNQ7VrXHxU2f1DJpu+fmBMLED71awZ1KflA4qwTJKiBSas9I9+Tbq1lwEVBG35Fck
xaMB8PyVf4MfWzzwP712xVkSYG+jxA3F2iPEXR1iaXSBLzL3g3XP8D/+J+aHDPZ0kn35QIr4W8RI
2pJZYj3W24lZXJd3283zwAxbqWxX6U7S9asXLoOqzdzxOZLKcBUWdX8CTyGNHg5BK++Gtq5iGi+U
oYX+OI0SRtkdu4Ls2HlVjHhf2Z8ftiBXJUMmk5+FnBKpYGyVyIAoMICG1yZw+3PM9k4mImn1jDjM
qiRxavAKueb9BdghD1eyOT4ehJz9ZeVFo7CR2UtOb2K13rUIgOj9Vh7HuYbGQX7pCt2FGvMAoyKy
G99/Bx0zSyom0dkkRzCyP/fhRDcNQIYtkN2gmt27zv57rTXGnslRD7KyGwzCaRBl5SonxDbtyrzc
tuuijgbWHBf16u/fWWYTq6WLmlmrh+OTC0CIzsGqdC33P3bH1HFykHGLtQIgw6VHb6rxmScFywBC
++cRKoSVDLi2y9GnSAaefn48jjMttdMMRaqp4fPDyQUY8F90OipjDkcKaRr3W7dUMbfwqPAQ5Ajg
tk3UnBTA4Rwji7Ymxup3Uc4a8XBfcELFtMfPE4eubpypobZAaWU6uLkVfm6gk6b97g4qorEDkop8
h4RyecMVyDl85wz0i5DuedeWRRs0j2mF1kMEJvFkfTxH0RdCxM6feZdEtouL3up68O93gnUZu3Cq
Buv4aKwBtxAZb7p+IQgSsR58atCx5MfYX2BXMlvUEIh1T5zz5CDUDlv7Pkq8uowqvvk06XjzvSXd
dstGL3TZ8qJ7cWMfjK75g7Vn28nxeRxFbDGzSB8MCDJ7k+ahW0Ot1F+rJAOi5R4vlyYoS1FNQ8b2
90EPtfmhyvRMoPtwuUWFDjg5Zm4PcUIZYLEeFEkhZPuZUq32GwI9YLCoT/fbmvyN7Fap/CPlTfEo
8AjotPzi7DRqhKBf2jJ7hXe+77+TnC5SNS8t5lHM4V+q5lxbsUrRMOsDhnx5RMgaz7dwXiGy4N0z
LLldRsPMuMMn8oYAidTyJZo1FqS/xzNvZf4Gnr9Qnfh+yqS6tlkUqqDkRw9LcoDv7vmjZ1u0qTnl
ncOw23qOR/MWYSS2dB8yi6D1O7aevHzZ1JFZPSNavL0b7L57wo++X37/hz8G8SO/7yptE+5qqipt
SnDyvyaH7Ycit88wAEIjcriZhMnZAgGTPKtayzx/naXRVqJ/xAx2O6Ye7ciPrwXB0a9k/2bUPoJI
bpc+AJFUD9Ric4DYWrBUuqoQQuY1dtSqGbZOkAKGU54Sr7RLWiK5fXLm4BYmg1RFtGs4PbHH7iTe
DzaN3E1vbk0iukDaEM9fm7jalh60N94/CYygY+gDPhcG9CkxQfRAUMO4cZ9ooqbHI9NURVVfbJ8b
Fz8MUpgUY94mc1feardc8YkiICWVgPXyPkTXglK5frwQ8oWo3apizCRkpI9O2RPf5DjJzyFLm7IX
JTNfVSnOhxIz16clCJvHRJCIhYhLhW9Wdms/RAwpK7RVwumugmkAkXrlS6MkZ7FuMWeerhq4ihxx
5V+wEKT+UwFcbiE29sKmNpzTlbOlS38HU4Wb3FN8YZkjkH+BkXsdjysd8vR+FFjmfIUlRZQJtslj
lRr23uWkZzixAhXHkX1uS4jOX8s5BuYuaGe5Xe4ZZ8FsUQn12jP8dSdw7s7opDT14qg9un2UqXyI
SKCaOFc+WzAgX0azIPu1sy1pipYWyKXUugd80vt+WvdINVJR9rgGP/nR1qG2WShf5q+Cy0VMjQ9H
MI8PHux6rYJi/rQMpsHlWP+/qEToyRP5mTyRcaXGZiLJVoC9+XG96A4RxjuiSA30pqlFzu2wtZFG
8GmRmPPruDh1eTNSc18NZd1vMoim7iG/hTmt4mGD7zr3bYodjYKztK+I2SSsxXHIyWZqKf9m2wA6
J+cZakrzae3d+RdCZlajkNoINdGnjFtBMxU9BhXF2SYjhNt0kjfeJVDO3nSQukc/HYXXYE5HyL/N
icKYz1vt/maMyT1rH/0+K77fM5pfUt3a3PdXSeYSsEkZ0F+cTXo535DR76M2pcY4MQ7lu8GmNSJb
V6wR07/qU0bYBCfBvyd4Kahdp3XD1mhXHyDu+CAjdsmkLZ5IYDGvhAa9LzHMy9fQteDmGQL6OEs6
tfulpt+ZSR8ccZ2yTfCXV4v7ZrN1QsGhMceEUOryvoMjQTr6TLT+5FVCFK3fB8SE/cIKv1Tmfooh
9yeXPRqsoweprjByMc8PX/9LMEK5LD/+OWerttDzUSZhlalPgFQQq8OdQ5FfiCPbFrI14vRncRfP
H4qusM36VQFbnYS8oALyCezWqBWCNYT4qTpSw0u8/05qbastF2PDXOUmRbHA5NGUlAnoWsigCwUR
RHGr8A2OzzTQryR3uJoD/E5AtA05u+PssOMqhMIstDr70KZg9IsOsgo/M02gffVSB8AINtCdGDli
hKfcXUL+8gx3ERDj7FdPxuVMc1OOPFOb7Wz8FaBRIgEmr/iocs13Yh8w9I8QYXztsmWNW+rsZCRL
yRja83qM4IeMdlIHeh/OGXg1kwdbBrMZWEqUTxN1iQsljdIf4bSVUWKNn1tWZV0RehTqh7K5nP85
CrRiE3c4nuYKXHgmpjUWqwkrtvQkbd5IFznzUiJFKD2JVRqKOJW9UFNs8fO64BQ+fmBMiqZdkW6V
5iPtPr8ops7qb6SB4n4KygnjCDJJ68TQj+3Y8SvjZIruIIcpNIetJNlvNpps9Z14Yxz0yzzWTwcZ
Edu2EWFdHVaRVzzJmhcgy0EZcZTRD5qo3JaLBKw0eeqjrjGqw8IM8DivUDGMxu1aZW1BmOBb5v+7
9ggyKhVeqsEOCl8RrZE/7M/MUWiXa+G9p1EEFbCI1TkgjCYQG2dm6TqDIX2T4HO0TxZB80QlGFq3
jfaNIZ72crq5Ourxcu+0VxLqzwPfDc5LsxwIMjCi/ULX0GNa5dshMu7r7HEOqBZRfi0LK+sKpfGq
tpEOdF6JNh65mIaXBZ+oNHlDCKzfRAvxKgtSUWydgDmrDBCniyJH/gQ1+siq+cmVgqLc8u/SCL96
1kg0a/3DcLQt/YDwvVH+hSANcYtKCLorThqCo7EfuTxoPWQLxdpK+vVCbuwZXuk2KSk17vsPfx7T
ZoCFh60J/Co4vpKeBqCzZBUzeO7jX5cNbPPkaK9Sq6G7BfAOLRShop2rqpVo7Q4zRIa+a3pg2uuF
xPpBaiEgYbKlsezV3ZQZcbM+MyZGJQfSrKfkpdb40cAlWMNBHOV4pHc9aN1k/3S+sgpucjB/DGhj
9g0KWkP6LGtfiUjODzaj5K9XIZzBErR2g5yaYusR6/2XfiZEpSWQz/kOnwOUyucLK4M4k7AgJa/i
00YD5ccitaUm7Skm7L0+9EII/ABTPO3Vz7xKT+N4hHxgmpXV8GeOwONqJUmkndrUWFLWa4cV2W17
Kee6zi6h3cKCXT3ZECNmVR9Z7k2CRVLq0wu//n7LZ09UUG5PDV9ZExGQanIfGSH/5NKyhfcjM3Zq
iJCEabWNOiJ53vFZ8EyUFwpx8ZO83Wq/YecHn43RNmbep2ZgyzYv4SeVbuiM9g5vZ2vKU6+eWwJL
JuV27cCAaIGRcS8FKehUA6hwPS87KfmLfEIC4arMF11+fxaRCmXKqmAuBSRtfx/FpT8qCgbmpoYL
nvFZ+eCh+462VZBtOb6YqlycjfLkv1shcEI9Z8QaERsjtvyG2A4Ez9v/yHPt3aq+LA4qrp1ZX2Rs
bfo78u0aR6hTbXdxSwpHXYEDQjZiVgGSX/Beib4JDKgdJNFGPRvOCcL9P8Zx9tDbUGkh8SfPcH+j
5QMzJJigjA+cclCGoK82FBO1BlLiMXDnfA+EjOJBh7KDc5KF1vywC63kpa/OCpdLBcrFxEZN1HnI
f35ujhwrYcF3WC9oJS8OMcenYwkQMv4OIEn+PN5kczSeRc0x9wVLxWVBmuhnzCQhzjrZ3vLYTSQL
aZPml4Rb1RB1dOxXROrlZYuk/YHPbXGBkNKIKFgiuPQojVZoBkKY6FoeKXh/tZav/4zYoxRKcn9u
Go5CCY7yjFmwBilBo7pwmZgFTMx5gtEUvi3uxrNYWkgXd4Yhz2dkbP7gsHFLa9gisABvxz07ohi6
r5EcNLHBpSXTL/3CHc1BZNrJOvqItgMdoILFrzb7h/Re6lKa2ld5cmJUv4M7Dl3i76wgUbIOe7vA
sCuZ7HbKfBkIYPCUEkGzblMI2Ya5D3bJ/RIGJabrGuKgPhTdol1SaHaht6bVu8ikBZvT1ZkSKyu8
Gks+4ktsgRvhpv+F4M5ni4bSiQO2HqAmBYhxsF2K+9CagdS2Do1r6WrhksRSoxO5i3pnBy1jYNMn
NMgxdF3b02Fm9LSXnvuw44DSrvn65wjE2dUI6C9P31u3xaQVhGqXcwPDKfcst0qGWkk50s3Z3tUP
7T8HX2hILu6B+wcLRMcv0XhPsNJP9xWjz6b2wZvoLq57yr+ezczzSw4g6MQ3L8ETVqNwvfcYrsEo
imnpNVrOeeuAtX4JQj+dJ5RvpgddwN9gUMFuvDrLQGEu2/E7BkqN6WlvEiR7zzKczpA44beR1xoL
3ktsaa54/4KKVHMmn8LdMjy4bLzdn6nsH9yzxckSdvABIAB8PJX9xtsgIHss2Ynk6p3WqMMjgsEU
wSX/BlIBZxXINmDWqZinFgl24OUvZF+g7odriBYA8v1EcDSeWDA2vvaIlyD0N8Mwz4JHEefZDL+2
3ADOCufyXYFQmj66Bh56Cfi8rpgiy6Lb4v1sMBQK9tJfA9UBSR67ulZaVjr2KZp92cB6vWxvvd3E
13kBu1EqayF6sCHalUpuWjyhIh0VkEY25/RuJXk9sej4bor2hrxF2kP/0o8P/FGhS4uqBbspAr/g
T+2EScFZi9+ZfJ3Y9fctzgAUT2s25ilZ+GMhybTk6OMR0dbsl3hcs9IUhPx+GYJTZRBxdaFflmQe
Yp0S4CQLbZi9scvMEacAmLgXw/0jAM0eagKlCfgUqgPGEXacW+bwMJWf9YLGov48QWvLALEx8Ha2
6NvbPDrQqVpWNyqGfY+u74ctH6IkGtOhOh32ZHzLViVWPobyJY/WkBmMFvJxzOwMYoj52g9oax1v
kA3d6kH2bSp25rTTDAvPi4PS1JSaKe0rbltOLiz7xtgFhHE33xDO1jKxz0IqS1FlHgKWn+8uBwvw
Byr/3kx4xwJvY+HKAlY4oBgeG0iaEnw+v56a7Vfj0HuxxfeDb/6sYpOm5TFbTSLcvDsA+AL5FV1m
IcEOElPPYtPCCIvw6ZuN/BGT/9mbsBfQqOZS3KWTDkXOlvsqgxRThG1TPhPXn3GtUTH9J6PeaWb0
b4UmLGXb0Xco851N62tmH94XOZ2bPUhOA46HXd7nJqSdNXflxG1L221+E/GmLSH2mka4w1T4PgCK
CDTvhX5c7i2OuSV+Zk6CltBDCNvmMH0rq8loV+EcnQE08leQLjYGhUpCO+4CPna5Yq9xHdx8MZWh
3LZmGBePH2chSd2YhY2FLEjjGcZhfZDR2huWIZvRUBRQVxuJ0IdhUw4esn80nkY2WhaLZL08cN0m
4ZGBh9PEFPcFzS8/NPPFCtEDi9jEAPSS76SRz2pXiFd7uczADxvr6Sr4csowFas2DkSyNaQM/5aw
UpK76aLAZE3xnP+cnu9AurDzLA15a1fEABUPcx9DXrx6Q5HmDIxKtqbVYbuS1LU0ZxgAbWOHAf0U
YDwe3wOjWuqcPuAmfyB+39qNLIF8ujmB9UbF3ZoBL1CqX7vGOB0Wi+GOAQNecMBHVDtle+f9wiKj
hIbEF9p6of00VVoXLAkwREkGLflZuYWf5FKVsJJHuZRVckHoPP+1yvgTNargl2ZofeAVgdnWcUEV
VMu1vtEzDhjdp7hu/K/lWyUbQR7f1TyEMniYX/k4gGi59hMPV83y/1RMEvE3yIweOu2C2yDy5+et
bZjhyk/9Ed7b5yRNW8K+lBTfV4ICvqUKLgIcY28GjQWU15KZvqO5hKVNMAh/o3+nktL01qzv+ZAS
fvbrdK9QmxrJrmlkzJQDtz07iJcYEsELint3QEia0PVvCddA1MzOTj3fWxYInQLWaSczbeweo4eg
EyYwbm1GVWhVjXPCLT329FkqK1woRNoAsbTOLcjQTWZjV+PLEVgz/7Ab+7WMIUTRvr8ENY/psE+O
H/7OqAr6fLv6V47BiBAHbvrWfvrgGICedpnUgwpNyc3shBV/vm7SAfhHrTBV+YSQn9UzbM78hZb/
hUTe/cYreWpvmVBrsHH2zjWYDGyXInFLvkfMhBI5mNESR4oP7sTfsxM4+J0hoq4pDU8fzSu6YOUT
6avn13JLsI4Ezbs5TctDsnqsk6VEN4ho8RXNhDSeKUz6hucOKicDyJmAnm84njAKGYh4tdW9n0gg
OqxwADsU3EszeF7hQ123ujhK5Ka+PrloLLGEdk4zUKm+rkWOn2gQF3mz5aA97IgbvUSk6BsMPvZx
16ps3JpR8sOsrnKeGWDj5IkYysgm1vOTZi7HNtrAzqXX5CqfJYk1EFOSTMtCwGL4lg6ZJGmCeQLW
ZvKb35lmpfcZlUd1h6YShTO8xsKUv7G7+HGx0yOr4axuD7tQIENDfE/HRvlVac8H2kPcv60kC6dG
HRYzCWJpxgLo9/3GEzUP32uMR/QlhrAmABirE1Gmmd+aNyKanSTymJ8emwUASRP3AiGz68a7+dzk
GTyi87pjiB3fF5SrFpeSj+xsrXRfFcrS6j1qe5QiAtYHHJmadMyxv3x0kz1R0+84Kbh1ny+cqOw9
D8DgTLEdKPyWz2GG8q+JaLx6Co1qazdWosWerIIHzLf2c4nMr9pv60VhjCR6BBnnp5zI2sxIQuF/
tclG6NZxMncJwV8XHXI6Kikcnq0YufNNBcyJM/O9RHH7HzpfUntiPyBz/CoCbMQK5ggLhuKoDeDK
HDwPps6Jxp4EwoY6ZzuY/7fKAGZ9gbvY1ltuM3l6L9F1yj3j0WplxW0rclZru04rRaLnqU3WVSM/
U2LamkKEsN/lNWow7dLubgPS5QanrCzD3vNtxZrcKkR+EwVdvX0wYsnRk2D4EDdtq+0IsNFmJMAP
lyDP40nsm0534FqRy3kqt52TjAZDjysDVLvj+mF2pey0HaQNpebJTq8FzBzcn0hwhalEBp3Rrwr0
A9SNE0r5XOMYIzGJM+pzejJf5eH0MI8gBJKE7kNiEzwSKe2fP9SWktR4GNJO7UUPUeXHx5Bol3/b
XqwD9WeWqo+boDul8bvC9vxHxSQNMfaMBVWwQh8zW/hXvTTnDbpQpXwsnTQcBDLCxYASiKD/lvVC
rHo9QuieHSzeRZBcuizYA4KSxIwNJXk2EjxiVY/B+HNK9v4Wq44SVFIUm4pfrY3hFM9CEWnqi3Mf
mcsupB8/pojeS/wCtSzQ7q/vq6JtvrzgnJ6PizgP+UMUNs4J1sFO2+PhzjhPVjaazVedhacn9zDw
YbDG88lBN6qTLDzx16Kvxme9r9Zslf7+9OMA5yOcN1qLUqBkvgKd44zeZhbsF2Er9J0nKpA1vTnL
ZBWInv9ulc5Y98g5JQ0PB7Svpkue2HlNZGyctIfi/7258eRpsUJ+5HGO7Cf37RzXDfebGK1R2ch4
0w2uINpAF4Snn6mEZjrYnpqOurXdYat/0W71BFcHSukIjV8bK8/pIdRqeLhXYGgfNoJwpOMai1+b
cC+Xd1zpN2zVG31zuNGeHYBZMF6c530q4I7ZBhLPlTuEvm+No764gmqgtBDmBseYrfv1SwAbGQyz
5x9zMnKKZ5YHbSlP+Hz2enzK9bn+pEzOmV9uzjC08YpUDhfP2xyK7JQ5kx4K+jgIcJQuyP63KBIW
wCQKmqIJYPmPBmU0PdZgGNDRDjxLimmGHXyHjTNY9CwAqKewXOJ1WzrjubaR5Nsy/yyUtXfM57f/
FWp/0MH/MT6PFOt3TqQqOFKlu1zBe+WCOp37jDY3ELTtID7hzETawHnp9GRB5fCCy50kap6j2lwz
09yEACayB0uiWqnXPZod2luFw0ruRDTZUMUsJD3gtWFmZWEBgKJWVK5xuO1gZKF/i3K5Up8XJ613
GduJjdRvE2mCX7jwb1zMVcCMff9yXgw+AeIuj4rXix9oVbgMsFMSqSVUN7Brd8naEOv5wvoErxZk
77Bx2QTgF6HZRT9wl4kKvlpSy/iYiH63/fmCgNUZu4c3s40meysouX1o8nzcLxwzxMu6WRBN02Eu
36N2PZdWAOwq56mwcrKg7HKlJrRnJAxLJ68ojcZmbzwSfkDWSdYS5a6ZVFFC8JxZ5M/Oa2WU8dSH
64t8r39VKIomcfDaUWasKALqWhIHieDqKkod6xBTF+ndWbgWHejLs5Fmo33cFmt0TGB2VJHaHv1g
pA63kRqA8oq2E2nD4EgJit/yfiD6O0vaPH1Jb4e4VLXicUfoHbUQqz518rai8wjet+T0RXbsmPIJ
OX4ZNolqO2+CoJrEvbXUiMvvzIrV6NULgK4pIWkbsrM24N9PACMwEenE6G0SZTlrhAvNknLl2gga
PKIygknVbo+XQMDxXFtLo+QGODFxBPgR8IISnZSo9WbmxNh7IjLPZmCs9njFg75HQT/yT3M4U8+b
MKbZLoZtUHs3F8iViFOFC8dOkaDGBBgxFs+vIuUSux/zNvF2GatV8eYt4UsuByutWyTNVEcQg/8a
rLSfmhILrcifYR1cZhpkj4MX0APSMCYEXVzw1r99CdBBANpwFA+yl1lg2v85bcJuSYfC6XSVtPqY
U2tq/F1Gf1AuYPFqka2slr8VXUMXsmVHXvwmVNCTsXu0xGTyzgjm+TrHTznE9X6QjPh6sewySZBf
TkXPccETKlQmDOSK6XsueVvlH7qv8l00PU49XmLcMOrx1KEej7UyxVdh2QrFpkE0jeW6yM9kISO7
qDe8oCcsOgWd+O73uIlHCIikzAyGe2WTmbb3f/BJdz3Xjmp69TGAYNx9n8Lx41PW9cOLPlxVdEM2
9pNNy8cuorKVMtf2jbcKOq8r7bh/LdMbp3RBJ4gwP1Y3ZD6fRns9psy9wV8O3vk/Duqw3WVjsp59
8m5F7M1EAxJpsWNNCHZfO11gDkENHXepOFexXh8xnbbkJ4zD3I9MoEhQJPyqllyoRXzv7Cfc2CVg
Se8SxdaiWLQlTKOVzXxzlIn4ml3+WsAcid9yweb4bWc3Uaw84ZZmoF7s+fU88ilirQomgZX7+l47
bMEbaViY3K6gSJTZIJexFix+NwsivlNE3/0SlUIdXBIQmd4KhqVO6OMxG9NcJzKRtEWJ0hf7rpV6
G/iN8SXZ1djEYm+sIVtCdbQCvigSjd3kYefqXZDUGhGeGiAmY/D2AXPApTPFZaK7gHiOnhQ4WyI9
iTScOaxxAGFChiQYK4rG0skeiAVO6zUsI+TOtwCkBKabNCgFPFWnC1J9Mmx+ffBrrj8NocazA25G
nxali254h9TNwSs9sx1uMv29k720OADfo1mjSQ9fGECsm9sgScfLaVwQE+IDweIL/ndXltsU86Ty
ZaRoqT2Zny4/OQEcV2sbBkfh+vJpQOYiCDUcOxXibrAd6JcsTsjbYcu0wyy5UScpU3QRBW/XpmOD
cf9Z8PXSD9Jq10H+OsaiGEvw9NjlgO/xolGsEQviJVWsqqUds+6619BUIc/SbtltXmj7xjkxu2fD
0LKYJF5zkQJXlnZZ20cTPqyXZ9ynKlV9oDhSr5mI6i5y6bFZjZ5ZLur3G3hAlDSwOpPdVcdGq2py
rYNfRY521A2cqNWd/9gSGrOmwOxI/4rLi0RaeDZbAYwxJiVHIYwTemEgz8OqsdEaMoWM6xxXVYrl
TeJ1lzOb3iYPiqPiKLMk2EZJw1q7H4PxmH39WMWrkb8LnQaTIXg/rXLYsI7vWKpWktcZ7X1vZp1E
ksONISAo5clW9SuIfHllVT3x6Z7KVz8dAA//qgOFVZU35uoiDgR9nfdr8hvftoGHpE75aGTXK0GL
L/Lxwhp72gsmYTZz2pkRJtlHmoyEBYPIYwdiXZfNsWnhVDUYYZlrPgXwzSNqMb85RGyrSR9Uf2yk
AlGjM3yK4o2lN9FvTt62jbHQli3hxxyEPJXX5JzN0o1OszMn0zVqepqC8FV6hckq7cNX1UjBBakH
POz5TVJ1aI5p8JX+keJCzGlMHVwnZ4bmYWQxLXwlfHZkKR8WO4ET8xKuc4uDtTy5Mn3t4leszkfK
UYfTaKkkLp2t1FHxArVi2L+lgVKjH19ZXWNd3yTy5ooaIOlZNtDVm3YFA3CORrKsAhCJDFb9Wus4
oU4jaejaBXyOcp7plE5slwSYoQZqw8n3y6lA/z/9wBZLjawRLc67nmpAjNyl3uZdjPljQivIQ1kw
0v2bfAoCd8DpowPzt4ld7teOmEsHj0pkFUGxxPhlVD396KtotRaIbgaxVA7a9CH4UouFiNwzAKcA
ic3IVY8jJd2k+fKS11ZDfbP7pe+L/sMDyDQrzwLlS0p4g0K45dIc7rCBnXxTrHoFjOELN6pe2aEb
EpqURHpoHjf2f2YgTbx2bgRmgB0rJANXEWeuRyhJhGskh+IIdJA8d1RtXww/HyFNiah+15p0HIWN
k+mxnxfXc1Gx7mmgdzI8t92QG4myif57HLKGgkmcAGFxWt53r7yPzOFmNJlATE1W8Urj4itrPAYv
ffdXHsmZVel3bJ2ccumFlO+gQB0MMexGS2stdJUCyZkVuq4it8+sBcAU1ACruWil9/XGJzTqDIMj
4Js4i7dFYGDL76u/qpeD4PC41fBdXnw4Pq9WMTDooO0nHzUx4EGe7IMBW2jVMqLPXV0Zo/i6CPnT
L4Zc02npzgjSnRhRWIF2plhTBI6gO9OYafYyoILCdCtXOUitjA23qd/zIRpjkRJu4OUfWJG+m8ZI
BLAsOvaW2FIB6hwz00lAZx5GqGfXqbenvRchrZ0v4Abql4bEprvYdUCG8+W/LdknnnPP9Td4Rd2T
nQC11NWXGNtqqqd9JTVNqN4xt2ab7CuYgjC4MjNL7TJ1QlvzlhG4U5hyhEc5pAZBnVBU+WDNEEwu
KogA/6ZNskgdZNfDIhXdmyyglLQWh2B5iQqV7ZqAhTjB4rIMFFnRp/E7OE3SEPOwszC7KE8vyWLB
qe1lU/ZiH4OrLJeiU4MtokCqKhf1FL+Z4M30T9rDoyn+wHdl0bTfuwbR6SbGjrKZIg61cmFGmCng
h3YYy/nZ43oJ6APiyvPQ/sYoPck4sqWFiT0BUe6bdQwTDdhQEXmk+GDi+x6W0ghPfkUp7fG1O3Ec
Ph5exufrfPBk9r0EhCch7k7kli0z996PTL5tp4w1yNP6Awr/QI3eeOvnS3jjJ7OvKOS8sSHvinNh
5NE/r+D6tnrzaokFpTA8vqOLuuP4c7ifEtqhpccVy3+Idop3YcsEDNijNZcgUJ6yoSEAhMWYCzCl
T1SoE3OMM67pDI8KX793+zstvEO2dkv7n+TPJmpM6N2KQDRc+hfnrBU7e5BQWYDojKYWw7klYwsP
B4uP0rnHF2tvQ1Tn3Vn52JfJTFIt2GGpfM6yKRTrjuymZ3SGWVYUWg9m5+IRCspDqI+RriBIjeBQ
PGP3S2WbeXKSpeBhy8ptQewhnN0juTYcpvmHQzX9K6gtYHs8ptWTfivqwk+KKpCH8dYkjuoaAK7B
USr1xplYqASIeE98Ki9lnbF+9rtYMFUgGrkSY6pbzsZ+903yFYeNIAe0TX9LKjn0fpNmedsPTKpq
0GhRh2wzH3QR4sgVaW3sS4j+sZ9YmxOw60pvkWLsShSkXAlAV79MG6iuowQqv7u5EjaVUDZYV9wy
yoLidXQnBG6tLVxR9L2/eaLoe+qcFnVr6e+VB0ZRCNs8S1os7DEPPhc93BhkraEeDrQK9TxP+M//
94QcHePz7uYBy3YqE98qq4eCj0xwff0dV2KFOlpZ+bna4tWyqLf1w070xdWxbPZfoH4pdCdHieqJ
3+MjBrt3XI0v695jj+w0l3zDyeKrzL+XIrDIoOUOBnFl3aJ0+0+hiB4hB4jN+gf7ftPsZ/kakRlm
t8KVm/eGa9IsH4YGZ+AUpLpGuxxnKbtHS9O5REuOf7Q28Q0bTt/4zLPKYzz4gl4EMiZos+S0ADFX
eieEKNk+s9GUldlY6DNPrRfCRXxUalqfTm65GMiQNWmLfsAJq9cMxBZXlyrjXm4IMOlxRIKFIeo+
5NU7QGgdI2usC7mVImvqELmBSJ7U9wKNJH0H7MFMsZClZsHcVpS9Lmd1xESb6KKaFgO4hNkiRcZT
UOhPBg5sWMKWRRhww/7fxHySD2gniSYYTNMHRvG0IEybydtW6SYccJpmDVqK0YwQwZ+ELTCZpp+F
5388gOkp3m3mUzh8VOaQVGZiv3oxK5u4Enl8oOzinA5H6QFn4mDOWU9NwnF3VifPcJ6tUCKUThqx
qBemDPt4g374ghla+71HPAFpAHW2LPnFqA6Ajv+oBHmmYGFFaR3g6B0Rl91kobhV05ucUdnPXWuR
P74Ol/XSgjBfje58R/+SWXNGVw170DfnceyqCA1yGu6Lb7+SyaeyhPJ46ldAJbYAJORYQ/7Hp7fd
Hm4Qz1jb8wRGSRWRTccTdVy2yO4bXE5fgj1p7AgrPgfwSvKO6kI3BOFVGJrR16gYpdCVawJ/bTpf
lyeA/dDkhNBT7WF/sOlE5J/H/a4ZqKlu7yyQxp08nd70ySmm7hDGQB+VRvfabMNp3KxBqdCv5AlG
Jt8n3i5dP+cG2CvG8q78kIdEKqp2jJneZPr6IwCH+dfexhNOuLaWecsfcJAiKYyxOxg0Dw/cSmKu
JwkMhY+MtFXdPRu0IdmInqyOKQHELDXhOco06bam7lKIoyjUks6hkh/OABiGnHsVwoEPTELI240L
dAFbGcMpKHZ19SgXxnaXYkvui22wfIeFFcms6PopgQzm/AYy/+7meHYtx7yBzxJX4s15FEZcZTO1
A5gLwrpz6d2b3QnRH4imfBnyey69GpRtpNeQ0Q6Vywm+247zcxAyWrYxSutiwr2jyX5uTqU2ZAVv
rS6fuzpqGRw6a6qW4bTNhc9l05FNPenKsy33qRRFtud8fJIVXJoxk/dp63zWes18u4LshfjICFWq
Z6LL8Owxs89CRu8EkTSLsXDh0fkDVzeFztGZwE7454dIpE9+afJs7VONuip3vJwcxGtQQ8WZ4qY+
Ko6mVPPN7TqidMyjJ/GUzhfFsZiQWO+H/abG7vvSITRdB2kyUXgYwRElanngb9SoOOvGAuCdYwIT
siWGyt0cLHIFDFmfI90hP4eSqvUsTyj7kUaZVR0rO1daz8kIPN8QXCVUhCuhKviw/rQg9SMyZ6of
F8JouCK8IqAdRka/I3Dg9PM/ff762BnsxIr8e8vwBtCi8XtlF8N7VyhPJWPUY30uVic08gDSqttb
ZEp2kksa/RYiLWI/AXbrl9dLArRGDKkfAHVycV51IMpGchwKGVIovRTnMlGSRy1IqBT7DNopD84H
AMIrsIjjJ1pXo5JSm6H/aH1X44zu3QPJdtRAjnLz50E4E2E740QLjZ0rgDBN52TNdC4Ls5w2Lfqx
NKOZELLaA3sLrfI/jR04CEqGvR9a0yHgsOYFa1OSLsCrCFRhNvPgD+wNFM0Mt4Z0VkEUSm75c9QC
PWiv9FyuJb8Jk+yng7H93CLrx+oqdzC4yG1hpcvfHlHNsQDU4u+cOsSNbhd7/naoRwE8e95fBtIN
YjtnG18Ip+8BnzzM+2AR9cPYOnBa8RAbav2fieeVMHQIbPMYrGbNGyCc1lWFcG4hdBycJmp5c0jJ
rqtS30sArraXwVjil+KzE0l54MiaJdp8YH0KWPtfYZHEYFamPPqNEFdVuw3j8ZcdsuFazAEw0CWy
FM5ijAXF72/Czg81Dm38wz5iHikpntVQob02hIIJw3xV81APe2H325iJvlvkurQsW2GeXptOr1sf
OwMyR2L2PQVtCTubkpGnsZZSnvdYl8K79ICtwrPO3uVnMDAwuDDH+yDSfziQJ+phbFcG8OD1lnEq
FGdMuS3QV8LHdcb5vD1WH25WctncpRvFmc+HxXGeMyHSTiR3SAmSM3QJqjjI+Pp/6TFFcgWWu446
ILWOmn1aFsTTRdORXYjm8ETnmgmy8N70vemLbuESQTIXiKj+NL9yaTS0Q12UCMv/MJaLkDq9aGIW
aT2BRy4CsWakyMXMayHVX44cSMnX5griPDpf4sb6lXN0nOWGosPlRgQDipTSb0ZlZE77visYcRrE
kGkZzA+FF/1rV8NoYt4RqLJeTSDbQckEsyUoIBO0IyD7Zr7sG3B3IO6TakhYENNACZ7PNo3RDdXX
KffgIU6d5JhNOLXPrdxhLbKTLXh3DoxjsALb4MoflyBmYRKMhXbtuV6MigkyH/evjgqC266o1r8z
Lw2O6b14MKM1ya4Zz2RV8lrnSoSjRQduOpF3J7ijuAx8cUp+SJsMQhnsIQqX4nxUurFWkEaw+koD
InGGpBeA1KHMI/bpQrB9HeB3L5bYjEczjk2Phqb/WOFCmEMEay58vlWczaG/xcrfXc0FM4M9ChUO
E0goxqKbf20ngGR2VFIfeQJIMt4NsmVHdzEgk5S72h/J1kRkyvuH0bwOqdHofRsdO7/jz+MsmrMu
ZlNDi773zDP/sn8A8mXvNEY2DjvrXf3x6+Gcg+Ez5pkr2n+4Eqp6YsYfQ9CMc6I6FcAdYKbQevQI
fp1/jpyTyA0eNMEX+Fv2z3ZfdliEdUyOa4mvvD2SoRfchaD2SWrzBLxYmCbf+ZZVX+Qz020OsV/v
L0TDN1ZMPeTT4k7o57DQcfQs6oX2F9ImV09sGOSG/oRFDvkB1bRvxWZ67Ux8kopXMT84tidE4Mbg
HiPNU28Gu9BOaPoCwdcZifC5vmMKiGAN1nL8Cz4Xs8jE1i0K9OClEMnwSf6JAVNQ9GvvHiJ2NJFQ
hdUmfw1+H5CzwaYYGS33NsbtFfR+KJu7q1XWUnlDtlcL1V3Bwn1iUtus72lPPBUHnjRLrOxEznpL
zkCX2Ejq2AsLmqTMB6LJF7pE27TjAVGJgDy18BzFJKmioRe+d3GgtMACwDV4dO9zJdbvIwQJ7Nft
HMp5odcWZFvs3tYFtpEgDt3DG7FrHM+dcM54PNrn9g4zFPXbKXLT0tFNCqOve094nVLhOgUU8Alm
aOhniYbzvBhVXCuOjhP4F2vec4bLIwn+JYnQCkYqZwsu4M/YddBK5jZEUQURAQrnLbHU9toBHguh
/tbhK2V0GYi4cp3XG9/koo6YB3b8ih8Q4on2NkVKQFSP4E1+JxpvInFEdbU1yxuIaA7EgCu4/A/y
4MRsNL9qkfGyuatpvwOdAlYzomXaMLdQLZ254WN7c5hNoZaBUtvQK0VAeXW4fWKpBfdfiCqvei7+
zvzqdgMdaKHccaiKRDqnjil1Dlx92L9KZQHQymF7OE+zpDe0v51uWkny7oCVVOblT8yYpYad5iNK
MtdZ/TabwkS74kiZFGr2tTTYtemex1IbqjB2AytCF98IsH1NgqFIA3DhJcI2JmA1tnGH7n9QJzk+
GpR5VVjgTLjX7i4HvSutJOGzieAZv2vmFxn+Y5EOdA2ZYC0m5V+SsPEgT4wCpi+5G+DaxKe5gU/P
QBj/09wLl3dRFVqp82kn05gtUXuw/MvLTfBkD9YMtpMOUv3tzNskfjEpX/qKUnaQJuu5M59TBesm
/08jX1q5KlEMMWWWQUUUoeSdr5kvtbYNxi5+SyvzFC7iabDjC1sXn14EH5tUDiosp4doEHo65fjT
2kwtRLj87vFI0W3e1ZOKIBenj+8xGmc+RCT2ZGxMw6G+dLRBaxXrJOVBcdMniS0ORb8rxdxzRZ6/
bn9LOVoQrk+Fm4OcnyU9CnsUQKfI0cdfLEhHo3srGcd7llZa1L1MdaMGj9WKpKWoJjxffjjih69D
XzgJc5lgHRhC9Rpzn2t5l+yD3qw/ZdigpmtVb/2hucg5Wu/h3vPBf9yFJ9bvy4SW66MdwFTIUfaC
hqfXRng5plqL6e9U3MXj++rKTSdLQiJRnM94QsNYUHSXK/pC/QStjnY/vC6K+6Mj+4Bn6c5mMG2W
PY38epMb1zBO+B8VZTWAySxZRMclIxnI1PFmvQ6DtDTlYalAwa97eCxctoEf2lFAheO8Yh0DZOn1
iQWdR0wFKdUKGbW4ioCZLF8JyMJk0LNZut7xKFfQQfalh60c1DaZdHWCnRat2n4pgZw4E9K3sf/z
5aW2dXRw2DJBphVNVsT//EfBMlQR4ndQ/2R2qOrUrWbmsS3FW6++L5x7X96VxhYQyVkacUPHVcKU
/zrlQEDvcgWhwmhvXOGOwNH8wpnAo/4RFa5zM1vLODz0A6fsuBf71tIGS2REPmLa+xZW/wdh+HvY
DPviGZDFUKJrM1UaRIbuRsfZ/gW2kqn8UB0M9xo8Jwj41U8Nr+MkG1dvFEUHlZIEw4SaJ5i8Gx/o
0K3wmW8/q57ky8gBsFFK4Ces3yFZmov2DQqHBxfw4okM32syMqPQTm3zQKLS38Wkgc/vWEPNwo8g
QYrpmkb19SdkAZdasXiD3X9nnra1djr25ZvHn4SPggctW4wwe7dWHkHtZaTucJCMv5hhG6waHDbg
QCs2M/v8+lQpt2yZs6yaLdL3nMlkjy7ruyyKVZd1fF/2gxu0/2AiAPnCJTHlhE1G2MOsgu/t/uPT
0ncUJVLkSYucCtLtbbTJBGphG08Cf1PjJl6/Sov8JdC22KtNHZka54MQ5eJEKyAjms9DoeS393/3
kDaANAuRYZsq82fL/fwDiEHlvyWFAlNmHvcVdbHbFl87l3wQ7gCc205XAF8nSxmwi60SCRrcXIrq
xNxslq7gRMjEXgURWNyHhK17OpJ0ffoDSi9Qbqp2r9ADWu1eRkhFvOXRgZlBGL3QtLIwq4Z6oREr
FxpcGj15ZtFTYICqzeDGB3WesmZz/aMOmhAzYvpW3w8y5qHLilTa7VHuFENKVQH2NwVy2TdrWQB8
qWnMehBcPYFnwCyoOYhTzJX5WOf/pyYmgSwvf5sYF8OS+LL/ynFQyLeTPzKS74ISX9V7fD7UX9fw
WYd6x+CHESmSfcJaBkkLzuuo3WxOUuY112GKVQsAoyOi17hiToYwmmHzPCOhzMnjNOTLBOMBHL5/
DiKRH4w2mxUQNogQV20SqNf0AZhN34/xwcCRzAUJyU3t9dQV+wgk4uKJFBLmrMOy7D2WcxU8Zxkz
WX+EyPb1dBXsrtWPNqLDfWJDVfa9RmeAe1kSAzt3GarQv/GKD942SxuNfSpyW5l/ybjRUvkp5fP1
FOOarLGg1fkse73vBDd32mN2vQ76fCed2cGZk5rXopKxx0ZK0rFjXK04RtOs6CBect8YrcrPegJs
iJPanVoGS9ozbkVolk+FnOB5ZizBOBkxxFjzquJJlgJD0w0Wp6qA7JLIDgQSLGLRfm6gg/qDpoRn
47seT6DgxZ91pVvxDU280CLz2pbRf4MDz21De21G1LUOIBAa+bqTN4rlrtLiw+utNVRuUh2znFze
wUUl4IQ2c1s00myC9tNSlCToxyiUmHjMRgRJx7v7xreE7RAkFYdxyDywzA5bXyKuutYaYFo7xLwf
Tf8E9uzraNm4oBr7kFc9+RBOCJ3+u+oNFarU1AmmMMEH2I4RInv+yc96ej005Gks4Cx/uW6OqaP1
DoWhHIpvJ9rQ+CHdc0GNwWayla3YGC+XUYwiB0WY6vTD3Tnd7ZgXwW6aIZ3J3vrYgd2wSPeJ3aV9
/s4eR9etnj6VORJVpCa3Z7cx8YjSCjMgRxlG5TW8gwKDv+/qsKjVbYp48NZtAkTJJnSNoXDf6uZO
Q6P3FQKbZ9HnM2Yp8J3e8INcmWxzT+MDkjERQUYbgugCTlAMo2s3+6aAO2N2c7jlzTJzqLWNmT/I
nV8owFEpmhBnZKW4li6Bf2BimONrkJIziiDzbe68qU1gMqgIQvJylelp1vlZqLHMLBSVLRC90PbE
UFw+d7XTosWKLB/jg0qshNGWAeEwgyuEpdpZt8k3RsJL/3r0Hc23TXyk2zvbbtLExDHJWi1RzMqu
0OqfGWZPTMHnW9YHsQFrE+safwXBQmyPoRLozk/4quNU9vVcXiNlQ/VL+PUE6zxblP3FYqDTzSyL
5tO/OzelnwfcTvFjv2MdlAjHoffs/3dsZEbpDgMIGuA2odJy3y4z2kz9w/NIev+OX9OtxO0h9g8j
XUnGs8fMchwdFg9j1Odj0ErrBZyEeuPpesdHYy5Pkg9apNKQf8HRm/Po/1Ij6lfWWiCCIpXeZbbR
hNSRhi3L8HhFKbO7ZiJt+EW91liUQKo822kZqYnpPfibSx9u4PSA/LOsz6BRhtYB/szprAL32rye
bLS7bYxWNi6Jz8MoUo+P+vvIoB1B2SSVUXHlx1iMKm9wuarydY+Bo89cHtloriaXMu2Yq/YBJRBA
s7q3kHQIuphBQTNrPZrkyMU3oh61+jcjMfqVWj/ErapHSk49Dv54OC5y5J6jG5Mw2YjJUcQw1IQR
w9mNjaaSKXLq/O67cCFpa4sOwfmw2zv8afiBn7IPSNieXYchY7hVlVl0ZFy8MaCdYHgtP/n7sAns
HAD5nGOoQ7cwwCKOFcfYmmGXaKSs9JCUopuD89dr3/GZ216bLLT5b8BEjJypsPC2KzVJ+RCW17zt
zPVoiO3lLE0GaevUsXaptcbjuLv5ju8pFgV+gjntAXotShsmkeIHdz4wPtJd17mw5RK1fkdCzBKc
uKHIGFnZgvOvvvPFT+Yin3HO7mMz9XLUOe7GM+J6y2hQFiFifqxcLB2yYMc03n+tyUHubJlqNTd8
4UkqOStA1iMB9Zc4vf8L0Tepyxsn2hGxmV5IWcHL8StSmRKHdqsaA4VOy2N8oB2ZyJWtu2xMnejI
C7B/e/ashiH77eFlg0k1mY0fslGGZ3IGLIG0IVgevjUXTwuySX4gEV84MV5u4dc6VN4HSb3TKd5M
BPkT7oc1YJeZCrGE2VrapkqoZNDwQxYkVanM0vJZuHr3UWa7m+YpN703xtqURkX6Nh3I8+XDafRR
EQN01MOcj9EXG0/PIcSGJHhWxWYrDzOkWHQW4vC9R+PSm0jr3W2Z5F7ojRtNMj9LHp38cWuEX9F1
l5T9WSDYwmLeZX3XS3iuIGqGbakz3jmXTWK+EWE+TPQmzt9i3jfjprcfyyOzCByc0SMJennW/p1m
jsLEgu+qFJyKfJ5NHMvup8D9nEfL750FDOGDp3JnT1qXkJO83XrnLkp+UkigrumD5IU4zIBEvTwD
lmeBH3bbDfUM61TvBKO0K+H4fjEu5XQm5scAqXbD5YeRTdpH4b/4Wx5NmHhHscfj6nXefciFHBoH
CtjZ2U+Z46Qc5LL/9qqPmVZd8LapfMwIJ1o5u4pz14ltV9Gg0l4YBvvewXiS2UB012ge+wkpfy35
oZ3IVsKZY2Zpe0yvuKhZFKGutwrWKYlKOFctP1Q+dRSDy8zY4h1rHanFoFgRf9uI2rra9UlyMDfD
mUFZDrH2/rhp7lFQzK4iqx6ZO858xFpvGIT51nebIaoCXYpMc/7qa4oxCN+T4f+/fEMSr2spyoFZ
VkLNBYfmkvFRge7lAoKgoRG7bdsMSxXYecGkmcLXt7p0hcvwm7MpUvfhvafn8S0UyUe8C2xEBhG3
G9+lR9r8OsHIZ9XFIcINb9dYtaM8uf15xYC8b+8lwkj2Q6hH8XiSIGBqEJwEyYtLi5IZ+1xEavHx
LPjmMozWxx8zcdwnEAHngzLPcRH7iZxb/GlEeMvVZZdfqsqvafBpHbGInalhDgoTOhqvaGGhT4oO
4he52RORBHSjbZiTDqlZsMBXnSgTVT62NnqsLcehFXxGuHcFohDpOflLloq1juIryc1Af/rRDmMA
PTjrdoNYVnnkF36ODF8oRvwoOYEAHjUay6fB4cA1Dg4aBBFbR0/NP8indV5ufwV87Mt8IZXuenEr
IkXmF2fl/bB+f02eASu0BMY19jR+xuqf2MxeESeib95L94bC1ZYX9NiZay2wTzz1KKKAsInqmNiW
GFotmdDad6d4MCXySvHB8pGvmggfoKVkz2oY8Ve2fYL/Y1TK0cVuDoiPZw8bRfevIcnAry1iOMsT
XZMbBAYH9kamqAVmIwTwNqHzBjf5QmgyvmzH21ciUaK06l9rM1GleKzUYNo3X3uyaLJjXPyCV5ho
Z+clHIzgIjzvCBRP8cw0wqSwmw0kSU2N0Tdx44AwyxwjEYK532qhFYx0mzzsh00aadFhy2Rt6/PJ
ouS55IZVP4DNl20N+tQqzDj7f9NscX6o0wWjTE4H1g/CFlJlNBbsweydbiP/hf7WMPQU2EdDokJg
uocszUnOsRsCg6YD316rHGsG/7gLsWSo3h6S+lCB/Sfjfi3vwfUIvP/Si6VFrN+dB/p1FHNltthz
6lNza55Cyx2O8cvphWFPxSGJCEOs9HWlVAdTzauaffjOocb1Yg1gR5qbcQAbT/x+BWM2EteW0ZEU
UCCNUji/FeBWVknHDH+iy/oDVLX0NK6LAAcEarmaNO1Sv5tNjZNsZ41/M4+Cj9piZGezJ9Bw8BmD
Zo37dm8RxywjjN8JI0A6IUWryxCR9h0nM0Wc9RpqALZRwwsNrozHgU3yiTtU1JCd0ZaBgVdr0wn6
cwiFHk6qgXhwLnVyNEVAObbMDqggtojmnoycYxYBmJCtvgPGf9QqfPXu/BzbV7ebB5ObFhOwZK/8
99RCAh3bdGKYVrWaxMWc23Y3voT/FVw1ANKW5KYGCGUcBwaHoPW/2/fWNe9b0chhAEgNPDjYaV7l
Gf/raXF2dZXr1i1fZCyDXmu4rYKv5yHRanNdchRLQR+ZOns4Jr8Ry+LymG9nscjVFZXysSNfj8bv
AONroV2dNVDAUmIq28mrQCjL4wo97fMw8JPgM2zxZPOQiheePNBv+bAojh85W1vxz/FDI3+vuqYi
ifKfncZs12QyUBLRvpSxnkTEkoHlA7SnSMDG9FK2xkx6ZwQEsFVqqXXoAdNKqEBoK7Db+lHGTuAO
osAJdqTarWvxBwx4J+3vs5PvQsxud/kOND6i78PijJb2vqfd/GfQzptowbR4NVARgH0MQM124V/v
N8IcbOMz6nLYjqJi5jk2jelnIOd6sLej3r12etEgRIdFKqb9YtoLBohP+YMbVHZUrURudNYhTvbo
5sH/D0/Ohq6kKRHnnVpjfEeLz9uWbu34fS2z5xV+DH8uJAWkf1VTWn7qCOa8P78jU7f51SMp4Qw/
9k1E85K/4eT55etzudqBk15/sRyQnmNlwWaWkP2WUvP4HkjIy3SofPQp6sIoE6qo5GFyWrVW88K5
DLV7gP2GbcyXkT3HYpjN3fG2Afl4U2c1PFCgUqGVT5vuiMGETw8Mb2KiZfJw7roOrd5iVuh+Obo5
Ne4YBMW6di7/WOXL9LVJPOjYsX19XoIGsuKDotsqj1lVset0na3G6VqIpczzmd+xfV2UheTX7yqm
tz728yXNgEm3150oq/MxweCus/SU01pyerXJVSy53ULvcwXpr7pW4CAuumRIxftOCkepUZmrg2eX
TeJ5E5ImAOamE6Ae8xKjZp9cPx9X0BPdphMrEOzNPWQfIlD3stiHz9rW3K6h3rr6U/IT5XdYSp9g
apo8m1alWItp/ofFrQzopL1UcAn0xAqN1Z4MhrwkWfqEHMe0oCIBkNIGM2AmauFWAoRvEppBFC1i
AIabNhuTWCR/po8SSH4tds32Rtf2SRMf+oMh4Cs6/1cXNmkg/LBZ8PXClp7gaOfyZKXSmB20Uaos
A3ebf6TKil2WuYtHKfQBo69PWo58iDC4r5n2f2+mECTIcgQf4S5+yF9izHdI3vCdpiUNcHEqhcoB
CKV5XI8ENHCJWbMk9gRZm1v93ItHTOV0FbkotcVf6H6xLtw5mhgxl+n5UaTEzWq8+ycljE+a33m8
lZNMkFkOBscvMRZFy1CmsGmqQ6rgj2ESmthb6kcBOS3XDtj6O9YR7Ll+oSoLagmYtQxiLdsGmGrp
CENlWxrUpsfZ6OQ4TRzT89zuIAlgVRYYkGLF4F4mU3ThW1AjBFpZ9SMROpxtDrefB3WPxILFDXNX
uswbe24RMvgWRinHjWX8P6utbx/LJ63FVITFX3YLPquZ78XAbLrlj4v7WZLG1D7JOiDyF65H9+Fi
yTnOMKQour3Xkh7MMJhKGnEiqH9PmWYDe2UwfM45rKwoUTcvg+e9paVgY9RAr4EqMhCL4GtZ5Iys
mORaMWb9A8Z9Cs8Y+OvKeen+yOcE3B2FOQTxRVUwC937GdvyznVhnhK/mKaDdo0A+5IEKMOdm4++
PuMNXlvIhuUGwdjRMaQh5opPJLVrOoBaScm6NHnhagyC9qA9aTiXaeokdnWGORBMHDdmTQQF5oKO
SbY51XDYipCRP64PHh11bZ43NDp2W2j+ecPP4PkfKcKr9VTZdCUR9EOoy8/znbZ+TZnacAjXk+5W
LqjrefTgZxOr1mV6MjHg/mrJqLx5j5j2oc+//9JLjb+L6HMVu3TLTJ0LLWodQXEaCP/0Ar7+vt9v
pHvTUpv3tBK96UtH+DvL7pYeK8MDSVAz6UO3l3m9+RPkpHLFEcbECGHXkWdZYgG+NpmjJJooaN5H
+T/3/nVcSr2vu4/jQlP0RpdXoWGj7ViWQMhYRp9COkJ9/3B4PuhNq1pt76+VPMRF00O+KvY6Odh8
ofAaVNmxlSWPs77oqiXMnH5bmcuAtbtaoywEggYqXwX9hrizU17iW/vKUTDkaY6y5fBflpTg5ewv
jc/F/ydetooNccoc793Dd5sp3OpQWYxibpVv0/i+MdFytT+4eBx7R67fSIHvGM6Ww7RRIBp+TMRK
gzKsHjJ9mF1UCEyuCTFZARnf6R4hT/td1PYbxfyVmiBGZWetG+qpDp6RnWxElOGVznGa+kDrnpq4
kblDSc6HQujNPPVL3FTvVzzqHFQX26ypExavCrhfiAV5ack9WEfO86SoSOEx+QvQO5h4SqmIiO2W
/zoHcoKYQmUZuyqN+jxCCKsaifUftvzQN73X6tNygWyBTtjjYIfNp3Vu80DCgUmzSo6Ydu0EP0S0
EJfpiEB1KJY/dmJ+aTi3sIUTP/xxsr+9IEcwzjHxZe1rL785IASn1wDzNsIxWQTJe5Ec5OfTQJfr
0EZ3nqKhcHoV0hbNqH13XzfhjQ3Hz5dM1w8nds//bo2ilh+hA3Bc42RMI2ibbbaPXhB7Wx9mGVVR
seB4Kzdqa0A2wirwzIYvZDk5tWXb/HTr8YJR8QNiGYiaTs5ZR1/Tf+bDWhbEb6flmT9KwOR8cOcN
ntYHZEh4WslDAi17KPv/GXoTBhmSNgwIbIBOlYLVxRRq3ziRS9F6xNWfp0qIVPP2WqeSB4KRkk97
AIFbAUMj3wNAHI9WknLY41MswZeQ8mBAsNtdytgBDxKnsc/ex3XvC3EwBcGEKUKTiJeP9O5t5GiN
v1sRm85A/oVFzjyfKbVNkj+Rvb4OTtvYq+U7zuw6ziYi48Ab5Qdl0hlQELjqx75O4oLnrDeJasd8
TovTgjnkNvFxeILYUPl393iyp0vZeG7q+Gx3nGTeQxxiQUuS98VHoVU9IRPHIZIAkxXsZKozF6wB
cWYAUXqL0G4oszg2/1/pkWru6v7sHBA88smapyaHoiK24Vryva3ZDjdvbgkcQxUeuNhcn86jsGDS
TJe4nNwKJLvj5iGlS4W+yapahAtGvg77VxGONulnrRwL2Dgm/Uo/9KOEGJ6YKcHRSAg83N5oZj00
fgbtPUJnIIj+COy19dK1xwNZ7qReMclwqvbhD/5Go4e1+6vXyikss6qjRxfqCQNOFL7r5OVQrH6I
Bz5U776acsDYjA7Yv2G4j7N9L2dG1khi3B1bsNnjMGZMdNkREFDeD7WBlByAIsmIrwyExNMvocdg
x+2hz3hxcFc5VpJW85F3iXfpc5EnOuUEFDrisUsYNAoB4huGOYHVI5hK+SlqzxB3iYLNtpdF5ZS/
t/O+mn7pccA0AgQQBKtWTlTKs6x61VN8xRf/hlsvmq0wbiZnx6BeVdMVWjHMJE1wu6CHd+l63qwj
C/+/X+kBiHo1uZJe70PicqVBbh9hWjcLqGdlzms7E5D9g+3fnGKWJAfcKrsnfg05DAp9tcBrPauY
klai0ebDfqRD6mSFddHHxTRgnRWQlBD5wW1Zxhgtw4jOx75nwuFGDH0Pwa6IUKvwRoiQShpDqVEa
coaFGh4qEDElgaiGNrWbON46VVo2Uw434ZpjO26NWU5bTTUz8GhNj+NQ8cM5LgsgqJx7QwURmaXJ
IbcNMjIHLbKuhz2Ldq28Qgst+eXDAEOErHEI7DJ4hcP/0VEnLmmX12GUx4haj7vJ4xdphUI0tduP
Btv7W/Wvx1FprS9Ul/Fuft4g2nWsF7sbPj4X5fRNQXxwfqbZAIlawsFrGesj1zl6tC1IvwuaOd1X
re1iUvLaihLrS+99+vl+4Mat7uDisnMNarynDnh4fUnP4cvO8jSGAmzkQDT/UYY3XYWVO+l/Le4E
8+lVIlzt2/hg1tuyv+qC8cOq7pkaQN0j55dshlTpRsqOjl2vZ1RJbJPHC2Ln6BBB0Izg+Du17vBT
3xU4BsJqO9YveBNA9kmEt9+qMyuNUesCTOQVsPfPhotH/t6XJWb2v5AFXpa9Mz8K4HXgAlAuUfh6
KXVgW2B2oOni9eH5Omk5s2+TtrEeIGgcdOM6PMnrKyLR1KBmzeEghZCwb7kJGrOKSPWeiNzobrzo
4nGC7x+09MRJ1BlbievwMzCAye2s8XwTXsznMbmIs1oOkRz3PJZkKYDSbfAyZ1r9MWQOp6mnnATE
zz1RpIr8nwPSqJZuHDYgi1VE1tta0dwcPy1DgfuFmkyJUFouu3NwtPDrKshDL2h1VHvTkmJTmnni
mLhtCjMZHUp2lansRAF51wEqxzAEkTslXTFQPm3EnaUsHU2aDcdUmvSkChlIk1w3hdDHQVJGEuXj
V06snBo7UZRmMJFFUpFfJqDjkWpuK60SKbPhqchYB3RVk1BnRHRyu8DS6D85m/rhSJ2TkTHlOanR
bEC5+/iJ/A9Xlh1Z15cCfthPcJsRUpf4toYEikz9RT5KbDpOLYJZ4uOyVcSHb7dAyGvD/uPOWMaI
BIHDbnbx9iICfHcqwiTgFpLTgDIUPo1KBZfK+VVD7r3EEmPnXW0Us3jj2lzZwQVT5cU2Tskk/jzw
ieZHyL57KHq8RVRyJbneeO/3rDJR+yXdlEaePfxSs8k3pt/7aDz7MUYFKTT7FbqtAeYhq3yrFoyy
6qlwVloKXBBKnB094YtRlx/ced0QwfLHGIYF4pwIy7wBIPiFlTAIfehjWKs52LG1vW01YTdJjZbP
1rO3c8FmxQ6PH6iUEFv0F5kGbft4EZHk6hbyMrmMt+R3j/87R+i7Kv9puGVdHEMfpPetesB9oMIv
dhnSegGDBqmVqCThgyezzabIl6PUgqON9vYAV2AdcmszMv8XA1febH/C7If/ObCI1lH3JrzXg+Zr
Db0e0awH5OiC3LiCXzEGiBMZrtRb8kesJTD57RPCRHc8iYRRwb+gpK4U4aCGyZ9GEZ86R/UZF8Al
iredwKarMyt98BoMOUWAWSu8FEI3OGk5gGs9Kzh6plyMifehBQnXm1VvfYsW0MnPWwehugDxgw5k
YYnoRaXO4ZD5xoKNtr58ErwTLAI4+HkXbQtNfDQ9+cG5XZxx2kcHlpgAUPlFIraf4CmDDuIV0Bi7
NCxkQkNMQhIabiZmoepkcjbgP/7/x48cvV/J9NDi6Gd4YC+RQ/sjE2L0IJ+OK8JJjUKaFHLdTBWT
Du/qrNTL4NCgX6C1R3wu0DY0SIwl0G11MszAP1F9e7OTB6swNm5Eo6Fm9FBULLoWs3PMLHuJ+AaS
qQB/HeYxI6jTzz6Sn0PegAYMFjAQU6mgwxb8m+bT3eDlsGyhZ9nohlXooZLilhsfy79c0HFKabx9
1mZleXW5SaHjPfeOC78e0kyroT5SZ+P+8AIkEEbttFGw6LELW5DSRHWJ5KTTQqv7Xg1PD4qbvsSc
F7godzQmJC4BR95dPEhRNooqM1qu2lWVI1piGZlLS77D/NsHPfORy5p+bzOg6+l2nZyjO4eugbLJ
OrNZU1+S5W/uUvyixb08Fq6qAQMAE5A1qQh4PQzRcYK2YpEGxNV/nODSG6DImZ8iOo0rHy6+e2+k
nWwTAhwb6EtgVWFq2RTvvYlMNPv+cUQH3X9wSzKHoFyvESKJJHjLJXOKgSe2dse6KbLVgdGab7f1
jUlYTl5N2gz8Hu9u2EZabWnDz5qJbQEec3mHtcK9pK4/5G82hT8OiC1MfXXmh8izjyVVv/lBO4Qw
0xQKioP9gNlHYb1nOe1IW3fDLBfMOrqJ2PFEGuICjIt4qPlR7C0DlfubmmB23J3eScdgaiwTKscB
Jl4TrkfbPg02q7vDpnu1XI/pap6SOmTnI5/6I+0YxbhGBEXVEXJwViYmmoaWqe6NNhfFWp0rM7M7
CBa9LQPD27KX3ugAQzcVpREtZrw9e/4x56FFnVux4EmG9I5jwEoCbDAvSSmqkHAG4qBiHx4d285d
kNviyUu7u+ibbmS1TiQwFxLh/1PXIH2DiAGsfkfUX1gZfEhHdOa8NdWRfh5UmQsgGE7cCnsNn+0m
K9B4x6rBRJEeGGSMB5GXQqK9clwWp37qZtJjeE/SZK32psB/C/QUXXjR+7k39bBELVLJZxwtwCUX
XLallZt/NkOqvmezj5qAog6FqdJ5B6xICb8iC/3AXAi/X1pTRfaZ9KZMrAJoiD0zzfjKetbu87fG
UwvcdE+4iaVIJcatyukv+leV6p1tdRYaRSUr7ceJaebcGpKSVkNBjgcu1kklqQ5C7SwsQtqbf+R/
qvu1gv5Z4VmIwg1kKaoVssGx+xpUVClmw/Hz5w0CsacuS8E2O23DY9HFHN4bX02Ae1V0IAn8BklP
WFq4fB5OEW3MiW+q57BuVEne7JUIvP8iJRXg5olErUvHkEEYIXyqXdAA5h6zEMa6gSX41vIUuW2Y
5zVV7tMGMJ9vuoC4VTVwPYFncBrYXPKTtM0EfDEO1fNBIiL16irkYiOd0CzRfNPuGwq3VEdYM2lP
Dw4oBvSbi2+WA4IsRn659kk7s7Z756WQ+4qR6OFRgSLuvLhwpFvWPgPjfu18yRDGp8KJNVgNwlHe
CTECLAF9GOxpuwgv3CR1SO4wuRCZvVj4KF9dcg+2msveR6sj4fkpGVb4B9P23UpA72aEpXXnlkbI
6D5ra5ABf9iJVXrJHPR/DY9rW5l+XOKcLed1aqaxe2LbKoUVTud6LLWLVSMRMMTqng4oW1vUh5VT
39bZKq8KK52FfmgwzCVrR+CzHdcrZ686GSgPsKLIr1PGWYvgBkRQUEomy8qoWXQxLa2xMoQ97OaY
SCRsBm6Ul+wIppTxUPilqU9s5W2ajJbNRREYSAo39Il3+d5BaXAUfVX5CrD1KR+prucKviiGsAjq
z8wxGBNACA5IsWKwOx0eTTpXSUOL6f4xAXFcNpQypGL232Sb+MHcCyXrsgmK8ul2l1RNlaItQ+vu
h3KnYoOrucZx3N2u/ChnCr6qjN/zqZco967hc1AhypMZ9DDiyphQS0l/7YPSV0LIr8IMyyt4wp+n
3cIfugxDKkjRwZPV9f8eXMJVa1R/LkModf72sI9ijSGJMHX/GT1vaw6CJapSy0c+g7+NqvFHtE9e
9cWVZUfI/KNWQ/1hEcTSjW9mV30rTjaIVO2oBkMwnwFBoynPsD08BFcEWqWzLlIdADN7/399g/9a
q9uGivcNBszzXOvcw0jOFHXW7dHl6aXI0t48HU3SYEsb5To3ioJKMAdu2bslozoLQlQbhf85eM2Z
iF0ukrn104W3EYY3ns9XkUS/Fn4L7zPJMaza9azwNlMeOHnuTk3Ny1USOUuIeFmszdVEcK/dhqRO
r3G5TV8HTM0pr2AJ9xhj5PlrbTCkClQn/KvCDx3lB0iGl0jAdfj8Lyf0Nwo31tWJc8ARJrF3kDj8
w0TOyR5z/0Rw5T8I4fPu0D5+srEd1DVhmolN4RiFj+3x43Bn7jTphp5F3ppwqLsYRNp8D2f3zvw1
VU6VxkQhDcjbAdO+Yz5T4sZ9OiyVb+funuzHkWjh54IBv2hFBDdYjt32ZtRH5pt73E5HdPLSASBH
9Qg7Y6U/PPjlilzgfjz/tIHD6y9HXx0ITRVK6jdapUqSpYzz0x7slnelymjJ3y36/OO42Aeq3YRi
2576TNQyaqTmuafAHr+12d44KunuwPtbWH13jY0AV1XYE6ZrKQ==
`pragma protect end_protected
