// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
iEmPESvCbcdwoc5ZOHjkngS0Zg/iABEIdDsp8N4jNt11QVz802iHphsvMd9QEN6s
ShmoBELFpAEHT+V+FQQf2/Lx0aHhANNIMRGzKKanWVqbfr+d9w93xHIiit0kEPRK
SL2BE2WjfyGkdE6wrKEItqezD3YJCZkYsY9KUN7N2qsf8fcBmh4IWw==
//pragma protect end_key_block
//pragma protect digest_block
XsVlBpGSKc8pWm6NIiXt3YC7sRY=
//pragma protect end_digest_block
//pragma protect data_block
6QdEvlLLtSn8l8kci3JSlRT0eqwpR0+gM0E66oy0LhYUb+csFmjRzR+XWf2i47Xe
XDo17yYfQHMycz67NqW3i3RtaskpmQ5Or/cN9G29XNBZCY4tf0RUx58IzkRy2Tzy
AD0tIXtEARZX5OzaY9qLHNZpKjg461Rjl/9C2FdL2NUptNYASWIrzlo0/B5URICA
FGLchrhRUUxPUR5/mMOVY29NhEM+9OER4L55/r9F4OIewIF0FRvVFCEaC7JQ6XzC
rVAsoC0OWM41iozlG1V3y5iKNBO9v8zIYcuzqVXnbuOxGZMTFED7iQ5ShY8bZ1D5
CP7dJdipsOOFD3CFeLRrcr3TiTCchG7loCCSsuSnGfioMoKR3ZDpfsjHpZcrZzAf
8X/fzMURYwp9Ds5SrKmpZUMRcE2uDLtzwQ8JsesYNoZe4FczuF297Us5RBg8ZwWp
B8Vxo5Yqw/1ioTdYXAbOQVQoq+bxEDVZdyBlL38KMJahFA/CiqmPnjW6PsFL7DWt
63Zk8uhyleWxcMwoWAo0GyhRR7EoTLd0xt4FM9FUAHtgr+p5P1JuNkS6/usvDmVv
Xh09WJMKAl8lv6PKMNX6hIJqfpjMWtFX6ovJSiBVfiPz8emod9xuVqka9JPEKcrG
Iv+vpt8luNcInKHbAwEwtzf1peDr15+kcUn83R1qgq9QxjwZ8srwhP3QzsWfbxXe
ks/eall9V26cTl+9PRLjyk3INCXwRqZo3m6ViOw1zcHSKGBa0cqB/zp6QCBhfBKu
oB/0VG4mGpK3/FiaibCUtOQbcr2Pz1TY2phZFyOKDVLnBDXi551S5kPDW3itw9mH
vV9L89lnJjcS3q8R2whoitBNuwE9MfXoRbo/kqAtEfPCBTU9wQ0R800TWBhD2xao
uwAm9aRj/R2xKUoKeLA5ylgtOykvuGsLu9kIHHzBE7RsprWfvI0rCaR2JSDojhGT
jBnGasTMwCzQmxd9xARgc01XCr83bTZz1OGzcU51/+b77THo7aVUoDjOPjRY80xb
PnVqlhPm/EI8B8HzXsKmVAAtOTEnSY036tQbyS6ile8Qr9aAkNcneGxZ2LChD50Y
J1eL4iqhtnsYCBopfufGMLyr5UKmhCO8WGyoAkXu+XWXpntif0xOw6bHCgZvVTqW
jbPmxkK2/UIS7Me64+iNDTPtQ+ZXvDrQBMStHQHXWO5KWh19/cjM3AybaTGWHVuy
jrBkPebJQ0wCle2T/uHSk4YHb27ZxAjGohZDXcx+mqP9GN6RWSa4FGtys5xT+N+a
9ChbjpyK5nXdY4GONDv4uEAALhUxkhor38/zbHuh0mZDu7eNKPgMyKnmA4C10sw0
80dMN6522QZVkszK6dGsGDIHKYOy2rTbrhISyBcBSCbYOy9li4pwBP/w8JYB7nzo
V55JNXWpTgmwZDSznC+Rig31xAPaF0db9R8nhCHNIdzz9W/hiwZ66Tc1GlKVGnUC
7+0LyTpjvW/bo/gmJc9oWQz8xd1XwOSK1M/kppLRAAfqZ17+r7bywL9FkIbaMtHa
ZmUGqZ+F2LNVPylAuhMPBS4YsTtsRip23b910fv8XyTidWejCrkiMEuPBQwc8Tu1
Zuj8N9anGtHVqDIMLbcEzJMrZYdJ7GiHA7BlC++6EahvY7cwLBsMnLTRLc1wpYbz
pHSWVYXiUzULBbZMEgAFKWv9e5CRWdvLwpgzIDYYI9iNIbeA0uRtkXBGhy7V3pFm
EJ+ZsYPtYZvzAa464xhT1lVxsENiRJqs0TmphBlL09jwefNQzip3Um/0zao5dYY/
l04bI5HJRpS6DX2s4q2D9IZUJ+JvGGOVai7yyuhnymLn1gV1Sv8YinTxCFBkP4Nx
SIld01Pdx3oJRAw1Ssn7ij2Tnk98NYYZbCHmLAL+JtmhIRPDCnBsFX9H8jShztlZ
LuEhAGdGUmswzUETCUQVxM3q5MxRryVNOSip+TF0YHhGxlJNYFeE5BeHgBWJV975
ZrH9UrqIsKKKhOI8Qeyx0IwgjR9F9YzJD2C6RQL6NdhgK9tJpA/4f6szKv5ZpLxW
oDrp3d4ArGRHyv91SWEmN1LrimMwVqx25GhNUp/QzClbO3uudoIwuxSVBq4rrlyu
xAQCWdxdC9aAUXTfhDFcdRewHRNspPNSwNSMgZBfHSxelrpri3YNRvlGeh55MUrB
nwod8LSIYcQg7IOikq541dEYz32t3zTnZgc0nnM6DwYuXaSV1BgTsq86PmmYhy8U
0+8HSQrF//I8GFzZDCVMUsFIdW3mUpu8AIJ3UPVfmseyf2s+pl1aiPPQmCb+A6V3
afBQzLjo5fwHZ2e80vqAf/RGbMrH84//cztDnowrhTMBJIatBMKir8ingLpbE2OZ
YH/u65xqQnk1KZxnmtJuj2z09oUrE6LlY3lzGg37B1JubW4f7XsSCvReEfam9xqu
/3dZvw0UAd4004/rlEkF6DhS0tXTE4D1+VbELE4qWNcWov82isx8JRk2cfPU7oPX
GWxXnMJIZGTtiPRgmHqw7NwkftxL0J45uxY3Vu58gH1ZoqF08hzekIVN9QIHfUz2
5Ym3GLX2b6ubUMipklgEENDkWLToX9Xv8YeAtfMfzvzEYMORiM0eoEMMqPGQ8NqU
RzKtlR0MQ8i6rcYDri9DVHrQh/K87mNEvWkhLDAKkvE2/gbq47Js6EEoi8fjha9z
+j/QQh8Lc2nu1/ZOa6HWdL5XC6hXv3F3iDXFpFy6x2xtXjaDdKSr/mIDuc7R3TM0
+IgI4n9o4WBTrAam9vc7xyZL8/JJzSR/AQ3onsXhvW5PixP8b95dgLJxj8FkPrGS
y6RMeA6VqqEs2VJ3TMVRWIh3VCaOCQ6h4umCxu8ED0gnA+z9NIY+iJ2C/3Orl7Yi
gm4qzUxM9S4mYM3F/iEW1yA0ZWft75J31wvmfj8iSM1h6tSLpljYSwxlZL0QE9NF
ylkL06k1IJ2rEORR9Y0Z+S+kw7C6zgI5zPmo7dz2JE/VCuPiS3baRpb+dqRr+Haq
sHjnP52Iid4vRHZfwxw0vQ==
//pragma protect end_data_block
//pragma protect digest_block
UW5eTSmAuZ/WUCl3mvqZstB7gXk=
//pragma protect end_digest_block
//pragma protect end_protected
