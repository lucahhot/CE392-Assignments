��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�a�ȝ똵�Sm�5ϟ�nb�<(����1��Ԓ�F5��I��(�^q�n$G+s��q]��``�+v�~�i"Y���1������ziE���Y.gڊ�8�ke�W�i8u�{v�)kV^]��g�=_�!�E������W��ZjJ��0/��y{ŗ��%Xq��G<7����u@�kc�8�P��̚�w�䔈�_��;r���ly� ":�I�:��`û�8I��G�}�.h�����G�s��a��3���:=��sפ��$��(-��rD���v"�LPm��:^��?��b5����Z��ҖWJ�=3-v\�{$�Tnҵ����i��?nE�m�l��^�t�*�Y2&h�6Lr��z8L0Y��{ֱ����n:����$Y�؏xߘ-bW�c:"�,�0{(��	:�����`�Bx����(	J�y��{޶,�+��پla9�]ˍ���,��I�
������G�M��J��yёPڇ��l5<�m�^	Z5@�iw!>y�Tg��)��;IX�k AեЄ���01п҃���2M����I�R��ۦ�W]|l�N-�H+���}��b(�u���`#����n���� ǡ�po2�r>V�>w�|o�8�Β$} ��&J��ajUj<�{� ��������5@g�(cCԆΞ���}��rg�c}��� SB�,9��V}���]��v8�mB�X� V����AE��i�+�^�)m `Ea�Ц1d�m�e�.�;�Z/8X}�6���Kנ��Xr�LqQ#��nceV=C<�ݨ�a��pfJ����f%|Q ����5O�����7�Gъ�p���t��?E��U�:�C0��ƾ����k�/�BȐ�����%����w(AO2��	A�5T5�D#�^�����
�P�SB��Hi[3D#�W�0k�B�J����Qa۠J��P�S��\ x�h��EzO�\��ӭ!
g:�\����Kx�C<�~����h���.TW��7��ax���+ Hc�� 2�G��Zy�g|Sq��c��e�MA`A���"$�{�'?��ܷ�*
�YݨA��`f������H࣪B���Z��vTlG��ѻ-��)6p]����8���[^^�x�L1�@�恘��p0�U����+�g�, �ި�|���bMˠg=h�?\�2�:�5�.8}��'n�����f��4]�/��чʔ�Xb��a��p	*D�aA����q1���e�Gh�#��\���_�N'�ICGs�IOly�3zG��1��V�c(�OXhD�rl)�6��<b�b�4*�ο��ER��~� ���!�^�&�t$wTߞ��Tc��1Z�S>�x�tq��a�k��$L1¦b�=�Jρj� �w���$%'�ֹ��9�r>�����X�_�~>��I7<{��t}�rh.G*Z:�)����f�Z
���te�;��t����4D����n�?���n����F���N��{Lĵ���a�K��CJ���EZ�E�,�W�B�s�?�|Ƶ��FHd���Y@���K���j�[��A�Q�y5%*>O�BM�����:s˿�%"�!F��]��p�	E|W�u�Z�m�<Y����hWg!z`�!�p�� FK/�A�R�Ʉ��tU��!17z�A/�`k��G����=������3�ͷ�0Gʏ�_�ÓW�^�S�?p��D/�S�v A�[j�e��(� ͺ|�#���2!�5�7�)��d�Kb�bWeYø^a�������Gh
�s,t
���� �����������Y�en���yn�U�Nh���ˬ	�-̨���ԦU�5��7#����ت΄[�`��]�[Mw�5���q1 ��ܹy�W�!$�|�� ��[�FT�HE�1XC1�G�NQ+�9A`��n�r99�BT�}h�O)CvV����1�~�պ��hU>7��A5?$��K+g�ds�;�"��i�Kj%_�,�}���H"Z�'���q�r����E��c�M�r��s�,�Z���vPE��l�<�gwL��}���Y�甥���G�#�N������J7 ��H&"��O����q#�N�xY������m�]����hI�y�_�� ֞v^��}�8�d��XBh4lx�CbAm�M5�%��m� ��V"3� �T�Se�(�J�A����,x��V�+�oH��Ⱦ�^3�T����5�����@[H�-J���5�T�Z������1:�|j1x�H�lg8������k�\\�;{� ۇ���OS�!jadyu��qI����pb��js+v�؋�����ţ����(J�D� Fӄ|o�~�١e�.�H�'u�ā_,%`Հi�b��\wa��W��{��Dm6Z~�m�+i�U��a���[��fh1�g���i�ݲ
�I����jX����&����h�nu�A�_^ԱWN:"*f4q�= �����En98�Η2{��_FK�tw�[��S���,^`�R�}M�w��%7aw��,�]۹oչ�~�)��;�2��Af��+�c `�k�I����(w�� �i���v2�G�aڻ�d��y�����We��i��O��o�.��V��D(���%�"�2�̉�U��b$��U��lP�c��=�X��j��@k�L�MJtm��]dΥ���b.N�)�-�O�>jFڽ
�q��R��v8�0Q�vKa>![Ds���L���*V{}���CT7���!/�g��!F0[W�I��8�Hm�a������8#ǆ��ywBD��Ɉ������W�])���e�����4��,m�dߙy� �T7w�5k��W�!����mj2w�� �j���c�L�5^�ש�h��t�IS-nR�:����P�D��6+LG�^��x�C�D�/mއN�p���l.�Ŏ$H�-X�����9^����P���V�c�P��{�I1�>�蛪�"�$��?�]��ȍ2p�Œ_#-�n�T.���ŋxw2X�-Z�ãvf�C���d��BA��*���Vi@�
,��@l������ �Q�� ��0FR2�o�:l���6-[WdI�F�����m��X<0z����f�M<Z�敳.�e�/�鶖�Q�p_�='f5���Q|����N๏p�jq�J����,<;�~H�^��0�ڂ	$�?yru���(���%�2׾o�u�h�&4ǰ� �Bd�7\/q�p><��P�������]��~ފ������-���s>y��7￳?�3�p�����RE��Ad��"CL��\5�U+�1�!P�_H���v�6�����ě$�_�j�(��J=��m݃֡;�����P��tVN�^�T��/�c��ܗ�y�Sqe����)��o���B/'o��y;GHͼ�f��08�?�WTg��f�R���/G�+�0����8�ڇGl��}��(F�V���̗�v��!�@��	��7��	�Ԝ��>��dg$�'Յ&MO��v3Qͮ6*��|;J�|��ʌ�S�6�ψ�$��ҳ+�.�,>P��|���� ��UR��v��7{��������-�m�ӈ���f,�8UXђ뽟[
��<+ݠA�(�W�[.,8�lB�\�������rܪ�ϩۢ`�@,nv�GŔ��L��_CعF0��݋�D�Z���ߍ/��Fhh�e"e��`B�A竇�]�^��[")��'��+�z�'�6�t^�����>�cg@-�)`�:1�{�_�Ǽ��fF<��|
��Y[ħ�k��]V1R�ڄNՇǾy;�*@	�^������<�i�5�Ӌ��5�e'��{�ߕ6�71lÑ�l�A���2W�bP��mLh�u�H"�j�9&O<W�|n����Y�����r�ז�
D-!l��:3����#mt]O$@���>�Zk�k���c*6v����j�O��߻�F&!;���P�ho���*��v �|=����2_�O�>#.]�q����G���[��ܠ(}���G�|�?��kb��Q��l��U���I^'��Q<@���>N:���(����P�?����Cd4�k�Vֹl�����
�ME�?�k,7_DϤ(崐P�ѳ� �ΒZ3ٝ��3j��ēԏ���}c'�^ǥP
���sO������S5��A�ϝn�w�e��<H*�M؁�>�������A.� Di.�C"�0�S�����a�s��+@O]"hV���_�d��e��������N<�c�;N��	T�u�����������Coڟ�J�<�Ǳ �f�d@y���H_�-d��������~��G.��t�m�\*�6�l�@jO�� �L#�������e|y��x� r�����9)�B������%䊍m���1����1=�P&y��@K�y� �zf}m[�1�z�T�3^�	���X{W��{l��h�M��d(�k-��5B�"��սI���}Y��v��U�h����-�>B�!��*�Us���hM�o����m��:����{L�x������hids��՞]��o#���I���	�9����_�DB�ˋ��3<��S�n�):�K�R��**�iZB25�
a�ߘ��GJS`��f���]ޛb���EKdY;�����Y]-��&𒨺`+�z: ȷ�mn���)F���}*3 UP�|MÚx� Y���+�������Wq���j��b��W���R�01iZ^1?5"�����M�aJz���̈�e�Ȅ��#�a�C�Hqǘ�2*���9 <;ͫt��O�vl�ݯ�X�R���k��
�y�G��=������H[�dj��H����F9�a�A� Um*I��z.�����[�@����d_��;�/+���wۇ�ּ��T�v�9������(��g<ڟ��}N�(�X�hj���U�?��학DO��/k�f�L�m�����=u;���F�y�0�E�M�^ߓ���,��ԗZr���5�n�J8`�,<1�:i�=�$�PY���*��4�y�PFty8�G|u4w�Ko/���9�U:i���Z�賅��`�gGz��R�T�d���O�9��FGra�
)�ev���v�����ӕ���$O/C���b+~�H�/'�˳w�z�vZ�%T�?h�[��;�v}�Gr#�\�f%Rd&���$V�_yO ��ve/�NV��'��X��"C�=�M����kH��O�V���.�"�P�ua`h/m �.w��_�ۍ�M�z$�^lJ%^��I��N�{�#�w�'ZE	h�}�:i��M��5�8�%��J��)��*B��������͞׬dQfV��WR�k,�I�<P`ͥ�X���Tf[�2�{c��:� �����n( �vJ���}��(I��	ɑ��:�@y��i�Q&u��^��6&���xv��r]ѧ�%����6ŏ|�v�cԈ (-rڨ�J@V�]g\�)�&�
�@i��ls�4?�O�F!�e� 
���t �|�u�)׿�$���u+��K-����0���(�6��F��d�/s�O��M�o�iz��RR4�6J��23$�%8^��*&��l��Gv���to2�y�ՀGY�j��Q�[�I�ү�Q����J3�`#��� ��~�Ł��;�բ*��*���P�>�zn��f�u1���[����͖�u�M���u�zH;y
R�!���b���9����E��p���W&�UY?�ɞ��cy���Xw�P�:8+�΍<��u�+x�S�����6�� ��٨W�n �y"��,�R�y}�7>�s. \,���y�Lu��Y#�g�~x}�e97Ft�.��Y>���G�]U'���4����2WT�����8jATO�g����)U��bF��Ǩ0bc��k�#� �^E�;�̗��h?���p,���v����z��h`?xO�t��6�������[��"����6hі��[��[E`n�Х>RV[3��-Ms �Q��"V��\�DL-L��t>j������U$����{�Z#��*�lL��ֽ��k`����E���oA���S;��M�?��R�lQŌ�KȒ���}���XA\Q�
'%�r�`@���g$����4������\��M�\���x.��=�60?0ewE�yZ��Di���y��Q������~6Ώ\��π$~������;8���#0G�oUނ�3U�i�7����,x����7K�� ���2ۧ���H�r���%�ʷ�9:�L]�+ �:D��G�_��=w����6�ݳ�}\���Aɦ�8�zFu�3�6��7�7���Jؚ��^~��4õ�I���t6��X2�J��e鹬�z��گ����^ez�ܜy}q�v��8�%�U��I��- ��cUX�E������e�v��P�@K��?U4-,3���J����jj.� 8Le�"��׼ov�$x�����~��+�����������.��<��AA"�c`�\OL�δ�	'Ϋ1���L����-�L��Ed��67��a�%����9^�(.p��p:w6�#�!<.b��k���l��hk����k-���f��WR�b���DUW����|>�&�%,Ԑ���u�x��TÝ�6�嫺ՈEA?'��pW����*9��XYpOE� ��!�F��X��l�'�i�^s�PW���O$��3�S#ߒ؈
:9�מ�p���5R�i�P�=c��fkXyX:�{R�ږ��^�T��As����lj�����UK�F�jS�3V�Oجˉj\K�䖃'�)��֏FGn����0ưG≸�qy��t.��qM��_*����x��"
��N���>z�A~6W�_�#�D������T4�B�]n�B�Z����x����.���'3wj�E���dR�r�t.YF��|�R�MK;����Ըo���0o��U �cl����3��#~�U��EWy��"�~����xOq�0q��z�	q��7��x�4X��I��
AC��Ç��$��i'���@龅y`�B��Ʒ'a(cx6�yd>ZrO=CS� n�,(e�C��1��LGC�߉4P��{l�Y"G�⑘NW�$2���C�B��$���h�2G�`�D۲���6{�\>�mB�F�����}��V��ix�<l��E��&C�+�y;������F�(L���MZ�y<�S0i���͑"��1ba�0,쀚�ÙPI50�\nڭ�R��YN�y�8Z��,���W��uT+���o},��3a��� *�v
0���?��𙬀0�c��tGx�SV�V��X��<�fP����Yr�7~Br��Z���Z�q�#9u1���K��t'��3~�IbL�j��6e�u�#��#$���i��O����p{�|��-���C��ԲsEr@��Q�%3j\t7�>�b�)[Ȱ0�mZ�c� :�����M_)B<����w饻+�-��պc$䝿U��r��D�Ã��PFy�����i�q�D�h�v	,��㕽�v�^�ERSQJ�\���Ru��Y�a�U�{ 7����n>�"��}����Ex�Ů�Q�[΄��,+Å)~�l��8^Y� ���L��ugA��q���T���5��iV>����5�9Z�t�Gut��-� Qz�m��Y#v�~E<��b5D�-�֗D&"�tj>.�z�n�=a�0<7�
B��X��9 �N<��Z$d��F��-v3���i���`_2gj[D�jPJg֞�
NAj�M�r��ip�N��KY����v��w��k�J�;�&/��=��v�%�E*�I�y�����F L��l�P0\Q1��^�}�������}�ɍ�{K�G�k1D��c:��>g0�@4�A�*.��w�����2I���a�f��Z�t��$��i�^��gjH��h�έ�� P���$ ��i�6�:��=���ĸ�qk>��,��ǜxi*�ק�1&`d�LD~O7���"%���	�ؖ��H�W�6U�A� E�C�j�����X��R��쒃,^i}���$ຮ�Qg���=W�Dg�09,6.א�ֶ�o"`k��+sIP��k��/<1�C�~�H̙	Y@�?�yK����{��F1R����z ������~y!��L~ۦ���1�wC�w�(H�v��QwX:�M�.m8В.Gp�8֖ٵ�*�Q	�3�%\��JVGe�8�|oFģ�1� �-eӟ���*�¿�3���x�!!@�����J��|�5��1y��\�y��0���ߡS��w�Y���)gv�U��oh�dƌy�3�{�CO�~X���������´*�t���1�E�jX� 8qhI�~�� �B9u&��:�}����sv��2����-ng?���n����"e�������?���`���&��T	�wJP0ę�9S��͔������0H^N�ցǹ��B�>�UK�N�29}ſrs��#cH09�,�+�6S�}�����X��rI�6��`��"
�X�DJo3J�f��*�����!�`Y�<�\V��G`��ui^�3�.7�����W_�����b�3*�7J�;����yQO�BM�ō�O��h�Z��sU�4�!�>x(U�W���kg%tu���מb�_w��&���c^io�K�p������c�M��:)F\ S�����i����3G��,,��n�Jk��@ǃ�|�_s�|�Y�G��su_A� ��v5תɉ�h�s+���?~9�ߝ	�H\,$� ��~�η/1�w[m��n����g��b�K�zȄ=#����RH��+9NQ^+(w������m5���ٛ�Z�2���>?��Z�5��4���^�$�VИ�c���c�r��캏*��'E_�jw��/
C��2S�ϵ^�KY�m��G�*5Vl�.u�C/���6mW �\{�`�;�.Hݫ���pO�%Z�wϼ0awJO�^��@����s)����m����ևtM�p#��7��d�k�C�p��<?���!���AC�2�J��!ߨo�-�h�O�������);̐*S��9��	�����}R�B`����^���v`�U�Ȁ0�e��<s����b���T���)�~@G�B�
��w}�C� r��v���o��M5�����TYAC|�g!��W\d:5�o�s�hY���A�8��U�g�$i�&N�M��+ZX56I��|	�(��Ν[�^q|H$�e�8��*
ock��n6���I�1���z�e��VI�n��з��l��ğ-<7�����A�����	�ϻ^�?K����#B*X����Ou��qG�V�,V�c��e�C�S�!@P�?� �޿J��p`%sS�%r���~&'��^�j���"���Ȫ������[�D��A|����IZ=��}�ޣ4��L�[U��CMh�t�~�}2���y`9�I$`�m��G6o��u~g�5i���|�3y���Ɩ��X�U%��@��m�p�$:����Er�o����!(��&5�����~������-����R�i��Im��C	m��A�����e�r�LjA��	���^�g���jf�ڢg8�)^?� �Drxj�l���KF�2b�%|�1��k����K[dM!� wҶp��#h� ��c�m��[��M�;��L�|��y>B����CCE,>�>�?�����~5b��O�W���c��\��T�,	X�C��(�8/�1�q/6M[o8����>WŬA��,����������'Z��M�M��rŹ�*�Ffl�*+��6�ٌo��[h`Ɩ��
�: ypocL*�[zfEJ��ƪ�w �mx����bg�����r�ϛ�g�m޵؆}�OmM�L�*.r{<�s���I⻎��}p�ؗ����"�:��a�ڬm�$�]x�� 4F.B��|`?7�]iƨt�`�a.����d���[�[h��|�+��42���[�˅���$���'��?����$�d��>��n����ڡ��1:J�]i}B>�����T�������kF0,�)	L��d�p%O�Ԉ(�%����,��d|�"�}v ����(�����G��@�L9����%�l��%��a��(�a�9���	�'����j}IE��/#mB����$d	E�������s��<H�Q	`�e+��O|>��wR�U�ܖ�����[���cg�6�a/�cM/˙�666=��@w���UT��pe�0�L��C��4@a�b�H+^���Մ��r��o&��H���g��� �ˇ���Y^� �1=�R�T^r����l��S�G(��@�>�˳�gm:��i�@%��>��^/� ��]��1(��=�(}�ӽ����9S�T#��� R�K`x������ޱUoB�%�"͗IK�PSC����P�7�O6�$6 ��p�X$1����>���U[u���(XX���[lb{*M�}��S����^����OoS�K~&����m����+{�dBF����7k�c�[�XD5�B/yӎIذ�̧@����G�@�wՇ`/-t����^����� 2܃?� ���,ͣ���3kG�5��44���24�}K�����,z|��"���;��Я�Ń���P��}\kY�̼��޻�L,�N]�ׇ:��H+�Z
dҥ�0KՂw��m��e���SlX�ߴ��b���b��䳟�,A�*1�D��d2�-���D">�J�,����I�{��V�F��N�r��t���B�XaS�����k��7�!��HQ��cw}�۾1<`��$1`9�aS�'�EUuWE�r0xorj�4u@�2=ɦ.! ��jG91�X%�]b$�� q�ɘ-��Ru3��3 ����з��̮�{0����(F�~
�����\�ॶV3h��i�!�rql��=��c�#d��j�͢Ɗ�qio[��p���H�K�.��-@#j�R=�n��F�W��f<�X�;�H��v��옛榰	�=(ۤ8W0�[q�,R �a���Đ���|ۜ�!|�\��I�����[lk������'!Q�Sn�t�션j��:�	4�/&�G�l,�;���w���v�r�������#[�qI�N�sX��Q/�NU�1�����{'�/�h��
�|MU'&�E�f[�=��%��>�:�zc"�G�ޜd�{0�Xn��P��rN���Y��4�e_s��*�C��iU7�����n`�W4İ>���"�fpA���΃th���:�v��<Φw�_��2�9Xw)#�T��b�3+ۡv�岄̭�M��n�|H.�ܓݍ�z�yH�dQ�> ��? A뉞R1Y}�����Ɗ}���r��i�3}��vL0LwU�Y���̘ŻB��Bm'gH��)� ���y�2PN��B���� )��*��\�%_��l���P�NI5S�#Mfv�W����<�H�ʔ�(~B��GFܒ�/�k��I��^�^2���l3�A��͠!�����i57 �
u�yy�E#~>𤫬�%91<\]�(��W#���Y�N��'��y�t<dF-��-��씞���qq�G@g�D(`�+Q)�i�(_A��0��O�8%�t����o[�kE�<�3�#��2ܳ� fU�S�����woW��t�i���f�7W�+�շSշ��GW�G��nx��d!��?v����0�����Ɂ����f����KC��+��?�'"��%��)�����l�?��A�7�n�~�xѻR�0�9�;v5��=x��pu��2���eYk��)���)nd�#YR������7*h���u6�I<m|V�}
�r��B7?3�A^��[�>�$��A�,i�����׏��\�Y`��J
X��'��W6��"�ئ�̔U|��шp�о��]%YL[�Wʅ��+-��C5�ɡ��u`�{�Y�g����*����4�*�Hs%�����1Ϻ�8�O^X����&�����f&�\�Q;���~zj����nK%�0�B����Vh���n~�(k��pü$#�����|��W�i�g��,���ZvlL~x\��i�4�;F��缲`�n�O�N[^oZ~�@��i��L�s��q��,I��*4a*��F�if*�ۉ�"��d��?�L�������NB�c�ܡ����Ǟ*�=�cDU4 
��	eC�Lt����e�2l��@F�Hq��/�6{�w_pO7��=-���w3(w$���X�s�5�wQ�H�D"X�2J��np\�`�y_fwR�f>$�7���x�,���5�=���wum���tG����4�M1���AT���m�g�I^9������g����ѱ���.�����L����_X�d3��]���Yԫ�L'�  ���e��A�yR�s`{��o����@^kg��d�&�>((%Ѩ�&��TYk�|~�\��>�v[Q���I­JP�߸��<���	4L;ܶ�]�8�(5���gBF���[�x���ӵ�X́�& ��|�h�A�v60��?���Ī�ܧư� b���	�g3kw���G��ϩ{e�Rԫ���2<V���!ߖ���h��"q<�,�nV촍���Q3%�e�J��UA�d�Z��)�����j`	%�V���)�L�l�d�rG����8Z��C��ۮ�S�tI��ÕcyvOi�.���%oc��%��x7B��MN�cq��UK��E]!�uj�~T�/�WQ-�q_����h$ܤT\{� ��H�n�O$�s��X$���A�7�=!I�i�?c��)�@���3�֯���8j.�T����A���<�u������^�ö$���9'������>j�9!۷k�:amo�i��2$��<��s���Q�^k1O��κ�DY$S��/ �����<�a9@��0*�>ͿM��2�¶髍�E�RڦO^Y��޹���8��/�erU�¾,� ����Ř�[���xß�=��������0A�E��k0���9��vw�����w��MfT����)���pF�
�*E��V�Ta;��^��!4�)���f�/W��:7F��m�@��l��Oa��W��"˔��\�v���dSʂ�`�m�h՟�T�����&K/���kϽ����$D��y���ۇ�"�F	����T3v�!� ����rj��k�X�4�`J���0t�����9>�PDlf'&p��|��y�x.�T�/�oPqK��a�\T����niP���\
�|�@}�h
���;/B�����8N^i�->�Ѷ�Jո��rf�JAMf���:�G}V�����A2!��v��Wtka:�Ǭ���<�U�>ؾ���n�EfN!����}����:<7st�Qv��粬�OF෮����������rk�r*�'jFV����f{�e��)n�|��(�CK&f
��0�g?���B�����0�Kۍ�	��V�
���;,$��i�ld���ۛ}��%������gf�{�:��2����bC��]At'�ݰn49�5M$>�h�@�U��+xE��8���*LA��\� �2���o��I��