// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
X6lDLEJGQlhp4sTWCFjYaBa7yFm5igsiMegkTkl65maCPDvyP0wDYt2I5w+PYBZPUFB1LgbMEy4/
hgtgtqgCgGhX+yU93r23Iri07bQZwiE4VebyVHmVIPDTZ3eAebdA2vf8IEs7V8Pzby7d2B26iLDl
7KFyu9bQIBwG3K8FY5VnJfMIV9KgnSlpp9KkKj0lsXNmNmjuuwzShlvIqJ9stC54ySvmDzbsvy7w
vHijbXC9xY0w5FdbVMSnTUTeJj+m1U69SzqnCJAbF9eE1gvo5zNT5AwXDgqabJuWaXP3ARcrKGDn
MbgHNqdqO7GVCHq81t1tdBy1B9DGdHoasIkhnA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 98688)
pJRvXsmR3WGJIaiJsXaY6XnZfRcHh2Dm9QUfCBH/OigNn5sm8h/JzqIDomFpHEt+2db4a4fXNKmp
2gfqTjH+YhwtJTIXJ03jFpMR9QH3lmko/wrSHG8+9E4ACIwfE+UZZzHf5si7blczkjpdH5sKuK4q
zuPLX/6blBUuh/x69LpPmf7uwkRPqCHxEFANFF+fwOsPAb0kJ/vefc+tvv1BVJr8sq3iniK05jjc
BdXhDYSE4SkHYXDPzsMFc4JuK60WCt6ZcdGl3+8zyyTNaA6X5gJoLTnPvdParwlWU+RFm09XN7Ct
hKVCDNtypB+XSwtLjU2Csid6Xfjn98X/HPR+HvIQwLBALVJGq2q5e3/Ky0vUPVPyiUiv3WXqwodq
QL6dArP5QP3ntygeyiItR9YPR71NzXO3CaiG3jb3tNUeHU21jwNyWNf5p1nFPFRdSIGJw4loYaX5
NFFhbmXNL++iQRIsxxEsZaJGEQXcdGC2+N0Z3FY/HHJAGgDafcrFsHJbnwRMcyfu9BnBrNRgsSj4
5qzBuLJRlOfmY8B7kcVHW7/WjcirIuDDV+UPtZl3pEsFpevVcuNtZo2B/cqWIR6DRLxScnPtwtBT
nJbr0lftZ4xuXu5/gTFaesPhQUjTZckAazJVKmgbWXqUALTEqVof+6z0g4NTdu+rjc5XeOYUhymH
mFHCrahaBLBjgHHtw/EXCEh6FksDe/VE8yQqyMKWf4OMSU80RcDdSnavJMlpKg/rrfripN3WpfFv
/apQZEQlsomadP3dE4vc/MS9bxUI3980C058xQFXX3NclSDLI2eLktgly0ZOAh75B10KB/JjyaAZ
RldAJt/TIgOMXv2MvXwBOF9ZeuCL1mcVVvejEqSPDs3+E34cHe5V7CIRdikYbsVINICOwBhrw+Vx
sMDYsxABggvW/MaCy5CN5lxM2VgH+6vAQfrcgrxDwz6ow/2UfuWixXwuVvjYqAN2hoMzaWRMnwgo
lyrWrFJ+b8KpxaDfHcqWAeRolAtVDOu3mBHwBisxWMyB0nuzW6ay/qWhQKziz+7dABJe6MMg40P1
vdDWJVfSoGGIsECH3iMkHTc+th/A6SmlAa+rT1R+/vW1Zw7/+Nv3GJTD1Ql0OLIONbsxulajDhKa
PjH+LUO6VLvlfr3wRp4kPPyBvYRs16/lPJE+eckWjp7hlMBCHgzvmzPLnZWORlh3twTJy5VE8gud
yEnHJlTaK5+hf+ugfaU9AGo/clTE8BaPdJbfMreYjGCJj+KPsaJII7DS965IUH8QUYO5lbTmMp2/
3rS51SvtArIks0pRo/mvyehzicsEe1jXKnsd7gggZjzL/PR7bdIbzJR8L4MoWZq5NeoryhUXZx08
e115QLkd9CaTLjqeqiTaYCnztX5ctUwAMmfQo8SbOmxXfy8nmku1IAKoOVZPRPuA84etJDuMZKMo
ZjAffIEFsJiyaLHW9Somf9ApmwZy17Dcl4GjharNM1XJYcZu/QqZIwtIj6XUJEGFY4jc4BsFytVt
eH7Ji/l1Bc05exFgZ7jjQR5ovIH144RCAZcO9U4A/xZRzlZ0envYY+Eyk+7auY+jZ6vosXTw029g
CooByrfnqLS9hC1lpAMnR8bwiG1bEBrp97zCYw8BzD40Uo2/lcdtbENdFDZKtGM8TO3hbS8QkXFI
d0MGtlg28XlB4MNQBRW+/Rup6Jo/krAAd+JskRj+5cZnDa1dWsdUaqrb6lmmKWiuBYAtjiwJMeLa
ftf3d4MeQM6ccLr1NXAd9I7lhR5hhtx4BYnFqBx4CCXkqRxkxpbaYAjKcSQnmLfDwX/UjCWMVk0o
0oLFaLmj5YIneitYn3u7l9rlmDWjgmlcaXgQrX3JfcPPuoVOFFmr87/V3Ksu97+ed3ecm08UxZTK
Ib7p6xTzFBp60Ipxvv0wiofQexBhfRQcIT7eriKTZSaSN2lZhJ94McF2ENvBNYZz8rC/KnN9A86w
hYQd7NJGarnxAjUhhoXIPP/+JkBJJseVag+MyWAnkyNhAMoXqygqv6UZQ7FUNVSWk7oatGXVuFf7
Edd77vWf5+mQi988nHjjY/CHz6hRucN29+QVZyQ3n1XSSZ/DsnQloBV9BmCXTyEb73fNU9plRgyc
h09ABfz0MxEf4qR3YRK/MRQG/Y7SM8B0wwLNJWhGoiqSOCFsQc7JOHYJmNeHepq4XEnlowx3AQAw
7EqArI2m5TsKerXUYXgs1R4CTdKseTcSVgBGOEK2O2WEfKogA2tRxiXmjCmqadXApQkwKcTyttjH
tZKEwn+OTlDxnwqWXMEZ3sQF0u9nJ9O9HNEEp4PqQ7yhvg6uEzzEAnEiG2FSOP0VzABWR49truOn
On+VlIpvyLgJQQfUeqfwTnLUjKBXdaGjczFDCu76uuaPCsV/Mlat9g2dswNg+OkEDIo3Tkt0Gc1E
+pWyL8Wkl7e7a91Agmvvwv+DIgGQH7MTrAzUUnNztqLjdg43TG99JmAZSMFtsP7xTVN0rfusV7iW
Wsg/Vh2qzq8EIw7RmgH7voawS3cWGAffDKuRwDeFft9a0+4OPj9v+T3StNCeUZoiFVVsl4Ze9B6X
hmkPZel3L2chQ9uGgpTKyBeYxnIi/CIZeKxE4Zxyp1KElLp+PLx910DthzFsbotdQgyvY/qOlx9O
SArK1e/ztB+6MHKZC7fmQyCn/RkZr60GQNDdrJ3e6J+4YOtjebGi+4HtMDigrO+gd+N1+FAnE7HJ
zgkdcPeqRdWnI1mF/i3v1fqQekBBUMYS4LQ3tYkpQgUD5ASNTOxqAsM4HrTzZ7VXpdOarZ9Stydz
9nm7O9DPtUpbWa915ejA6l3/j1fh2U+Wh3gZM0uCCIM0tRjmFm0onennP02yMhvOq2RPQGaEcUeP
iX8YiGIgjPtZaoZ3JOtEjABF4Y2cjw4WBetGlnnhj07YDxMAxKRGporBSa/kQbmrsDlA5EBPAIo7
ID58Zc+kRYsZ3/75cMXzIw54It1dUC8IXbRD3yVj3DUmsx1L7LIT9bR9rv0pNZv7hpS3GwYB+DpP
viECp55KC21/qJ90soOEGiyd8yevodGYQrtL7tHeiz7ujHDTXmZ3GIq6MRLamnFVlwbr8RIbB0lH
vGHRK+4wn1AKPV8yiW00n/tEHHsYCugZBCvo0NEBAg7DnVby4+kKbfFxVTtNT5hKcDcryDImMrTs
vafaM2x8Lc2sFKdMikmHFEIWdS2XIRhnJNvjUNeexVxJ12SvAk+zK74qrUvrFt/Et2ZvMtQYSjt1
aYSoOXkgn3LAW2ThNi3fCau+qe/f9VixmkQUD2pzI8ZwqxVfM65GFEm3SSgOnk2WruxAL2Q00fip
0ojqHtsWXnl/YxxjlzfJNVvpbKFTwOh58FB1BtnIejOC+gQkDzZrXIGsahE3FXehJ0yyxmYB5Dhm
IvDmxj9NxU9gRM9nMvFc5VD+uxxV8omhzlvs832DtjVeObQENfNZ7AGMgZUzwDVo9W5OPefZ6yyG
6yPHS77dwFZaiFBkTGH6ZXlGhHrNd4GYGjyprzbOqA1qMgGmnxjccpoI1585NfnlgQaTzS5moLB3
fTahY/0lTPeXr2q9NhTQ4d7ERi1SXG80xnfOdm2KIJ4X9hGnMyJ1hH/NUcV+5js3ax9fWGJGWLzu
7MAGNPhqn5xMu9uvOuOTq5J4lmT7Ka6hPcu1afIdxpGVlsW+ba2czroDVLjjrWOO307g8w6eEUep
Bw5C6TDN0mFpUgvTRqn8Lpg/71q8///5qVj0SEkAlZELmPYhf7p6Fu4TXr8qz8hL8gJdMHLACwmg
yO54nkmXA7KOlusbf8/gO2jEql3d0HSJ/IDHYDKlVA7b3r8T8K+/4M9wyeCX5l6nwlEX85mReEpN
9pEIxj3Do26pkd6q+t1FkrHA63p2LHwhcfMNL5fk80CtYs6oneKGt020je/gtXRj4eh8efQ/iFKH
sww9StFJUC9oisIfYLI5ak6DL719xep/yK3dPHHxUiRu4KtsI3iGnT/B3sfKEYsPKS0jmAUXhVj0
eiajvpx3zdzf0lVLqiLftPO65Veaq7+hOospPVzko2dp/4I3A5gqXnTiKTNYn0OG5Lelu8k+wIT7
lNQnF0f7sHIVGcPj2RCCWXjnEYkiN7m8dCZFa+4Iskdn3VDNw4mFiU8HZ3sIum+5iCKWf4GdH5Ix
+RtWTL3z+R1BjgJWVQ7jOauxjTi182C7AQuPJVarMOjhU2ZYEY7R/HHMpStwyLNcMRblemnGTvVd
fRuIyAR8Mg0bZESyND/K6L1QS8HQgp81T2B+PfTV42CLyuxcRlNS1Rpvz101WUI7xrFFu8MQa6Lg
BUm8eqOq355QfNHhCBwIDLIjgQzR8yFFW0d1i9xtMGxkjrVGz1YBw3Y93KIhlxGfOu5ZhLM15HiG
k+TmnGK0WrtOpP51kLLqY2LGQj3cHjovNgff1GMrP0dOtdkTArLRTgN20zda0pXdLz463aE4W2sD
qUbnGgXbASFsNGz5fQgvChdStk8AOktkYJay7RVlhYqfVETDJ8/ZBq7SdwAtxw/J2kNl/75/IHJk
YpxbGygsfrIK6NZSAuT425ngAn8kxqB4+blhD7wc+ScCAH6YgALeQpWD48Zgrj7wKIX9I363QdFG
qcgWwWVMJMFAAWu6Qisgyu08rSPl8dHW5wzuC0Xowsyuh0kgZ12LOWmKFtYLRQpHZdffEzTg2DrF
eqLYaB9ZdxlVeLqiCJkpjGDHcu8glmdnhhoSPc1BcI+sHYdMqCI0lh3MH/SVoTKo834JqJGssFwC
GXqncifk1982FUPbwDfsnbZji3+bewyaoPdOGi+h/80qBB6cbD58RRNkemCemm2TmtVLkvko7MZI
GJRJGZUOUoIdSiozB9ogtlosNoY4Am1CdiRGLJFhCKx5C3N1HI2fdvHMNA1jkgYD5k6nI5+OFB4m
FZs9282G/xW95rrNc1O0SxEWQAEErRfswLTv9wya58MCkzANNcPHQTnn7u6s5A7Rjq6SJKZOGTuS
S4sweawbz7xfNZhmpfokXxS9WSIuz7Px2eLgKtevXyiMZ8DEMY8XWro3fA11jUysV3OBOQbWTAcE
U1zzFuCnlHeYCu+ofbRPKtIeoTZC33AsBPh8me3tf2WH9Tzjr2+QpidRG8gKcwRlmvIKPRCYIKsh
SVfqUEqMly3NerzYSrwnnK7wOxSiqf/mVbq/FKtyiRMBTDKWPctU8Hi6ny8gAB5dNsPOGW2uMbnB
FldXteZsdwqJSF5M7CJqCDtSt2MjUbcPtSbk8nxJfLNXR5+tYsT2wflwKK2tHcQtRU6ZjrpKxfag
PakG26YUVwuDaeYocSTmsyP7XDVixaHKiQfmt6VbcZxGX+Jvai/bU5l5hmz5r8DUvLV6m41d40YG
zd00qzpyFb91VeGXSnIEifK/V9XsskEp53XhIz0QT2VUVD5/Tg1YxsRzJgAvR8RCoHFR0BGgEW13
ZpD1aBr+D2w9AdPFn1qqIvxXf62asxb7EgUmRUg5gVsg2dS8WQd2rnr3wXwmxLXp0st8GdAfr01Q
vA3j0Hby3k+4lm6vM7ZY7K6np2yFBd1gNeDyE2CFyPxBCEiyWsJK60nhFiqCkzKSH8PTy3oP48Vp
l5lafyWutvmlxRvySBmp6NuwOTFRR8p2nixm9vipieULBOtA+QwbGw0LDmyKjsKxcTGjte5Yz86P
8Q9314mMjj5SodmnqUCZIp2Mcp5lsVGLQ0LydBBdq0k/9TvR88+wTF4i/gtX0jKa4ZHq71C4Wcxe
sZjdODoKA61hCBttzV695zYBSpCaiRsci3l97Zey/G8BjRzdzMrIUWWsHFo59S6RQOYKIwaPZK1i
ffNS9tjpCULnh9zxAR4f7gOfXbzshKwEEZyiDSnMtvKp5O24DxGDyVH0K6vJnApSlVvERIp/XT4q
TQWbeIkc9xWUzCRe7RVb+ZrbUO9aJrbJcGE+newG7GaxiLT8920lnIwqDohy4kgTxl1nWT+G64D6
Ofu3WFjeLTwWXEToIcKWJslOmEgCH403kOrm7HaticRb6WAfJkwenvfkF3zcbVUvXzI/jMF46JNc
LNySeCgu5Mh+cFliX5ia+IooZuSzDTgCphX9yrhqLxP4Nl9iSoI4+GEA/fFJt71TdVDtCZGfkYag
/ZkYuH0nkT0LOCj58mC96rT1OKYEv5YAJ+CeJq31pAe26Za8uAXE1Lc1qtTgEeQtQF5lh3XJ0GmS
s4WdzWJ9uFhX20Pa+zoWxgENPBte8LnnTBDSAkIjZd1srsEwWHSAStb6VdDtdWYz1ldEUxvl5SpG
l4SvS7a0FLOWv5E3RKMlLvL4OpYjq09K7n5c0tQSlzkNDsoB3Co3dUBxt2feNwyMXus/Jo4zx+Al
Xyu0H2bQw3mwNWWv0WdZAUjYLb0m2xh5+Pd88xFFtIWu7IzcIk9ouCm+DlVvBKZV1Q5XsaofS7gu
DvQZWPfdBI1ziLm1ehxRgaoSWik1eJzV93niilidrzJow1V3Q9yMqNDTqV0/qg7yfo4OEizuY9h+
nD13GthmV67jjBqVblXOpshPW8u2+At4is4SoIft/erSmw+FVjZqaEh89yu3M2gPqeRgUgJapO/U
pES3T5fg80rB+eRYVfkRRmdPNTlxcajrvecWeuPkddyY5zwgNgCFPIiABXGLRy+METeFHC924wED
qHtu9wJ36aFUS89yDRfpNvB16oQ0eHeJzgNAqz/1p5UY17EWgkHzObW5qpzNRpcF3bNy570zsmmU
etV4witBHJnOtVNx+LzCDz0oK7AR7qIT4bc1CyXGc8XHVcZp+MupzziGKWwNa6Z5oePcJQmmqvmC
3iELEt68ESPfl5huc+adxMnzLx+wDO+qxB1Z7Jrm4iclqEZ245FciPl/wVhEEf3nqyIvv/Z865HN
SlFatrb9oSonptPKuJhE/uz3sJYRRQvRHD9lL+TWSkDnB2TJwa0ArxcJqbimjqd1F0ECaHlW7gd7
y+6ayoVq8kE0/jf0fpev0yXC9CdKJIGhysliiC1qbzyVmZU1PEnPbzdL90r9Dah312Tz+uKBJyGP
GCrZJsGpH+3mwod3pn4sBiYhyzVkiWglwCSMV+lHjLBV4Pa5/LSyM4jzssCznNC8Rk0BLa6dSn6V
1oggZPRo0CxU2HUt2g3KbReNQ9QWHcP1vKBVnBum2lFcnvGxDhSO/mI4+ogAeRryHbqB6oIhKkGf
KYahT6hEMFsKkqdu3xYsSdUlhlf7ldyoDkhfppT9Tu0vldyY1mde64oN0/Vll+PmhbeB1bowuqhT
MUc0NgsEn9sqISAvfXYUXTEKBvRD9Mkc2U1i2srZDf7YA5/NXRPuss/3JBDV9iTpy5o0MbfRrAyY
PD6Yj7/zpO6QLK+jmPuMfAJyc35mgI2GlRp8XWVrDTZErtGNkZi33IcQGggYKXzYujIx8R+07Kun
j9rC48g1ieivq5WGQUIbWHTq7DCkE6fgAO8/QEIz6p18oCmUez9xLsOdq7FPNiyIan6Skn2FdSZw
UQ6tDOb+OLbzmuQHQTp+8EJIpGYm95ouW3VE/kO993y5dQyFIuKiBB2D+ezUf5SMnSV+IRE36StI
LlIJ0P2ZkBYgDA6TympKt41nz/PSP/Z/97iSixS0LVy8gS6DkW60QvijoStZYkPXaguVCN02cjm4
J9y3frm2YVzcowS8b8nfQ2jx53HvDy79T11305FeVvDKwVpTZ6yowshOKbqkJf7DXC+G3wvGM3TK
t7G+8YGTiKC5yE3g4FPhcoLdGjwLJUrOY+riqelVhpFNjzR/55Tz2smX77KvbqcohJxpH6gusUoT
Bkqmbo9W70IPOkDtg2Gp5ZcaHAo3rrQk2Dj8Gk5ajf0OUOnCUNqLhdQI52lFxyBIPPhyFAwJtswk
eTo7oc5PcRt+nhFGSptaN5lpRcBVcm6r3gPhTy2lUGY+fhxhwdeAK/SG2z3LaIdiRRr8p8n6hG3s
FQejCIpPQkpwigvKaA84bq0vvfC1DIvjUyhdjHjEFd40WXmBK96rUpJfshvwH8sdJGkKm5HrhhT+
guwuZfsEyjbcWBTxkB5e+/tBBccT5cSuUR+7pZ5PIqEn93IhuFW8JjmdUjIGGE4nT2cthY9QPEjR
sAEjM3aYH7o0Qa8HQ7HTfCd6xXjntyRa5M2EfrxdjfkvUAXI2NmXMRi5XaKNzxizWqqLyYAA5OUv
btECkkISAWHeYoRTJt55rXUDTiJKEboJQJZ0lMSAgjk23MNdPz1TP/S01vAFF3uSj+sicOdv7c8K
LL8uwx4BKNENJsXgRm6SIqUgImD4SshUoKLp2H68NzK5ri4wDwNx/6bTh6oJCKTzmoglCVevj6X/
7lkBvEvhFsr3h49k3D01reyr/32g20HiMxCrFFk+aNz32tN+/h9qsX66ONtz/L7UxrD5pugN9n7y
wBMjRv4SvP1zFaYHsj16wXMm3EZa48KT2TAsn7zUFSXWlSbFgdB5RekV9UOiCQ5XdlgSy8b9c/b+
y3gtQVDxHagDJpAok0WkvKox/vIulKdo6pRAMBigGxGZGeUUx5BDH9m3uQKQLqj2qlJ7MlCTf7+T
bPVvbH8T1OsrmhKBdaLTc2OHyp9nh7kTWEqzV7JGlZckUNc0kAG94lCPGBh5LMOzF9LefGOGt2ZJ
cWbBJyec9uK/DrajekXQaAXx1tvSJV0BI4NwKIIVdDtEdJOpdZfCzjOnZ/oP5FnMyAumvZbw7fAh
AeZKRHBywaYqOXFLsrEADYwi3JoRriuM4Mt+BZjrxHtWtJJDFtIOxZoqgT2k1Zc60bvfcPAHJWvU
237fO7AkTJ3HXjJq0j6W998zkzPnQu1lQT7QXdEeXueCj/QuKYu/Ilz8EwfIY+b8n4RNaWMWw0d1
0p4PrcJziziAiv+h2OjLbaeLe+ITOz6TwjTBDDSmONr92Ka0RQrM8VpZptchR4OWaaJHj8zuqJo+
XMtxjvkhGnJQM9B63HBIuGq3LnKyMbGJr1391o6pOx2j0f3lhbn8MyXXU1nMbeVwFY9tcPGLnUTz
qGXv1exmN5X/ojpvQlBTXnKdW99bcZSieYePMNa3MMhHY/cNzcrB43MjKXd5dDr/4kt1/X4Cd0Af
98iW0lScjwulzLGu3wsiCJLVmcx2YSWM82TxRXBzaq31fSD5KLjhZaMzi5K+h2czT/3ZvL0oerOc
PJr0jnJ5QRjO2OxUA6s5N/3I8fGnHiYR2XtI2BwJO8GkQ7vY7sOEeavrRIRf08QTbtGKyhSQaVP9
1vTNclfa69gYE50PV+HVyYfdZdRfcfF0ouvbnLbIUUqPhSAYJR97uO1bCFC9vbSTKNodvaFEIu2W
EOAadnQoMuvE3K1NeR4I/+u+Vbt5GZLLt5y4z7JXH3leNuZb0JKt1P71CFOJ497bKc52QWL5yyhT
V5uHyq18eOy3kcEcwVY13lZTKQjO+z5N6m3Ry09uQquI9YegZGRUMjxMNlGYmhLLdZKmFa4DQ+ZC
t7h/v7mWDp8LioRr7sW9nwxKrHL6MG9kOFgkWexONSK6CsHpp9QxASQdP0LHwVhcrmuXkc5N/QZB
Nc41AexhLiMPqvtVZ6DANRLEjRKX1DiH2Ca7g3fBIX2blP2dA2rl7CrlIMmNugIBaNoK8reRCCLt
56roIc6ZD4Ysko8lWtsx4voVwr+YRHPOl/9MckPLVGEcJMsdjaRM+8tu4rNdJMv/TLr5pZFPTEVp
O+61Ea0q6jnH5o5AUqn7h1vjziOt2byEYsd22EwM14miyKjORv1R6fPviZ9Y+D2vPQc1MwoF558a
b29kLgRfX+y89aZ2Ztq9sDbG2z4rM7maNi5rmz3sQfDf/tKjSJlqWZX2ifJPWXNgWzsRpzGyRKGa
dEM2fyYiCV2fs1lR1q9w6HjUJxYC6dO4hg+eO3DlqTdBeectIXp7BDqVt3qYbn5LZTN6BNjfjASr
rt+5AB5LdF3X7tUhTi5+QNfeJJbAcZY/vr+o++2JDH2ygYRqE0lW9SQrd5fXXE/h5bpxTKJW8rWI
uNIBmpw89E/oRHcn0V2wxpqgJdWtkFoAOHCHDjDdqxZk/26VIOkFAuVifCXjuftycPwN5+Yx/rUg
tIxMpTSB8ZDoc5j7LYSYAnpPIyF1fXzP7M6nscALH3uXiUZRxcJ6CoR0X4WyNtUi3cT/MVqv6BYb
W4bbduC+GAPMyrbKAFrTTdfOnfK2Iss9sWG0lidMjh9+lTEZk+ZGIpNi/wHVsJ/WBG3spBEp6pte
xoqp/zl9C8cXBHlnib5AU7OInSijty+r8JMMSS2ZF6Avh0Y4Kpoh26rBBWheLQBplLn7IWupzxBN
nxg6tBTMMaVXAy3eD8zkwkEHoZAMrfcw6HX7UdLzW30VLkEcSFOjFIUenUKk54WQY3QyTY3Qd1Mf
VJV+jnef6qf3Qu8lflO9QmbwPUKaIRMW72SyrhR87+AP9xqG1uCw4OLeQW9XcpFhjyG81OO+29xf
xJXa9Y8a7OXCr23KeVeLJv6pGBAC27unySRGmGPd5t89LbRMHEP/Ay+4IHA4NoW3W2qUetPcUDw5
MWRE8dMknzxAlhr1v+zeslNm5DfoMQdbesOSNjxVmiVN/8XMjUbNwwJOxRL1c1MjkLcmxgc9W+el
UgJZeSzJ1D1xufuNOnVRg0ioDT77yAtYiBcgwMcHbloa5n9v2Ctnk0GuhwJs344blCpZq8XZWGD2
PsX8KqAzsYnXryVSceaUYj3FUo+vnX8Tl4zDhbANfjdhGTL/puN/Acw0FtnIOh94IgssWofxHOET
1zBkQVrlS8oN+iOgndJ5f3wAgcZFn8IsI5Wnk7MwcitFgp/hD4kbPONcGIiE4fjp8qh/fY56m5s9
3eDKIuHnjoXNPcF4Nw0SFoewb5fDq9eX+manfV+lKQjtybSMdBCdxYohhwW9OANQ7L91F0ep3mYR
CKqXKpQMtdjZQjFi8Eqp490je5T95BAbvmo2xROa+zEf81m4sQgdZs07ycvWNJiesB6T9vfh28bX
M8LDIy1d0BBqutZcwH5xeOYQIuVlXnkx3yl2dS+x63lL7S9O3lcmwdCO9t2uk5VsiB1ZnkyUUWaO
0MT2145Bzv2SMBSuca3VJeKVRQkDaiGO792LRYnYrNOrILEeR7QyxF3GeP2miUEG4jDY4Xa/JXBw
j6d7FXiy86lx4wnkciAb/ygodk2XMEigpS3KOKuUvoL+271mcaO/ka9Oangc1CqYzB2Yie08ZTlV
xiZ4DttmcGLhxsO7/sA6jFSU8AxRcG/cCgDSNjWfZiyW6s+osOFzAPPnSsoRQfyJjkYOyW+JFVbM
RFWyVRb6WzNrwU/qbMdfbysm+0NtHyp7YAHgLVRWmbAhxxed9Lp7ZIntcIqf9AjgR4bNs/7T780r
qIyfSygoY/NNq9gIPSkbd9UDuHF7634TOy4jg1snFcJvfg7DTul5xe4PjS3A1P9m6dk5DGrxbYcd
5oT73H9iTQs+kv+dLr6hFg22kVSd2900BauMLmKwA+icYxSYizIOr4i2m2olFJGzKmkAhi2a9zUm
B5B4JMOHvt5BGVu81g8f9LoCDDsdOzV4lq8RTqgbULy7ifn6Epo2uHdtvJMsrqJMPbjyds+zH9gr
r0CT9pEqXMtO4Q7ND64giwo+Nxvsf1B7DnwDkCpkq1BWidH5u1HsC3eTXfmX7gVE1Iy21qVwyAsF
b/Wc7Y8haAV5VdqhPm/7oq9BqnutLqxN9jeDv2HvwpkQcfmL/5Ymq02D4w8G4aJtVGpR4c7nLXAt
cGqdnDxWlwT1xlhEwT4RcfXrSvtfhtEPK71Qu7vknpR1YDyNrf+PTn+bfviYq3Nh70epEdrEl9J8
nCfEJmd/25j35hJfxfI/iXUuNpv2wIFLQrE62ps9B2qILDd4eGg5exmb3lHvUyoXdvGaiXyxi7fO
frbHH3yrlwlLlaFH8SBavSRur+DwKAPzpd372PHbJgGKKG8ZFqGcl70TIo0QGBQjVarO46bHfchc
xKaMrpsAg1Ooh5FD+psv6wrGVGRNrVpVY6DMRUsqMJAlBLC3hBBf6JoPNRLBB4HKb5uEHcuyDEOP
JMsxrzgdl4hy2/zMe88Zz84F6qVV/9G7UDA43fJVns2AVTGHHSCTSVykAleaGu8GnCArwFpP6itU
hnlifScel5EVJspzzL8vVZ9GLJDQ4ZJttyMKLcMQ1HZI9JbzbjrM9wxs1YNYEzHEN3EIhN+Kex0W
x4juLMtm9f/F4lyrDvdaVUq9MzQHSY6xfDtvl8du7JnpDkCrFw1ZVveyPrc+uAolQm0Fv63ynED/
+vPZfL304VsFXftBKX0Up8sygyGr3uiuyuBTDPOkuC63+sulFEe01kgZtGlFuIYnqUmEAUK1fFzV
LBTdkT/9eWB7N9YaxCi1iq4cHpHsf+cvcSFZWgYurkFy7AXrf/y+RIC2eIDOZpMFCg9S+o4FBjp1
/GVzl74hXdpQXbT05EEfu7phSabI045uUkDb9AJgID2mJG7DBETonDBRtNkOZIKeOI9ZwPGaFtzt
yBy+nFXWqjbQOhunMyTgPQi0yLYr5sZlwZQhgeFluvng01bBLQvbEBe7NTVLtB1R/Ue01EI6CgzU
DIjCsbVnNMywxEm7eYhtG+YUFttKB0DxwRgt5uzblKs5ZZoF2FaBisMhXigqluTh5eoZ5TXU+y+K
AXZtgYkzrz8eteGGxgLKvsspEbvKt172xObwRXzThlW+0xId56czXQm/J5IJkto96trGma9qHgX6
2OE7mzj28cpFXDYhXSe0ftMnmjP9Mv9JcxpD7N7cjvUnLT3YGaRz/dkv1xPY0wrbDgYbc8LhGY7m
kpw/R1fV39b4hVtsduONMjPwVFkJ7J2cKpQBC3vtqOSbR7ZhBxWNXbUcWOrBL0APmQ1bPDMJaRV1
7L04S0DmKDSf7RiBosCsJbnDjSUSbLHJOvnF4QloAvx2fx4MP6q5Mx5IyBJhM6PPkqt95UpCgTBb
r2O4QAUGbmvE95zGRAoiuIqAM8e0tAINNwdemE/L1rTE79KJPfMvxnTCoR4S8nfp2SSro6lcQxjN
nU+LAHbvw5lPET/iOeZUITeWX77D2jCKfL9JfmCGpppfrHBWGXQhJ7bQS0iCZaKl9qLCL5QEjjSs
EjRGdG1VCpywm3gyny5t5ledaB/wP4kMqhsyFc45yzkTE3mhou3EJQbv+OdRtGQYwWWBe1MIoGr8
8jJpAjc4z1s3787X3oFpx/BhffJYggBgOEpcU3R8B54TDIs/VREszMG6d0+24FGEn6qVTON3f/BS
ukUZrKXPu0aW8rNnIcc7lseobVP7KKIA+Klmg/YGZFZeS3pIDmtIuE7uHBBaaqpLD/GBjC4BHQoC
ftoHrRHq9438BQdplgW05/dQXv7RUjeKdt4hKGJWrqy6x4Ngt4BfDQE++6FxgN33sQRu44AMMbmH
h0Jp5ooPzN2dOEcPVormUB9xatbqRWdiC4ef0Wq1wxICyQSc83OF9wB6i0rAEOKeEfgkKaJsmWe4
q55SFaSCSHTyYafx7zyDTg/sYP43DpASwTqofZoWvu9Z06Dnp1Vu8byLLwuArGTt0kHYV5QrfWN4
qYcdYGL2bTTem8C2dXwsujHI/YT8r/Kb/M9DTv9VEhWeh1YP+MXez5gJaCscoDMido5dBoS8AEfm
DQW36xlZEHa54HnXRYCTHkToSx469TXCxWScFnN1IczxKIiXoH3Zw2/97uO7aYNrsD3Ny+cM1D1o
7UyIpeMbReSqHf8iPVXGIqq03af3s4HPhdMHC+VdXJhlz97gjdAyFP8COBIm1TnxKdqqkVDoa6Fd
/37WmI3so/C2KjpLdxuOlA5EFozpzliyjwZp4TL8Z2Si2MXLxZQov9e81/1pr3QrE3ifoXBjH8Td
WshLX+A8bZGgDNDgFWYHdwXiuY2i6uj2vAT2bhbKGx0tZEqN1a3mD9hyeDQHeAwHTDHVlXPD9LLh
9FyuroGj9rz8hZvElEObqYfEj9LVgFiy0KZaoGz/BjM/BsZSiRc5Bek+Di94kPx7DjoqlhqlDOP2
wDDBJKNQtFzhDvO5ec4fRWzwqOPbluNkAnLwfiywM4H6SHwm9wK2gRuv05GuFvaB3gXQi053zTII
Y6OPFlYgApttqMQFcLs84Bs4zlMMNvI0g69JtVNUStNmB/VJiu12b6T7ZbxDiNjreQq6MwOB7/X7
MAvebpLofhDR0RxHFt5pLdGseo8+j7vqlPsndTzqchB7ZFZXT8ne+5EUt4YRLK1dlAqDI2Ls53oC
4+1ZCPBMRgJWIbeHOT8kliwOhoRA/N19tGIwWsa0O23dwYm+d1dmwtL0ZejPat6swjNrzqdRN3VV
AR7ltmqacP0y8/LAb+x9qzB/s6ubll8vjYMe2Pz71fzvPumzJJqdxJmVfXc99FvvCrGE432J5/NB
ef2HpnhyqeAIXyb3p2WOVUKmOMJ/kX+dbP8raTDH9fDkMk2uJ86Z9OWaLQ62enXr09sxLNUei///
tBT55AHUXhvYjNwUMaoGXcvGHVwn08v4WN3GrWU8erccnGJq/S9MX+11R/c6d/fkiUHEnMgtKSuW
hd0CPeMDMjLbvlEkbNLiPn7l/XPX6VffDwwv7efczljhIQN7uPRPg00fVUt8yL+MaLvejeD4RDyx
CL6tKyL33ds7f1b6Wek37lxrNle/LMdO02ePDAyO1R1+iwuabbS9l0jQnVoaBeaxHP1SI7Q0H2Od
f1K36gWVsh5QakeWOrSYHNZHNJRf6vF9Q0Q/i6uS/mKot9O7QLua/T67dexHpFMyRc81NQyoagrw
WF/O1L30rRfseXgDTI1qI6r8TyIYGMSTuAD7uulTryKsiXL/DHdKL8xNpgNArQilr1FAmVe8lNdi
YiPRz/TARGOIkOw+M1NFrOv6Ji/sH5IH5HxTyrAowekN47VbWo3PX43y2tgyl0jJKnZ4LYnNkYvz
X84Xza2fx5d0f6iqDU0V0Dc9e/JpNRXir4ASVknKjHANl9/CsDTTfVayOATeN7y/sU9yVzpNOtpu
9yK+H+NGghezJjHPZebSficmVVzjtg0jIxPLnUW1kXQuqq+QUC9b+SlmnHEqbnP3YpFNGAWfD+di
764daX+hpZdtACVdyhm5IKZDTLXrmQnDLU/F6u/BHKpwxep5R9uGONpCNKNfdszJp11kXWV7vGDF
y3LWJDiIYK0RDaQdSHJFx1RYBEXoFlVuRBQI48JX2HoZlSyQpr9NJ5MAFk2CX7DJz28ZWAVeDn3e
IA3jN8Qa5rL/pMafE85pjwlye2r7WYWuiSS6jrrfuf/J2fIR4XQFT5PRd11fWbrpPIBjpm/5OCxW
ZFFHRLpqtsjrxS86SUwH/G3NBjeksPKPZnTnkQ/RRnKwENt4Xa2KEDUa5ajg5pak7qmCWpbzXir7
hXbdhkA7N6AM+VB78z2YgyjA9uibZD/go1H4B5l/JnvPifupQsKYbtkDjoMXuc9HQcXYDf/TxO6O
hw6F+MqP2SPPXq99gX/tw4FqfBOpwWC76hio6GWlnTrc9RDiFa1Fv58V0jSJRFiGnZeIafUpexeW
730KsehYTqFm+04LgcTG71gt2OshpwEW+jsGS2gYdYZ0q4bi9mtNjyEZ7hnyW3Z8uQluyG3FeW4C
fimWbqZy8IqkNwW5a40PADxiIYoOV67W2IKh+MmZmqN+4YpQS0UHmf7djNP00euMmxpIR/P01kTP
f7c7nbN0bFPNxpx6zs4kQzWg7d5AGY/6L4a0E+RxUS3pCas2/vAfQmoKjXxdJNi8HggneXi8/SxV
SVvlZeTtsTkdCuaBNJX8l/DR5fYmUpOmq7wuUaL12YWYMdhHCR7N5ADY2RUY5jPZzgnYUdU9QqrH
GwMaL9TUGRohKHA8GffNYK4WWJpSvxuFVGRfVqfijnuOIMbbaUP7nBCv8A8cW42qHec4eM37/iZg
xOIY7hxOXFfAxrLdvZHRcGzqcEvWK4aJDukvs7rBXrgdL1s96pHCrX17nqgVSMCxW8oJoWhPE5e5
3GELNp1JN0W5ySumJ/56+0lI20bf2T9utZPyVtUaSjdpMp9rE2tHyDcVMJmBlwt7pSKbSOduDJoo
8Ks0kIOUQKWSBTdnHnY8ve2wFMgVaa1uwZbhhn37hKEkBLleijuzDuS49BFtOULmKHyNhI2hlz2D
QYVzccqonMGCOS1jXHx5cDMGhl+Q2N/Kll0DXGAEGp4krEHeEu8hFABY+BPcgJW49DMIMqKcWTz4
NKDv/bKMXM8Y+Aphjye7l0JDMWKNI11GHIlz8QhfrXyISIaSJrXXMgIUkGmcl/XouwjmEOrPSGKy
6640UaI1WeUumclUCaC2O7kS2pODRwdWbJFhOGsDAkiDTNrzjtHUagzp0oZbFK9pgXWtSZDmMjOg
kKOr1KOCCFjFRKdnj4Bmw28/fFIATCDozonFbXR9/tP9Hx8CWyW+ghnPCY+gCMvDBwt0mvchSuJR
cccBI/+J1GwoVMF3+qX9HtRjUASncwSeUSQjpuH4OKuMm5IjP4XsI+Uvb5ZAKBS1MSjj4lR+gwJR
luolIYVpydu+BB5X98ldjxumbI2ntfyVaH7mX2zEKtF8Sm8F5+JHeOFydYF4Wy5F93s+T2bznH21
ut8cIhpkvQbX9WRRAc5QRlDXc4BADN7MDcQO58SpR3F2YqVBrCpYnya+VVgif2QW9JLhswVVCDU7
2etB5/L8rpXD4iW22+98rA6SOALsZqMMfBeHrtUp663AL3YhR7FoErBDT1edx+SLF9lkqiyEhj5p
vdu3y2Mu5tnhKLioep96BWY+5zdpU8Rr9YNgXJupwspvX+Vx7fSrGeEr+nKFBq0ZiMj1EvBSiC7H
gGggXjM60y9PWTz9bvMQ7ESfRTMolNLWUKI3ayYuoFG90U5QESZ20uHanz43wIELFEg8AU0ChHfE
YjTPgxhKAoLWNeCq7ndFsnvQuAJViaFPVJ0K3RijhFDUgp+gQAIl29hKKg5pvcN/sBcqa0P8/B6P
/8Dhd4qY4bs4kqb1ZTlCaVYLrp63QJK5kdFVWZWaXFdv4gyTWMlyaSMWNWLq3jQqfOdAB9LJ557i
DYC1tLUacbz3RthB0tHg1f3loQlUSFpK9pt4XaNeB4Il357GiEzUebM68PjPjOAq52U+w//gslnN
4D83qBHwXe56NCJlTMghFrS5qw1fh/QEFNLVa7mB99LLqbbiiJyA6pqPTtOv6Fc+gWm2ZS5pOlbt
ASQq8frkyhKFYqOZLhg47LrP7k6XKL694qcgOKaPkyrXq+HhdDxhR7+UXy/BqPlmTi4uDtWnreaT
+DlLuo4QVfhHcSblWOrcdA+2xrkbMMiK2/mEaA7BqVpiLen2keYyTZQXR+++vh4kYFd1kIIEO7xt
DIQHYsQ5p4LTcFQBK4cWxQ+oBGukRdnMTYm8+pDhlATz+M3v/FxUQEbHJQH2ToiY2d6cyvKUQnfU
4Pu/b+Kao8N7CSmQnaFb+4aCpIbVJs3ZO5QHbAHoePoHERnDzGD9nhuHBebXsp2VO2LUBj3siLj5
f1X7mjZuTazTCieGRveBD14x9mvS3v+8GyQ9ZQnro8mgGh24fkXVPJncUXRgq0bcRPlcfkXDqofY
ipaFWxJyNhOkjpYadZsUQlu4hdz08q8XqWjhmb6eQFIxW6cFvi4s6rsTmaNjPu6hLjSsZQX1jbIy
uuIa2sajADJpMRwCNtAo2t4HblNBJdczmky1ucN/11kSEyQsVENiJ1y/4QPiZtyvZf4BAWPpElA5
satMNwPCtshVFRnN24/lnQZOPF1BjufQhqRRcCREg4TwpsHpIkvyri8BXQiK23m+nh/1G73tNxCR
9yj+8iqmMbujzUba7XVTG85VYSfxZ8NPNd/bXSSsbMadkM26Yf1L2nCfGUhY0pKyrJxePX+XOyu/
LcQqb61Xd8Ru74qMPcIiLGjUx92Mte3NbLzVy57f9uALOLwN8fpxzTulwwhye/YD3FotzBdMDVFO
/XhkjL82XY676lhNNr3yaP4ZtzQUZy1gOgNEqZexsrH5IAyHErcSuNXFiHFoynIfaMyTwmg4ECc0
tuVckGIvxEcXmohu4q0oVpblw2E0Fi/6R6u/54D4sjlLGBJO0oG0Xmpw7uwzpv260oSq+RjZ9j6e
L/EzNOAhrq3+tYFzlklkAtFqxFvH0Joqg2xPQtIZjfL+JAnIZimFjMaQNvzRCPwpJejBbd0MKpl4
aSeSRR5Y69llgOOEpA33TWR01OelwdUH7DSlLJfGOb/TM7AIVeRst3a8TGM2NkDkLFcrzdsSFpWX
EaLkAZgLOTs/rNp12ybHNcd9C/QRltw4R+FMMDaUxVakttovaDwSoyIg/PV6tyIp6oa4Q8oEZUfJ
VIR2z8voWLYtaQoWTvrlQmzokGIYloTK8wcUiAEhxUNpUQ7GvHm5gdgD0bzOrN7w4paeOtVMlEA7
7vcGlVSsoXZwz8VH8pkDTJbWaUL6arv/ReQLkwHxX2fYoo8zp6RHAIxf1eMnda6mYX3AXIpCGf/6
RN6dvFJPrBobf9PVto1eyBO9upwuZgh12JPl0iTS/UrRnpWuA0bDESsbAsutBDJ6nVvyMgFXibUM
eHuMvB19DnCMj6Yl1QcU9IGgvb54QPvCb6r1maSj7XZ8KkW9w7F4RhwKXwM2byZxaSyUBGXvom64
yGdIBuTlORiwZD+xcooOh9d+AEz86NAzCenNeeTHktvvQllB+ML4jDtj3y/YMfm0uRTEFhLpqNOa
T3IVYhwd2sHSggOaXgf7kp3Hf7QYCUC6B/kvRYJt3ckxJ+vtrX1eaEnnLHOGl7zeSik2pm6EIQLk
VC1t2fePK+u8hLUJJCq0N/K2bEnxKI+H5OrW3EV8l1R4R0YVJRrRwIWjjx/7OoUOzZ7cVsW8STX2
xoT3SMyg2CG6zFcssCmcrSqKW39cCjDpTfxL5jy8xlHgn2gpJeluBcEdL/7Ng1uVUEwxm8M6y1kh
lbYVTn0KB/CgoJmtjuBIGhusqdk6U/7xgmijtW+J1bjkotzofvpFEBXqsZs3nJ/4VVgZrDzAHn7U
MQpC4/k1sF0PK5dQPweMFP2agceyYets79qe8RqCpwILXpzaepeuJwZzRolpdm3YQGZWWzh3O7la
/g6qZ55WTaTC/xmTZP8IuGOt8zD9AitCjbJaVnvpIgsx1DKI94MydKczmHj+47mH6AghFuvQ5bno
3ZWsoS66U+IlOxnI8tdUIAE8UkwCrfPHQv8+yewx/pUr/uKzHaX9iXga7lTHaMJ9wLlxXhoGx4Mp
wM4WKpkoYTNGb5vwxLfdcxxXjrvnFk9pNc42QXVz8Ri5E4ODLnVf049jcivRiplz6niX/fJvqBb/
QVwjVF8+P+WTqwuFi/xNMB6E81d7aGUnX5mhXarIThpFyDaIh1oO7I1Xtv9JFI9g3PonN2ebgQJ8
Wdh7mClLUSlUBa9f8Mb1BSUj6sDZCCMis0AJ2ka7YIw/NjiKnUeHVWeFpcaG4zfut6urpOKmiMPY
ioPuPaz8l8gKA1NdQz6lQfdd5kLd6nzieHdVf6ri2yYAXU/wm4giLgpsj0t9IxipJZJqQSAf6AcH
TH4VRFGWEo3EKl8jbvNqvb0f9i/LRV4AfI7Omndhi1MnAcmWxYqMM8/Wf4pJhZHBYQJJ4/B6xm/H
lOo4x/FcK2PtHj02aTZk/HXwv5vsahTqllgFjKShDhvaNDu8rw+h9sbF5RtUhK4AJK9crqVHuZhX
5eytxRIYZyDcIxASncZ7Lp2pWL5oEkvzggTLdI2GM8+nNm93/D+nphvCT6ucc8NiH2+TBUwC8Beh
dsAD+GQFIBi8hiaaJrYXuDMBWtiQVA0Sg3DiAw+OO6cwobQnJhEtIwCBFEJKn8mTUzVpgbTS3GSn
qk5/l4Tuo6/6IvMxZItc8XDTo3rD2u5rq/0RCehwWY7in6Yys8nUfYcpMVVsuG06BU4GHdJDABTU
WG+7oRg2LHnK8EF3JtIHQ1FMl3CU+0uu6JDD2VGknhuzNQ+kfpL4h3MKk8ux+3sjHVAsoWcevx2E
uZqV2D7pr8iqkWF/lv4zVMLIRcdpNf9ZAMiGfl8K8dznzcm1/ENaT7DjoBsxisi6Wqc4bQ1FnSNv
mqa87Eh1tl90lU9/7VH8jKzm3N+nZKB16aHiOb9lL+Jg2ETHfiWb6JHVLCwe3DLa3yrHKu/Wws8r
THRonA0Qm7Q5+botLI2asjdG34F3wv3lbcTF85QP/jDgr3x0RcLGN9dKaLvjWJtPM3ZDHuk0v/MT
B/s2P+NcbYCmOS5Yv3ctn5EbLnsuK1y4pOtkDMl0/G7NTkMVLbskENd6eosCv+1X8v1xCmlP0Xqa
MJ2BN1ISzzptHlR9rdf3LTB1+to0HTP+Qo5HI5Ypfj263iwdBDJs/vP0j4ia7PxaBh1KtnyyAUIp
3vXYLSRKQwavNQlF3BbaqWU5i6+UvX3t6v2jqP+tAHRAJwj3roJDz4K7EhwEF5ZjnnMWJ0DaJElK
uggF4cvJHXOhSt28WcQWjF/a1Xamw/wuqMQW8VGYtEjrna6CWzyjq7cgoa2HUqb26Bzf4hZHbBLL
kcbxkX/Q6gGflG1MLJXA6Etd7qYY1vm7AzGrV0gN3aJ58MBHfJ7M0Xscl0DB8iJfq9Jdg5aIXL5L
3vCpaLoODTA932S9SOv3JVnC1qlmlrjYgup0nKedW8mffxNymdHe+eP0wDOnwF4x4fl/MDSL3dc+
9ZCH7teOD31HZlBaEpRLK37ZtSdjizJktKkxn5xyiskohegNQCeoxGAp85BGKKqItvbEr3rf8Sq5
moxhXq+Lh6aQDTIzuH5/dSJAA2kYPdnva85ZF0ukMvQ9kVD9SkCrJljXN+cnIAT37SUv57tDQW9G
nwfLNhi1wtc8SRA2sswqYuJVRCBnQkxQ4TpaPkpnrFC5/3JmZD4aMKdBtUHkj0JcUMrcZitnYWLV
+o9O4S6F4mWUgwexsftrleL7VCdDV3Plw1mJTWobFHVqNxP8rD1tGcutnRyn7SU9MdfKPbSRWuMZ
ziD1PJb1vCBfDDEK4ztOBerSM59pdEOAqF+JcQZH1Ras21x38OUK7gyWFpUTXhMJ7639rTbf5WQq
wlzanlXkuxwIH2gAVMhcoTCyOEhiVJ7q1NmKEc9J146fHgNLm7bIWgO69UCegBwsr2TkpmXODZqE
vI0a/n9Skv+N0o1xxY/yN62FxUr1Enpb9UBgO2df833aw/4wl/pBCYxkOQOly9emofSjM2E+8/TS
SeyTwVW1s7MN2hwVOKxOZgQcau3dpyX6nojo0jm0CWwwKLbm9gic6qcBFMMQR/ZQy2WxcgQzMeTl
BBHkSl2HvBBxtPuOA2tMyOwAtPyQz6xYXO3oTiSWuy0c1q1CMu1RNfRRqj/vDi7YFCTHMeVc/54K
035hnI4WhOSEqAyttm0fTzsixEyqiDydft4HROkemcu30LTh9UBg94QOReLJYVc5tsubnzqzqLzY
9GI6+5wR77B0Yo+EuRHmZ1LrOGPCtj977brGn4IqTH7eAcXCpi60A3o3NbWoVRH1NBS5t2pChbWZ
p8a1dVi0dxECnyIVvXiNtAU6/fhqIjdaNM6eTSuwoiBECIiHcJp0eubkUcJZqKlPZOiGaHQgzeaD
sJHwlgEdmefqkBzsbNxINM5TaSigA3NQ36eqb/ohCBzLTws5Dm1M5AEeIjTLbcFUmpS2zmPLU/hb
qXTng3h1uoJ/3AYWyR8ci/e0H1gklsk0K17bkQEKkS6txP7D9jPkU8q172jOD/C5zZAQ2n3/SKIU
Zhb7lvF7/CsP6g6TIT2Vlm+9KPeWKMr6gEL4pKx6D8y3xia8cfACUkf2FwT4DuIvfpO4L6uW+GRq
Yk36JbsH1ls49b8fbPK4IhGPZPK+9XemLDR0a3Eo+15TpZzAV3+dXR+pMIZ/ZxEEUlrClk4sYj2N
ikCsPAJ0Pn1+pYXn2eN8MAYfbENGBE6E6opf0HXkF/vM3j8ilCRhiTw0l1EkVtjsAgOwAdJwLMK4
5I+aRF7uD3ev04KDngsrc9DYumiVrDCZ4M7Rk3HER5AKO4HFY3rGXs4t3NSgG4FgdkX8va7ccIHq
tzJCe/UJjJLHhkuEWokR6ywE0A/d6X6kHiHWKjLDG7f0XBPSFV0Kn5vRS31WrYPLHpLaFp/0dZLD
vA8OCLXvYHNE6s+RqzTtbLa2APIsSQTYNF73a8Ggrx6AKTaQjliEw4Zj4YGMgbgmo6L6VhU3uNC4
xpwelJklWHoik0tNy7vxcZe8W8bjeoBUc9GevcKWC3KZL/xkxGOk2+g5VuLWEswEvKo7mBJNq74v
fn6bN+qVijdO6Sk03nVIR7M2eo1auKzD6twyYuB7fk6hby1tOgh/Kb2VIajrbzxGptQdzNd6SU2e
6J4CTM6e2b6gp5K4Nz/1wz97i02GWUv3H8YIkSjIP+aOymTIw0O8P4yY1BYmgUXXfM8ZAO02nUlZ
8lgL+G0g56/c/qm++eBTmC54s5tM9UFlDweVFQloakQAJVXRtI6JNky8rpLvC0IXFAduyFOcJsqu
ZW/Te1sXQJdJ2HCj2FotH0a78mSikLyS/wOsX79+L/RMwC0FDteZr8f5MnSJAbEL1AHdCo0Qg8og
5s2b5522Yy6pVmf3ilxrk2KrKy9eYJI6lu5HQ0g71r62mpPZCdb41rCEaS94VG2QiF+VmU0+9B2g
bvB+Zye8nTAnRhc66Q2Il10ZRYvso/y2Kj8zN9nS3yIlG7NhvAJ7zB1G/DhxN5m/k8qDKLrVQFwE
g8KMcrqptsa1pQ3OeUYMRriKcXfvfNa6SUmc50RgmzSwkMXeLDua+bRJbnNyAJrdSf1de4AravWy
q6IUC6bNDKkrY58OvD39upybqwnlfK8dr+pzYfXHRR53FwMe7n1Gcslx2zKq70G3LtIcM7OebJ60
g8sL9+DFJT8CjpDareUPuoqoAzq8Ii2WDPBKPEfSsqlQnBv+iO6DJxFNuuXSuZz1lM1e4lq3KWfQ
+PSYJgXO2gYnNvPmcaiXuB2FadFPySKEdsXH/0pKEjbR4XVXh8IvutRHi1Dvx1Ki35uduFYct9ID
qLn0ufr/KQyd5ehfhzQbUtpgD6vGvC+R9W54xliMARKWkU4l2+0nMq0NHlos5HoOaJpxNpSt8t0Z
8uUoo/zg5RDD5n0SxqZlZJ15rYmFVUI4OjxTbiHx1yTwBvSeGTZKkH2cniRcJ4207MstvpxtU3+6
Osx3YE6Akz3pnSXHMoHCWleSCqYOnD1ZGKKxZD3YXkcZRoKGXrDrvrqSHl3guO2rlh8VAXEbskx9
rzNXOnin/6zDkszkWk3Hc5V4L5W9jlL/CXbMfLzWKEiQsjdRdcPLyQq4VxdojjZZ5qA55YIDX5T6
bRztaEA7L4jxpu0aBtxPtdaCtgV/RI30Mu59GKEQuGD015ZBoLluSBYGpnBd5u4r+bmptZMnLqyj
2CRkA2gCG4dYT7IvZSpTbmKVTnvFDFhYUPjiEQvZIPc6HXKTTbWQL8BY5D9bskUK+W3NBmwd6cQg
0BoJ4w8a4Ogd+YO5kuV96D2kOtPmZhar7oc/D7a72srDrPDKYffuRfe4PM292v6yYL6iNYiumexG
/SFuqlkOw6tdC/+G6v72gWMAOIJmoBV2oI9waiON5dtENWltDfyJXB4E44MB3rhii0XAlZbCQcOC
EFYRLLfjbtR761q8ACLrwZBUdKYgaSsL9QfxXNmAJBCE3wCiiZ/3Hqt2cyCHgXC6WfGVBFGnRu3T
YkSgbInInzygS7RxSPqMffCdy4r3wYpBLHLdGbnvLfXLtEt6xAtoPIRBM/VxY2Va5SgihbViYC+8
HhbG0D2cV+wgL+svccjCFfozMN8mRog5L0qDatzqIy8SDFpbQXLtQy/1LjkNbivlozKy7HAJljJY
X9cfaJNLR1R1RMklqKSB1x3FJO7Idb5KoC4Aj64w5SgqpoqpvIdk99PczhJahu1jTtKWRP9/o5P8
EEGwRHx6HPJDYY3vBWNy2llUokXHpEv6E5qnQoAAx4wbMrqNKRkkKvGxXDPZ6FggjKZjVo/av3L6
UyBdyMId1ByJ2I1hvn5JHZEVXqWEQ6xX4udLMSXJt0DVbWPo+88a18UsiDyw+Bj6dKVq5+//Vr+P
OCCkaZANFzOAKPPxaa3RopFnv5XGD1ZbqghLO5mfjAenw7xv5+iui+qmzPayEHGWDcpjuhbT5lVG
P1twYNE9mmWsfNmTmPGY7inyUEeklFKWirMMurpOBZHcmtf4s8f9/H1hJpG9RZFpT8FO+7m15kKI
a7LcSjQTD/vTQpo9Ygfrafb2lA+XIOyx9+sfrVNLNO1TCFmz+xRyycbIMVLLgaeP1fFymoZrotOl
0a7DL+a/eHJ0teWLRTVfKv/qXWReGA/+C086XUfQWk3sGJIYfKSat3Zkmxd0P4hzKHaJWglOen1b
4k3OCrhjuTlJU7Wpx1EFb16dXRnaf1Z+leVI7H3wc3BUZur5Fx5c2YQZJw7kIbJ6OSadCsU8fMDw
4B54ZTi1OF/EaURbKuYZTFf5tPHLuyoSsVuFRetrhXqAqK0jH32EJX0pDOzMptVgXIEXQDRMkle9
evSDKtaK3ImOyX0rWfXXeHBwQzKoZ7lMTyUYkscjGRG/4DiyAy+2gb3faNOdBonc7l4OCHY3uvi0
sZz1GbZ/5yVUlxa6kUyWqWNWW53+CgYQTVyGHmKeGNgHq6Y5Yf5voyD28RioXl7og/2DyZgXumHx
3+Zg1xWXwUl1XqAvNcRxp0aV8pUZDYtSdOuROAUQFA5Jz2+xnsP5XGchADY8n0vDNPMc/bCt/iNw
L0ojpqFqY/5yLMLE79LCOPjJf0PJOB8QGOruZsuBeETJ2EuzKbN4OaquGMCk82ICZpIi90T/i9Oy
VvFLOJsHJjOQ4Lp2EvE+cZ23ynu/UH/8Shrl9xVA8IwslqGStlKbAsis3+wNWU1k4GWnLpbbUwh0
gGhaH29FeD66OahE9jo+qQ9iZy62/GZrcuHE7Dx0bFhEqq9ACsbjPgu2YLR34Ru5QHNaoY2B6e58
Slb//8gJukMMcxbLPE8Z/bnc4v1aDc06UmQtCLp48ITMIa+VveL8Nsw8elzLtrLnmy0vzgm8zWGg
lKktf3YBLgMQKzjvHPcQqzjtH1HXiLzQQjqQOYHDHklrMEXQz57wMVaMt2DTMzOdmH/JR09igjzK
tz122FuOY1xiyTzCJXieU7eo+GEslhn7elhNAsIELe/setmb5KJigg7Hr0joF1/eQUJrkAvNQFF5
ry6/VGCxI0F26q5zJKJl3LWcEz8uEiKyszTIdSjiUO6WvhhfCpyt3y9gzfGXe8Wp/KJXOBMMi7tq
oYFyTNir4Ma5LOOnqxdLQt6gruI4dJ91OLFmJ1c+Mb+RWz+SjJALEqq7gIg0/7p7lcIpSSF4wyN+
WT5ALzOz7VyPrIgpSNOWj6U5j03bXOvROHeOQ8CPi3tz4tnL7jidGdpX4eHq4ldVzz4d1n2HDU1O
hSrxnvSSEm9eB8R3sUhRihtaCRHR8evo1wSmewihWLXZ7kAutsZP0/r61QyjYPkoV6TdICS/e4Pa
NX+RjuyWAu5vaisSUe8Fp7CgxtJon95fhZsmi8YcxVxtWi/p+JWNGPYTPTT7PsaeUWwRzNDr8IfV
v+c8PTzaCSD4dUYHNKI+HRQokm2pyyeyEAzJr/4x/5lSwNs24QKga4TfsPpm9JcZ9dF03kVal3qT
nl9jslZNQ/PSPclS5AdnIQVoGenZ1rjMUMId9JRthCm91/5OEqU3/mAjkdMKNdrlZT+ngTABHwee
gRYzitoegdsNO+2/K09dk+RZoZltlQP5TjINBl6BYEPJ/oAwqrgG35wKIy2V80QSWEgZQMnId1i+
psCyRaLu+lNIAifnz7Sbm55Cy1TcxzgHKBmpktGgcRLPXMs9aHVEVNm4zjpocj/kJZNBmjXF7bsF
Vh3ojDyBWg3ZnZuJCPycgdgS6XBa78iuaJJyqS9E+y1aEkuVBH34u4/25qta5txwG9n6CSGYJCw1
c9wdApHpuhcs8UNNPlTHrERE6OWXNa/384Ji7Z8holEUKjp0aiXpeCeWNn7sBXvwXNpysrK9Z9wm
nNTCKYCn/YdU244ogGb9ph46OX1duwH2SYbPIywtAW61sik88kQNztf/EhP3TVMIPCoLe0QmBjAE
nj2m7SBili0AS6HQhlsLwZmNo1nMmIIfmFrNYebQsd60o2C6DAgOuaa2JybK1PhMFjonTwPAmRus
4pmHWgxEBJw6YtNG6T4PUshEad6036Ow6cEkgyKnDKmW8TikSpPKqLzTV+CD4OuUzyASlLoHGbQn
h7xeykBDsBev/R9Id27nhNrWMSRYK+Xd37vYukqdyTe1VihMAaORGdcAj/Z6UQmbFawo/xgeurQo
gcb/CwOaPSiphOSPd9FdfUzpPZFd52iok7mvwvwSbDHV5KQ1/1rs4JxTaS0lVobor+QnsY3EoiAk
Qc7PnfeJ3OEq+mJHGmmVC/BIdsn1MTgFVJu6c6vzSrCPdV9+/i9F4rlZTJX3PfiEw79BilW04R2W
Lw2ei9z2QKuEgt4oQPijYS1yX+ZCduZ11w5iYK6oFvcLQzzPOTtYMWNptxwZKvIP9SmEABbgnWoo
lSSasjWJ4SkZW1nBz2K0O1rwBvrM/ci/YO68Pe2aVHqDmarmFEWSBG5TmLpz9h32D4wtItJ5HXjr
HD/uyPIG6egq4mMZGc/emZ5A2On9cxjbiusEwNp3160uOXz9vuDUSzeb26J23ObPwMaJR5b+5q+v
aEghcUBnER4pKDhI9NGUxgUpmA8Akq/rDfVe0wkWcJzo9q04J2LgtYBSlwCCf7boImFpmuVAANS7
uKmaS3Bb+Et9uVBzvDATmCwOHiQLfUaEI+gqPzJubnGP09KMLVS0RFuUJ5uvn2EOSLywxEy/obrU
92sS+2WOef5YyiV6q8gIYraCElEG8VpwV4bZw4zAF8eZAGStPAgWQFzUeCT9ogKgOyYlot/ba8oe
XCTb7RBX3105wBoKFYC8+DUurgOvK4742scZN0jS6GXtAi03jbw97KKQAHzKASMBNdKqWFW6KkQt
8V5ao7momL1xn5SUu0TuUNevIF362Ezi6/vaxKNeZrKUtd+AM5v6n1/s31eefHr7hZx14OU5VYqW
t01wdIEfJ7P4YesE9jWnVwR7NKF47OKDQjkxsRLtkq01KBp9BADbMnxLqo6Hju2zEO/U9XQ+wpvF
i+qOuvvZJ362Z/vmzpJQndWBcC8yjXFUBxnGO9nILkZzexmEz2iS9uLBqBzP7ESP7wmbzLoCA7/u
WA4EiA72AXmGXwqjXo2MdtYIa26R5IanGfp2tnS++h5PbyyMX+7ZwhT6M8aVtAqgnXSKFXm/L5/Z
tSXW1uP8P4r2JIBrMlH9e5QW6KYEcEKSedOByR4kse4alWyYX667lHOCcdZVIGHwxBeqaq30rEVx
kjrK80E2huFttatzmqZfDO+JqWnCmxeR6hFgT009chCAMXNYJlIURdkNdFOQIFAmmpvtbQRqBwjW
3WlyruTVN45pQxIVTUlgONODqGHxJuq3mD+rH/6F//Jfaj41mwCVqDuKktWiI7nrXC0glcFCC+vq
RKsFNd2v2SNtto4WJwIyE2b86povdifkJpfcwqLwT2sz7zO1EvqHrs06VPyk4v4O0Uk5xl17E0IS
N03qLnUWbiZAhbyoGzmJ+JiQvUNhxOEsnN/1vGcWe4kF+CJmWpaRlbRj5VvzEH95VEP6R/G+d+ux
oDBqQP0am7FDtftWQ2LdkQryy33VZawHWp4+9ZEFfdYqMvXYFJOnOB8ArV2q9eJ1Y8AxZ971yt6K
gtYsOLyEMtdDjkIOFV/snFc8Errtz/WYHp6gFk5U1WhjEHfiVv9YbQfG0VQ5t38CeqBJbLRP4ggH
REt8SVVGIaecw5mAyQakn+MHFAj4I1b8aS1iTn4EiDSrMH3+yQou1UCFXJf1JeBlLDu1Z4KvplTS
xdOWjOkwK//VDB4VASjzzcubidpyM7WvBzSmXz5N4m3GK5sPWVmfW1vNVCleLjiLkw6Mdlkjch87
5Acy3SOHzvGOcIvvht3SWOEJqj4aFEkpa0dQUlvc95NdbsvZuq+RbNf7g76ik83SdP14G3vDQPXK
l5HvhTFHIGpGWhcQhqGx5GnroXubzcJs8CyCaTIZnbhxkP9EtVG59fhM9pvF1x9OqSoV1Q6rCE/a
YYPYdpl590YenwaQ0ml7ydUHWohyALrcdyJS4if8P80NhOmCkBKL7W4YXsrHVC6jxYhg3Xg9GPIE
aLBomXokB+QguvUtAA2bgOFnJk0tyNTaCjnd6cD99xGOZiR1P4FGAR3w4U1BcN9C2wQFJVnzbfZe
Ezhae3EbNJbbXTsiNbrAI5VrxeBJ+JIEPlnZmK/pR7VLupzoKqLYb2Jswp+QwL7MEmoUpRp3uvDj
Zy9UuIkc0pinfAcNGa4LHbvfLwh8JM6+k8BgmJ0/xVyg5Z7HX3vPFH68sp1/5bTvuGV2ALUcK3sK
WeadmdCLw41CmKiFJp5Q/rrbumPHbk2OxJBSkFS35gxriq1X4h3R4Op7O9JoUt8yVZeiNivL/YhM
VUjiJ31UvvmICuOWTrAHj5K2LAF2+R4zka694C3Qx83olKVwnlG7Kv/jH1QH4lAvw1gHnxRctDJp
EdwZuhc+zufrLlZSQnIrwwMveWEzP8Xe2nQlYRq1pBeWmSmWzPw1vMpJ7FmMgMzLUWn7axWitAY5
nQa3rJ3F/3xB4eTaKitXNA8/H9MV1ym0frq+FQWkvOdpiv+G6+wozZmqs5lt2j6Kav/RIlZTFJcL
cXnEp2eXpiRQJNbIKVj14GLnL0rd6U/RYUZY8MhF9XL9sFQ4ZG3w9wVukoPZ4vwdTkuy8ISm0CoJ
r2d7exXWv9P646pc6EPfIuFsXHic0z+ls2NIUSlihoxGe9xpl3IPNLpqqlhqxP9O+OP9tOcMWSS2
MdK9wM8QFA+xhTtzNSBZrSAEYPO+WQ0wR7tMJJyGTPGymRvn+hRySj2RTBlKYz3muj/AhN86DnlF
0TJixONJZIFb7Jdsyu3Ez/e3eET42lU2o5vVqVfAB3oHPcaCwx+2m5qIcq41X5egVkwq6Y4dyubR
lyAw4ISwkg8VXP5XNOowjmA0PpbyfOftxHhIeJT8ZPROXrholrBuxMOdQSz4x+s8y5SYGMywqewJ
G1TH6VhjyWhgoa4pCZQnoLwurVMbEC55tu7fsk3Tdo/icBrZjBo9qdQ5iGWPTxzJdOY/GrCC4PPg
f1o26EHA43yb/3NEJSv8lP4AGurMNGfbZWFwruN1lej7i9gEmU+aNGSPpE+GMJO+7sGIAur7fsV5
ktbZ6mVzz2wO6ItpiJBXzK+PY7SJWbO3qOZCaEYpOrQZxZBRbibsjkEmvmEFkXURl2/oJtvEuYQN
fJ08guSuJzQS7ze/9k54b9u918J96NdtkBt7KN03pWGgxUpRBx6MQDqkrud3//NO5MdRDo1ARE89
Yd1sTLG27Tagefk4RDmdag12glQgWTRXtBKjRQszG631PvfTr9xcONR2pENCMWM3OmE2I4AO+tgJ
2fiNtqI5ulensLZDnV5tEKoVvh05pY4OoJKnvS4laC55h1KywDhroNB/McU4Rhrn9bRXFCq/kG5p
21ouMApdTdYT171ixZvai7+fQIBjwrXDpXvwFdl/hXt8mipw1Vohm5vvIOmKM0fXHlsk2cdturAA
8TtZEoJB8WNLidIUNwLnkfP+Cr0M89yLZySVj54kfXX/cuCxZAIAkWrSh2O7hmse8I5Mbj6hxsge
eKiY9XQZqlILEMZ36GzgKtFF84+2Sh3IByfUB5S72ezsxXbuQ/cbhdtoB0PrHNJLpjGvqW9aO+Fb
EkgWuZu1RQmojzN2c6uxUiqX1vbGYRRVxxB6/y8JE2KsR/cwGmkWaJrtBJNU8J6JOGjujaCh3Rtu
MbwHn7ZdpbA51rT7DyV6r7ORGhmxRTWGs7Hpn+ig8bSkRqCEaVq110OybCOsNOjmDx2VloxyzIw4
tVt5Z6UnD/pLQ3WR0AaD8YvkSYTJriKTO/7zra0kFY2BrdtyvUocumrWaLTXDZipFGv1fOEChtAT
SGSg3g2UlSvc0+eBpRxyx0QfCBUTQiPWa7nGz1bs6TXdzwpGzD0ypqNgYlOcE0gevHU//ZoSp/9D
nLT/iLtav0pIYWv5KvWN2zZ4lNmrIe32Ql8KVmFGKBTifESYGLA/hDnkOXejHACPh+vKGh59sn3i
rAAvq6DoPxutjdsl3Bd/HjX/5qyavJ21HC3Q9mS4CNSgBJUsp/wVmkRTD13Qj0vz37C52FEtPaE1
iBnrNLERY8jSSnYD1Pva7pA8mloxh477ycvnIlBzQTgudl8sHPif4a2w2wgpk2+6Kcp0u+aOYxwr
vQfPddzZd+IHmGbqI4VGpRaOXIBpDNv2D7NxsTI3bS5f0Lq2nFYpC2ccWlLbgMxGX+1J74kOrfBY
0o3AnFMdVQFmB3m9ID5sU7Dufbxpd2Z9NtcC121JJlLjOQVc9olk6Esww8HXF35KlfR0Z/8j3phX
RzMubPac4gXrIgd7n1hFV+VxKOsShY3oA1p80rqMc2PXbJKwe7ilBq0bNh4rYTOZpjdokF+MwAVh
1PZBNzXVmoDukK2pS2ZJidBzNZEvo9/7sFZS6nRPYdjAcqW2cu067h+IkssrJLL7yTu7egd9hAYB
3UuMi9gnqVrUo0sYjnlk62PmHjYQiZC/5fnGezeDIHSBkI4hWu4LCehcajNCWOd8cgm+lNAWpKnn
QvoWnl3pIAqG8ayEfo3zpgLZR7ZoaKzjqLt9+2cpUoC6+7ReMBLOlVqBzDazWp+cU5+lAhPCUtF6
kVUlnWKnPAoRQpH5017PuJJh6OuW5auTS3X8Blp039fpR6zXti0Co3OxGdci5fJx/o0InSTu7n1Y
hefxw31XW1CPg1Jn1DLf0zrGqzHbSwvKTkmfc/K3MZIUgpLMP2fmCFlqINDtbUSAYr64vwt0H4eO
D/k4QvLxrwfnyaVfL15TuXvJ3GTx8Hii8hFsroOMi9Su+LBkURrl3cxpCHKn9UWaSaJXwkfvEGXb
nC7eIva4QmxrVmXKuwUbuqPuNP0G+v7EoqIbf044KJXW//JrA3PLKlNjVXG/GgrbqPZS/KSkdf0Y
Kb5Epg+Ze8ofWoqI3F7o1/BmlnCp5NqzjrH08LrPDwmuOmg0btp4sdRE4PqpKjY0BZB9+PtvgxyF
DlwXF5svQeV06EE7GFJUHszpezAyCWziz5RlaDsfEeZS0CY5xhiq0LUu6StllVtQCn6a4AIq/gjk
pa7WN80f01fEmHoMalaVRHG6d50O+E/cdekMsDTQ5CaRar4EM+Ntkqx6d0r/AFYpf1vEYGrahuWq
TnvRw42LMnDNjMMLOpbI3U3DCgjG2FJ3cKZt59187ll9QwPLY3PviOI2AlPY9Y0SzKSYs8Aro31H
i7YyLlGRmYWMJE632YtElwaWx+fHguuGez94qhLqryRVYhlu5Ad6MLwZPkqXB6uKYXbChYitQcXw
Xd3VRglEgvVmFBGvNtICF7tzECSPdZNyP6bbyQE6WAE3lBdy4D/1Sly9FJaJwr0E4NseTPB0rbLk
3wJXH/6Exr4w9rtiuJUmasXlkcOfXT/dmE3M1LeqmQGnWOzGLBRf2efS0PazNHgLxCBI5iZVy9rV
HIXecRrRpth1A1ROlYVf30mEgJV+NrJ0Th1iT1Rhn+Po+PC2O0SNF4VrVjdPXtyiX2P/sjGcY3mH
PRLAaTmkRPBD8rpzbZopHJc7AVgxPMx4rKLgHrkWYpM6SmUalJ6WPWkpoH/vHcSKfsatT+3V9lrF
YiaEcMTEUtPli+CZmd2PtNswOB58roXsmwqIhnreY1bHiQrSTPFdTgOSgURusx6YAKoj6uBMHvII
hGtfhRQ/r/OXA9lDM3oa2vyTUK5Zgzmp0mIsYEsqqOHuJUEM6hwhyT+2HV02Cl6vpEBZ7dYgsYfU
9GW8rHQnAaptqgeM95FRB2UQsQoRSj8qvzMkWWXkM5INt+YzA7HDEol4vzTsHXZuXRWEZqj9Y3M/
z/HMOlTETPEUY9/DDMBZN8q2GVRpiu+hTK24J/ZHpzBoe+jmzt0ik67lDVchexAVtRVdC7q66KH7
T5YYEqiN/4xaTBpOaMqBO5QkeCTJij/3nQcUf2xK8W2QDHj3W26klbjwJSHY12E/6KNews0p5FTx
bOi6Hkbx6AthVrYeTjOCL/y1qHFNdJ5MTzlNAbKrO5Hdy27LP5yxjyO8DmbTFNNbU3FgjZzV+afI
9YUiAnVq35AnvWmTQ7ayKBgp63aquL3bCXk3DQh+Jp1KzQcSjOIWJG1PxE2DlnCi+JW1C53PlYvr
8p9n5Kqku/KuF0/L4LHWQzfhZZBgd4g4galN6sl2lyj2GzASevNbCfmwmcEqOMZHbMsgKCo4m042
9Q6mz57qyVGdND9H4cPzySXfU/wN9LVMiDiWXlpsqNYp5/OSSP9Ne7tO850yThqETQaUalzqFJbu
AbeBgAUhOmg58Sm1j22tP5F4lJubCqE52SLZA8QBZIGS58p+Uleija8mzu06TqG8p8wM7cFYLkz5
uqNH2GwjtCM+TUCEpS10arwmADH1zTDN9PEiDoDL8qj3xIWEBCGsQ2ODnDJxPuEIAzE30gnsTDJ3
ALDMDw70xg0kfX3jDydi3LqY+ocZSU1HzNXH+1MUlvH7u2JGyuFfIk+wjdCWv3X7BcFhb1/9FAUi
rkQ9OiUCJplJhY/b4Ijw2eReAtKXxjf7ZWqRX5IoR//rdsWJ13lm1hcXF0OwIZdLydPowNDI0J/l
W4VtbxO3A1bsSGRhqU7+4jWBM8xRx0M1bs5De7M/0h3ihFC40QQhONbmj6g/fvQyC+KdrACTofsw
4BKrS+d3T4xZJyLQnDFcrrt0LR1qBgkX+mRkw1BGL0kyI8CcRkVNMhLDOX17tU35Dw7tDJ/b5IAK
40Xy63ef4UmFQF20S8H5JXGyFPxRrRqt8XkoleQX0FsuwwWjFwr2Y+ic6wNH+hfAtyRc7pYuJK4P
oRgCtTa/0CvXrwTwA12sw12a4zxNuNGk8xSehKC72QERTugQ/nNHzdcyMbyBB/6nAdekBKI0vhra
4Lf48pcPTOp5leCZBmuQ3WuHl93GsaEcrPazSCN/pzscDB1DnGo5quqUx6VCD6zKILh9NVHkz7vT
/QDKwTu8BxiPNAQ+5l1ZZQ9H95+BqdjQJHnyUsiIpSrHGbBrYQ+qLprnDnmXbea7MYsecJdw3ESZ
vejNmIZU/Gs0GYzO3q5A6yfj2CPzAw9t6dMdTzj0AjePe/uAq+uhfnUpVQ0TLsaXP+PTfvkfxgt1
xE44doW+NHaa/gkT+caXEKqe+5fbqOQ0Yj7ZFXCbJTKpQGpqcPibeoeU5IFu2aOwawupyqyTNNKR
lgeQFZpARh9ADtms3hSN01wCtTYovpeZMOoSgM0PpaTciTh0zxw9gF901ZT3Vb1ZfbQyHvFXnVlE
wZiBmGmybbiuW0mg6OFbcAcAxOKy52BxAxTJ+td2UxZwc7FxhsnhLNVGkDWULg4mwa0ZQMUQoCLI
KKcx2eJLkbLTSeUhUjI4v8pvkq5+ZSUKksKZPUuEKd7Ni3doxHiQi4bS4wAETSOfrr6+hUiVbG7X
8Qk96JH5hIGBV38N8AmiK4nEgv20aFYQtYLn9yZlbHCE+ULehDMk1n9H2XUmUvUJ/8uJ0hWlU6ba
eUwcy/tOPO41hCJUr3/VS2kgdf8NoZ9ILu1k+qI6RcX4WZhVRunMJplwYF/uCa/jUmNhYvLFCHcJ
MwErUY4bOaqjjlubHUP0oZ9e8Q9mfvyUd1GP0b0bEq0tBR7f1oG63Ae7RDc/EkPLJuDOt7JHqrp6
WGz4z5TAGZLqttyMjW3SBA6bUnWT5vsnLsTRgd1bu6G0FthuKLYnGF+lIyiMbOhwhmv8YA6Kn+tB
Uns992Vep5wGMI2luzJ1P8sybE6gysi2DkRguUXmtpfTV4+36OszJQYcgzI24pBeWWOTdCa1KWo3
92Ex2PYlrgjKS2JAZxF59jYjec+PFAE6t4RJHETVUdb25VbqV4QEXFdM1V7iqfOcPUgpFN7i4vtB
t5WQKdGHVbopTIKvhSGdP7+5plb5dO/E4xfGLlyu05mWhexqFH4qMMC210MbjzIfAm0A+6MQ1qPA
pGVwkLwjiKlMx1Y91yXzFnULptJdH0RycUKskhBq2lJ2ue9GAp+jrQd0a5VHvgmuNo2RT7spVyBg
72ogRgJFlaN2Suodu4Lp402j7Dil7b0sgOedOmO2l8GXAZtC4zjSkEJJBQJFHHiSMHEbhsaDSlv3
tnkNy44MWkciINYK2NMICnNWUc6bN+SVRWZiY1MTf+g2uJMmwYr8EzoP4pE9lGU9YPiR1n9iPYbD
mU8UvGDmDcLU5dkQli0v1ch9OjZ7Hq0wo7+jX88bxPXWFimRRPZsBRmTuwNXzWnT6CGYkaTPfx4o
DR+XX3YocUpehkPbgQBkTFbeBUvzFKnMDzlwsgUH8aQ8ibnvl+HDhXP6D5ogAzAsDw+zrzIijTxc
UEOhOrXajGxyKM6MKn6p9xTmrp1I6MM5dnS38g1KgqFTS2xSomhg5UdIbpq+V1kbP7F0IhWNMjSw
vMSoJRxSfwOW/JLJf48r/ro43qqUFDLCEerCDWNcwkUayjdzeKCYYuh6tjBFkJbJfCQN8ewujQQF
b5U9COgwuMT7s+jg+WHMO3OhwzT/al97ugG/C5fLEKHog10qHAN3SzkuMrVWCEXRXkQTWGb+x5lc
tJNI0Cs46ZxTv9WZxPG7qgmDc80kAUtNsSu5ZBvwF+Q2bsJgD6avoy0VDCxiiKkiJymFbd0ja8QI
ozyeVXtxWT6UyLK5o8PC55d+KFQ9ocKQxTaI8im73OTxVyawSKaqkiBjaCMLm4Y6N1yd/ArwBAmA
Uj08cjsry7UModW459yNtPwKrdF7A07xP//A2kMs3rZqRS/O68oauTU7iAd/0E+Y1bL1QhT4NZsm
E02gn/pBdXYjC8LVIBSeDXhZ/OPNMxqBXmgzXQBBGw81nOwCJ7Si+mg6aGWZzMHgqOB472nfrpf5
wavunLBUOVpoaz3vfUs95KpDdiTLOY5QNTwsJmV9wzRHrGHhiwwc9Qdyoxa0eLGpymrh2rTlgjZH
2mVAjdfa3Y5Hb2B8VIT8XX6T82gPdRd1yYmYDT75uF20lnFkheOQPNitVcEZHvtA6c7kEbVxIa9G
4ZK8JlOje5NZ8WWXPPGYHDLg5mhqaRn7v96IN4fcftRlhwtOF4TnLVAinrFh4XwdDFUY/4k8CDqw
4lWiz/dJoafP9s/JhnGkyyITRkYLiiLxvloQjmGGa//dXI3++BiPMIDTJb3HiMIaAkJx95VAmtiJ
b1tokcwOk13FLnLODwtfGgVX90xHRhye9R73yq0A/qt7GsisM5w6nunwmvdpq0kzEBzTKx2o/xUp
MvpCaxfWFEOSpy63JbrlrKViiCp2VnDRaxMgMnH324N24L+0/uiD72eNIFqAppSIJoDY+GCg46XQ
y/dXNw7ifq3NnqUIRLigUqmIGAnjdCBGe1MeomJWVU1nXv45xleOl62wwu4v5HkWrCMZD5EBT+TU
eknY19eTAZigY0zOF+07YXOc4ptbn9THVa6kBE81EHLJ0Gsvh6Pmre3AJnOMxG+q1f5hNFgTesxo
9PQEX4mA2qqawSPH2L5yaCWdRLCK+ai66AL5Tp5m6+DtX96rmjuwcDQKJGdiwWCSCrqujTD0kaTv
QR96nnCuhbwNyrbIt6ngjvz77zvcL5nru4YynYmgj3Bf/AKmd1SAyX8oIqrTDgjTgghAqi0iEbYB
nwrhoRZBgBa1SlmqgdpfO5w6slE37dz+UCEfD42iYNTNk45pVWUBYIq3GK0F1wj4sTlbcZbODotE
oHanb91lvYk09Dnn2uig2WrSrrYCU86KD2TfCr3AThKdqK81/Qy32vYftvR9p9z3DI5AlT1qY3s0
L0HL8Y0+igMZe6nJUAN4gXRksjV/GTZzufpMkJqSzvozZSIdAgcNz/0XcOcIUeftx9huXBeYPCvz
GPikOPu3j/R+ov7dKtJLEfNYDDl3NlcBQEqxg5fp7DQhHtIGMbwd6JosykSCDHj6HyHk1Gapgn1i
hGYUPUn6PRCNmOXmzN1wAMNsNDRBvA85gQjBIoXnSSJSB0DKtKMPQiBQQ9GFXFjeBwH8PKbV1xM9
MRUejggRNf9FcYcOaVPwZbDIr6hz9izMObbgA+p4yKtTnuDMJGX2WtrwLHVftUKP5kaagwJBpQpZ
nTLAnbfAQaE4sS4OI6wsLjWS65hFLc/hmFqsIsFFhqYUkdx8MkLZa0qGNguWBSzORr1+v2HXiLUV
SMQVUUxDDOTQzYhB5mCuBTbESUfeSOAcMvpdgKRO2SWkbdWsXuY8xnBzrcMn2EP34jd93UKYyT2E
DoGYXKnSAGeiqgOaruhnAwrvBoQUmgipgCrgqXBdxua+17oZGbb98EmOycf1MztDKmSInffIau/a
2Etpn0Kg/L1mE2i4NGfWZBcM4zS81Ov6g/vTecbP3aijtKYAu+ogNb/ysz0sMGtcm12P7vZRfdf5
337YycCx2fKwsxvUCsU/1aTJ8AjJtAHFkU1wFKiRNKjIhncdU5w2BkCpmdSKSv233NFP8SNjGQJg
IOMafrzOC1WOaHqIqoh3zDHETnmICwlMziwjaDK8Lm2RXjQYAgvymlFxBtyFgskuUQl4mx91zoFt
xbzNezL4v29ulBcxfjxXYeLmdj2oFKhjNW9uQgiFo9WoWSDq1+tVP8nkNjj5a8ZY/OxBUcexgGjT
ucsF3O9ORqyb66MeXFMfCpw6Q4HLXDTDLjqdvDiA7OlUywQkOkw16QMyZ7mdTg4lMJ6Lv0/Qjezu
NChIYV01MLOTsc53ekwb9SaxwuGHDqqeSkWaB+0aSAS71AViI02IQlG8GsPkEjmq6eIDMNiedhMA
11EtfMgBKqRVsOP81BGFLB11LYVe4ch3u/9XWd7H3Wf6XHtHe1Reg9d/klpa0pUIc/7Rq+WKfIK2
sb6+gyH/tmvH8Py1zP8oNWyurjK3N5BQKWf7VsP980WZjy/NGW8FfSsraX2epakXYn5Dfe0l1nEy
bRIK8N5snWXs+NxRo3XRjnJX5QXcnkhIw23rvxCCkMgP77Dyrf+Ot+YkJBapg5gSGLIY4JP4wLb5
QGTpFyNSziUPPLhtDHhMekIQ+4VR1RSsW1Bf8OqOzLv82GmpBNuUBj9+6g5okQTUBYVyOcm4ueFN
8jCpuwdL+AOJH321TqlO0ViPzgLkpWyBk7gjjMZBpk26RCvTcY5Ftn2O4K9CNv/n2pLdieIQJspu
etjMqBBUPlYd0kFJDLQJFexw4xZN/AsbdltprBvBDHfNh11jOh3exjhXRcd3RT30QjEtljm8Y3zq
3ZAyQ6aIUsHNtHPiqD5KNOYq/JY/TDQKny3PUAZtrYDu8QNHrS1xc4ilxfS2DQ3vEpHovH0ODM8J
9Utol8OPyJuGUS4NWSupsjizWXyJNI9a1PSEJ1ESXWhLd5yhtyjJ3bMnEMAS/uvg/LX7Z5NTw5uC
W0fs8QOeitD/OTo/WvnsNofDXSz5BRRvINCXd5oVIBVYwZLP3pDqbyIHbvYLn49g6PtuzwlXjn++
NRDcJhGlKJB/6Z8C7eZu9h8M6efh1dmgKQh4lRO3MkkNA8oN4yciMw6Te2lDtUcxg6c0V/vXWoko
UQMviJ8AORSym8BfOLy2p9Vw1PdJsGw3svj9v4u5ua7J1Oady1TxncxYYgRVZOFwi8JQzTMaW9nA
TsNQLnIvIXfSdN8kMWfWIKUdXG/k03rabe3jonkmkj8TP2jkQb7FXEHRnjtIB4vzw+T+RFgsHw+9
ZYyz2itNEH3tNJ0zcULRDzCtvAXCiCPUYsUWwp/r3wiStMtG3YY5uUtU55JMUtVQ9bEKwG06jZbZ
Z2/GVZT9HfsjZTp7nGuXyKhLOAEdEviNfl9EGwXZSt5IAqw6eZ2Y0yyY+GZ48Q8wmDqedZXg3p7Y
d9CPreQ9xL8uvrvGrlnauuEwjKCTOUXUhUUX2uNnzqCCLT83aBud2hz6fEDfx/demPeIVRb4nmUk
IXxdqaS7R+HN3vbZteqEWe2peyAhSpCiLwAugJEg3+MGwrFlzvNHAf6lqNCexJu1zqgQNDyH+Ksz
cbEDOBuyjjN77R/bbbUItlVk25iCzt+jCNkB9kVpSNb0Gq8XTnHjHWxpgMxM92FsoNMCI5eO1GBd
6reBsviTX/XpvGMO6fXzY29dBPTQOOFVopisTIykmmEVBmaixM7L9QaRHI332WHig/iKkRaBKv4e
wNQKjgKHobLl2iyfTi9YK/6jL0Y0N5Q/JuhXLUW7p9T/WqoG+Y1jdUHUbBcOVhSVeO5/2jOb3BSd
dIjzZicIBLdtvgh8HnoV2qz9kD7dDTxY3eVItYukYwVvE3KHCEWlSXsqfjDBAw3h3QsoU5XV4iqp
F5xPxW1u+ZQOvuU+Szq+MJtAoEpdiwmqv7h/UVGX1/vs77qKZEUdU8cOc6KJrme9i6zabFl8xIij
H7OFoMskLVLP+0dC9H5BjeAC8YgCu8/6yEeUcfF6NFkQRWBBK+1tX9Hgz2M8fsi6XURezHniKIJy
jfCbPaKCV61iH7mjbzDUR+uRQNedt0zmyRKN/X0pU03oUiZ7US/zC/VK9fswcxFnl9a19jjed0jG
N9x6JYbwAXZTm2zWgyIpOHWhzr5/Dd3+ufxJ7Ptgy61WDzIKz68sZyBdiiteub9W7dRHyy+tt3zk
rUj9fjFJgbMk2wEeAru3wZVt3a/lsojzUf7VPWMVQW79tdhdN1a/kLauHYtcOaup9LGApEj4ED4h
nIFpFJo02YZGk7HoLtxLBZqHhHV3NxBcP+DeU8zobOoYZoNea2FbZhKgcXtDzl1BL02tmKixSpCv
q7d2OAKBl6aRv77SD0LvBesJjaHXQQSbHdmKYG7W/lLa6mnyJRRJWQpAUjB3sSb39W5n3qupte4w
VETfXnNtZCM1xFRjyLtwhKisaocxSGPTbE1IJMto026qKlzrcbgbqpB5K4ZWF0s4XpZF65h0hpgb
O4oR/ISEuqaOcTkRC4VOt8PmqGHLZKRRZXv5587vnRBmSmFSB7WieKReXv4nRA3VRRij3NYm8uCR
f3cq7vDp8bnRufMDlr825hkIo5UkO3vfARLuz6WjdKLRXs4ZSDCYnWw9/TKztm/Vmh9zU+oJyHFh
hgYAvKZiwIw8zrSkiDSPoJZImiem7g5ERMZqFznv21CO7A1S+DIOz1cGKH+EaW4XKieTopnDkOC8
YspD1xxYdvyvG+J764vMUkfV9jWTfD123NIwp/KGe8lbKN+Mg+RqupJJUY8le+N+WmisHqJFZEXx
JyOozimATjJ4fCQ+kEBBXBoWqBIgTLeYKu2TLJAuKbuENHrzQSF8ZoIc4W3ReeO+G2Kb9vZDEo1o
5WeeIoD9aKbxpJg4P81Y4QBPQghqQnOmjbFXWiJAEShZRUdTf7/LQBioBK2GOqp+z+pLT2X9CmWp
p14bebhFrwICK+zE6IpECU3J2M0vNQvjYI+JRWGlfRrnS3/vXLcmPgmFue2XshYqh+tfIYTbr/f5
b9XTfzL2EjDXGsdPF/r3SoJA7VCRwIxFUVKfYpaJfCnttuUsl1QqUKqSaPsBMdv6R2BkhodSOveF
xNt0Cvf2vjRYpTyIa4zkY2OUUni0rulA6wKnZfegMcG+NZWTnQbdqKU/nC24XcRGoDImnv2qsFxL
usyStknuayXUJndTqx8u0ETwpeK/BqO608wqJQP0HN6nCc+24JNlKqhGNhKU8zlxE4zRwJ7HBTj2
XJto6PwMihdTIlBBcawx736GeedHaByWbJBCYdOr0SDE26DypdT9WF0R8Buj9pXumMiX8PFE7RDa
uwyf4v44UFyg0QZnZgYWYxIkez2Y+B1cHvedsSsAn/+xKz0lxnlvLcFd9GKevrurRamvy1radFaL
fJPeTG+ssR1EEQ+YI2umoKT+uZlocFLY9OA3S772pfDLmw5RH3vX3AjFMDx8O42SeDPVDTPlaI3V
uWq/Ha3O83aMimTOLj4OTOP50Z5oUcTYRugU/LAV+9pEYamlJlUfwERqw2EMJUZc2FOdZg/Z0RH3
BYLOW/+VYiHH3a8vfeD6A7xf9vBu5vXGWQvnwGZd8fG41dRsjN6bnUb40kK+lGOYAoUXhxzqugoa
a2yeTncEDXdUTtrUXOURS/a0Xq/D+JLPUXg5m82jOlFYX57CndZb9gl+Qa+11MuyFi+6DY8YKJFj
SDPWJw3QxXafK2Pnb6ns+p+kNP5gQRaIp0wz5I7R51xGHgbguuC8PoP9BJ6wN0Wak93hfHPGKr1s
OImzbV9k22mwuCwlD0XNrVCnPC8OmPagzrcO+rUC1zkqRNzmm3wryr5LDlXXT3U+uKmEmS5N456c
5ngcLN3OFoaU8J+d4xnkS4Hs2zgpeFR9IZFGKpYBHF4HmuKForakibGb+OlhO6GbyP/TOqpXgXMi
N23CTqoHlb2hh64dZ3TFUM4ZTN/rkwK0tDTNvIxZqRT/xfMsEZLBjVg96lvrTdRafXLFMkcNI1B7
Bjan1AIT2Rm8kcsE0Ir8ykTUkQ9/qnL2Etd6alMpskEUzrVtmYtSVqhPjMDFj7Fk66gl7Bh9NzEg
Xg1pTebEspo4uqjnjK5MMgdprq0TmouFbf+FGWHCT9tHcG+OczdTtHspb6rmTMlX2U7HYYddjVJv
2D19C95QDqlMrvlIEmI0VRKiv9ZWvSuzr7SwLe+l043LI+rhuKXMXJ1xXD8Gc7K/sG/UCF4logjI
WiIkxK/r2veU06U4zi0n2D7JlmwjR3uqVCSFrUgLoDjAOB8Q9/sRN+2Vffrj/CDHF2WVXa8hTYlQ
cugojebe45r89sW20qsQX0OWAkKV1gdxLBzPAIS1i+4GqetERJS35WXHlNveZNeKEEGzzfMpBhSa
Z5Vg60vWXFtZlhC7JldXgBT0nSRojnFKwtN/ywi/eARTTpTqSIELPsSlp20memqEDi3iqA6PdLXf
jRKy4A3qjkKQE3Zom8NLY54Efs+lwseIe4CUGST2RdTJvhWfjXlm8QqtYmS9TZ0vQSJHqxA1JcN+
wnh8b4ah8/jrKuiXM4PL2Jz+9jTbdYwsX23IJQepWgEZ+MLzhcCnMn9IGMOwg5wft+5xrAvSY7As
VsANxDl26uXZZtrFKPVxPOo2nbo1HYIkD9hMG01bMkumDXu75jBh8LWOXer5UMVv8U1svtZKJNwe
BK8H3x+eivt1JBqSdhzSp47+1JzdCBkUja3HViBbhU/LVTBTdjnt9/hCqir22kFUl7igNzSNQcTv
e9qkeP6CANYdp7SXHygnlOxpeIzY/x2UxPrTlmf4mc6Xr5G0F9bisuXPaWbdt8zJRmo8mMyl7Zka
5I5CLPIaTOZDFJI5p7oFjOsrRSKhfbHjgLupE73giOp/x2U2VG+de+fCPDy0uQkc4pBtzsojUMK1
w54vOw/ba8S2L8RifNWimQgqow7bniuQaqV6IdRlm+t2BCyCZvzlqjAFNI5qVx8mOA0ym/t1hzft
pAbM9mh5AeW9UpxQGXE2oXmIz1BQ0PBKav7HZAmk1qznxl9DTE/ys3/wsCQmo/bE1whpKzIW5Io1
tOIUBLe2T7wWmKoW3mm0HN3mqqsMTdpl4JswDR9qJ677psWTYmWP9zwGRlie1XUviTHxmvyAYivI
9IlxtTGJHr7U9f1F7ZcFr3ceeKdXCaieo45w33CqFCsVuUI+RVXxhlFnIefYkfLZT0kxR4C3WpJ/
XjwflpJ+TDySYA5xMKfFea98fDJDTmPpkwSlNY3o7hgGPXoXzEc5rIVWMAFIQkv9AingN+45wFnV
P5M94sklFYg9/CGdpFAT3/dNk0Z3DAeJqkWk9p/1RyUDUn26IIRDYAcfO79lBi19tZtoG0pjKNVn
8iiXRv2A6pYXh1k3Wf9MKX+mH6IuxXvg1CrBZfENX4EL66HbFDoK+e/+i02Ozw/qNXAIi3c5g8Nu
iy894pFyxepqt2G0mR2oAWa1jauSTGgq1w2Y9531o5C3VuMnljULfT2YfZLeqtbXHQrSOXAMaMNL
V4gEE/k1UL061eF942QYX2d+iKyaGNpinbpQjd/ls+HItoHNpwAO0q9McWVp7g56rqWsOopM3hSZ
2+xg8TWRv9RRnkdEDCMs1XdIg/pdJA3tgaahlBHNO5o7knbmW+4khMx8oACQMoNQ0gcB8INj4z6A
XQpoJZjA9udoTlxSNHEmcKOS2aX0lqgXtAB4Yb/bQTCBs3MVEH9YVqIEfrm+gUaG4HKaaCv40zg7
bcB25o107vDFzRYKWJwtMyyRC7T98Wi50cIKZh4c7McqLhJ0RdMmUwg9QcCIMXcdmYDFYqYWHL5M
YNvuU1oP5r0U+CcCDyZJ93le2Hnzzt5XXnli0FAFprwHUDGqsIFv67PnIcMRVc+mhooQ1kwzWFeD
G9WgbTpctGXlr8NjQE1sXULS43pDJ2YVBsGMbFIa6XFIRK+UNZlS9flU/UrL5NwMuK0fASf2hrTS
xUZkfWnVFwei2Q0cwVI3FEgDLpqzXYBaJOjeDvX6Cg3zskyDebTilvGxJqVD6/M9/+vW2fXLhhG6
pC11/AeFcKBBE5PCD4m3nrV+MOkc+3FHRIWbw3HFXNEdG6QLoq7GjTF60UfB7c4adu+JzgFjRhmD
lqHwTnmlYaNLsboUb9hXkqa46qCMA4VsDZ11wW9W6mfmmTqfvN6DXQjwGFNjAE+XZtOKzE7U4Kll
KQOwbMvdZGrIsWO1fsEznmNypog964W7+frCdVoREGlx9ekZW2Z4a1gv9nHSl0MYaaUxS5fFWepA
yNJobpDbNFMnFbzvU7OmAeADjXPNMu+K5cRObiAhPicjCiLgFNJlQxbCw2Mzu8TObqMEwYE8Dr3C
C+V7FttSnpQFKMhy59WqtYJRHXt+9esXP90QvnH2UrbEqk1P4ji72CZc+xo4y/lpxiTJMCiscUEF
23mPUPr1RJnEHgVcESUN/h9dCQzM23gFDClI4EX+qS3F1XyHQvM0uFONuy+nTbo22OrXAT3lz884
cvCIYkOby3DUefPQWY24K1/6OTThlcz7x9gYGZxBMfzU6WtOVCRjXFjyWpNa/xo96VVBkomchMrD
f5VloXErVXEH3BYeTHsVMuCA06rwUHvhayGVcTNPbQxYdUAUOUwXNPzqQNtfXEheVBw24LUuBvPj
qbueFeGdfo0XRdky4kSINqptlQ2oE8SL+jP/U7fMBUfhx9WvOgNOcTgK/6rAQZFXIpdPMTFGY16q
Fpn0oZ5aaj0LnUArpgC0ACkK1f/rv3DPGRIIxROHrtfns82CyJU5kTfPJI+eQ2rlW2RHFaF/Rr2R
dLIEVYxUueUJuFojf/clpI1IXcr3HKgQpyHnhNLpPxOJRDTx24VZmfuviY7oTauwAkn1d1ZceqCK
cccEKlecmJnSlesHlxpztAc9oRrgQ9uZtSGzsNq6N0qTLPDHUREF7HBVNqsaY+hb7zrgEKDeviQN
B84/7v7o7RixS2OjjxYPJvsnawQv9bMg/dJ6K16hBzShWtRxlPZ09tzM/kBo3OjZKgBYdalWN+aa
wtxUX3ukvfd7k0AbTt7o1a65nVRo0KMkJyrTUPw6Kcnmvk9Ot7xEosdJRphn9MCl/YNe2PgyA/Gs
TmhfkvfBvDfQycNCpm12DLqRlE8ic7GM4L6AFOTuyjxJh68KGTaA8H2T0Uh+RVJ5L1wyQcsjSIVb
adyjpvTUxBg1xBJdZ2LJNOwnfceyx2Iu7yuYCwzWNWOy0pDwzyf6msDhk8qz+2O2emcqu6e4lV7m
rmhY1w5x9fNCZR+AiFK94FQ3iik4SX05p3JVUsFoxwQS3d9sXZw+KH3Oj+cRd2nQSbEsO7Eeh/wT
PrjI8EvkWWblf5gBIlqQx0yjbTED0sBhr1VgsQyA2W2aHjvUHCryswtVeYQser7eV+rJj1vy92r2
7ppA/L6rFFMyGlnH2EYBXj8pCg2CDVsJxyaCE1qKNc7qe79+PxVHOHExtCDEVBw0uSqPBx2AntUY
068aXm3gQ7OhcByCKIDNIkVxKb9H5rxfLDiLkCFOHw0Lyvl5VPeRp24JaHD2pNjAm6XAapNAhARD
1odvk1uCfPKatpjwKYlQmzc/xqK7mauSwHvrOSwXQMwQHhlPiEckFNnUyyQyP35IqVEbngXiHtnS
w84o/e6NeJWdkWyysajdPAFYcn8E/LayUPErFUCBN6A8VU5BjeaOJFfJyay0xGjSURrRzAxTHKoe
ey9XN97MpIERDqzFMthS8118RMoPr2baiJYRyWor58SalsZlLbmbFvSZyZoLEFxMoPPhaBIbZopl
pwFkxOPGSB+/rILYFxDZrCklznuTLPozUqfqkpBxCQamTXL2YtWNn97T+cDj1PQG3P/ri50gZ6m0
RiwsEDwP7DV8jjq8mXV8oak6LJMAxIQ9dh4cU1k9ZpQZ2dzvc1/wnlnmeBg5M8g92AWZIqRBZZqr
CttXtoyddSETySvvPKa9b2T3NJgX0sL5AgyNZXjjb8YFJONjE4Uz+upgSDqo5z9Q7Q5b/bsRGqqh
P3VO3uOh5Di206aIuwQI27l5BdoIZ7lKspm9lVILTc4qm46H97dB9VqEKfWDmRqsU218QCbSQnzd
4+ZH/NabF30Rb4B8uNS0p0LTfH1nmv1mqFwyX2I82gtSNi+avp3XcYJkdlJAQIcAF9Xb0DhyVZJX
sH4UuXKTopve+sX6byLK/sNvJoJMH8ENv/7mme0hS9ltExyLt1z89CPXn/otzEZlbRbPR+3elXpl
iwImfuUutlPmH2iK5NI3sw2VjEACp8W9BBNKp9w6NRVOILTGAoQNAqWvXW5NgWiPbg6h9/M4OwpL
R7OMT83vtU1FMiXHxPQhPiaoHxZeSJIY6cwwJYTGRUJMtXPuMX7kxDYh8gY4Z3pEBSQOb3MPEex1
rf6A0mqAYx2rYJHfqb0RtHBcsAelu5OTaQ47RfZYe95t+q/LdG9358P6sfEDmd0HYlKwfxXAORMN
ZYFV/s37uPfJt4rdSUkpMj44/sGSgYKiPmJaCjD5RXfvVyScSMbo/7wrYa2+avGc4VeJcQskdckZ
xgPpWtHdPXg3hiWSs6JeTb0LhBrzSdbvhBrCjotxx/I7h/uPX5PLnmcaEKsUZULftyZn+WnpjRn2
PcldNezoXZzmE6loVpw+MjVvf95MK8SO6DPJFQPbyoYXy6DjGCnc2j9TEPH/B0MQmVSOBDa0Cjmv
jTOc8koLt4IRV0UORRoyvvrwfp1YGyvxwJyWboe7S83sycjhVaL18LYtmC/wtTHi7yzrnK2LpWmX
BWyM0aKJtyl4XDOSNW7aIqiJ4IEeYAI21Z7+L2R3R8JBA96munpKJ6QC9D5PwuDh4AqU7HvO6HxW
5lEjpFH7nD28AgAleORi9SSQ5hOKB8BXGS7Oba2fWt01XoQ4Gv76d49VmuIFB5oW25bPqbmbntOy
ORYXDH6pIRMfiuEvSM7byjwwqs94ZOaUc8lSVkQQ7es0MUYqdrWZEm8Cpe4tLWYLktI7iMSJeJiv
8WZpT3oa5hA1CKrVr4fHZDXLR0OJjxiyML/UqCzehGl+w9AuW9TuaqYk3MOPWczwDWK1hd6Ge/b1
MdPM3b6Uppj9lF7Z2J5gcPQ/K6C3qNr5u1t0ciSLph85xVFuL4d07231sCLGqaD9Kw8temELY3Q8
cnENSMBoT+3SAIe91VGBIiDeElV/erEylB/d7N7v/gOCNrn72Tk1/Zj7mtBDI95TfhEm260sbp2R
jIQ02lRv0YUTUMpPRM+gV2C3IVKK71DAFTxmEgz01F/ykQ4eeiCDI/z4GV5mareRWIE7SYH66LGX
3e9A/WyLoEtwq1vlwa3Lu6DsOKdACh06TszKT+g4Uc/mROM8WmXCsuLuhrF401oGDqz6UmiAlcCA
B/h1uJiJ5DxWL83xW/Ilh77JG7PwxfaYtAItzAvTWQC9sjBMpY4FQFWF/5kxInp6282JOESdEMxf
ET9tXLVHElKnItoCEitOWnHzcciTGK416G7uW4C2w4F+hOgxX5O6oxCXmLbnrH+zB6KKjSSH1pdg
TTZQqGMmpLRsYN8IIliYp0tnnwFAsgruPpS796yTDWCQJCn3pBN6dvCftX4rM0Nv+b2RLIA3KCls
5nXwB7LsYHJv+k7VrxVBvYjbZAGEHZpMCfGBnIBdoSqVT2QgAnjk2mdsrCU6TWYLdThCCSOUzjIq
z0xs5nI+Cz1Hu9ac1vMGYG83BwQt8Xkh8rfcQ52MXx3J9pytMIalONa7fFyyoqqY2iTegJckLfE/
lKCcfRNXe7J+azM5uvOd0tQ1ztuYzL1Ztd1b9T+Fj9QgTkgB4g77zXBqMaPC/Ttg5VNnhNJxlOU9
G2cxwfTNi1nW/zheqvkXV/W8f9WSCh3PdfVARkwlMmj6hz1/KXdH2veWpyTFD2nwrinpCJOlF9Qg
x7mRCKUdW8X+bSH4FtZKbbuqUzHkEQu3kP8FHCSwbxxmdhwOIArjbZVzqpeinhCzzTfpCYuk7uVU
KLVXmPFF2p1BCi8+hpMEi8B0fMFvU/7ZhET7z2DL1hV9GK+asrZy8fwAhotyXaBl6itu8Z0KQgSX
pcPsvzQLf+0elItM1ewVNmZD0BI5bAodvFMk79T2/Jx2O1qcy0SATGC/H5oZafEWpxA9M69x8bjK
M0i33YTsJa7T3RuRuQTkHjW2MMAL2pdbUac9KcIqAALYEo9x8mP2fR+3eoRkxOLM6uYewjrm4u0D
bgp/9IXEn4uN9zH3xF2yR5+/xO2Afr0mrm+Xhj00tJO5eJqT30wVCEID/NZ7H36SfnhBTdEBCrkj
IQD4qwQHYK8g1o14mmBfBIGEnRr273qay7O88UBUeHuiPSMrxqGAJwh5SZHSm+lPxa4vy6jve3UH
NJdTsf+PlV1ruoQ8jOV7q4wWoISoP04Rdro0cmFPn/nLDRJVuRWe3jBN7XlKXWzN4U1FIIeoKwTv
NU4DIfKJ/UHV3z63lMTMhzkV13YaeiQuzGC28Kqgm6l1gu1/oi50iABeIa+jxZElITZOhB299n7k
k5CV310sNK7/zy8F2WgTca6B36lKf8HjzbIkDCjZ0xLWm1d3n4iYgjXBXZEv6aQedEdxQ6vzVJa4
Oim0WYgwW/OFLAK47sDuF4u0ud0vUWdiwKNDpTm0wVYsfr+NdTnm7iaZlq9VCb8ulTfevzqnczI9
1813j37RGoKJdMM8F5b6LaLlJRvckguXD95QLAzDT+lJ02n4Ik2YdHKhiRjrkL/PqJsJBfMGna/n
5+uyusKaSk1mvjW+K5qViGtf6l9EmfjZf4vVEafBKynM+jN3oORp1q8xYdldYnss4W1hKJH1c4/3
71rQXbk7vUFKh7vzceFxqjN8Hy31YqpuAb4mrEz0f3tTDIC7rba1BLpmlk3JRqxNruZb/4ZgNb+G
wasPElVgKjqfamxDECQzaLA9ZdzidwWGdyCG3CpvW5a5DECqvPP/UyCGw96uSUHZ9HjYzdglDG0r
Hc7cUPUDOGr0K/Hpc7GQfhjs2OeAtz5kcnbq2cyg0sxWmu0K56xJSiG6iNbclwits1upw59OLnI2
hA7Mp9yCWCa8zHh7mqKMC5P3Cc0pveQdxv5SotysPMXHQDA8erxRzjlNL9tlIjiFDflMSmP+vCSP
kJbMpzYkAnfC9FdzvrZ7UmFhOSA1JwcwwITp2H2clix14mWNGbDo1m4hat0xXmMES7JygyHWyMvw
fYb6K11u3a0LeJiUgFLW/22bG4W1u4TvjCE10YD08mnsdlu4JpjNLwI/NPfP21BBH+gTu13IL51p
07vEY+PI6rAhjeDhdZktHfRZrrkRyH6BdNKrSNkQ/vRtqRb994rCmosK3yM/0vXaiK5PIJHw5cUK
eNVI6V+joYAN+o+oMhxmBgdDgmYF6MNCd9+VGAMTBvWOZhu+gr1cWg2Jwg4z1FwgmDJN6uRxr9iy
h8H+Cur7NUwxZC2lyIcVP3HIQeCeah9hHF7gYw1p2SKKks92j76nMzdkhnY5lSBnqYX5rxzdLCJe
S6tQRd+OShvmqfly43npnVAXV7VZx3slNsZ5spDOODQJB9QVRXnWH/N3m6aWVxK/Zw6NlsaRDjFr
3XQRpMPgSqNQyMTwwshQEucfxg81AWXzXzEhmnRzy9AdYvqiVZDnstnAyPU0p+l91YFYKu5wdJ5N
Q/2pbBPcpRCCvkSLDK3PiDX06uKcpFVGTnsnqUIGFB6+mv/K4+1rOv8hzzSxCWQKlmqa65On5sz+
74kRebvDcX8p//dnDA/GPMyYcfHhZY8y7jdU1GktoM3pgTjp8VaiFHpMTNiYFAQewAK+y7XFExqU
v+OCneX8IA7ly0PToaySZsz5XMWBishEaHyIw7gPgrnhDith1txoDHw0DsFG/Y9JRGt1+fOk0xmI
N1rCzpx6fWj/ED71FesR3Z0VixI8oGMijjj7OhBzMGQtdpoPLnyfG/a2rgY7S4wlF8+jlScrYcPZ
7j9aaxOif9jtc366P1gYWmL0CQUaKLAyDYYOebAmDARZ/H0xf/a560i9Ux3vPMX2dOoFT4Iy6JUy
hMrx5h2tv+2MBbzrRe+nV59Ys8RefzfAF7J7BwFY0AgqdBS8NjtzKJTtsLU6Uoos+FQGWjTsoN0Q
MAjWQWDrv4M2B2L/oxBecdQAHBh9Yuj/ZiPR56QKT6lPdLKBVGmDxrMDYDpilyTnVa8vliZY0cZl
feyOeeQ0knzUVsxUbJC6CP0KHVwAVi7yff7G1BE6GtZo4qNjTULs/+R2y8FAiw+lT+ECl6k2z6EM
YTNNpZJ08bXQ/GQeXLxcrdqIoq+EQjZ4mDL6ZwRt3JzrJzosWlna5RV17CU28St8aAaymLT8jv+K
7YoNtREB8h03AKjoL9C79m7RdnkNJqHSjjbc0L+eXPrbF39aMeQrRqwYM/nUaM5fpFaAPUA48rJ9
SiTqkZIebaX96XAekpB0Yf+64u6VhfDKC/izozJsaSHMEzA3vlgXBUYk3lVr/JEM5gv6FLrTveFr
BwP7Q2UoI5lnaPPUHcZcaFktrggk50ibtEUy2hl8/sQHGpJY9q/IG6wTSC58h74YA6cVwdndyI5N
mQuW2tRU6fIvUuNvXma8tljt3DgpJtFGz72M8CsgM+Tm5FYR0aRzyW6VSv1HkZHMJFyrcJ+lFSsg
HxZ1j41gex0MK3OB9buiR0AUgEFIRfNvFF2sQt2dlWr4EBxtbOg0tBe3K4zhPR9XNn/3EiEYXKSz
363hAkZWsr9yMykYthJuln1EIocXM2n1Po4gzMbQ3APqyy/K+7gMkXgyuhNna4eZMO9rNj7KNzIT
DsHdmnJS7irufeUTTtYJxlrDmFmRcHWAUpqq9f8GE+BPooQ56KIDeV6jDp13IppYhTDe04u+wWSR
T32762oxGHj2edHKIu/suO/q7hjHV/W/GcFstv18u0CwPZ4pVS5OzK2U3FhVCi8PYnt4P6CnvamR
JN4Oqg6d4mxVMZ5Fe6sFWKsvT6kx/LNQ5VZKn0DVAXSdoMluBdon/AcNRAfOHtSRnnU0zpBht5WZ
afj+nDrqRwXRZZHCCFU0uIAo/ybEA0cLKHzLOQ30UFbl0YvL0Wka4ZClX8Ik3L28yyhXIe72CJPv
n3GVRHvVXMYn6GquxF8tZNZY9FtwgaK2WQH65Nz62aUX1qbmHM6O+7ZV43C133ZyeVS9VY8Ust/x
HbLyIzNNsTpoJONxGbTG2i0mDO8q7K4v2A142SqA9vH4Wn8BJwxK2wjg1ulU+mXls7ZNMyypSw8M
r2D1enr3/ghdR8iNCOI4Qmz63jxEEk28AKEEHq6nKSlue4+Ali+ltml1HK14Tug/EZonXFSTmQ1R
YDHwKyfy8AKMqEXm8zbOH+CzNdy9eMzKQkfzteN2Y5nKxmUv0qs7uP3Yat6soq5WET0IveHIjrec
yrNAebBiNfo+hEYzka0OORcHkDl+MptvYuA88H1C0EAiQQ17i7dMP1q1Ysq/HCNbs4WVd3lre0KT
ecEcs5zEevPlSUBaYEuDe4I4TV0S15Tn1PyRaKmKdaToAN46ZubBlATtiPQFWxep6k/LbCLXSusc
YLz/aIuXEl+ARJE66xeVyVz9Zh98xyRnrg6LA+EWmzne2bpraPEI28pKIEX5n6KggEdQYiV5Auc7
FK9QtqVvLx+XfUBZ/RktS6ML3ZGYCwEeBsNdWET0+fuuCZZt6BO/Gx4O1QBEBik8UeNSX6SWUccD
xR8bVaTFwGIiqJXjr7ZCU/TACHNhASu6ON/UYoyWVs6S4LYEbXOnHaoLKXWfbm0oF6/VloQ4V1pY
Lo39W4LmMzWYhGu9rgf9sSN6cQw9F35xX+aCLNEp5h+OyPr3NqYQy0O/FQCt0nSif+1a+AwuYV20
Vqv4wLmQI73hVzli3qmj3GtUOLn8fi8UI86P1LzvlurSNpFbPoRYW+Dja1/oiZKvgWt165zAsTPt
4qQn7521jrP7gc2+FGXsFNYG8HO53Uofwo3Aizx/pD7kOeXzFsVjrcWe8pUlrDIg03LFGCCYoIC/
DM3Bgj+O4pB8iU6VOcHP7XrSkm9f9BoqvhFES1o/Uze6XRU/7BAdzWhCukSVDRDAuYBQzqlp6rmm
OTMMFAz7D+T88b5/3YsxawW4xGb8acNRqro0Lurgoi/i9JEKdH0J5ZbRDjK06kNDubqOrpyvv6oM
jRuaqY9NoI/yDbDhCgyANwG+9ETJBGY/ZeRZQjxoBvsiNex3KLNKP+WN0boil/IurnVFjNm8gsbj
PY/XC3NEiDtV7fDebdvFUlIrsKeTZVPwUxa2q0Sp9vKzi8B/5GuvrzxMCsw9ygDOMadIH1AfzVf0
Eth7sChqQ2Z5cvc3cR3sQCHaxZuc8fGKOxfQzeAYlabe78g3+4087G3N7nzQokx16Dfls9KBLDNs
J6B2dep9MOaQlAWbbiksHdNB4YTZc0bDYN7i2crgPaCHA5XR0RJrQsbNCfh+Zz0V7xG6/Br4V9RI
PxczbV3+koCUmDZIU8KU6Cpsbo+6JcXpG+04UItehA+iN8OLdDuAwoTNEJgQdfcbGHWKnz5NleBP
FTF5N3MICp6CGFA9CBtxw1v0ZPNenNF1YoO77AUKKT2HHKT3xcC54Wu9XaPHUGtOKTPsn64ee+Ye
GRCDy8f8x08xjx0bl5osBMwuLLt+cDZNNgW+cZMU7Up2CNj+JLrOYX22sMEvux+tMyAG0WMibLQb
4nqRK8LYfN2OcNU6cTOxSpK+11bYfUK6l1pFhGLzZn7ytNlER49QechrvBJHqLh7PbwfAR4of7KX
UxJvt2py4ipSIgdgMnaFP6TZVP4u+Qlv8Jrd13FQUf7Y8PFwhwDYwaZI/+4tyRedWaoYT03ZYmM9
gsefrEv5sQfY5FkvJVfn2Cw8cd7hQSRKTK/xdAAv+z7s7/vWZ/6U7c62vTCx0IlorHW7tPdUz8H/
M1gvsqVJ2uR7U56V4AkSNUsZHLM10eDuC5EPHm7DRQb6k75RIRw1FA10RIUchhMYBTDrK2P9Drcv
Teq4Hu9wZsma0vzpBut0uUdHOmg2/1izefgDvWdsPfBC0kg7E2WGN+VIft32F9LmiYwNjf7SIykG
mZNE/p5HROlsCxcYPkP4UmWVfIXEyRaS+GbkQfwALeI7pamSiyIwcD0Wk4wQkmGLLKNJQQMNSrEn
OXHpua2q64E0LdhKGkCTQELJjFiKkfGcwfx3T+l1EnjTNE26Il8lyUUzSQgdU1pZFQ5XPWJWvZVE
/6kTSHuTsT2DqiURhR8oNKjnpP00XSfua1myF4m5oUxApgGsxB9bUqW5CYkZJPb98/T24eds4Nyv
0CY2F1oNHOTLSJQpi8nlHkh4jr1rTkzwUXQv8e6wqjlYONGNXvG2lkKPnmzc6X0Mv3sPSO+nr2dY
47rSN75GqJ2Rmk6mGcjIL2G6pl1cuIdSfOoV6U6JVGXcVt2v+Y7MMCj+7HaHIwJwtJupducQUhGK
SagOeZ7lm40AQBW2z8GpRgCpxYvxyNCMI5EeqK2O74iy0KRZG9v/P/erz9HmfEzaeZCOnKSRWOUa
DV9K1IfYaE6lrWyk7WX7r59rT8hlPpUFOff3++3vMmpE/Rrk8RIH8tUjJO3b5rZzhUUDZBqyBAeI
w5wOFfy0E3GpwuJjSYvb0G/51ZZopDICdRfeKl+A3uhtx3yg7dNxR/PXcifoUcchxyq6/AI75GYh
mFZG4CyKzsmYlI/e3uKwmZEFqOqDMsz+mOhJDG5slNAFCRyZDlLau82yxUicNz6lEqFNLiZnLemo
8cvbbG7zBKfpgSYo/vqjT81mm6WscA7weP2k0jNxiezgwaT+PpltVDWh32LRGmK4ZSBM6K9p2NWe
qhk4ppKfW8tCOl3fnnxgGG6p4kLftQybYIkg9qNSUAehpB6x9e6cfY8CLe3YHUzswwKvt5zRuD1u
nXlvPU0xovvMBBMVDApcjs/uAdAI1TKhaHr4guTTv5bxADW13u3KvC3W4cHRPGlL2U+rw3U56/GZ
6ccVhC6PKCUurhwFdLRn4YVeegG+UKJnWFHTkCf1x0J4eCBAsflapK2PX1mV9d8/DRco5ErMO7o1
BYhbn8PHhnBhQsXY00vUG3bbsAzm0BqA76RTK7xykaneybGmksgPE0lc4PYuUfMsKL2AcWCTvBw7
VpfMwfJxxLfQ3n0+6e4OR4ZZv7AwLGnHF8elDQvxS4m2JJ9I0okNUglmPZSYu9YOchr0KV+0VnbD
aYX+9+2gQvmlGl2dUrPaJtzlAD7SyhSJ0sNT/Ay2iH1v/yXrRoEp5NHTG4kNkofmSfmKfD3CTgio
aVqpOJ5BOCi1zY66uDqV5v6YiFU40MxqOBhFdErtlCSsE4yJXxYBjHeB+oW3pMMg9iGP1o8EKIYi
Ki7Z7lE6pTQjOBjbyShFRxoSuFEzgs/6XrO836LCw3Qwqmlyk9MAYndqYnBBW70pyuXR00q2qWeC
hlfj5A+PlwWZpGf2w98StJMUlC14WPvikJIjpPSnXd+5VGprlcAetaZqBMgNGu8ucKcccY9oZMSm
KdPZAOafk7PgRXe3xh/YCd4R0vMf9WjoiO7vdRrXprBQf/9fh9Xm5eXttZejy+z9PNXXb3t43rz4
psp/qbgKCFm56HQLnU8EvYMHibcBC9SU7oZ+0ndGU70NaIMWLRbCeTeO4z3f+i5iTGqxDY+5tSyS
EZK6E/KO9L66StlPgCO0KIRr88bHDCLZ8HutMmFnV4ZdcuIbDDofReq/PfOzXdB7iAEEl5OvL0Pm
ldt81tecksuRybvyJozPO8ijdlYzn8LPxpts+D04ILbZP6ngtlbHa8wypdzo9+sPNIjZr+KQmAaK
3g3ZM3EJsSxCkmtyWPmhtwOTf0yAyywbrFbOwsNOKA1peCQkc/eTngGxXTQeVfu3tYI4IlyKeOQi
/2ex3RK4JNRWjI4YUfRsYoN2UhtWZU+dNZ8bTI6naq3zgFFoo9C9zDgKxK5W8oGVRojgCtNSm5Qq
iHXW0zla11EpudTXSyR664+huaSlneJklwO7Aq1a6d3deGg5BPEeWKhba1VYTEggMILPLjkR4+M1
05sIc1zYHdK0pf3CJYLZMwSciL5VqoRkwBkR0yNVvtW2CIvtr1R/sgwKAddMYap9N4IO+5l3aTbi
LUlTYlAO2ypWXNywmW86YvgkBuxZUyoF0Vn6/fW2Qmd/NZ7Q0Hj0d8m4ysNzAlaYc+crzfCvtPM+
8sXvyrZO8sme1gL59p/uGtBmRfqxr7CkBFzBtowW3hDg4kdfbQW5T4xKkUujN0k1ly/47dDq+RLI
gK8IL3Uy6oFKaTks7Srxn0HWxt34dK5IqWG+noeD8SHusHpu5Cv+2YHxiNhTDAGew4/exZccsmbI
g9WhcNz56HQ+1wlL8sFkeipQ36L/F4L77zMRhw50azoRl0ukpRhU6IkQ9kLQypR0U+psaph4aK9K
z+8FEEkQ3V/PVdCdmCaDrWuSSWa0k9Fct60uueWTDd4Zx9MADBaK2TNiHsDv/PbfN/8FNwe3kLj0
jU7nfaTZXyZbF0OFM9valcDkox5v41xo0GWrNBmwURteHztobuZ/oEGkao3YGBt6t4M+wrzMjTKq
1SN0aKr8O3xDKKaICHQyrhA8nvszFcLz9qvrYd3p8No1H//27KmiEBDEnoQpNmRjvYyz/Eocn/kx
KaBWJjdiMO8Yv+sQgAWzMMRKlZe7+LmZ6YYMAIWHlRrxbLE/DYln0sYASYGP1XCoDNsSRguAQjWq
rFJ+zvu3ekXAy3zLq9wHNVp9KHW3BAcKlgHRfrNSWd75oJdV3fjgGhSAba7vV+e52/5AIVLFNsdb
mLQM6I1MI8ODUdwPY8eowRdVCgcWAhzzQy07hrvZFfbLTlRw1njY6Kx5vkgnu7zQBc7lE5ws4fkJ
Zcm2ER+lQmG4RjkUeo6KPLKKIB2q4iZ9qMaGwcPE1Tk3Rzkboy4LMoogFwrwKkz470x6h+X3D2Hd
TxtkXJr2u6EpjJUox3iv1qieKC6XiFhR+iB0uCLhkuL6kWtRryryAWX5alRONtYKO3JQ5s4lvFvW
31i0PMu6GNXn1BBR4A/3jUSySy15tes2q/8oDK1eYsIg37ADTyNKR7dASy58w9kCNpWgKnuuJxzo
qkJMAiFH/r8wIpmnpyB2/oEVYXbs5fr2N7F7T1Dd44OjT+KaL0xOksn4uqf+vgliUOX81hZf3LVf
v5UrmYODIZ6Kcrn9Ey1jliPf33o7W0CWvYIWM+XchzHG7BMUp/sxflIxwk0myr8NtphBwtQTTtn7
Sr8mk0YVgT8Ala3P4OcppNapn0Lez+49KxlC85lyKTuup6+jpBBYw0lbuqKUnSzLZzTDJcKN6w35
vVaJ5GvCnX1Io41gTnULcQuUi+xi4Gs+EENnNvKCYYqEnNCTtLyKni38xZLH79mPBDvL2HDrnIGR
rfwn2dHpA9idji1iefGSpbgH7v92A6VwTV5AqKYRZuGEQ6gn/ogp73UagKgJg/yvqh7OwZKRKDQ9
YQvviWBXt6/rRdj/fSOWqx7RDfuHJ3vzUH6cDj6aKLqczCJONt27LpitN+7ZBZ6aWr3VLi5n/BMB
9wXSs/8w6leEtYdEi6sLciY99X7IDb2ZBZ3OR+3uIvbWBcNpfF8Vy3UMb0jeQHH/e4ROc76NGvpY
YTyVd88X++4DJ+i1ugf9OUEIsGdYYIGTXs9Y+npVL6UwhueElNh6pGH4IxMujcgWQZSoXSEHo/7p
lKyj3p9jzc80GXqqitkySClcAXThnubVCw3HCvPx63rjWyUhdHRY+/ma8+HjxpyzeG1vL3hAPITr
la1HNCf+mDZZ8CD704lfKrnhqsnibKTH5DCGM2UB/57lXGX1kEOWmij+XlHqEJGFMRXzHt7EwmMV
+dWHfiB1dTJUVCuJUdiJEGWaVazsXnqrrLgQWMPsyuSJVHiDMpPsK+L7rkL6bXDibwescxM2uHez
uUBslb3Hahs2vpdzVNd7/UGITl3eMAlVgVzbntsaVLovQfSFkOya04d7BMk6BRmlJM3XGxThKIYU
B0gmKqXXVzFAI/AQB+PXrYYjUr08MRGe8XvBWjhbcXPCkw3MeVknuJlIPvEb+ueVtntymZ0arVrR
5S33cQFkyiPomPZxIbAgS/QCTErfj6P8oRviQnXNx76ee7BwaWDdhEWUnXFh7VCHUd9ZxG7/7PzJ
7uBiz/Z13hAwieyh2KK3nYNKbojZZmsWQG7XLst+2SMqi1ufRmfxlEuP4JqZ9xlrcwYDlHvivTK3
otjcBPdBjB8stnXgVomkh0qLQ4u6UJoCBUdTQJhM0Ke8HiFcWOYk27v08ESlwCujxPSO4BawAtzW
mtdirvGamLI9VR08Vj34uucTvu1OjEABKQZ0+Weda1Mjar2FE2fZyhVvRKjGSMQwCZGdaQUYfGzn
6f+FuliP7dvD0jPLLVmgg+HSsLrl0OJs/yLlywVg+BvOnjR1+UZksTTghb96mLHnuWYNSe26AWT5
vntbjWd4EnFbMXGVuwYb/RsgtCBlolD71+CqvaQ/zp+3ROilOroVT+1g7qnVu+SeUVzay9Nwgj8s
+4m0hifhYStgslywfvj2a8EE+J33HoO1XSZv6mY7A0N4OIbaDV0HD+gZEGXYF5rOCNtoKC615A9Z
vWhDSw1CNu0vOf32OdpYYPismOBjftfdsoQ9mDvgbaBPA76k6JZprpkNVJlxl30UqFE5xhjUbQ6n
sxuXT5htpop9pmSUTFU/3IN8dOLHnJBSz3MEmoS4Hp7ozCkzeZXh+vQucJSUNDytAV+vHv8fjpgN
Alvjp4KqwvDQ8HMFiC0JGDOHO/xOsqLMI8/8PU8t8x9lNS5mfw4wChWB1WP2zSJmgXBfKFixfiDv
mg3gAJGVGoEkzZ0wpHLmzeG4b/UdB3BWjJW/panMxb7sB7o+ekX/+q5s8tIhrnugkXVRN2X1bSX8
oacyBBrLf22Nw5hiSLFIRd2oSzpPm/+01qqvD3cyFJb6ysIcCpBIneQLAimp3G/u9RTAeOLTCLGH
e8qCEFAwVVusKC1o6xRUX/Ed4hlOjoCooCGvGxb+TT9Flvz7MFSBqmIZo5NzIUt/d8ujvQI0Aff9
HDdWaoEOK0XDnI/VoU2J+8upIq4IkQwhNpCng6X3AqARh3+obT4rT2Frc75mcmow6Mal13mVN8o5
reHHGw8FTNPz+RF0Hd9fkqzfxxwvk9W9LMls9v88E5C8vTg/6C4u/Ctcd4FOSpz+eKf0ywwgn0YE
AYNJlIebRSDkBoZTuewtz8dartYiwF09M1l0puVikrgfJvrxmlanA3WBmRALXh70FDhbUvpbMVvT
cEpTym2kBp+8chhxkBpduu9wLRyflgjIbGhyNyklamVyTy71MS9UGzodryrOA7aYmUcu0EzXNfB5
xqlLmfAMeSS2tvrwrxMViSvexOHLUyiPQARSALIKlqsF3WJ7A2Uq2NGjzqUZasVG95hnBFFcV1fm
d/EdDAbELgIG69iCKk50CKhf9mjHSbtfpcdnnIe8linHH14WGe3b79TpLG6W+KDCvRI6WT4CtzC/
1xwkkKC9Vzgz1bL2nuJRTyeun16mD4hu1o8AK9bG8dam42IDmTqnhQKc6G45Z7NATJOVCtybdFul
2w0fM7ADiN22/K/XPOn4LQT8md5ygGJKumaz4eeFmUtcYC0TbW8Nf4gdk7j8gudwcfeU6/QfkvL7
jveEMXTHDHfGdcY0XfxQoXDLn6A8HihvMsQ3fE2RcZXIKkN7dC5SqIQKoVRUsnjmMwVH5Z7GfbXs
pEqndB02vAl84aK7kTPtVC7MwiTgeABTbU/birGbJMCxNoREOrI5kSw8svi9QQtKOxJX32G2EQA0
Ep8GTjyeNNl0Pj2hS+TTo0oxzXEc7xP/gJdYFnVHciPQk5B4DqkiBCIyau21rrfVPbURglXD5Hbe
Elb4mXkuFrJhkFXMHN93L6n5Y/kjxxkOQFa+fRrV5PpAiLsF1CDwEKzaO8BSV3CKgf+CZ7FD/bS/
KjWCKBUvEVXgwTG0naOannm83UQ7zltiyvL2R/P37Cst6l2l4p6r+GX60pfDO3BI2SOCT8HSpMiH
pp4cive9u48xuaU0DyydQ3PLhop2RJ0aZROEqyWNRitibhzs3YsBiL5OUekp0n918r2nfgi+HKf7
aKrmE5vhRjjL0A41oQLXUcAZckNRm5rmbRafwlA68AGpG7t9/L52i29tGZei0abvLZ6zfk3wxlMy
65VdoQ2XHbgkC6CYpXgt5Bc0hssAedJ6uq/Ffh3tf6UKDfvD2SsZN+HM72oUgbIrosMP8yVljygn
IGDCKZ+prYh1JZqVnnjJw3mOQxc0+PPlZWGR4P2lpdU6UqARY5+OBRAfQdz03JMqlQ8pjT8KKYFF
7us/B+TFFhPyFnZWEELzKGLF6Yt9X+O8gsI+ovxbpusY5IyO3g5qtisOTgCt2X7920JDAXnE5ny+
BFBXQy7pcYfINKVvtPI7IceZO01m7a3sGeidN3hFEQjgw+CV8HyV9OEQGS95VhHUI+XZz8IcS0Jg
walinHjkrCZGVkf9csNFQWebuKsmXzSA7mJfOyiyO89JasPW9b1SB8wHSzH/uaReLgAsuPpy4cS6
3B6tn9JKHI5httZZxgq1m4HpTG+9jiDuEuMUez/a8e1bU0QBXLFnEmweBBvKBC/wViJkLX7LWHT0
09fTxl3sFRjhmqMs/AW2aKpF5lSA+9XlLNcgSGWYd7gHcVAm711lZQfIl8wbzbKCTgDkaD2Qs/FS
P/aVs1Im31G9St0qhO9J4GJlKrlYy23K+JhnAtpdckBs0Tn5amHmpCc4gc23+toPO4qGcZ7Vm3Nr
XV0eV1yq/p26rpVk02ACWJXKE8/V0tR9NnC0xqYkOl8mZbH+jwFuyFerI6Y6U30ZOXHwvuLtQPjv
nVRsJhN0yUH63Xfyema0+mzQTem8yo9BqP7K9NypXV6oIg4hrT0FkC3BzCONGeuwEuT9h7KgK1Dw
egrTU3GcNJDRcLAU3UUncBSNiInsoME3d4CNE/wu4+Ap/km59XWmqqgJf7eusQGvYqZzucQaMKEA
bUUSiQqJPE6hFK3Q8Mry5h4jRq6hh9ZMadjUoU0ITNuM2WjqFIfKaEz5P6kEeOg7pzbC9Zoh2W89
OF/8ZXMWmpgs5tyOa1jVOYti21EzfPP+jMDmVKOpET7MEO0ndqunCa5wxUXrigMXWy8yKUJxOnVR
HZgehAiCUEKSgwvO55HwGB5G8W1g1gsrUyR6eFfyCVnt8g5X3QW342rT3Qhq80cnjOqNSkPmuRh0
VxBMw0oJb3KqEvenckL9T/khCnJRGixrLSkLmB5NkfHZXc5EU7hedMFQJRdgSAzV2o1Y50oGIqXo
dOgAJC4RXH9Q0XCvVcAjOMzWOHNZUxpVs8zmnKl78evpptw4q9LL+xRDf1YOq83hRQ+OHbYbD4DZ
OXxMrYpRu74D/vPXVT0EZsxZA3PDtrapmt6ednzTV58rQZ7+aP7CxAGjItk8uY6Gh+wPKGAYxKZQ
gczVQC6cCvzU4RYF9szO/dE8e1iIiPExCrfMS8/gHtZMOguh//T8Acc1jX2El4T7C4lWlaKnVy6S
YpD100AKTom1MTjEWu3czFIoEDQb3aW0FAjtkaKpVd1UToxx1HXJrfMn0szaG2g20vkKOcSBdccw
Ru45FtNFbOFLZltSoM9eaJxyQ2XcNVuku2wQccx2dTmPyL7A2ggJ9ldwgk9zH5whVUAcdhXfil/y
Mt7kaR1o7s886i4wagXCi9R5ICb4pcXcj9lHYv4wxaFfhRTmYV4BiFrpu2If/HDLxOuJvjYVDPhk
bcz6PrgbVPglOn9bTO8IgGDYN2QxplevrDz8vkvAti78koFhGlPC842Qz6RKkUahIcOmYo7uN+LN
si1MFlIXAshFpqQKDeHl2xP2gPZd2qo88DNidVTjpx8MFg9tpL+1PoF7ezFp6iaNMPNH8w1QA16N
GzmCcqbWZsJ3WP6V9KoHtq7h5WuqXpfhCrAZvZ6lrAbE1F+NJlEfP07f+IPQ8nPyNklW2uy7FX97
h9lnHPHTZzE5EcBt49+lpbxia1GAdZbRh+F9Rbc8WH1W2LMom599qf8xgDqanG1cencAcSnw/MRN
4HA0Kx+xeO4u/kFd+Dk4I9MolJIrClBljfWGnzeAwZCGZrEvtY3nD6BIuRrrvZVqPDZRRLeXZVwF
xMctVgxFs4aJ3EcxoNJIHpF2pBsL9Ni4l7wua6x4REuiG4o4q8fzA5fLCjDwvldolN57FJqNyEUs
/h26d+klW2WYhTudA6erIQ3ExTnoH2dhCKqiNqOUtf/Pl4BSa7vRCRt/MwyZtC+3t31JvVUYPJiZ
Yg0aE8RcTyzh4cTZ1zYNB4PZM8mY/5eP6uBnGZfi9mGCTZ5vquOyp6utW52n05k9IOMhoKE7eXge
yrxYxFAxhUhNvLYGs3suao3daQOrqWjGJ/hcPjbtZwLNu7zKmGpkC2wL9yQcFLZfkTDc0av1HVkQ
nB+3RZ10BA2ritCp9MzaH9B9vceBPICQWJ83a2ceOMT048pymhLOydR/g4a+sTfXY70MoG6+yWkX
5E/9Gmgr5w55T3PezRCsCKzaEVf463QDZ3p7vV4TDhZ2qalCkF5XT0pMryNa5h+Ry5FbSyTYjQP4
eR/e158FK/I1h0bzK5O1CO8BzS2u6uQ7kAQMKPe4yfjZ+VM0IZ7nJYxZUxzDMtfNr7yRJzA5iC+3
KdZmEONWTYygz4mdQmaczhG6JjTUxLg4m7lVyU096+qLmOiApzS9xEWRrJRw2RcUA/3+oCnr4yVz
Cn+iJZaEO6be0/WUzAlMb1z1Mmp9TN3O/XwKr2RgK+Zgr+2iAlpBI70aneEk84FBLJjorWJtG6nj
zuQ1xiaAqCLGW94/LJvr7PQZVKOn5W8zr7H27Q8jQfH5+I9xPtb4GEIm4ZoP6MUarO6o/vg0ejUQ
YydfW3HRfdDTMxngMFSEf7d0Ytj4PpUiE3kH06On1JKuy8V7nqSf6KYoH30qAFt4rUfmPE/LZo4m
aWZy+xUzrDI9+JhQz2AL2Mu0nwTr2GH9j8eXqkPQExM8vwUWv3qFudICJH2v3mbjfML1D713Rj4u
fnMQoQiS4P/vqHtCvY6KrIVqGNelKsxPM01hQ+WMpI9zdNXkqcuN+N5Pz9g572ENO4aHd8upjFF8
QD2Nd/2/OsloxWYhD66vqeVtGM1h/4H04MPKXZjgqZeoVfwTA1WbqSXgtufDUxQVEGxWeg6Uh4cP
5ErOVDeU+QbJMk+/uu4Nu2kUvntVhFnODKhTTTGFcPPxRTXHFDNOeXWdIv1QH8eCFkHHAF+u9N0y
xlXB0AvF7fxruMEiANhAwM5nB4445rYWKWKrdKbo0xqaty8KFkEcrf8Yr/N4Jj7+ECGWqaXldQQs
ZDGvVQVc5Fu4CLWQuSi6BQNmxwaqpI6ri1zQJ0G3kfVSrqGXzAyg6Sb+TPFne1ezDmUc3ZIGfNG6
170kxWIy7NCQpLDrTwOSCWm5lDZKDepdA0TMLK+pv0BWQPb2Sj6KfbIpRVP7IKWyplhAYA27UTuw
cHNSI3RDJKabKJVJ69BYWG3asnxHiVoKynVO78HwnbuDKLWsLM+kVusaTzFANW/Yod4cY5Kt0A+c
gfODJRATx/fahO4w1PFy4Szdldl08+6R64DqslYdr1iBtGmZJuYbPXxMs9yPopH+VyPsQEW/S/WH
5bcjSbtKfxO1lY9B1hgJ4x2UI8MyPnykHUrB7q4gnQXkrOU01tStqcNuNFrlJ3JJwUEWLf2LAzqM
SCXAZ5sGK/WVwGeMmLP9tslShV/kCudiD4KmIxtANkq3eu+fn1SEYc0FRQXW1WJc+dkn5liTSbAX
7Hipw9RPOwzw/aBQ+WV7OFNSoa8ZfI2COJ5BSXYjpjr9MSVNVPq7yxznLlCUi5RQ4/VVaWwvyY/1
NefKBO46AHmW1kjqXrpDoava2ny2tJ/6zBPy0YE/jUlVotJM53Yr5bvr0155cvlaeZimpRkCovg1
geM+/z/l8UozL+yq/nJxHhBkbBaeDc3Mhcj67GvDNFymwBJa5LO2aZtkxPbcFPDrW7KiM0fez/x+
EhVjPu5vtV9y5gJl+MugHDnDd5nE7qga7kL7z7ROdf61EFgZcL80YMsmDbffXlJwBcTaEnCqnRY5
3D+fCVSGlH30v9iCAYhXY2HNjw+5guumtFLxqCAtepCh6Bu6PL8MGshLzPv3scb3vX6fTWKSIerJ
1Xm+gC9VT+EmFwlCkXiWhD6Fetr2Bqub4Gr0Zq9jQni3k/OD8JtXp/2ioh9ZXod/0b2YbJsQywe4
LhPCUFEyJxcN7hiPNSQ6ejK2aH5KRCJnjfLZc8hGjcSq0m2IAITSiP8jgNsHFl5Gz0+bkfnK7kME
b/cMymtmKnCIBLdbNPsqSpiPcZFjTT+bLv0jh41CxBczUFRd2Kgk5zlvBcsQvC09Jk4ibWWE+Wgn
jWpqOGA5sd3djc3UfTJdHiMbFZlIxQr+rEEiUMuJyjgvtObYWhWrGea8ixpZL9tjLed8MSlkRn6V
A5gLUjMizdpOqXZg1LcFksEGzSH3sZVMWc0PPMkCQFFv+NwsXND05eg7fd1hZZvfCQW8dhQSZgM0
RdpR1CgzUIbPYskIGms9vBIf6FzcgCnLG6mWAI5JK4tBNDBXcdzxIEQpxd16GTbiP+HOG3EINerC
31hpPR/flsC312jTDnDZBJqcgckhI1YYcVobwQdi7E/fDUohFFOXV1oRZERrrMskayUDWTln8PM8
BuJJuNTK4omH95TllA0QD7wN8vKqqGaYF0D/mAVQ6TS0cJ4RXjMCTcTdwB2K4OVYB1L2thTfBrp1
1Jlg2SWeoSWqOTsS1pot8PfF5JLc1f0eAaL4xJbk/Gf5Gfi2b93Z/k9xA0z3wgrIP0VE1XtYu1pL
6rTu0lnNa2jjmIs1VhvxzuV8nZiaHBGgOkTfz2gM4lZZp6y1O9KPZImXF7bvJ4DcXVjHWQ4I29gO
XaMJgWpurzdeXdFa9ZWnaKqOoYFbOkBWQkXVXUdE3UIjry1eald8k4EwHghvLZH99SfyelcKCsnD
yFS9+GZaohjXD04zcEaplMh8srlzyaen6rW1CWwxM2KCV6VQSt47mt4jc8Bp625WHYwZexx6Q01Y
OJLo3TX082dqLSS/etKiksCq6dBYYyT/815G6CuW1zftZvXx7z2wq9MhPDo3KjXW9Muu4ORioPw+
AKENOxXDafLBjPbrRwYw81WIBn23QMPKK98fpzrLo8mZXhBMQJ+Hin95dgKA8atVvgg+mgFe8DVA
YZ7PjZlOJDOf2tNdHfr+z+hyar34aQiJJq/cQp3xyHu+BR5n7q6WrAi/Kgs2b1Fy8qOJ3++VoJDm
k5fzSnuqfb95WAPVQD/qEJ7ncYuoU/bLyg/P7A1BOJ/hm4R7y4kaIGqGC8tDskOlnCTugd8NkGgm
KH37ul78kasd9ReHi7FNMVcNaIokXgwalt6bK+OxIgnQSyRCGE9IUvdZ1YLlQF0i9OAUVPwo+xam
UNEUI57TNtk1j8LaqgcsOf4AFtKY70Uc1rDZcIp3U7L0O6UM/ItJ4lcUVPmMqakAuUPljmSWQ+OS
eq7TzHRXl7V5qzb0hRG6V5/vegFYGRq8s/87FdPEB4FTEaDFcckYfC3MhIwSr82XHIN7uBpKHFT+
RgLf4yV49zjky0hiIJf7892vRjwyjF0q34EKwyTQeUxb9r5Y3x6ObHDtXX5yFEC2bfV1W3uzKm2j
NiUyohZHBiLkFKtyzXLMajBcrvVXknf+u0VvFbANrfML2sa6solNYxDrImzqoYdiUyS+bGYZwJfV
n5KDXExJTTGMtS2lDDO2JzmJRfl+KpnHPK0B+U8tVktp5GcOhrhoLY/sKJrZuI7YRLmWUB/U144T
Xvs4Urf1y/75rWYO24h7h8VzTxU9H7qx286h5rHGwt/56ZjWilJqmFQo/Oo0pdGKODhd1CCAHABb
150BTkJYHyzxAJj5mgEQCfpcUM7R1Khct5ioGIAts4kI1xksfOTXEWEGtoqvy/+xwplK0Eyx4vqh
OOycTs/PyQhc3oEGCu/lNVq+UVXUDhrDhYSF9dFLOHk+vN1xxLCMFhNV78CU8GpquHbCUPdB4mg+
YuKWnYqbLhBMti6b7L+WX5JN0dC0gK6/XV3D2G5uv7wHGtNd7Bir20e2oDbamXLZ83Ao4zh9Ev+a
9B/78hetEByyUyXY4/CkZQmYAv/JW0JZKWVmnkxePlkaeUn+90oFGefxhlKDOReKXPRhAE5uoGxi
kW0VQuSun9Y5O4I01ti7M3si0am5ADghpEHaDtHBVzmeCfCt6pnPobzmp0CSy0B3cxBElddn5GFa
uWhMj+6k/6g7p/OSoxD+vC3e0c8rLnYpTZ2zbklfaUeJqdB6vmTC7GWzISUJyk0sdL2s7Wtmf2c7
rEE02EtvBraAw7BeXaJRephSajFKqKrFk5EZWsqRgX5wWmfuth7kkdAFgp9c599RQiriGolzql3S
GYbdmrLmEeU7caBH8SyajKA9eGqHSO4RcogchGkonfs9pStdJCGU17Py8Ms1kVv2FNI1GTShK76e
JzeFFdWTjEfIDkM0+jSviN1O3+XAONRAnxgcgdpWAv/n6KjaNTJ5shhCvVsA835eoMqBuC3O9Gv2
/ww6U3CRl9wZXgeqm7b7oDQmNNsYfD/Rq96WO/JDMq3pSkNszUicM2JZoi1P/dysS4+69WWLYsXa
051GtzbyCMAPrR+p/AP4UjBlApgnUCiowUROz3Gisq81cv42y/qzaK1EjmNg7Cy+AP8sXHl2KkLR
ykaQnLZ2wSERdRseUTHWUsNA8+13tqhT5Xi3o5+RSh2Hw6hNrMvCKLczpvW8COajUZAmWBWvI8Mp
StvBNHLPkevtzr3gPWHOCLedq8k19xpykQSpdAFK2jOsR1dyZWnSj+CMwwItWp5J8YKLj9QvRoFO
a5Qkfisw7C6NUWZSDSrXZSac9Wur/+1l6IEmXAstZ+dPV7FJuX/9lX4wpdC6gnLDVEqy/FyxzzUC
Qy0i1eDQcWM4Ly6ErhO/FW+iC6lkXUO/g21GBODp6Xunb80jA2R1D1xgt4z73PvOhFz6TbpYjhVF
qY8vfeLOPL6rzGsDVV95x6qxlOkcl2cavA8MYDCiY3qO/C8s2nerQM40dqUTSn3sJz1y5Uke2CuY
GzVA9uS37vKMChUCMGIS77bMFbQ1OFAd53/mDzzeOobIu6MKAxErITsVIKfvfWvljVKZq32DNlSO
+cQSpicbNTyRrQxNMAqwAMWnvZslqwtUvotKk3+M90w+W9OSiy/9/z/MZUZYCCkGVVIXTjbCJY4i
+5cLPM+XbQxErp6h4Djok6nQPzuUSOdFyBhGfVwjzU90mIE1F/dPfxefMX5hbabKBGOvgoFuBBDw
vE8CW4Mm1XSC0NwRm8JWeP7HyeAzGPB4raWH3wSDuaVhWhl+eXgpozpntNbDbZu9S8+uU9hpTubw
BMiOBOD5XiGbf0vMqEzAdSdvXdY5IIbiv69lyS+XQjm5Frd/7/7abmtwBOv4kd1V1xga94stz4cJ
uq1noOLx66nyQSjhQDkHID4IQbBVb5RQnWJObF+XhHfPf9VsRoxpMbqq5dJQ1ZxMeYwqtZ+WSFvH
Z8W/tLlPZF1kMUw0d1M8STkEDLjhEfOtilHaxRafKYq6dpWXd3bD1hl5QoqbsElPo2h65SISkV3H
3oP23kHa6SWqABijBYb+AvX4ufRCdYQ1QRPmEbg0zbDrIToXa20L5ge25VCs1EWhQ1vazGL/dUHh
RNZZXue4ssi2BmAf6x7x2uQvKvyPGJ9UY7zhvF2JxIPgJNg7BOYeMqbp1IApnnFql8QFJGv3Hnep
E6mKZ0DDKAXrV76E/pTvxsHk4RUWjEgXpBLgKb8R64MIoPufkhLVx3XSOj2B/TXSxfhfzi/Au/zW
V3sVwl+kuCzMVEuvKmpCb2JL1VoWNYmJHnnTNy9tS9MEkYgqvfaXyj0VtVfMX1unT5FeuwtHvaZS
FfERNkKUAJVzPSTy/l7DvkkYyck7N/ot4sjBSQtBZ31sMb166oRLMYfquOLOXS7cCrafzN05KbJS
J6OIkEHlZMl8/ufVK+KzxI82DoI3CWHENekjG2kcKg6NTkFxmjN8UKkSQln2zxVLZHmqpxEPrtwk
EjleOluUhnv0dXcv/hdc5yN8QfITdEjUbXgGbNl1VTc3zeuiN5sKMQlBrmpN6GsOrHQkfIb1a62M
Chc7m5Q5tWc+w7u7a77bfWV8XrxArt7/kmpj+QOhL68CD7Wh5AWBpb4CgiCfkzld7cAwraB4xQS7
/bjql0f9ApFS2cfowXCTRmapFZhtDleBUXcOucDkvkDrytrl7fmfe1+bpF9ujIWyzzXFUUIfOIR6
6h2Q21PDZZjL1k/FPcgR7ZQdtBXzwydvXuMg+qGWMZOEKK9n9t4aO3tV7QtI2SluQ/AYRVIYQWwl
gp7BUUE1fvF0VYsjoZYIWN10tBDLy1UkmT2X4wOn6PuDkITT/g+WXGrz3y8ISGjlHriBrG70U+lF
g4WbEtVBY/QdFm68xzEYlGKcgnQ18BmbLPwfWO8VlOeB+5NXWXImcEj+29lkkKklB4L1yBtdSir1
BOcdELF1iZDuprJrimlp1U9dX1vRgFLPZ2j7xYYWzpG3zSNkptCkOt1W3J7HiB8Sc/j346RdWgCC
sLtwuVzvuswdJe6ohaFhLa5taxTB2w+b90vsk35cNW/4VaGbQ2vYhQE5+ruapUIK4zk95QgxaDJ1
eRJ5O/YkAMOo8CP9FzWUCiG5puLbWsofBDH0frd3gr6Q1HRYuiPhv0BuVjwrDU8qeA4H9xqPiS3y
EyssDn8bcOjTC07lCGCj5kFTDQsH7L2Qi+Z/wl5pcnGOrlpj+cGCSjjWP4r4G4z6LeeEGhgVKx6u
hrQVwyJdMYCcEnYYZg3roqcdjGDxQwj9apARqVjHmipQ+ssAlmZVVO8Ke433HOHvtGCgO1lJBXnX
xKnLL70ZxN/p0jiBIKmK3lBEj9Zd3AfIVJdy+gG6zZKZevhOkVAVqj8G4Q1GApEtjYp66TQ9LOjL
LCFmXb4xRx383gWDO8ux54K1y4RYS2iV62rHwmqyaD1EFMPeyEban/wDAqUdStftdjJ23k8ktT6B
0QVl2tWP8WooTRgSClEfL4MGrsiFM1xr8Iwn1LimTyesGlvfYc9WDSfhNEPn1gDFoHoO1yigxLd8
h+1HxXnLkL3bh5Gw8h6foFIm5ufph5rpgsufS9jbYVt0piiKluwQDa9pgoa6rAw8KH6dBV8isTlJ
BNnLPmgZKfbqd6QrMK9dcNxIqe4O3OlSIrRIyHTEPLXNH/2rAUWrV5UmKsoZ+HkoQO37nkHYFEpB
vE1ulhrhOLs3GD14P4nGSbhFn2NgogB48Vr+MFa//dVtmnsrLbJlT5NQP4fIMnkx5nOt5S5QjQy3
po3a97UfvHkp4s69dWsosfc58YfOJVy4TKbHbg0cS4vLcfAiQJkmlSQfZQVJQDw0I9Yidj6X3OE7
YkH+/DpfzXVwBn0q566WorlvCqm3TxOxhuI3ZLG4LKrNQtf4bSB/nUx73vnPk8/jOmwONDQf/U8f
mNRSnGTUmQIuebeVqzKP+79SLfrQ/uB9DQj3E9MUTpO6QZnr7S1v+pl0LJ3Av1VlgvyLIsxcKt+k
GclHikKjiEn7Xv4EmY0Losu6Ap2dDdpWtnP46RO0LpB3Fwkbp8R/6JxVW9mDgDucaBtE/xFDlSna
RmyimncWjq8DrvfMAVKqCrAUlCRhPhWxU6M2v8AywJ5iVhVYrSppEhMenMPL6Ov0MGxLtsGP3ZZg
KDOu2qpf1tr4tGBP6t3u9Es36HF//L6fG9Dtw0ZSlLzuiFPH5nSn+TvS//z87QKYoSN2JEiGs16e
DfNNHVdq8HV1IQzACueNN8YTWX6pZCfOnQHSskaA6G01SwdRAIfMSuEZJvqv+iuvp3ThZJ4g+Hm+
TMjaG/u9yxIDTdOHSAvReSrUk8MNOxFkXFpIb/3UMek9ynIQlEz8qN6Rvu3Q6ApBXSWMAuVEaQud
RhouQikQEE+/yY5ot0uXwB/MVxoCVTMic34DVSNUma9wulhq7OvB5vmCshwTQOb4NxFpc44KG8yS
EEoVX+SHOoH6Hvu5GHIJyI/DX/ZnghD1ZVsqkhfwniJjTPwFVTvcAFermRRvHqM3Fc2t17tpZHge
2MNIXfdFUBnTh3tWeoMX6QRHTLxddcK9QlnMrEjP2YI8ynyBsIGUqBnYAmaOOuCVnXCgtg4Zq0Eo
Cb8lLox5OwfT9Msm1ochR7OEi82PkSbI770ZYYvbrfswelVpABnWAKaEIO0DsgwkNXf9CcDDqq3M
ok7DwhPtnhrp8tL9l8BMsvMYcFz4jmrRy5VWJpaMs9nb3LmHhOO+caZL6rZI8Qr8qj4O+xZAz/fF
CH5x4X3NV6hgh9gXlAC3OE/cmaraRrgrYAAMutoBI5tphsk4v8mUbB5GkvxWsaAXzeBrRarmPJgq
XXl3UHG7WeAAsduT9sC56rhMz3BcyDm8uq6iAXR0pPElfSWOJzJO+DDfg7hC8WNqQ2kp1+JylTAP
onQEBkevD7mi27/qps+DbnJKxbzPHGXfEH3v4ciPCkSla5ZPmjgytAMpebqdtD6OwAh1sY+nWIH8
/Do//uCoVeGN7v2qD8hH0YXlwutfaxr9gbWdiztVzBAZfm/HvRRMExHgrXW2BRKpdVq05cdQa4UM
UwD898/RAdlWEpg9+G9nsMGJI2aZ09OonWzwAm2mWO2NdVsPNmtpRb5RcpTyHg++F9kRuXdRBzrw
ZFJLWS/1zwyliZIQUrzBFXQ+kGdO4CNQoK1Rj9YbGzWU2tLkSMjsSfaXBgoJYnF27ymswVMArJik
B1hhU1s+bv77Vcte/fzl0k6OAekkHrQSk74QRNqFUGkpL70K0oE1foKtHgOc6UZ1SYiAQ80Vq4Qo
N1NaY6j9Yvyh5+rjscdouw+CW4fospmbcc7Len1UZ1tn2DIcDi25irQgx5U2vgU7fVpT3pN8mHK0
MMByvREoXOtYJI5F4AQIfymLuXza339CSpVqsHvNw8IwOnZOIH9/mxywbP3nUAtBwAC+VmfjoZCv
ZQvqV0g7Ujv8SpJ5RU7DDrKduLy53L9j6dhBfQpcwKx528VyfUFKVpgEuOkPbSKYKDnOOSfTPhxw
IDbxcf+ZkTy7nTf66lporwrQf2fa4M9TeQtKULOdZvrvtOO8oNFs7uAP6ST9AicwQppFSn7Bejdx
3LCU+Jq+vIOqfpX09bNU+IzYWP3NdTQZNO3D13GVHbTrmNBmS70p2EyIDtvRhuV04FFvghc+gcMt
W386gDcHxHUaI4A144oObdP+YrnfDJeZLuqzsIY/3IG+OOPpEAnOhA5iGMnbKcmBt7iOIU6a03u0
TlLNVJ2oJlzaSRAueVYpQaljrNCNcVg5kgS+Fo0vpskCgtxP5ypj/kzK12Z208E9JW9x8eb8yFo8
xggDIYYv6bnsOFxMqFaTndhjBysMIAjRLu3nqGCRQiKi7LGxXNHVwa9PRLJxSO0Uu1jqQOf0tyBy
xtj6jEZSbAdR1g3nakdS/g54m+co8o+U0blQ6rXh8xKEmKY8EBlfFJiDibDJ8nwaLEUIH4PUxrkT
9ocGyWX59FR02dhmdhNIJ7m697GUootbzb7YJJ519eCW4KKL8e8dInxBhu/nMFIUu3tgA47k3TVP
gL32pWUKmq10r80Dq/6s/mT6gR1YxMdISIIq9PP6cbS1I0h5/cKQyhOy+g2pVgqCZg+INlesueqD
iyFe961PHBecgmnBYm2jtAowkt40tKjEjjI4kFJqMMbq8dMT6bFyCnCqCCZuZQTIMpIkmZ8MmtKD
TI9GUb+vqLCpH7Jp1ogzD+ZLO2zpQpQ/ZkjMa/OMdhp/dUb5+S10mltqRw1La1ScZcYGXmp8XlNF
7anQoewy0batqr+C1JCo8tjMUaXqExA/NM9BJyWju/99BMAkBi6qJjDcGhGx+IDfHiS1McekANKv
/vXHg4/AeuqdjQw/vAtwHo0k7NszQIY5YAQSv6GKnL902ygICWLQo0nOe692+R6ZO09BndhifxI8
pOgXANdgZW8K//8vKGUOADYxkHvGvQ7YEWMQUUDEQeoGZzO1ZchhTiFQOr7bM4TgWiqeg1aPLtos
QZXj1Jiny1KHZ90L1n3eax3vV1xwbXHQS/KQt/DEa7/+v4BBFfPx9gIZyOOw1XtBjdDsu/y97dvc
GbhwY5puhZCNeydSV2MVNEztMUc3QMWdnzJmMq8XbDmJPpEQPVWbQkOo9fAzJHULs1tMBeOQNabe
7sJDAPAWSiulaQLKEN1dzAmEyGwIyIumPXQS2NQusyDklr6DKMPF/wcCr03eXlkMAaTW6IRcjuhW
xOHiG1ptVGOCYVDD2+cHSH5B/mrBoMgLHxqhzgUqN3WTiUHZ7z0hdRdIoTcgRh9RGjoefEZa9ZPF
X81FStCV2kNzy2vwEATOEvoCSy40jjdhlm7BnSbVbvs3MCB8rIH6APeOCUh131jny2RnIrRBvHV4
OU0mt98W1AtxC9kZg0fFTDuxqF+nuG4PyHFoUqe3THfBt2o3WZSJ4RFCvviuSabEQIahacXrpqO1
3Z5IaKyzERwNUDP1sJH5C23sO4Zt8eAQAQgUZoRRlykFCl0TI/EZSbstcl9qWHieIeViYNZbwsM4
VzjaIb0EJP5YKfGR/hTID4/DX4Z31JUCWW41vQb1qqyz0/C9flS46w3syrydj538gByUZfg508u/
WzTUyFJKT+AtI/q8fHfmSQhIQ56TZt6fXs8xstZgTnrsbkaxKK4X/noMIE15PSZrbORy4tbC2NAV
ctI4vtMj6c4Ig5Oju9fXqdEutH6KJYa7dMMsnBLRNdoXKA2SDYqdsR+UfoaehzvQjGAmoA/u/44c
wZNWz2ICwbVOiE+B14VNa0lgoZMwad8Q2fAha8VBlvBgGsjHvJcgY1QDG2/B6PO0Fo2or3DMJJv6
hXt3C0j+MY4budrMmDzIzp0RshjQ8/49XNN4rdDMkBFL49EJT1Ru3kfbskkQCeMpzqfTXEVZB9Mk
qA3Bgh70efnkAOI6HrYTm1ClVh4VeM598x40FPpvZSJ/jjMgcPXzMobBNHdsqiXhxijdOOYGsKLP
3ovb2cjEP0dRGUsqU3VlrABvQpEghDr4i00FBzShrSsThL0Gi0jlWL4Q3ptXpHIdxF9IdyZFfY9n
x0inogbxXY/NMmGdsHiHWv9vIi/ABSA6Wwy0CHeN08Xlody4QRL2xiOJCFvILgJylvWfgx8PYNtP
ZniK3xF1cSLAdRr/juWqz76QJvrpKLH1TKFhfLuk1f0btm0cF4TpA3nbAmoVuFOO5CwvsQaRkuQW
0JhpoWJYKFVecz+l4ccJqs8CdWjVTvKeeracFft6D6B97UnJGpa83R2PyBUarVpgO5Gi84zOHlYR
Hgm6wtLCSUHywW1s6zJYs9U/rsqyttgsrHGm3NSiurqK6JjwWarwIsl80TZAAAe3v4H14E6cUYqD
r/AlyB722AxNrk3zIfpB/TJHAbXf+MiPS+gGoLr01ceB2VP2w+UT9FD+dpcrjg5BgEJr0+By1d+N
KsrNUne3wgQPQpVLW5bw8ncv8MpR9kHascMEgZp7yP+YzFT/IgYxGOmDCdzjZp2oS7sK6Lz+hAxs
0KA38lG+qQqSwI0ty/m+OA2Hvr7vshn+BV03/ivB2T4HNg0NE8IAClheyxqPUNRJisJaQf/Evd7C
ZL+zYDTdlI9GMEMjVjm3o1KB5RhoZ6UVtwsuNVR1m+adJll9BOjfXfduqbG+CajY3IjT6WzXDHXA
vP7yVGqHSq4DKAmpDG/I7Fq9H00fOBdOli0mllDB+m/E6jLwnJPdqT8WaM38rhytHBzL/G5Nr6zG
hrUtJTmQw0dfawpwaJPvCOWn0Mq21Nd288YURZ8HgMhcTUF5nxr/vMZ/hEhytUatOgTSKAVR4ldt
F8HWNo0EzcxQ/Gy5BrfkbHjcfl0F6MmsKu6iQ0VcpFTbB7j+Y/Ep4Lo6UlfmiKtyLuWW8yQvJ3Me
nMFmZ4OVi8GDO3xIOBKkANPnbCgOahqV3EB7dn2tHdteiOuOZeWHXZ6WyfAgqSBsKjFAmAz5pBjb
o74e2LNiOCh24by+2WiuJQome4uVpDjzkWrPPNFXcE5KdMCiwdriVnJoO/loEhVoywRwT7RY5/+4
BpPDQEBetUAIMpxSIirj6b1DC18PusR+JGXjwy07LVB7SBFMrRVcn/vXH+5vAxVQ8ftlouZSaYYl
mKDjFj23/2toitrOYgk6AKuesF8+tJNqdKuZ2nzWxm0PUv1P9515eRTrKi/CREOTqvsjujRvE45h
RrGGjvf656JxkcNWeqhsIg5n0UyvnRU9geDZs/j9en5DJDTlvsMwcH85zy+8EcycGx56VxYw59Q/
ZPhatwSYkvJOOM07b11kqHXSiwEIh3R60ISoHS4E+0coxE8lCU0wdctEUp5FgXrQkJcOZgwyHO/O
4kTEiuZnF/73avqoia1vlCTR11M7L4OTNzCdOijA1d4wvu5UYqaWAutkT0Rc/7i/sWN591E3D+L4
DLwm3rgh67CRY+R02A5JB2s00tvpiLULBGRCKtsn9LVPBTaytL0xOCSajmTJPO7d3Koz44+osFOB
KmsWmYn8MXXmIS69jW5mkvTTwMR8dVy40IyNmV5VL56rRGXNNLJbI6XgXMrPhvkX2SFmpfJyVs98
+JMsBo5YeXSFrNy6zvQ7sgy1xN9TeHf2tSzGrBNlkgWKhFto7BorHoQJRYqydaR2/7Kq3j7yMfB+
EJc0ovK3ssEqrduFFGeTPE617xmhLZNQAPMEoXzVfTnLwsQVeZz4ukQPTcHEPVz4IWqknSjJWfup
MMy7vSV4TtXqRQRfzMxKyAjUJnoYFF2b6Fi+8c8KY7bZNJ3aI68WakXKg01Ft+gi4qfTDfIV9V7o
SQMdrCsTI8FrOHQm5WpGy3WPXk8wNuBfqLjyufdv4t/ikuVrvWNokNMRYmt8MvNLX9dO/J5Aiwxd
nBgzNRQ80NRjm4Db2yOmeR6xqUVxvHzvd1Z30sQHbkPmGnym7HQAmqD+6u4q/VUjpZqcB0OAoEEK
Sa0Jf6EMhkuBziDqiFR9BxAPnH/tYTBrsWdiFvpgpcM62extDLA0L/Hhlz5iyCA1hH0+7wJQUYj9
cvtEPJs2lZ2Tu2rufFkvdehpN7vNyiWnN1EkPKsWik6neVIimh58mhtcD1wokVtSe2qypBwFyYvX
Sg6WOFzEYl2IPfCbA93TaFJUmhL6DVOIIDkQH50qjmvQRFQ28HFp0y1mQ/BThaseRnqeKSNoOc6H
mWwobzVng2t1XnQePtKd/mMt7ONGCvAzY6IAd1yRWbnd8eoGNF5w+uNrXpghzqrZJXdX/gintZPd
eQe5ZBwDU2cv5T3djjj+qLtRn9V/YTd2Rnw76/g56WiiD99xPnbsJY7YJcm9zuN/Nm9syghUlH3Y
kFm26+Q3h/ds5AJN6VL83loVYasqNh9TyxEbLYzQGkb1hVPGXKH1VCmKZLj9pDLUdqy0Bc4xKFEF
9vOsaD7mI20vqmgJsdkKDFpf/581/Nyiuq3dkDxpJyrjXz7VnkM1GU467+CnokRVQlj4sMqHZFeZ
Kz+v2GlZEkTnZMe9KVbow0PKWWHmN+b+Rh1j1aoBkYgUUI7RVXLhmUIJQZ5f97yg5NDDyywLtS/R
bGkW/Ebi3zNDJ20272WeBw068CPtZ557+1OW6kHuO9CmKq3fo7hSP0HdfMrm82jLZtE1drPGTPdj
bv7fpkiRZlyQGQwmBDB+qtkcuj0fp4WAknb6vaaBf5wG4lr1BACTTm5zoWDtfbgbdQT81WvWUh+Y
tSvoa09Z9NuJaKGgnPuZ5z+Kq7bFeAVWzCEec/eyr3pKQXyw2xK1MeeQ736UDM/TZKKwILRUCFym
FB9DEasEjfpL2/rYeiKmWlsQnXP3y8TLPo+//p5kHFmM4j2w4C5Gkgwf4QELLlrqwvzEpOE4JTlC
nJN7cIoTTuddDVPUV0G0pOTToz+PiRDrAJ9UElhsuGblOj+ByBtl3EzSuPGKnCiODuwq3f36C30l
vmofvL+APtR37Idqk8MlKCk81dszJCGNM++WUTmZ/CzAgEgs1xiEJUJBRl6tNHXs1vijRddOo390
Hx+hUqwOBTgSmZa3P5VTtSf7cIW/4uh5a0wA371/h3j5ZRH1AqP6q9CsHFT6IyEPyBaUN888upbl
RqhFv446q+kC4wfscfcio6sbSmOnhkQtG6sDMOf/9ZN5jIy3XDU0rSqbZnfKYoOjF+iD4WO6Iu/w
sMPZc0da5DSTeF3K4VPgF581qhwLURSaqi79M6XyoU57xYShjGjvlgeoerbNWdm3bUH27fHUhwjj
wA0s65zzf5VdeReO26oVsIeCNtQqEpG4bWcr67N27HWav3vPnCr2suwKwVxZsUG98U7+ygY+l83n
k71RE1yCCLte5VrW6TAVe6P6Jnzq8+wYch70BsPYPvSUs0PIILICHeHs9I3iYgS7kk1rp2grmDdI
nzkHt4/akr8ZzRPattNJ9ErDwI9AQ6WHKZ1Aci5RhiCpoywItE+uLp8PyjuHeT6Esn9hqYw3UZu9
AjmpWL/tt3IsiLoSjqfM6v2Dwu8BrZ7lVxCWmVWuf+VWfLOktZ0DVSb45TIP36U0ZDpyYoSnLbZ3
uGI8v/6jg1AR+3NJLSv7RUK2kYMWIt1wN9pcRjcIiGTIU0+oYFtCOBkwCWJdBLPKMQvs+8g7Uxoq
g6DaU1MQbccmpeEYdqtC5t27iebr9tH+2DxMS2oALL+JKgspvW4YrcVEf6cHHM5OA7BKbHWZowuP
9pfBpQsAKTl1FkHTL+DNtP/pnY+sXjOw3u4EPjNBZv0/DWCE3+wI+qpbTta88LmV96KHuF+nI+Jb
RufAWMPwBjt8tWjqrwdYPSqePfA2YnUHE3IzXpFDuXjAplMFLs0BXRaR+ItFx6rvHEmlPOP/Ryll
1EfPxYcj21UF+FvePSrF+4VkkoSyGggIClhasAfPUHiWRWAsLxyJx/Lrzm/bRYbVDyaYFhuyReII
6+EcNQPjdVS605SJJwk2CvKzghv3l8IfUKrcEDPXo/fvGw9ci3FeegNgHP7qKeiQBf/csssiW/xf
3xgcADOShUp+SfIKfRDxTLomGHbqEB6UawHAF6/n8digkXO7sap8o29fAH7h5OZuib0TURPucdcL
tSuz9ob2jYYt+bd4Msqex4IoG9lvHpNfHS1fdusi84nQTBphydlvMDoddl7GxVvPxA/1Sj6sRdCs
wD99m1sZ6pV33eSUXL0VVzFUplmefRfu++kZhfVAW9aLQMqcSFN6wePKunccWsodPk3YiI29gFYg
TZBZG52ZLO3IOdBerJxuR9N1f//7IanW74q+5Ce0Ot78fsSz9IPext4mHayhv4xNiog4d0zA5XTZ
gC10xK+aCV7OOyEIT/THF9ykfoxy0SutE+OLTw57Y5ASQ7c4XenAWAh0DmGIaMZjWLrNlsN3/YmD
8mkPiDHEFrkTGCHzFG2dNZVtDbP6osVy8Z2Z+IC67TY5OBBCGBH3jLoo9FXyd/e7uB5FDi0J9QCq
MFralSRB1NpvC9h7iv+Q9YdSLUcwVCkcaXcbnhivaiiC5KnMLwdJPCibdRgRqhxbtvoOjKhc3kkF
l2fueEhbiuMLLQV7c+dBAgYIb0MMYjqHhEsCnESNd/8l0EwoF+EgwC9P6nwss/nx4te8fFr+I2zX
5jNjllNE56tCR1T2x1+C6YHIIWVfSBNNVmiZgYBi+yufSBJmfpW70jNTxELYmx0MXpQyQdMNvm8T
aoHVRQh+1xo+UC7tdLoTjoqn0l9MCgCeW2/PgcFJr2wzrcceWAhNEMeURZnHLiLRZDd4QTXV4WPw
gb5JcxVat/1FOFtAQeIiv2WF5hnZDyfXH1XzJaRVBdMFB085+z0ejDRCCWiT3qN7lPvp0I1s5z5e
ZI4cCEMgDgIdTizvGuru8ThnxM7k7NEdhF99MNWP94mjtAQVwEcVxG5Be2Ug8nhUp3vS78+YX4I3
3fQLtxh7EG5RFfJFNM7yd4ZHcZgckzvdEzIGkhOXS0a8u7KJZpYqHy45mgdP5VA7/CnVrk5vWEHV
0k9vdo9wQFiNIyval84LQGpFh15Q+OGHV5bMGgQZKIbspEMacnJYH/Kdj/xgVXILT6rjke1Q3sUO
KM+whYmfCCAtm9vSPpfQqUX/pB+0VVKOq4dl51sB7Uf1xwvBRZ4TNZ72FPGQhS82LBulSY9ZCsel
pPlD4nIWqlJL9zYw4M8hzIJiUCOVdVCpuZKFlOWgxfe+gKJK65MWNmHrdvxGnBbxZ5R8s+hU/erM
SzkB1t4E1LP1+Ori0uhZXwm9cz9iL9lDymQA8gTzJoAVwKo+wVSNAGwgw2+caBPjfQev6qHnwBjf
liHliYRjk0Wei7B2gE0J2zK81uv8aRzIfiVdxaRKggkfJjm0vmi/FvskO57alpaz1B0RdwsWEdy0
jU6n2IkY3Ex9tUQsYKbOyGzS7PuhJUsHGnnbl0cnQv5Bqk60C5VFZweLs6eZumv1+bTD2SDbwTpC
8KjM+UtKUsJTDe+OqkVBCtyERemDGpiuTVXZ/1XmrpkC7XoM8ZMvfdi9CMQtnXuqgjLLzsx5xHSx
5MUy+MJdki6lNf8WcDSztorbz1FTPSByfJs6/oG1v6Hlg1DG62Ihv7iJIeTybr+ApIKDPF9gfKoL
mijNru0uNdGgwOnq98gAjuxOtna5Q1BURpSS6uSJK2ACFuuxGRCObS8W4N3TRBTy03t7YRSqBbTg
pr3NuLQwOMGROC1ExVP2ctv9tje1rAP3wHwkQrtQN3mR3HPX5VzeCXms3AJmaZD8y2y9y0smwiIn
+l6GhyiQLrYeIhbULOhRoRJDubqsiaKNMCVSWdRF0LIptpRd5oRbLVR6euuiq+cOotBklRlXqufU
4LtfUSWQ5TiOy+vYKft/vfd/5GuTHG5nX5WVUR0K4kLepULZJm06unX91/ulHkqngH4JtehI50H8
zIfX8BG66o2U/bkd1owoqiy4A6th9+SfibjKLy6JzphsaSaXDgEXXECLA+t7DVeZMq30Hc57oe2v
oYqxFnOCYMTfukJxK19GqI/wN1LjYGKeeLWcxUsLrJMNvNYX3zss42aMft2ej0V0yKZlcZVdOSfm
dT4eV6gURh21Vd+nAm2ji5NNDAkQAPaiVKV0Bt9eef2/atjOAX0X/JCRxL5OthwGfdNisB96XmC3
U5+LFQzq57CriOZ1KNzpGGAdmGxY+el6VcyasnFr1R1k2unT+Wf09Dw4seUvMNMjRhcba6ooQBrt
DyREErL1+naJ+wavcl/13cz7BVL+OfoOswoKpST2Duhaavgu32y7CAeXfVNUROn25bw8fmDmmafe
HiDRR3PtkDllU8W9EId9lCSRGQcBBjlxcQPICmj10xP97VNRCvTu8CEV9yRg/Vha+93I0WTiUoj3
nUrHqCWM9orJa1CJNE0wZlOQOseIYadJHCzV5sN7aHXfJeF551nlSWpxtT20rDi0X9romat3pNSf
HOPbthG3dqAtaoh9r9RJPZOVtWpoAue7Be8ral3r/p1c+XNwO2JUZVXkAufhkzlxm4Q6iHsnP9MR
Zi+9RKQG8f6X3u9XMGLRvpYQ6RDHZT0yPzyOMqdcco6vV30f82TrhcLqkODoe2/bG8qgkIVUBeJC
Ril2yYOnL2RP5fV4HjHbbQEaXk8ZRN+XTPHGnDvjWRNylmFGxqIpP5epPvsru7yt/uyLoP3ml/6t
FH7ir+5rmsf1kjDQZPfEhkCPOwPvar0+xU1sEOP2JIFj8cqFJ0OgrIraq99l1bk2kCwZdpc3zmIt
EisiJnP39p2kZLdKVHckBaiWmUzbdsO2VsRs4m6DAB3/oY62a3N2V0cNlQvC5SX5zSp8MLARH5/7
a6emlN9wNcEhg5iDvr6nDRxKarZ14xI7GrWNdcsc9rNt/cKhdbp4Ik1/pPEfdEWKX5SwAx37dI0i
GaWllLEMaGe2/fF+PHwvzok8aPmwLHckTZ7TlBBpmxMaJ8rBJlz39fzEnJRMOCXKXJ/RbLAVP6gj
tBUwDKeUVLDHovugCDTIXCxZXJ0soJQypXRpU5EHWED0LrV9wW0YqnZ77l/Pauf/dMq2jG2Nk3jS
aOmWsLXAPYo8WS+rEJaLDahFO/nlR5G2W/psH7rW4tOpu0+iukD14k6KyhivZtCpzLajjKZ3GOJZ
U5XITAL433MCogK2KnEwMmPdIKMaEN9c8Wsd2Q9785uOZItr3S9J/5JlRhn8Z/9QyFHR5qJeLco3
nzSFiU5eMVGVnJDolH2OvWMKUYsisp5FwkQuzK5UP9Y3/U8ZyZBcmxHTOEBJJFTa+VtXNFpvcAxR
na5iivNbCzoeJx4OWqnyZafZr24SpDMw/Kdzb4DeEaBJkD8cB4lyVx0hXFyx1AW9+QDcz+xSAPmw
UDuYlsc8xKkahzAOe5emFEK5FB7ickwTveoFpe9Ap0NpvIlxc8CpOjAMJwvTs+xYglnP/xGtQlwK
ybUbeNmPb7YvGpEIh42zNNgFl7o3PDX206JzOFMfLG2ASVGRj3vS8cy9lC3VqkgMA0d8okb394Ou
T353TDjO1gTHWCzEJgt59KdybGReVQYa+/EYSfZSfl7Co3zRXRFkeOfoo9GdzEkalfO+0tXM/cXt
c/g80ce2FAk8vECHZFQnYQVLCq8kSBz7MGzIR48NuVQeNNRvPm++Pv2ds1pOB6uYoIS7cy8mZoGR
GLLhK3pgOIYLimndNF24hscEL7mhqkIvghxA2oF8hmRX61TOca9/o/NBdkG99NofK8jZBEseFE0/
DeAnDWd5TDMJPgdnYyR6bSvtB3vKLcgVzoJzPcYNsITyNjJsdVMDN7lo0Lq3aSxAGUbtu0Q6ZGQM
b7kfgwbaBaax4G1Lja5dllAXU5JPV1qCMu4bL5hWd0FgjpsVDEBsWp2NtD1wJBULkz2SluXmgF3k
452GM+Nadj/PP1F+iPHAxITJpsSyLdJQEtvwHSimUhniDe/urG4ALGKuWKm/EgIN7+3WmPkse6ai
PxetTzH4G/tqv0sUcgSyFpCW8E5RUjTa6+B3/7LSPXgxykaXZeAhTtBvFR07ysmWQDKGQfhtzN0Y
1TjfGJD5Kb3LLcOuboVwkkjZpsDgLVblAZ2/+74Kpong8fWkefOiOvs0CF/YcdeO7E3CWJ+uEc8b
s81KfNRCypDgiptRMlowmiYDAvRhYh+vamTgqRz6pz2aFFREromIZEs9AbHOQP/aulLTKgy5+5mY
9ryBfSOTq9iKoP68RpCl44JBn9AM2Xj2CIkZUfk1wkyVEpOPRwEotJkLsLycNsXTMqxEuqLADNb8
g9H+LD6nzTLwaF3MZH1q9YCTb5HnIy6MjQoeRJzCVN993xR20BpCo/wE4wAj4PfgpKYSOn5kZGro
Fe0uvK+7M43cPytYvqFDJk1DfNL7V6qrne1KfuASZhbvw/DL4OF41jwNBOsquXy1/6+8eYpHGlNx
2ZdG75SZrCt7bXdljm3WWkzfLXbRDGC2ECjFEMNe42+MYlTI0CUayXjGd4rBwFYVfGMH/k+Vq/x9
KSVDltJbsXc851kSlsvo9kDW1avjDg9BAn8mCJiN9I8cvVqM7MHAkkRdkTkiysGZ4zREisAouKBn
uoDUHQn2GMycu7F5DNBStoeTWJZhu6UOCg/X1JjHq9ldNHUf9Kw3p/SYxcpKgIIZ93MnPBHyJsV0
HIbntPwNF1crBfQ+A3m8k5/Mt4rlhUX+KfHJ+ahtaNbPbO081iQUo3WKCh7tceuN63QY3Nz/rvUF
Lkkoh1X1kjzCTCcjpchByhntpI5U/D/lpFyiWvoowajKTGtIMCssLTEZ/RL9DrigOowUeRLCirYH
rvG5mgA5aUqzXLIFgFWBrJ01nH5/WrcVCsi86NmBMVagoNhQ+Z49BJVb1ASKN1EdtVjr4ln1Jd1+
3fRyi+M4oQubfZk4ITtZmno18NlUKSy/LEPBGbJk91IzMnqS892DaRRMyZ75yY3XfSjDQ8C99Xbe
ZyAeiOJlfmQ4uJHxmZW4kGKJ5IzEOlq+OwOXX+dVawzHBi/rw56Pjv1eB+ZbPYxprV38UX2r3Uc+
u8o6SjBKOw+FsoeCx71LUikC8As2cwpDs2Xomp711TRcSPv6kgW0bgp5/D9Ht7dbQziO2jHMHXW5
v9yeYyasWIzqcHoJh2aUSLtkPvuab5JVJ+4vFPcsYlo0D6cATY613yYgJk3jdcxCeR6UZGrS96BO
VoJM+CQ4dr44nNyLYMD7Mv4+s8Xf3WIArmg9psofVTSBkA3aWJFkkbd2SgapYCfPGIIuW+lNdrdl
1xAMGrnrWSEWVFxm4WXcY3QGwotymmY8vufRuTVcL3sgh/8EugwYskpyQbWi9s94yOLPHZVf2ONF
tGjfRI86DrTAQuNVIWq3EgPHPgeHZ3zE8g7qB8nTwU7zSbTSSE5cODBpPr1j2bPFRcxurQP/tt81
UTgl/qFNC0SztAoTbxUZVriu//dWOztldjAcAkkB1S0vyR970DQlu6u5fFLfXKjoS4vB+V//vJIZ
R9yYq/L/EtExJtas3/zr/3oIwd3DUIghu69hIudG/78MZJH01Og62uvCQYWAb1aqwRQHYdVZ/bEL
XwuC3ihYXJJGCf+249IvdJzh9rmSgA93DsRKB5FsBza2zVxHjOupjFYl/zajmf29/LZhDEwjw2OE
pwpEFEHAyw1aN1uOYdJDJOv/iuQEDX14W7sxdf0hVYaxrOpN/7YJSsdTe4S9Yf/pM/BQlKkoic7c
4HdlQ6GZ6Tb3Eznm696StzmxTbFx0tiviWVAb5lWKE/oBKoURE1PD3IT0gzClGQwbQb25oEHR02W
H08DmsoIZ+Ni8UhSQ/UXdCzK/pzrim5Ahe7oLPFbDjhZ+L43A/ym8itESuKlXMNTLDL3K6+0wnm7
I+gTh7iBhEoCf8wG2ocTuT5YkDma6k2OLcbLdPf1VA84B4mAvmL6ilHKw5aPVgXT80ONbzxAlK8Z
YddL1pICfme/b5LKv3P5CByjttVPyEAqW337C7U0T3dmnHNS8XWxdNOJaR796c8UB66jTqt1Hl0Y
IvciUxNOn91EkxF7M3s/TSITbcao2/zSYpbcdY8aRMtRg8i6+6uL7ZZnBrIHTIoDJg7xli/0uZwC
jqHUaaSJm7TlowxdPKGmg1JTaoI73aBhHSbUxLttNKYvnES5bqWWfPsTX5QWjv4DLNAE972+QzJq
lwxlyq4yIRZzxZC8Xx6KbRAJRKNiILRHDmmPoHlFK+w2EEAnzGoPpEWiaAbLK6dKhmsQ+3dM9VcQ
ianPrHh4nGDRXchfVUDC6aPFWD4y5EZmQ5hcJJlCGsNLdIi1D8l9lieyjy9jb6tgE/I+VoIzj1VA
op3BcBHxVv5eNy/8FjV4WZMLCWRSJ91GjeD5Jw9yHw9W95z3Fau2qy2b4uvgvsvPYf538zDMIbwT
0XJpT+b1uusiyeDasPPr+Bchr5RAtDIix9PVOX9XEjZFVhwB6IUEwKaEuEsy7PenZ3S/Cpl/Yba0
w1HYBWxAQzLycphAayhOSro0Ze0d8xvZbti1RIDYn5nhjMPzpAFbUWcw7NBCuZ1xLWKjhRrjaw7z
WocbSDhp5dbj1GppJtSI7rkEbQCheGHcppPKyIsuZsy8wY3EJ+kbuorAm8MSSECLl2XUZdjmUcwn
LcndcCyZ6Pwz+CUIq/O6FW74Qi6KOnqlLByNNn7zif0cya9t7zgl9pTTUsz0rieqeiGebC9a6ada
+uQ0pi6RXFyIIHiz1GMcQatozD+xa7l7fRujznulq4gW5pBCcd8aTbLrHJpQ3Ufj7xuWfrMuu4/E
DhyioCKNrcDPDACqMRy/Q/tqG4D+cmd1zacm6xXKHG8lSTVngbwww9DpdK4X1ck7EnX+8gI4Qpsa
XvlKuIZ4gBjUA1aFrRI2ry2BN1oWcglwZL3cxdfFcyvR4i4fEXHTvY9VH0OXI91ZTkuPD2cLUCjK
IjA8H05gl5AlLrl/nJQP6Ml7hqnzVKQP7WUXlZ2px/HyXS9GIB2GzxAox0xoKobkw4w9Jrn1FVo+
DBVrWjCXVPQbdU2wJ5q2zpFtrVPH02gaxUoLxcPElQw36+H0OFlEeC0E8htFix7p2sMtu2ai6UNx
ym1UEMHk03VVp4B4IYXAAlD4bmAdxA9ovp08B7kLILR5g3fQtEEbfS5c74c3OeZs7C81hbAfZhH1
RtfCOoV0oQpVJo9IH94J7puLr+rkL9AOxSV7HG+XCyg1tpc+E3PkXxH8BGwJk1ZZTmYAivvPZUZj
DBUGIjkHHsBBge+rmKjB8p6yauGwa8f+yBAcM8vEq2Fyh0hR6Abif7NbiBTXtR0ZNSZGKvWtOAWQ
ZGv8TIMTvryxd4LmP9pSygDx4JoNUECZfEmcPkkzDMLu54J2jRir46IGmOfv1HOFHvjKvgErt8rf
tOR7CMn89SeiSoOZ/knCMkV7NFMLwQZ90gJWEClhuV0stdKwlsnzgcNG4p2cBrNBwjga+vBkGkx0
IQM+cwZLmj3rbIlQHwYvS+JsX6uvv6dnf5d+241ZaUrs7gm2i29kPmQsTDbrHbkQKVVkuWooaVCe
NaQVY09smieh3LsirFxXnUAU/A7oV5p9UaRk9erFsCThJ2VMbxTHfmOov4ACWoA43rVFS8Yw1bv6
HEX+7Yn6xw5Oc9hPV5HyTGDCVz14d7fOEhxVlg6Mh4v/34CuZez20umsf0aAMeNjNb7OOd0lNVsE
X+B1XkVk/zbDKq6FOlCAchHUM74hADK7a75KsKjdrGspDmow/JixhUTkeI5nLbLVW0JSpr2zr2OT
alWgu2GnlujTy+JZZEwWSdadNIGF0Z2f7YNxOtI0eiwDpxsAdJsbxBYZh+Wu8o8DRZFCLpclXbZ3
PkITrKUsKaujJpHzsIzRp6xUJ32AQQ4REVZmYp+PjVSsvhiNn3vyDvWHAjMWDtcqCc8dF049o0hd
Zq1hhGgLhRcf6WIpk5c/6nsUl0OztAhDEnJk4i6cabTV8+EeIRr9OMZt6C+zt62gCK17Ns7ny9qE
P9vJ9ld1LPfuam/lsdyHjYNx8cmXkGT9lhT7u6t4bnfS46hbejI0wm1CTaEyQxztqL/KMyOxPyox
GMMGJCwQAWx3csYttb+JMccMmPdUWUdYAhAIxDYJSLiFq/9YtI+YvZRFi7a62I/VX4qH6Lq1fwqV
6IQ/XbNKx+vCLGxtJMvyvNI3aPVaG49l8OS69wB5fqiN1VMzaGjRIHgCeLXdPA90VnrhVrsgVQ2z
3QfVrvhEPOY0OHTBRFlrhq6VeUrLrBBaUlTo10acqMNQ9SdmwGdov+P4hAsVWofCELq1Cda3ojJ0
wF3cIdHDqhW1tzGObb56cXk05OVIWg6HEwT/aXVkS+JDglU5bTYyyAjlLzw2rvK48Na1z8CS0Bvt
eWFHcQwcCbB7TSTmKWwevkD/JBZaGXdGgJXwnVfpZvxAXaFYh8Iu6W02yXZHQbEKP9HKZjf67AB+
2OExqqSVs0pQMnLu0JkCH4d3Ge8jdZui5a9KYTKw5Cgl0tpcTmxCK5dGoiiFan/IZCRZH3VgvXXT
8sGoab8iNVQJhrdzGaNop+zROUGaFM0Fe3AQxlwDJAJyd2vxJFj8RPuk1y/QXFdwrQ5DqVw4piIb
Ll1ay/p8NMV8kL5BhEdV8RDNm3wZhU/XDR9Dpf4gSy1zwjZVoAJ63TUg1QaNxayBFWePD02QA+uE
9T7w1LOeqI4kM7hU7/EHnMKKfsnpW+fmk6V1QOlJf4pq3im5EMx5hkuc9CV0L0r/BhLBEN3uDhgs
tUze61DOmkTLbMqWBhoDeIS5U0xaWL6vuu3ulPP0ZXCqE3aXdWq1qu/MnzPOcie9w2mgW0xSqU0m
x9HlDG+H4es1MAvS3TnJZaQYdFkhCK8lUDec3OiHFp1UgY6vwHMD2LEYfItG9Bsc5+Lm19h0t+o6
q5SI+m5s5/ow5sxU8VcmcuaxDUTnj9ebcU0A56Q2LiSV82MUsyTxwKF24tVkf8oIBQY5diQZV6Wf
yOPXhwTHeAtqNhkJZ9fVTJG4dGj5Eu+OmwtL3eSRgfQ2BDJHXx//oiUL7iqlDvmc9f8Ml/tzPlVK
oPI37NWQPFpXjTVje05a10wgcSCZdL6girNnr4uNrSEYQ9RbAzmsLetoC7Lmu2UbxLu8XquXMs51
KAmgNDyWF/ObMDFnog2UgIZbv9aLnysHudv9vRtj/arBecHN//Glntk1GMDUSwQHCBhWcFCQn9sW
/ZPUM0HbN0N7crKqjoqaUpTficrOZAIwUOmwVVdOuHaUqmfsElSPuBYKOOE2ucyOXz5Cxql2y8lB
khVjsqVJe+PfA2aDPKnC7/ADoC4podE+Llh2B3ylwUXdWkOr4c8BwmomRRa0mGKADbjdY9pHLCPS
IIjMgNUwFUqXUuiPivakOze/kidnDlC/RYgTFmJdLQBhbj+oQNWJRZXbWCEm7DIe0RihjB/7dpYY
DQacZa0BDyQtOutUNf5BrpHpX2vl0de0FyPOPRabmOWfXyGasnfIGUZzkYG68DOwoXi6taQW4w2h
igXtAdDLAgo98vctM498ajr4EWctvzOdIO3MKTmis/+oCI2HNB4Qy2pZGWpwKDZvJYcrqzDCbkpo
tvr7LGmXuqS8BCXNcr8SEFb5Gl5RmVI+/HVkxdbCDcTUOZz0UV5IluEaw+H6kau4JU7VwV8oiO0X
exL8HTsZu/byZVbR4qlnpry1AJUadoA4lROatskYJIrsHxEMcAXOc5iKo+YQlIHpJHsJZNuO5iqh
xzRkuPpIadvfs5Y+M4DudgcwCMmSQr0eBsCpYrWzD0uXuNu+C+ZwOChVdr8CBapt/BuzyBxGaGAE
v9Yn4FOeKha1nGfc2rAfeAV+Hq6zTMjDriLewlLLanKymy8WpqYbsixlHFtAznoLqjc9jXrFTXBm
68sPXUT5aJ/2lF0YcJrL+glzl9UPeUXVqZ2dYVKHRprl4Cp+1npfRc77lDLj6w/M7d8qMKv2S/xv
Gy3aqn6WYZcY9FGgnSRjFcMawkG1LfJBsAFZchMsFSeaGbkVdP8jl/jTxW3J6kNxw+KT9lBtAwE3
Jde5SrXYZF1qnr8OIVHKGWc4kQXX1tcfv2KXx1vofHe/Io0taatGUoG9e9V0iU7+F1SGDe4X3mb4
gOxBRQEl7oSlgvXS2GUXwvrUziuDSGWLUMcCG7QFmAQKSELw/madYr1lFhtpnK73AVKZhCnRBQrb
VM3y6d8byu5QjTlOTGiHHRyXeYhKQ37uazk5CUDpOk10+0Ilhac2jH/NEFnfid64Sd6J9a/bDc4Y
WXfTcwm9gZ0nTHKkBpqyXBStFio47OesfkbcexuBcYY1jlppJkLsub3MOyJoNKDKpC5jp160QPCd
b5wy8yJnir/EPKeTH6dnkeZxREHbCY3/+ZeaQy67lpvXZeY3yMdsuklyqeQT0zu+un9N7JznRjMO
mdl++hq8o85D0R8N4nZVPMANA9a5E5otIFMS11G75Rr7rtpLcBMbPq7KMAZu2mx9UbSif/zPicJr
KMMjcfCQwYgJFFDgIByWNS4JZvscl+1nG2xNFEqD3MMRgBgysJwzmE6+DTNuA3VSlERTVMotgBvD
r9DNbQ0X09eZaZ5D5b/vrViy1FifnVhfNMQ2Saerv0oiN9BsUDQS5E+TiHzHQlchty4XsT/buX6h
K1cWMxXR0HoD6jeSdHrTcKoEKuXcowEJX07IcTpNH12OYFzSZ0zTKsG8sU3TuNEYg4R42kvSX71k
ZzaF+uGvABk5Tgk4QLaE9Njy+GxQJ+8fTSyfzws8CWiELF8j/slJMaXOxZkjIU72Lday2nxdZy3B
pgQlqMRTvalqzFvo6wMss5WnvFnA9Qh/dzKhJXWZ15taYSkrq1+tj8x+hajsEtJZf/mUG2n8xCLp
s4BaEB6gGlcdUY/relk/zbCRexXL4rdLi7CK/WVS0ugUQG76Gl1cbbKyl5gtUMbJ8M9s7NSGNBFh
n0gjyN/uJzB1hbl0Zogb5q6khaPpNAzivXbN4B+vZ0xPKf1fYCX0mF3rGZitoTtDwTq5pyu+fJGk
Te0n6BvHVSN8wn2IOhaJnomQrtrIe83fQmfqVuuRjPCBDXI9tSjN1bA34GgkSEe3tACaJM4hyfA4
7OYedaJBIA9sBDF6i732kxWpFTCOkXHpN7JGOHhf9WN0nI3aD4/Ut5ZzUA2JtZVdmtY1fzCohOXQ
V/oEvRZcz9FRdiL26nKMp3tj18BmgO1N2+hNJjnwsRML2vCvREgrUFsrvlXD+k3FCcQ79HdZg6RJ
/o4Z8qLG4v0A1bdLbaIX0IiTZz6mi4/pbZ9T+UtQ6POUDlRmJj68L1+HIxWiZTsDTA/9PYVBqDsa
ai4j2cffv5uiSxiW4f+wrDP01oRlHnP1SzRLjGYIWw7lHLIzl4uLjyrSOxn/gBOlJbV2zp0cTvtu
sec1f1ZfXIAPLY9wdRufo7XHi14P4dEuqO6I4XdM1AhdLJBXBmfNAB82OXy7XoJPoyzAYFnoBN46
FIaim4GDtowfKfF/grer3vkAzRlqkwTwk865UWTbnjsaTCwgqWOi8RwSnXM0N8g4pAeOk24P7gel
reg51a59AKVMTS5KOEUD7hfh+yqVl7BKvsLqe2WoodQc3g/SitM5cSF3xr5Eda4tYEjCfOlzEvjo
Pk1hvddDQBkD+S/9dKD1XO1QROsSTxDc7wPQcMOx6mZoMNeHus1xvhGlQXK0Dve+GzRFwwzpiBnk
nTd1o82YHzwRI70Sa1RBt7/wOiQOjrHRIkp7YNfCGTp23iIGa6+ufkSk3zw2gf1ZW9+fNIJlmdWA
Bs1VS21anSe0ZBj17bvZkHAT4ee9Nr+CGxCOhsIiMCI7bx78muDkEVUOw4ypK3R4BJp2I3nt/Wib
L7JhbR0fL6GNOXHm0cGA7xk/VnROWNBxBN3r2c9kSYXIlvkE1VxnqjJhvht0Ew2UbUqYPor8Br9A
hKhDW0y8xQv7GHtGVluOY7YGggLVTRPYUahK2HPv8MCwydpNxO0+YyKg6j2XMLbd76QoUzR7QEHp
sk1c2kPowKqnGpayeEmdC8Jhsa2BMa130C1dW9dffFCGGgv0ivrzoecDFBpvl16WGJuyu8cXlFfJ
2aM4veW6av7BhIJpQERF3Zee0KcSwS+rtKu92FyNIEuwkIJ6oOKJBYZr4uKEIhWPtdfQ2pUKKHhe
i9YJw+xdD1BJWRh3a/kM6y8CcjOzH4bKhMjuRxPulAyU2DUQtdCgLBS/T6p3wkSbqtT/FEMp6kts
q2/RacPc4haTilJwa16KM1/hF31ftW9CHS8+mWWNDc7MRCSeCiXnF2ij2+BEYbGDTNYG3BwY1llg
XdsQ5bm17Uwe3zfnvFgxmQx1RNRvBdnbujMDAmvnDbuByor79zxrVBhEhESVLohUbKhQ8M33Kc9Z
RssEO6/+UIB624ooXfefepaLlPLskAKWmLkjsRbuU7n0y5jHlsFteJnsanj6y1pEakJtaddyJGYM
b4lKH2S52Rr2p5yOHZ8vglFlgtXOqzIR+bcswlH6SmDOS/B4sJVhHwkliO9yLlo6QUcwM59X9/8c
PcEsvXh7c9S6L7GT5N6UvKklnGijtMuU8HFW3oaHYn8S8T0WKxr0SnlnChQAT8SJFsapeHPpYN0A
ifawNJSecXPQj5MrCIyJSqE2kjZn3moixbHHPUZ/hTNc+iiovpvP1EJ4UYpoYX1kRO6+5wJIk9YM
5qQdtalW0LiFWRI7GZkNjH74UYEumF6b9mnU367pCgvxiQloSXKXjNeRuOFtQyTGl7/P4yqh3qP9
PhTmVzLGp9im7gBRiHXJmz5y6vfPQa146U0w5jgH34mApHhnS6i86Vd0vUiM2aMq556W5560xlsM
O5cYkc7zv6rGtwld/YCCcMjWlekUHH0iLYj/62G46Ipop2Uvvj988x0EmZHPML3ac1sLy2CVPHdl
qmP0KFnIlaRGjHQ3JVq82DwbN629HLNdlucdTnU6zcDc3XwFwBNjUlCfzmyRGBNsXkHWctzZHto8
LBb9GhRbHqRs9Y+xPm0NTTxqq0f3F6Sco4EXwXiG866yo8kJ3B2Kh9JHIUVftiKDsm7cQbpPKoCl
9eDvXE3CM/D/NR4tX0bG7Emzr9+UsskaQHnz5w/q2/Klf+YHwnmn2nhMenNBbYDvc2RzIuzSrfXk
CwoZSwGY99gsIbZYn14CpQZ4rPNsmFDJPFcwaItp8Q+32OZLSeNovWc+0J9yNNjTxNr6cHP0S2ap
wMJwgF1zThbRJbtgx02rx6VS0vMY5TZ/5UrCYEgQ77YRN2eAsCNZy0UZJitowjd8kbhwZDaVz58o
ZETsKR6MScnqboPwXixIAi3WcnnF3AMxVTsmxMzeRi4JogJz6MArcv0RDck1gt6NEthbxDTKFKth
oIdajNIK8+zZ72gE0rVEt8TWWbNDAJ8T+i3Fbc+Kf2JaLp9x0anBHdqBLvJvegOMktAZe7oKBc09
GIsSn2O6hbYrsovnQxHuckk1DL+tCgJ4bY3zsM4jj+KJBbxSHL+w0TN/RBSqLwP6wdFWLuS8BcMJ
E5ILlEjkmKwgsCwxXtd8+5o2nBCOlgBifxL3sLVvpqvV2D8B06XZIavGNOtAad4xY5EyioO+9G+T
cBXPaKj1N4iXBs+wNSPrtWjK/qNEHxfZYI2i27Kix5svcMOGdRK5LZo9/LKEscKob5x/QHcmsUuf
3vy6mkbsUgZxrel02l8f8IXJR6vB8dqOxqQIcBKwBYALOkqb2rWsdnIqnqGCAaMkRt+eD5bXX1wJ
3H6si746vFh58PAMEKjypFrIkWBjve3F8RHHzrrGddMnxZgSRc0lDU2tOSYGd8EV9y6Onf3I8zWo
fp0skgRPjHqxxRXzxzNKeE4LezengNFLMEhBD1X4d1tmg+t9zOQp04Twb4NfTcASw9IX9S5bw0A2
yKK/UJPOm8A8naaUwO2nFC1H4xg5gRwjuIMGHnXIJWgqKiBnW9GNzLapQ3TtpI4SsvFm3eoNbKXX
AgIvIH/i4zQqBs1HW145tRbwydhf0nhex7IyxWBqh82xrgbZyWw0yLgqUIew/qmbQF+C76/kl00v
U51Z8GSgJcD8Ln0EMA0kCSJsUbfrm595oRX7S8p0XbPGR6SefYFLPGH0ZvzXjRnfsScsxYcVmVjc
R7VsoHjzjTz5LhZ0H1ogH7fJLUaJw4dHaaIH7V5VlbEI2yW+52JAf9uSfKCoNBwCD3cSbxjL+L1/
bVzw71gnZFOTF7BSsYCW3ZwLReqljJECEfwIilW76RZuNNqRUd5MO+g33AIE3p9lS+uKqv9AvMCE
/eLWY6KjbgUn5um2NMUr1SY4o9D9y8u2K4PrWmzasBXrvaML4UkGrBXJT9S79V3Yhl2wNNJJ4s0n
zdDgNxxjNicl5dgOwD+PkAu8jcSXn8LY+waWXbQFpS1pi23xK5PKcfcluMX60F76FQFUzGzgPJ1J
vKDkQzm8D2pflBgFGw0+Hs/rPUlhAFBXIVDc15qeJ77hl5n0Gy/vh5QBfM3oUbYKiW5bSOmlmuBG
4JF3Z8G1ycOatq6SGfdQf7ZyP/06LEMMSP8+5RcRB29nclBM51Yqd/lt+LxEWSrnYph4k4HggCZe
juOyDps99IzkY5oIOToPX/lcW6fWjlYAd4XYEJGvtOUo+ooXlWsGXYZ3Io22ZGKcaMbry4LvP4vv
JQrGhX1Eq8035NI6Y/CRzt+CmBmL3DALGfuhHeNOrEK0M8rokOSEkwVMOw5qXV48a+JmOFJzvneF
RDZGOe51/zcX3dv/+9ei5nA+nnR4AOn4CKZ67WYitp4otdBNDezMu7oqaSdH/VKkXAIY8PjyqKZd
bIeN5bZkhBBIlPzy2cAKLmBCANbZ+e8ZE5a/RopH0VUFkuElWU/brw10c9uDlshvO+nM5GayCYE7
wH0GNc83o+tByzTu5q0uKqIVv8bQc1xJVkK9P3J0bpQftEFZSyBKBfYHkS90qL6PvNpEizrJN9ZL
M6y30J/s4lij6fO0KR5oftE3Y/7hmNcwa3jprPMfXujdf74lmITzpvZC2RKqn/GjObQE4DToNlAt
ieH37YuXoU0jh1hT2OzkupDLvM+mWqK3k7bYh+EUwdgANHWNv1anUfWuKbNfXc4c8BhAzMkVnLf0
DvHIt5HZGX2N27ez8fBxGhxl6hzjixtfobdQgbjz5ZI1n3/QxIi2PjjlIOADhMnhFzEgzJhiVXsW
DRuF9jDZUeo51e6/vAvw5m2VzCbRB5wr9W7eX43Pz/JLXHRu7xbdjTBYqUsIe0G6+i+Yy7VvR1/X
o9KxhdG5LWJl7RvKqTKBvyXd1C1v/tSr3MP6WnVQLH2OmTgdd62uG84qhCjcWEWnUW6MR2wIjjFW
rK6pv7lR9XF7n0f8U8Y+jK27JV1vskDz+1qPsjzYUDvB+L8e+dIzYYglgzM/MhNVdZAmeqD82xtg
FGbmGEqlRJCP9izyqayMCcHn/7dPTTHxwRoI7OWos+QoBePcnpCHa6vCx1eVOv/2+LU6V3j+4eME
Ljs8H+37dd9YymHaTsXvNfy1Cq+4gXsCatmpzSuWGTv6wHaoVffXzkh4tH/uUNeK4nfGVmpSDGZW
ZmrI58wukwHMBPWZe2XPK+wfOrhprX0CUqD79ljGzIB/jKwK3VN6J/9+n5ayFKQ+/7449Jx1Ma1Y
tTaEHbyCc20m39Q0z7HIYe0N82LwqnfCDvW3zPytDhl9s754EoVChrLZdKzHVRhHUwxITv9DK3Lx
zhcxDfNpikeuCb7yt7ir+O4cP7HR6o4ovXfaFU3X4DzJitDMcIDK7nv6n0b9y41nDkGRu4umfnsy
9cZvAe1h29St7KOn4Nheecfc1KqxgKFM0Cen6Bd5hDScowgDAVQRPBqQIAIGnXmf4NhQ7ZfMob9J
X5LCglEvN8p4id3xQBw4FgMom+IB3cKJX7TelMBLVExHluzl+e2sgrlkac0RydXB2VtiPvDM44S/
Yx2c81VXeMAQrxiGdyc88M5CK4hit54Kb3+zYorzRPv1EPGvnGHhWVJgda+dSFd/teiCK/5Na8O1
bgka0Q/mw4bU5j3NDC6bZYkl3OCcg8z92DRI1r9t7kR8TY4PAQnrkACIYZs4dcvNkszcjMg2K9l7
UpBo3ldWgnqxOxHkbhlVK3tFklzQq6e7zOtl31nLv0wvA9VnIVR4azxyniQgS50LJe1Msxr4K8W4
kh2r8AW5qEZS9wuMILGdFUBkL8idlFgzvbzCWnxwr6zM9qhDZSqaBWx1mfiJK8fsFZlFV62ai7eU
mtq3gmeLtzm9q8hFlhiiH+5jMyt6PUjmnohpqHY0raeBwpQ28+7MhSax7PopFS19lovgEBf6qF5k
G6EypHxFQePnEhCByTFhaPeqbc41ZEsDnlSRmqRchgHPaQKGHYUeIk6vTr46LFrYSK/ea9Mwv4fq
xFLDqhTpXnxhSSR1TzI55WC/csZPD7UuuF4s13rSfwDk7fCXUxoD6d+uOAcXY/B8xBgXqszjmbzs
2+4aQD96o0wIX1bTuZZYDTTww3OB4zi61pGqgUAH31jWwmflwqfbEmPnWJo6eIQkSj1X9IqIMwDD
CZC6/b+IcS0rtmtmVUzLF5oWSGY6VAtDFBIgU9PpPu4KoWu0UsxCRDsT5InJ6baKvrpytGkHu3QG
EoZHn2bg3R9RY1Wq7JlyJPMv+bsqhFJrkt1ts6VpHtWEh+lGDqnvKMgho/tUwbiT8TbZU7CyS+Oa
6NEdqhqdfJvhStxb/5gQ1BoLRWZs1GmgJWGILlDhz+QhXw4C4XpCzJOx7Qsn3fNcIjhhTMjdg8Dh
9yUO1G9OOSLU1+gNF+8Htcd9qE1lEm/B/H63CiKQYwCshRBJWY0oc3JOtt0VM/FjXNeZeuc8jRP/
zW4BmDKr0SHjch0oeV7sm9GYvezeRVW2Za2nulXLnex6Pkfvm87GLvQYtCL2wFjTB8KxVe/8pJUg
olq4auq3NM4v0qyyru716bfzPtRpkeGCGexSwW+1C3ysOZgmbHIzZQN4B+GNM2eB93qerpzjpJ+k
yqvFFzT0xUEgZLnZJyIYdqHS/Zd7ydg0/6dIWkbhzYLE1FS2aWfgjOTMppK3irH7pWj7gGNiEljs
GDm1Kp0FAwJWG8/Z/nQAnFznfR73YXKInThXsRmVCfq3YGO+jECMB09j8PSjl2ZFy/B+xO7v8PUe
dgiIWfW/uermKajN+X5e5EYPiB/DawfUcWmvjo46zNeVey9CZq54msd0RrXtKpz//F2IGPKglwfB
ZJlfp2lcTkDwP1PdyuhHgAkbn73QC05wlCIk3f8BDP2CIW25wi3+uS5o3yM96khcASh5Z1J15Zos
2BO1RSsxUgJPrK9MwhN8exAKUNvgip2C+QXrMJPcsGpoXNP3Uw8ONlqnfZvh4NpVAbEiuGfoBdJd
szGybz4m0g9XvrPdJIKol9Um45GN4WyEsF7I6gpL5fVSEwtvFxLfKhqRYnLfqtXGNCNKF3SOdAFQ
gQD8gSsr76T2s8fYMBTFfDIY/hGJ5RetB064JLkDz+XkexmmtAF+wHhAY1E/ZWUOU7CjdjK/dv48
+jTWcnE3wlLuo3juORbbXg8VnebQBT9D3lkQqV6LdB6cjavEUrCJOQztb61oTQ1B8kUs1MlfqjYX
b1o3xeSU1VowHHrvj239L5xHAtxis+uCjuSjHQ9o51Y16u3rSaZAcyE9nIYG2g6FpaxDbNwD2Shc
AP2b2rNzb1dLHwen0101Izh7KuzFsPp9y2MzFZHGFmSIEpNJMyO4MPXBgplU/CSqiSDbjkXPpVS9
hOFLX+pR7d+CP7oivX5wwEWFFrMRCDZRSQij6lVu3GQBHnu61bRgrADrRx/h2u1QshlWgft3KGL4
bVcWo7+KdbAsRSPRTiPtS3kW/z3QarMyY17y3h2MCq3wmQR51Pad+lulTs5OnpmddUj64hd81UwY
NWWBDoBFA+y7JfYbCSESHso/P2oO5n1XL6HKrCckT8l2lUm+sA6Y4cjc3DjQf+K+ItQj6z9igDv8
wz6yHTSrhw7HMKqi4UI8PIHgII6a3wdmLlYB67wq8h+yUP6HVphI0s9RrIWxeDqf9tWbFLUVyxlK
gu19jRTV0H4dbZALOVBOiuJ6PiVZOi6tyo5xq/ZLwyf5NbejEpm5yeAsHJGyZK8319lW4IYC57C2
NEAtRGdpwWJtdXsJv0TV2L0ybypuXi0CZAx3J1HljLzV+OTTFeyXnQq/Y4OapQRbrDjlZBbcgnPD
ZS7d7INkuNfwIEfvHKEZ65jgdg4YPulqdFgAzIip9Qvgx9n4kUPEJS++/D082VHXwc7EJEyQM853
bUqXHaJqhzYtcBxDogBV6KHY4NbJP3PEkQOGrHm64iO2Dc0K7ht9dXqDeC92DMcgL3fygtktqFCO
E9VuhtpUct8vVCjk2TnVNmugl7SF+fUSYN1wkVOJdjcFqGX5uT2dA5qZ5vw4qZ2uDMNVulAx6KWQ
MQ5pf4EpwbjALCfr7swxl2GCmGqsQeHlmitKW+X5hy9Xu0zmqDfz0xCvNfQgjMx0hAbsLZMws6zu
GwqGZGbtuANmeQM3Nuwf9OOkLHHqXlq3spBinm4UatJTuW80MP0zb5L0Xjz1F8PFWAjCihrEHB2H
oOL3GeuyxPUhGjBKRAY07rr4uSDU412fKhMcczxrHgh83stzhnQc5UHeLnxcPV4oxlW8skovxQjp
j3dTtpiTm0DD4wKaBmosamObO5yEU2/Mx1ylMdytDdvHZ/UyKsLyorIvsQkb6+fvMF03/K+CkivC
Q/e2KauB3kWBPIUwuabT4vtGu5v1/EJh0w4JUYkf678Hzk9lwbRHJxQiBBlfspnPl4B6yyjo4wbo
hPB6XLj7wsJFkPYVXQdJr9Vwg3Z3iXHnNCmAmD1LWLdiuP4bD3aozWdrOsjrF7Rgz7X3/Y4FhDyW
piwdJnP1HeA4Au61KrB6n9ki+MozdZtC9C/R/PzNZRx2ca7v58zYOfgoylMjt2iWW+VkhQXS56Qi
qdhBi2qt9gEtUSkqZsyaTEnw+ncmjwiYO7VOqiEC4SnX3mHqkE7yh/6XcZOc2DA2vXdPdzvRD8js
FSnkv1saYswOZH2y5gS+UNVojbjZy3ICzTOTPLrDtAXBugNmuVEbOezeNKTooABeP4ioxlryi+6w
nRZyW/GP/Xui6VhyPkgmS+7Qq0KqqbldxufBYy0lqTPu6rP5HIeKfKna8M+Fu6h9Yj8EnTk74AfU
Heq30ZpEtsSJRIOEeb0fVczDhMSE2mx0sMpMzMEK7Qa/JV+o/S7IOgBpo6zlqfgVFfCV0QENpAc8
ANB9oZjcK7sKnE4uozxjZeJOfmvXk7BCkgRjMGFMwrFO5Gz2xoc042nR4kqspnSp1oImGtEbvxCm
G+8Xxp+rf0P/MOC5RIElyVgax2kof0k784X0jyKsYeoGobxatgwMjp1gW0kOYHmUMtSsYYSoQ3Ff
M6YoGovGZ2e73QN90rF+00o6kzyLiLAoK+hm+PUmgx5fVVPi3nMxsfay2Q9UAUOkKFqO1G3ipcBi
i4oXkwx3Q3vz/+4QuqVkKyk5aelO45+NLIUVLBU86E8uykeCSnG805fLpZ+2wzOvr4iJqVCjdKW3
ItzUCrQRxTguVd0YygfzufdtJocTQtbJT80iv5Ezcq1xHSkAp/hzm2R9Q2gU7c9yCYufflGPoKWG
aFuyPwZShrhfYB4igikkMHm2CfedpLX8T8ebaQCKhg4UF8Ze3sTSu9e1uo0uOOnabLpFiKdq4X17
brKk5kQNd6aOMgVV0NRi2qez8j6NcQlo3AJXdWCazX+oK4H3ktFwFhZ40CoMTdk1n0A8/cpL5HuA
NyxMv7q9pt8YDDjFD70j5h9s/BpKFhTATQzl36NWZAPz5V00uAh+RgQznoLKO9L8+BRWmEn8WBOV
22FwoYW+SkdiRXFz6JMcJMRT6AL6J+EKCAi358oMs4TQQUU3nQsLh+fmJfNTR4qLLdszb9AMlHs9
zh9JoCe0AR66lTSB4NGvfdcbBo3mhglBjjmsSo+c0cD1EfT9Jp0VHtC84dXXsHGEKj+Mp6VO0ILC
i7J4oNCH4NwDZ+f4o6cY4Kr3oSR6+a39ZKcTyan2b/CKhItLiODoHv5PuCt6hJJ8MwGjqS/lA4I/
euGnyrtP6vAff0jAk2nsgG5xcI9GPzMtHiz2yjOInFcI6Kteo8loBjCtKG3IHrbcrGonb3VzM35k
jMGmnfGr4Uyp93WcquZf6+LdlT8KgSObLZhUbjkTkmA9j6ruMvTpuT04edNt9XkYFyuPx8WeOj/W
zlBw/uwNpIBHeCKV1ZEhpPoHysUqTiyWXRVBmBhsfj6udH3ru2OBPOhK4WleIiusUTecml2e0l2P
jYoKX4B9um2dUaI8pDUwcdaCpOm7hcuGnRCxVKagDQ7yCmnpA+HfJk5jpV8ck1rwBsLzNf+xasQ7
eUH8wNNeR8nFD2hDp3Vk/jbNnyvivsiPeKwB2CKTGJZ8HTqsiZ2zGc/aqgrLPh/jkS/LIDlAxZ+o
d59DORXjwC3t6ibZyEHfI1RSc6RoByFPywcHSzxbsBhzsNbbsF1TGVUUvK1SIHJGLRjdpYTd9Ruz
blwJqP0OpESEe3pZN7iS2FRPVYNVW3nHiXcn3+G6edioaInO1AvdsFU2s54WXETweC9U5e3R7FfX
xODXpLkrtf5jlqzU43I4UB21z2G+jGxI1jda46hGTX8/gHt9EAObt8YnJYIr6Ad9L8N7NmvlhGv/
VNQepxFLOy2Yu2SP8/qHNp0VOnpxzrb/x8DNhi+OVkyAlype6WUPOuTU4FQYil3bQOwaXzro7TE4
9d3XVyrcyODAznzv4dY9tIzAgobqG9hHB2yOwoxUq9jIEpgIR5CDyoWQyMX1yB3uCvv7jzgJKVCF
HgGp3GshiaMn9wiqCCy9R3i4TdTpPqIz0oNv3gMb3C1fXf2hYY38YETYTFSkyoVUrMBVhUkaChaR
zxKYPz429IhWvK57Y1F3QPsjoua/VotRyGiyMyvVpIUs0Y08eawkBZBUOasy44YHLRkRwKLLtDRz
Oi3oEEK9lITmwhGioxHYe5KZpW/C1AzFML88gUgAECnGIZmVcvXhbBVRyqF+XKVdL0TTjvjpLpeo
LNOc/vJ4xb7tGNdPx4tJhj9ukwami7snk6Mi2DXekcT5S8xvx6EJXrl0TeS08YvEswlrY9XbEt1L
pbQeMGEYAAuflaDTfqgnLM687vR/1so5uQBKZHzQP0S7fJ2pXtljcJqhAi+v2HnBdZIrXf7GIJ4/
WJS0jZtDpEruG5fVY65Wmmwp2VnCRf5U52yerN4QQEqrMEl9AcA4tSdCiAlMzhIGmM2bXaEE0pcF
1JoncozWvjtkYzUc7XDSchRtBetd5LtL5vx6Tkxi3mNiFK9H3PSFRnxoetkLdhjyaU033ELbxF4v
sRUo8HaUvxEpHjo8+9WLoBDxvzHXwBTVtSAR3HtUhhFBZh5Ltu1/uStCzzPiB5E798ChOcvgdOn/
jdbXjAPlDSgXxMGW2S8EarNmBghc5xSE11oHHNcm+fmCZnt9lxaCtQxIfaLP061E9yyM0Oe/T9C2
2Q2mQaKFpUx5ZVvyJJPaUKQFKHXQkCx5eVSXj9PC2DcELLxJATtjcx095hyK0ngshcfiGHD1TA6Q
QAZUXmuJA042tZy+r9BSx4ilZBzR2PqtU6RnbVJhB8BTpy3yZyD08LvYZp1IUxKSeB+cFCY127mf
0NzTfvtsDz5MUmJAZcXzrtMmMHKeyr7Qeo1+ro2fk1Ja71QKa45ROIdq6NVguzDvK9cB9rRq0pUw
QGHjt6ANB7NDtaVsxzKV9AcmjIkrCsKP87xyetCKYlc76iey5/2nk5Tobafi3BlRjsd5R9wJsjK4
hgoUcGMBUvmxWVPIcyfZvPpVzAR8OzfeO5ePIAPN9iNJoranCE64ZT65loQACGUjE26DZuzwRbrQ
y+aHBIrc3SNcGYonLtqT5A7wekWCvpc6VBtMXEYvzW7nbCoShapguzjJqHnKS8i7t6w4ZJMIy7CJ
OIpNwFjzX2dYXXIDZ3M6QdetnTv8QVd09dSnZPJd8TKrsHAgQdZtrJB0b4ZCMV0ByRyEZpn0xqUO
EGtBbX4oPQiy3R13UAqwnT52i+BR6FQwJ7/DLCT5kA8+hRhX1qX8Xlj3awIZ+tvBIsLEcCMS4jGm
j1+AYCk0TU/v4YtCVn7+TOnIrHO8eoDkbjY+pn1a5LdEqG1IAwMnKuO7oxSxfBO5VpTuNos6Y5Mb
ShgGaiT3BiNWu4d3e1zuBtdvOozk/K/MqIz44Lna7NuQLXGgBYyEDlx8cxgEZSblsm2tTjH9VUOY
Xe0kVY740B5MRyBGCxKR8ilKR/GbQxEBludG21MHU4miSFl4oZvpVsIl9Z2TZwosIwZbn1HATsqZ
YKFt5Fxoj4FLVOtI1Mdi/5pWemw0nso+cV5yVN/6SyuUXmpJGPfx+9EWQvy2YHY7pYsAbJDad0Ts
1MRW5qzTsiAe1HTDA2xli+C03R7IRcfW3i92qD2rEmmnQIjtGXM1/qKWDtQJ917EPMhlyyYgeyUl
Mzb2S9lfHXGCTWNaXAqeNefoCTnL7n4SmUXF9iWHDm57S822npwZM/FQMLqu6NgxPcbC1Ykh96ah
keuGfY/sqlNf59ADRDTyVmqSTA8TgMUf7CN/NYk30PX/k0m+D5cFYxsu5aEjaKRYCAs84Cvr1kkA
RbiG5L51OLSqKO8jdeeN25MAYqpDQVNB4sdW8xExVdPopGjiuOweCjuIIu2FW8cM+kE9mS5ShbUi
6IU8nrcW3e5Y3YbnwY6nfDFhOkagLL/EnwORpEDVJaO1MiP7aTS+0bBmSuct/wG6lALO5ORT4zcX
23UROGEuHZ9qh4YBL3/fjTL74cRVyFWRmN0ap92KvG76PaQ4yFVJvpm94p33/dUlTdl7h/RIj7Wg
M79Q4dJ4nMBJJB0ebIvVbCvl0CXe2Q3rYTm429uJ1jjYZg28Kkqhn4e4ZT5WGnb0191EDBG+XKTG
RZUr7c+Fg9eyP/9wBMX2P06E8roiIfruuROKRQkXipKaB8RdUxfWEbso2HwkrWoHRqKxyPYRqc53
d5IzY/942hUqkArwdEq9WT+2rsK4VWRDE+fkTby0nN1n5eGtqfJIiCohFqYVGTnfKDa0OegTT+Tz
H+m3/8fk+Qr4VWGuv3TMEzjEHR6N79x6jpsd+LnVSKzxry+FvzPyOh9X5QDL6287YIHpwMpIX9p1
0T8rFAVm1jREiCHS+Sail7HWbbDRPUDe9CljWxmbFou4dlbf+rK3H4gEu4ekAeKuk7Zd5xV7CSNx
BR3Ow8xlizh50NVpSJJ13CSDOaftr1OVMJtoY+UB35kUiBn57BBHN0Q7afJmhmyBqgzhnX4lIld8
mdRvCxUT9J9BHknj/w55UFuTUMvXaXlkYLOngYLBr3tojtljIueihK86gR3zumZQy15AQ84LOaS1
XwSsqedZWoN3l7M5KQD/tU9WyqBZZMWnS/MQXNdXVXrMxlSy/S4pH3hnvkeFFCzxQFIujYrbC8IX
QPRvB5fbqwX7xLplpqPgu1vimHOcXMOG3w3UxhfPfHl0iydiYfyKt2p9q6AI2ugWV/54UQKALhP7
ZI0tX4XYXI96MCPjlDNrvFlQ2DDCI887uU+iImeCsiJiRd5ujpezqVtd+PCFmFCOjZghoVmSijsM
U/+qaZei+gDQUy9JupN+y3Feo3l6JpKiDZGHyv02fzGLjEaZ17w5aJliDbKGE53V3AXKGCrdxGD8
Wseo2IAeSi55rfAFPurH8LSKatNTM8NF/IGVyKjznbkQZN16plMKT8U/B+CyqWHPDNz1qLdVW71C
3ca8i23t8TEAbCDccxnd7PUiTccjBuPHd2bD+bLPydyIEiG0WaDz2saRgABEtbYnfUOaauENiN2d
x+29KJT8C7BwE2GMhTCyTcsCSFdfPCUmZF82FwpaQdrKJKWPKMuiamVfrJuO9nhLS/d0yIG7h6u/
1f7Pca9HEUOaiCdgTWoUVJsi4hfM+caJ57JdUg2We3eaS04H58icm1EVB5QK73mCBnkDlKJlPWil
kvq4DUFCM/0+3i7kpcFa0xBEWMZz2SRuJGxN0Oifejp9hT7Po+/gO5F1P8JlDQRm6eaUC3zj0tKc
ONllMZmKYYpVpfSYNPAH4zD6A1PhqtySOUvdzzZkQWR9KTyoa6P0F3jr3YZs86OR7mfst82hjSlZ
sBrCsodL7OWSfyJvVnpWjzl14M538rLBTMG3wI79ZJvb6VgnqM6+YWw4Qs/AwmU7H88hbRB9Gwou
v8RXValaxrSTQH/IW02VSXkIcvgJjkqfjSTQ+3YgVUgob2xfcxApn3DKTEvHYuon4a3DutuMSdsn
QXjMkzRBQqO15fHs9Q2k8xXBeCpJhPvNnqMlDLxwQI4oHbzblEggUy6PEFnfSGoPIVwSa9eT66sd
9UaV2yap/LoHJWqk5Y14c1YjYtROuvFngLIJnAerWoBgN18qsymWjU1OiASMajI0KKecMn7pL4i7
1AkaKfCE6rQ34MZW8L9C2jzEP7Hs0iSXIdYbGovRdYW+l2KScTE7bNUBVLbkGtnOVxa/vssXGOwd
x6ROgeLWqd9fi9a58Ls784HhTvRfttTJe9k63xZkz97dhtmWgTdQXCc4B7lY0BQwjQDGoTi7LheE
9Aj+P9r2W8TaOui/tTX9LUAvWoiJtj82kTucoFxnxTzh6F+y/Tk65fqcFJS+Vg3qSAm/a+JkhB4F
NggrZtaHw8VsXN73EGvTgnAXYthdHYBE5bI4DL79SBBJl48bqrg0esNri6jN7If1mkW7mBq4zt5i
ZF7lhDq01rB7eF/P0NV9q22zqTJJ5zcb5JywdzeGIrrmPm/yR1xEGG6X4be9UyfTOQsZ6CbdD1v+
0NpjJqJPoKxn1CXTV4tHu7//tMF4skFtjQUv66KDV3eDXF9GaBDEKYE8XJOPll1fUA/0fxxAOl+5
RPSfNmzv3aXk+AKnVqQGUbtkNOBclMIhzwXewVB6k+r6REBnA27h034yaxHo3km8CQaEOXLoKOAS
xfsQM0k2zx0+Ly/1AdHb5+pmfk0ZxsbRz9yXtnQaDhkiulfolHkNJSkkfCgHCMhpwc2R2jCv7Mb3
ecmePIDl2KscGm7ZQbIAeLnaALJTuDUJ0mPe/D4UKDwEDZizslt6AuGSzk4J91oIrs3qm+vukTa8
v49d+myWNOLPbYzgv5AmMUbboU4s+MTp8BA3cKxwy0zTlZPlag4y503eSDv1a45KkC21in2JyQZa
ZdoF6KJ1uVBCfZUawUbauhy3D/iMveVeRbsRg1GFN1GsglLyzdlAVwNKl5/M1JUbGrTeSnT38dFc
h+Ggr5yfIKhpAJniU1ZgMQJ6TOm9PAJrxbUhPhv7XTrzhRgxOLm7WnqJW4QBFIFXtJ2UdVcL3nZi
SbUkTneuaVXWvbCKOqP0j3DIC5a8CZ8M1joRfSTP/YUPCZ40Wcgx30+sCOLXWRrp9B9/Fuq6ss35
DAzvHI8WfwNZveqwe6y5Vb3mPA+rklU5EW20XGPGCleGDsfyxpv/uy9po4G4m+t039VyQ2vk/N3Y
Ykyfu9zNPvbSiD5rMDZVp3UcFH2Sj8ZMHtRULxKDwlbh0RN7Nf9eTogjifqvSlAqo9HIW9cBKfKI
K4CPsj/6RjZ0AhFB3oXnl4oapoqyCtnClsfz1mb0MhRVDc3eCHlD89Izqfcs3ESlnd7NqwyEFMMv
IkTRqN9TEGCqFtzYC6KlA0qBYwl7CtpnSUZBtyE3doF8JSDUZDPpELblo0RjB6kGGzZLS0SZLSYc
gXR1+nttt3nXOBzaiO/Sl/WQWIAg0kEnzByzgWux3WZC5FOORkyj8hUtM07ODNSd1+IlmGxUD+/W
ybJG2LZC9JGOP3gG7ILzaKkfCyK88b5qy1g2GG68HNKdU893huIw5aPJQyojsO7bZszbuyFhr7c9
Upa2NZyxm2Z6Uo9xRh7iN/ht5kDu22hd8CH/fT34JK37I3QzB4+qfVhnqJCS9/co62lmigaUB1kE
vQJwMRCt7dvDqgdbI1RN5J80adYJ3Xh48XTF5hCUJQFFA2u9zh8hVPemPTya0E4RSFzCzfyuJOU7
qtv0DDFWguSQEhCZis9BAJ/YqOPHNOWpnk8wqtI3dezgL9mIis2BTi/H5q7WWB2Yd9zXzyGTrArH
xQoqUJVzeWrurYbtOe7MuzQNk0tEGAGrpajX08MmXrJBa04rDqTX2Ggf0t3k2J4f50nDl4IfHuFx
YWQe+/FLYamG+ecowEsLw3nFrqpDk71WH19G6xYJYY/vifLAoe8ZAprtSA16/ozV7X5/LXWGYCXO
7ZiIS+0WllF3hNhOno64c8xpwEyCXQTzTl0ngP4+Rh4NN9ir/zi7WkXzenDU8HPy7ve0faMz3CpQ
84ZZMnCAMaDktNnOlY9E5nSsZzdgAJz/9zrh6zB7hw/bLEf1lJyAdVWwvVZa/fbsPFyIUDR2gKnv
hMARora//18Qp377TgExPr3fJAHF49fRystEL3VGcbtA02qPatjrYbpk14bjcmO/z/aeFOzra113
6bFP0S0Rkk59gEHvWKPBooyfsnhHXFTAqxjxO3dGeRYbX0ouH+9PLBPPLNB1w6Z6yBTO9DNOlKdE
oeIif2XyalO0KzwJplmNlhvPFVs0yiYc2sWG3mifkRPna/Xl9zhfXj09ie9iLShN73WtiCQQLakg
KTnssi+15b5/Yx0vYMDEFbEZGYLfhB963wqXWSxx2Zp7VdnAC3QLIOsl2v43Hpn+/cxQXCHDXI/n
GXQk+yxu1fF4J1VUJD7DBjO4McxpVKn200/+lW1fSdF7sYR+QPzKJW55d7qfxfMLU1pmkAUeR+0O
NsdJO31OYGKX4fZj4dud5j9zaiHFoWMzbz+AVyk6BB1Tue0RhwZIYk5KNd+TVHPcP/umhQet6+HC
P/vWwiEQQVshm3CjCzXHMR/pQY/bF9CnLPAK6GgQUdEl3f4DpgwGSqCxOuiFez8LBdhh4iWGiePD
fr5DAQILZ1oX1405+voQN1rgAJHFBOiM+ZxBOs0M0ywYU5Dxxq2LVUxyTxq8mJr+H5PaodI7hGMw
VQ+8Eh5zQCcObOKsvvZZ+QsmDeAEmcVSoU/mhdcR7k/DEQgToqwBKPKK2hqr7PQC92keh6KKLvrt
DGckorAX05Y2WEllluzzKgYb5M7uRSnoxAfuFamR5c04TmrkEEVwSAxWVfwnUKBRXx6s1006bAvp
zTAlvpVLOUC9qqGq+9rBDa37bFlOKJbvy0Ipn20IP78w3t6750SrebeWCqKGULb4C39eEeFO5+th
/8YeKSf4NQHoj2ItUX17UK0jcSNJ64bKch9wD7bAhPmznKVDdDuIjrDTUx53lmAyd7o+/SoJCs8J
2MJK+dv8vuMOjhVB5E9OrCGqxB5GkQCFdfiJd2oIsxuSand3S7NO18DU5oSn5czi5+XlJUpQdl7r
4D8CXy8oVPwpA9Jr048mR7fM+vu4uWVSGO1/WSSZkHAz6Ut7cwgw4sBfHi3LVpUT1yc58AE8xMYC
uWaikfczNL+Pf/85Pv2Hc4ptHSlGsIKbNhlXSnRirnQtnZvfSqnFzGnLvOiuQE310OkN+N5BU39B
hJGoipn31W2twBe0x6tC/3x65THKneX9XqTQOUXAyEbh9xUhGojqitFk2MGA9uwJdkGVJWxRqX7z
iYTTDN34UAOmDXojRqwRn63/feOFKNh7+CJjAxcLdVhDKAdI7uhYTC+SxO3dNGunLfzkJry6bdmR
D+3OlcF2HODo6yG/IreKy+8CEvg1zhFKGG4N4QIx6P4c5RK3dGN/FmSANz+ez8XLMTet++P0a8Gs
nmabb/mOxCsi1v1rW7R1Sx1FVqVi+noaRSwTRABT7DQQmfNNyn2Q0npQjHEdYRhq/r8Fd1+v0hOO
Gb6Z7APnGzlq9WciP+iScY4X2Q9pH7/oMQBd15qvcTCwjYjv08CWcZ2GMW6P0M5ict5xm77lPlL7
pNJmYGHWrRm9xUrMU12+03kOcpf4A1/yXaGDpK6ZK2Ve+jAJC3SW6vpeiPEUKig0PUDX05FpjO6g
KuyT4PO/+Qp/CE6pub+C53/2sI+uJTzdRG3ukTkjgGMzfm8vqCxQE05PvicQzwUmd8W7sa2K6y6/
FaxUxYedYrrPqCryMZKMPkUHJRfHLAFsAEeaGpZofW+lJvQ4vuNyyB8Wy7IUsv44Bvdv87cqDNq9
F1QiPs0rmIDcujcVL8u7Hnmx+prTNUOJzsD27PQlsgGV7cfWf2L0UVJe7TSSeEp4FSkXrRolzGBU
LsvII/Ho7w4z5gwXppdBhODWB6+9NxlyhICX5SJR6HUzZhPqFmO03IjEQJ+jlRcOdoWMY2t62xmT
kwsSENjtJrKu1dxB1iVddvgQtJ8yHMYPWADHCKBD5d8mJCPkSmn/g5RuGbvgPwZ2E7Gql8QDgxjZ
rEBa3MebXMeFmK6yU63//E3XlluR+w0yx7lMv7v8V3W9TMxiMAnN7IOts8/8XDKhSUG0HFEXnjCX
OPRE7GEORBCzuDP29PbkZPcDfUT+E9uZ0GQLGC4PnLSBaN4Ecd+1RFSsxdM1AytGIqN6Y5Sxyi0c
fTzEY7FUm/Rt1CAr81sviahCz6xaf40vqy3Bztk3lOZjsK2NNieuqsiMzSHfUWH25bNqdeJU59ho
saE7kEPB7nWERkRm+jQhwaoLQZ2f+xnOvxHmyZDcrnKIWEbSK+bzKdJ9MlTN7tehA2E2G6FCESt+
m5hPqizeFqGE/l9+Q3YirDtjySGUyzx+5ReXj6LK3U3WppQrmDOYJH2iNdvx2C7AETGD/l/Zno1b
ix1+8QEVmmBRU+OB54yRB8H7oJ+FnFqshGRepxcvId81qrI7W1b32s2ULj7PCTTXxFAu23Czbppu
oZinN1FWnpfjaV142PCDsR+I1F7IheAtN12UIIgacvAmKMCHCWitGLYPbiS80iDJWf5bVqTGj9qf
F1/2CyxCvH0vYGi9gVqvmV30DwjLVdTqurfjJe6AfGT18ehnLc06Fh9SKHzC3UFzd4+SEhbw46iX
uajONtgM+i7CeTXX5ZlH6oj6y5jz6uQGh9el0bLOKb3DCNLxLHqSmAqB3yM2Wu4DHEmxy5OpyVc1
NBo6vxlIZDm4MObffxqiW/3kZGnI4Jf9zpB9BpZ6OR6QY5z+6Bcp5TSO7sFn9So/M0ZYapAqLAHP
dCnx2dNcpyVMDu1kU9JAkLnuwvrNWessxwavdx5gkSyuRb1ndol44ofCAWK9Apg6atgwH6y7CI7X
WuXlDmTOmsxPQYmMvtNaQx4SSGvvlc1Ck7BqmCpHU9Wi0sDyQFDImAe1pCSZPjvJrQmVasSvcbUh
HDb0gtgDG3elhEHCSTHahNjCfIdT3U6Ah9LBOA7FC+bSNM0YisyalgRFnXn+agl7Gkx0DrSdHatJ
kEw9ZO5D5EsJCsEYELCnOq3dAEAct/itxFeyPqVXhe1P9Y0HZHwPg8rhNb3MWMpr4BKLwVl7wEDv
zxEK4rBNppGyvKJrtCM/jgYD8QhtqetLVzA1zt9T7LkQy+FRmV9bYysJ3C1Q9b6Cfdz5O5Je/Ivr
RBDn66+o0G2WMCk37AT4pPSQzph2jDBQWzdNkTA4O9jrRTHtokfrlidcolsIwTMkIib2YwL6duoH
ww4cJFPIEQLa94oc8mGfPZaxOGTwDKoSZ8eCKIEtPoiBQJrvGVh4wnm67/7T9QjXv3kBXeHatGz8
yNk0/SnUwdM18/199YpNZBRZ6O+M0KavjTx+QoZFqz11Z1ymeqqXNp6WeAWOhtacsQ1GsPoe9aPj
Gn+IFj9d/UuYlEd+cmj+HEdpf9BrS52epiHnOq7r8T+wCDaD8OTr2BPNY4pl+UM8DFJyQ3RJxS9x
j/qTa2m9MzLE2yXuVhFXsZSjDc6VDz4OSDAZGMK4424abITjopE7Uk3120JuGssyfp3gCj1rgi0M
OVfMmihyDhXE+xzk7ydBggD0EVX7vGR8KKRkfs7Q15Ph4UY4WkANqFUaAGFLIj+4fxJFMJzhr0Cr
jHHLMCO4zXpRZHMWcf8MibGdbhvGitak9JRD5lTHN+NtnfMHZCskSbSN+kPeGKzBwWqqyO2SltXr
kcxlPnx7qNHlBqeMXRELXJmazWzguQnhuDfhAOy+krvvs1eH1sCytJJ57hjiYah402ugfnEtx+Lb
UibZQtSlpLAcq6gu+J9VVReeq0twCiE44SJf2SJhtPs1RCd5VafarIEYDeSeNlvPRfXY1aYWjXTO
O87LQjTPmIIlwvWh/2GO7Nbimt+xb0HhZ4MLNzfLkPPRVkYQAGSCsrNPOGe1ohs7F9cm2TmGljAS
YGjX+dpyQ9FUEIjGp1wusEYJIgCS5g5NOyX4V9+FY6MX2FCHiPpIBH+cCL/IXvz/rPYkjxNDkwW0
H5tEceBTEcWkhj7ya9e7isD60P4YnCZjQDS2M19d1aMcLhmMfzhLPLO7TxFSSKPaCyKhlj+bcwZt
yXCWcuTBRfRw7MznAcTKXUZK+OOIVdyo9106hvUQcDVE4NgDSNpGmhYxfkJAod92brs/cmDy0hvW
FNTf9eGzXcVRCqLdwYzJAi6tZRDjOgsCYeG6zleyyld+/0TX+2JW52eaL45enAexJEYbzbh0M1mf
w62bQuJC/Da18ibOPfwJAVViMxOtW4rAEW8/2Py042OHjX5LS2gYxvVybKViGxlmT1d7xOYzzSP8
HA1UBaHDAhS1+RtjfvO8KouBheg1L+LOjbZZWZJswaNxhepXDM0kRP0x7bfGqsiPK+NFzAA1vddQ
maIkkmikgm3AKP9RL6OQ3obpldx9xkoTvozCLxf2z+zekgssCIH9EKxky/zRavOBLXDRMmC+iisj
hMBIp4PVDcgmh3ATQMo7ej93/FDjG0cVMkz8zJtl549qHOoMcmeBYgqxmJR939uDo9OsNQPLGUfL
VtIrTsuSgUj7S5+JKfVzQUkjLsqmuFv8rAKUWGFFoDJrNeegGUwRr88gARrJ/ZXCubsiIng7bg5z
AhdDjIBrxRaR9r8gBX9eQN3d4ln6wxJfdPOmWxSRNQCQFy5hK5XOEeigot5LYaT1xFRrNQeCS4AH
RjXnqEj6PrrToxR6JsFoZrfyaHVGfc2AdAC+8LWNuJPcqjdit4Vrw11twB04/Vz55kcxW0DIee4d
hafEG2qsF6T3pOe4MX/J2iwDinG/aW9zyIy1H7RhlAXGtgu6vUiBg88mY1yOBgCiCCDdk6TzSndT
5POCw3SmpXyakk68sEgbBKv2EkHPom02F7x/madfdO6jJ3Iw3we5o8c9qlUUj8dLXiT0yjfriYF8
FBjkYOzrYE4PH8TOqrs/8GqgMLRk6km1vgbZalu0SPjBOMRIIyb1S2EMuBckeWFctnW/h8DrwRdd
EdMiWopLyoqJdGX9bxhf6jNoLlEC3ZYAXAl8SZOT59pMJgrvCUmQrhX3Q+qVj14evamj9cI24I1H
gf7y4H0PE8S39c7P6D8jE8uOXpI52kNRKBVd88OQdAhpmHSo/YzCXgwDsdzYeaI03f1ZHUgH3JlV
FDKajDRTG21+jeg8Cql8iL7U9oA1vwUEeE8fqHs576I975MctzfloiNc8sdqwtu0qikkqvRs/A0J
ex2JIyed5Eki4ZqZh3mpzCvxJdh5uGipRsYrFFsiAsBVzNjxq/Pl8yhukrtEG8ATrAgx1zNurXli
QftFlP0HdcX9wsBfC7tBVuBj8TZ/vZCtVCAlv9GGfeDWDD/ycWyBEqFW9I8pemzvajf8a4okOX4G
CIwt4/RUGoVijcGGq+ps/EZUcg1It6tjACk67YjSVdaiYRq03pzPn0WhkK2vc4Y+ULoD0Ri0XVp3
rIC6pWDgLxfIXWmACSb1OQ6NAB689IbQCOFOzHA69OADVOwlnwvrKva2uB+z2CJkswYwgrfiTVz9
Jf4nuWCnRkKF8Qdf0uaSP8LhYNdH2OL6DtC9vP7f94GKRHdAQZU8Fvbldf+ADrX3m/9q8NWzEQ0P
Qvrc3mFLMqMz8Tc8dNWmFmYeWDPo2lpOpPzfxJcTkd9hfHQs5zNSyWe2dcWks01Hnbze5WoH6gUY
KXC0bMaX31b84MhX5uf8aFtQuedowkaesCqAo377FvcxlfXyooi2ZfZZL2VgIa54Y3yLt5Jma6Lw
N/rQyrkJ/Ia7YDke+h74YaTvm/1Qjc5av2sdxUxG0g4onrH1s2+V6gQB1CRS0rBEYhSHlQWH/A/U
QLVJ1TBDvvLdbSaP6FkZFj0SHMq2r+wrpW2AeQXg+NX1ttXfjTZaCczZghxNGezFLKiYoQxT9Ktm
o2oyVwbBvX5SfhYe1s3T+uuqsspaUXPJfuoYMjb7kgOrMDyBpSl2v5uos8TQ8R7gSWuA+B73eLNo
z36x0S1E+KTNJBq+IUy4YUODaS+S3VJJ3DKG6q5eJdYBIVS0lQn7rHAqCSC26dTTcG2vDeu6cRva
phx+mmm7/rgMgwt2dPFvu+Qk/QgFmAR5fR7H0Ab9GJWLhdL/ryUYnwVL8fpmcQaZqoJ/XVHlhFpf
g5IYURUmq5CVE6dYzZKHuS63qW/I+U3hs3I3+WiHhCXxgykRcr3Pl8SHqG4hAQTTSeVlph6jABEh
/zXES2nJJEApGzWB9CxXVj7Pro5luPk1C8TrqkuRXh3AQEEIQSyv1QG1NGTN7Cb1hCB64FxwPtXK
JE/+xuKvZxKiLeKWvYulXR9lqcRsiIw7eEu2kKTiVQnAXPbiABekguqTayWebDll/T05bZneLJy8
lQw//LNKgVB1GlTC2NxUJXZ80CfDFNWKbjRx+ChNGDr12LGfECdOD8a/7LOdbtk1AdZgqG49wPCG
ZVHLEHrgj1ADnjBliCHlXvx6kTwdaUTM4vl/tjKTlqFL+H8eVA+WC/jgBSIC2Y+REyUkH+frbkst
hxmP1nIubUai+AE2eWMrD7Y/oxISH36v+EJ0GvEc8zVEXKchiAemUn78pFnpoGjopts+MjF2AkTO
NRVjaOKVj1Sx8caeQVbDQRXAjRSp64GlP/V0DG0VJ4SxPp10tGU7DMGWYNcJMYwPq94q1BwIE7cx
XUQxkSTRIuMQhLfckznRqDjDosObwTWt8+uyLEWUaMUqlFADvtBf6xRlaDhx2eLocTiNQ6nw7Jem
xortWDX6nNOy+J36uCGDR2UKnongd8AKNb+YtYGKcYqhDOwRyxFjb1dsFLOqPOQ8kp86Y6QqnSLG
0RkuB5oi+Wb3EWqS7tXc1P9gCy+FzixJrgvMqhO3PPOHhXcYAO8QLOzuvJlfCozBeJMos1CndG1m
nOKAOdzAeuMGDDyLh1gqsCZwNxfJQE83/bNdLb9/u78MaPlqMjmNTGZ0tHMp7IZEZMIqvj+8SOL5
RkjyKO8jkQlP1hIi6qbyv2RevzHK0gyapJTxb440BUbmn5MDa52XeQXEJhybluvIPCCA9uUubkqa
oS7KhGOT5UbUwxr25LnhG0Fq4EFW2e7WlJiRPNP+wbFq2Po/PMwN1GgjAPL9fNqNXx9nq8S8MbG+
6wCDgM5PtcJwZa0j5WtmW9kbypZp8HDevQ67UpKpgHsSoDwcqeaq7gCzw8ldnmKAxJ/SnU9FXMnq
BS8EjOM+5SYgRD9/a0ulg0BHSxg1itAr3ewu7oHsQ8OAv3PvuD/P/tc1zQRHj/edwjpdHINRqZv2
KZexx8GRNf9KALUMTgj1xg7ZNvDibYcN7MwYAPB5xQR0Jnc3/OWBQCxQe53yI+0LjOs5kHKdQNUP
KR8tDsbXr+mf783U+H4wic9QE4kCru475Qz2nhcCSIue3ByL5NEcWTci5PH0p1zr3ogmAT7hORk4
3hVorDN/EZz7/t5u6SxzlmaAmwllX7XmWNyuX9Zo5V4BxPThbcr3FzelDnfSSMFcGeDTPGSd79TI
vuPZJRSvfrBNIsNlGXcqKNOvlIUZbT3i6Ex7wr9NrshxXb2JfT05UY1MkBR34KMTuHRDEeDl1EJ1
8LeuQnZfgozc92qCSwltMNiybzTKLpuQiecRJVWCPgk/wM2WGGeyzeEsrmrgISEKyeU7XOnf7hLB
eHPjZC88/tmEaOh7IeZNiJ+L+IOg+QVVnCcYDpWF9OLtt/WnK3XU8A4GkkGY+peZxyu1GGniBOPw
buzaoX7zg0EjCAzZgwwOoTaw0cyz1lReygb2Px4/qKGqnp3fw4wFQQ1F8i9xTIwadKvLRJeWADJl
9gevj+p/rJiLxzaWrUs4KCVNMw096LIqKRTRja8DAWrFZOkrJWM6YYdhpuggaCpHVLN5V3GkiJuD
BgQ2ELLTyl0XH7xjOt8AOy5zGTf3M5D5UkHVOBFBIYEqeJMSyU7HF0J3npWVKGXN+JLhs1E3osdc
DUvYtFTPlF0tMMuUb7n2LFePBlx8XmSFjEiicYy7JHpmuP+EPU/h5q/LMFArvT55HO162MQdeChN
qeQOCSmklYpaVimWUs+c46tgGVRPdiNuoJnbaM6V2d3f9MlwsaM9Nf0ZW/j6tEnyLe9sK/YFKDzO
443uBwlExM8MtWYRBMS1axCDHQyCDq3bODCuiDSuQuO2cEMhJ/jAhpXhAmmKW3xDFzHSt5+OLAZr
Jl3xsqwKbTXqSqtyRvWBfnpsvioj/XO7t7wpJ5hTVYGrY4zuDmw7RKwGuLyV6MH5cZrwEalmwUxz
aYofVdQsqcfYBK8daln/zh+lJVR9q5WnIczG2r8V9OZ48iffaOjzL1xSXvmZQUgk9Up+vKhYjaHx
2gzavUmJv/BaYIFtji8Xd+d1j/l/GzCUFMmh3AxdXivX/z5YrmWFBXVcmtlDG7nzK9lBGLVp5fc/
WE/9tqQGz1Vfv3eIQYbsckOL4BrtCCg3yS7ynESFyLN5i8EXe7C6MLS1ccboeMFzjezE5d3g3Svp
Yxa/cLsRVZtY9is/gQVS6LOuVq8B3rlWghzBi+yYLyDYAch8F/u4rQldtN+LgN1x1xE+AeBFMY/4
nN66Rg6giqAa3kz8YD9rMje5GyulpfNtDeOqykwWd2i2jg9a5ZVw0gUfwJBw4huhZMHvmysbq8cO
lY7Dd/p3S6vo4WQ48G+mgXdScSIlavA9K1movrGj/D1zq+WLUlbqTrwZ6ChHsIuikfvUN0YfUy57
sz8EPwPswgsh2vb07QB/RyhaxSZ/Bvg8i+ovSZfba6UXDh5FrqGIv7sA1juWhghGddVd8t+Zr3PV
Q2xA7nNJYOqZkGtCmCpvs2V8gYSZNsvM9+jox/uhMizsQ7W+jiDbtQBhyetis5NtDq3TBiXPmy0L
pub0WKcM1hpzKpSPNGjmJTv7Sivhh+zzehgN/uBQyz05oJUXaLjSV3+xJRxqILsFXHgVj4nTpsgs
Nb7FBRztW1dmPes1p9FztMg3AQNpRbe2HKpLsupOPOgbrNTwTulr1QrFGlz5wabpz1oReNR73Th/
sCYNQukexE+CSu7pGQOLWEgLaqcTzTVygsuyDFFZCBKYXQ7rQa9TWuG+hfKQjig/0Y3NiXUkoKF+
oqm4TIjV5rdCyFf+RWLu7YKW9EtFjd59ZD0BAvsSX9rZK5/tGFGylP21SDXeWYMFZe4pnYyj0kdi
0TRdg3rebaUlYgJFOi034O3HT1TA1YdK692tUXceOYi0nU9Vhl+TANCodsJhYa0fs+uhL0Ecogt2
yZIIKquRJBVcIv7bEB5BqhgU7E6KRwonAhSyDhXeUvHfL9Ntkjv8+ApvtIWW0FLJ0XLYrAnAzliw
FyTMVu+S9fCfEOEvrneZvaNVrqirQDXcnbelcbqQfl3qjq2cRk7HfAcxKt6ibwVlMXbj8WVzrj6T
bAe496UPNAIoVykcegwwl3gHKAPbsBOXg0ixUc/hxqkBTWT2Gbze1M8tC/OZ314h+ghjwRyfBqB7
thlF/QjEbWgdx4zmWr+zmOkRrpIHLn+cRorMb5YjNWWTj3uQnBz18BJpmiN2nA3PVpeb7pjpZLmh
WAsg8TgvhFsEp4e0VVeWYHE6frahm8Dv8T5IRidD9057J55/d8ZZ73DflPj+W9oALVh4xkL/R8i4
9/K5qFSeYzASsWq9mCcgk9RkRvufxXdQ+SHSUduYIsdatQsDP58BN5xj9NveCo+Cy/EFtArbbDlb
no6PZQv1CbyjlCPPUg4yKzyPf9Snkt8PNlKvVyP3HRhKrvGVbSkyrHqIzUfrLS3Z/TFZq/P84DED
D/M+lYlnF9i+u3vWY/0aDgvVHP77HQmELWuO9Uzscagn09ixwq26EV0gB4OpH39mPU+/tMQsrSdi
C9CWTaziHfzJLJhrQUv0oRTMlP3szYDiC6y6kSTenEWt3gMVj8FWUOPB91sGQect2pWln4P9wpax
q6bXeyd4BEhbGedW5Dlrvl9bOcMNTys/PFloYE4pUOkbN2/ysoRpfun70tDU8IEHPBQ75URLAEky
W9iD50WME5kRjPYZEdE8W8cYeNOBgLeXF/X9Mk4qi+tNKhP8TU2EE44DF5RsVx6Lftdmxp+cNn+e
a+VyYlveqktRKls4BJPDMFjrMaMlV31qTMlzEg/jizdLU4r5SjgVlIbu+Kku5bxIBc8Sxwtk+snM
e1fSkQGe8VWmyXxtB6qVC3byZbhvEeQmfce/5ZNuUNDjxTjnZ3ES6HmdjUzjRQmXjmUlY0z9l2hF
UPlVLlz4AOamfgfCNXEPua6fOqCVoQCHSlmt+B/QL2UON+qeVKmLz8qcXLj0cJPXqbR/4QeZsnVn
avVEt51fo1O+3vTW9BdRJwTwZfE4v1YnciH23tHsm/CJ+T8nOOb9Kf4WHCj6qYZALHjxpiI/Smlu
hH+mdcwosA6fLOG2iWndjxIGu25o0OnPMNPuJmGkJfYbVp0kacOGiVfqBJiAyqZKNZ/XMdRhNMVF
wHS5DPaEuvJLqY+KI6yYvHLP+sDzK6FPleTAwhLViVIB6faMRNZG/ibhLSY+DOjjxByaJ3YngSkE
IuJR8yr7R1bBT54Fm+prxOSViH3Xf5/68FeFpfTdnZOZNHvrJC/wFl6OKNwQmiIwrAIW1d6G/maF
ORvQStCwJPtahOIchs0qpIjVGu+Oq1gGzGOAJZHvoOMp4O1vuRwOlXddaWZPrzm4WNvAcl39UiUq
/ks873HrUEH9nMoYqTvEVUhK1RA6ykqkfTlWXQZ1N+fEm7lRVHkGzhuQG3pu87ruekMSPcnAaaqN
FZXfCe1gutWUqjtgzXj6BMQ5acFgwfh+VAvWyli/F7Z7Ucf1aUsH32WwWiWQMuRPb1v08RU1VF9g
8foObci50z0sy0Umn8C/QakwJsoZvNhv6VSQQrQEGkZ3QKHcTY4vvq/7rqViw7nYdXJQ2ScLrQgH
RHXWrZhIugp5+puzOKAHTiIt8psvlhacZr7ans8horFnUMd/wFjXMYIGi+0poX2s4bqM9nqycqyk
hQ8FVylyAMhH0wPxMoRAMxtY4A1toGILJ0Q/bg87It5EPPtDqn2eB7NPCocbVjqrD9GZ09JqsQSp
98o2LZC7q/UvWKhPf31e30JgyARDUIZ5ut+2OSmINC5/2pb0U0ZEpsVIHv2dir1WjPHa3zAzHjYN
KeNnxGckhqte5KoC++KvLhgM8RzdD0WeNKP2wb6dHmSV/x+0DN98j0leaQO+soUrzFmkRnhh1Mpc
JqWX8H3dZIGyUppbW/CihmnmGu8Ln8R4tQCw9BgyXGqyqoMerdhBVn5+mV+0UVW4eba8SBkTyksW
NPnNGBMHDiQTZK5olQK7cqvxmByHj4Agzn1am+dQZTtMaTHcYqYNzRRkddBeIAPn7iRTaGPaFD4a
meePzp9rDJH2jtvEYHGIVUFzG691vP2RY7Z38uHrhPwfaG4F4+ruGNkDBsnDBXoWnBP1ptFIrrM4
hHZ5haB93ZNxCmtJcfNuhhkychAuBuX5jcMK20D0fFsCYlWUZdUgmHb7CuJSOcPFzLx3skmxTb1p
qHAUD6IPS5MaQ7fI7vk4D2MvI4Ivikv3JB2NEWH41exzTbmITSF9q8Yi+JhCJI29K3meyWft+//X
3ewukw25q1l3mgEszTAyZScC0ICaYFMMz+UHzZ5pi/dehYY+vE2C3ET19va1uO6a9YIZE+hY2nop
yQs1thsNZEv+gbBR3dQd2nEflkPlWNZM9Ou2kO7NOyCvCE6BmmTZfwh2B/tVe/UjMZF/yrh3goVG
94+LpUYSL2fsnqOcxisHk6QlwrW8VNhbB4KsOS0nXB8jag6MP/b/XZw+seVSiISunBSYcQ6STRJP
2uSEvtquf3/0jiPq6a7hg3826MebDSe4FsQXlknNRfSdeUzolouJ/xCSnXoeiEkFxuVRALJ1PURW
OP580SpiWONhZevszVY2YnmJbH6zTyihe0eurX7sWPrkKu0tXNFRtpuFJ70qkXMRJVYkkMqcwSYz
FCGmpf5VgDp4PeHIqgSQUkTu2TszD07uXbmT6ZE0oNK1AIzJ6DQTymwIR0hwR8tyEMBrviePoTgS
g5lsYUDTP98amFnHTjq0cvJ3Ir6NzFiDWZFHWYC+DxTZIpzPaBbopJYAKVZoXvSVOWNythZRY0BK
NI+slYwARp3l4MR/ay4ZLePyPkfq1ecEasbyEtoCbfxdpLo2HvSLI5Vp0v+aPt7RnmUX8M1gw/c/
G+gOiVmHiIzYazfk88zMn1Lh5LaQtn9ly+TVloAnguwXorjk1JqQbrJWkSGRsg2NTCWC9ne3s+d5
fVBwNv2Z9wQt3lvmn+f2shHuJKC6i2RRPMY7JxANPEYalnjC02D3BWt8C9B0RxeOIxlMEoz0gMZQ
7ybxto1Qlutuzp8RU4OMYY7/IXfnzyvVuoKqjS5F0eDDokh7cNz+OGqy/5RrurRvxw2r6wGmRBhm
MHLp9ZPgm47GRHCJqBMLw52qxJ7ZHgSF+YwjK6AgBK1bH781yrza+HBISOqmzm3IXGAUCMsT1sTr
kJkJc6paXPWjTx7nqgj+ndY864lv6FWMbj73I/hbffpe03ZtV9kjyoZD+fzt/zKbrVTNyCyQVN++
yYQBwkLEx2d7Ewtsgt1HO6g9RRbHkTqOSWhukf+QbdYFc99kG069h/E9f+jOlWw5qaS2UbzIca0I
tmh74GaqnBHO46/uMyeHmEW6pyB4E20+QPmolfT585RcN9zMwy9YMPPK44CEd8N6WgAdyEgoCZZO
AUdDlX98vUycrWvlEYAMeTCCEiD4AAbwM23qP6YLqLuhStlDdBg1GWwJH0TiO5SwbPThkZhpDiFE
2tYJ1NxJtYpqdRVsF4FSrhPRMl829d9T03xSQVv8oMAwZ5UVarrWNcjm1SvnDaymQkyxNTGQB2AI
J37a7IbxmoKtl9SN/lfbMcW+W5gcCXi5AN+berN2SgbS8ALx+NJabOpa/km8fMN8RnvGCoUURYqP
kMAlftqUcJsc/L+MGXC1tDWFz4muih0PVtVA+hKioNDLJJHRFflWPteXwNbLFHg5kH/b2lCvKqUU
uUks/wBG+rKWC0aF2YbSxOWAahfrdb+WMfQvKe0zNFg822udbhJIaIcVhwBaWUcsBWMTK6zwqovp
GqhR3IzdlSzHex8iVu/Z4J7kCX2YyQSbj6xgpViQKgIwjYQCYmMQDRDZqzcsOpNgSNDQNyGenUVX
R0A7rxkpM896+X+WUjcpG61HvoR0qIB6wbWbpscuLI9JBJEPQ9y/2KgO/eBWpFr8y9Nqie3wfSCO
Oyj4yhP5ltzyNkxGk6UczJFyEPoH33+MjtKutir4GiQP2OTupriDT3w5vL038UE8Mnsqqjn3pA1Y
eUCrL57hKbdk8I2z4d9RluzKDt+64pj8HBnJhrKNgF043GtMtLIc5lvvXWX2zG20AUDTqhg47wN+
VHVzX3N2ZU6dq1+IhIb+x/kgF0td8tmOqzH0O2VRe6uWBjqHzNFgybMazRHrrDcGT8BpY6lXmrl3
vsn/jv6eLt3PZI29zm7ecMp//VtbrEXLNuz9wUVrQqMnPxtctD2u4LhrMqhcLN5WSu0ObLcTP3ZZ
KaE0wpZL0M+zhL2AzjUPB+EDRm69NVOCV00GBkV+padetjN/UUO/w72GSIitQCCln2evHOVbCdhC
DHqqhjpVKPk7lZuBs600sTFegcnV/l3CTwEOFOuB35rqf17VmQ+SnKL3u1EC9q4F6hTrZKPqhX49
fHpJXf+6d4arzIipuoMmmAwAFboEIqUQ34vXNRqOByQMmjfua2uu/qADVztAQKJTZ9bLr8H12siu
sYT3qU+2VldrXqWXRXsrz6SQ6VIiGQ8HLPR/TbEAZrrDcEfDl5TN2zJ5z41v1cQPdOuSoW4+KJZS
A9oCT0tCQjkpAT6baLyt1/P2hAlg61lrjrAzL04M02Iiam2IGuz/5KTAO8eiH9JfQDwYj/1sl1Wo
DCAdxmCkva4NKrKrMqe5U4/cBBNvGydbao4nWYMP/e2NI3yAIdB0rt3n2i0byq/nnosjWqnjLaSn
j5A7f8YweapjRjXbeHfQsm7NStX55DLSwPfUdLnyHzQO2nspYRJy6En3heoRSHgvuCDRsC5WjWR4
/GRa3+nnC+X1R0j5YZYj3fv0fvGgx4BlJU62igF/+5EN76QYbpjCPKH7K3UxoZdWyD1FZd4/QsZR
Fl8iZh5U0KdoyZ4Z35GSF3J1ein4BL5AcKYG08p5jmFaW0cl8A+DDwauu5+pB3dt2q3D2DrfKhRA
/Mkp8DzRgF1C2tjE4Ut3fzR88savkXjePSc3FCNjbSwVNb8WBe6CO7pd1NYoA7+2DeIe2DKaGBIw
MqtTiWuZu87BAbybOYgOMs7lpZhSjJY/Mq/AlXyPd1ubKWeAq1iw0kb95s4at8L/a3faQtuQxv64
9Erqo77jJK825uYoO7EjdDNI9zP3Cm6gv0Ioaso7vPAJKBisX1s7u9LIZz8WycTJHXYmaC2uZXst
rPROR2hTRjSe9vvveesnjGzUd9mgoTFHYLed6fyVra9lIKF3r5otQM3uD9OKjA/LyVmkKds7yzId
7CZ9aJbDJoEi9n4ogE6Jm4Wv7vjFYpbC6myYPh1U0aaGM50RDnunc2CZ7mbzqETaRHTykmuaCPPZ
EETxzZfPgKXzr+yz+gewkqh2voazj4biqJ/Tg1xUmXGRi/i6NzbrBhRkulvLyE+7GNMICTcX6hqG
3WZDxzBWHq9LYFWWRY10E59m0/mwMaXbFrxH/2LeCWk7JA9SuMjiu4AszM5n7dLqzSBWTv86Z6T2
M88R2sOt9Cdiv1yRbcvXfsUsQ4mHS1zAS8k6lJHxuqoVfltO6TA7WCEVBZo40BZCKau8EG7IWfoi
2tB9UfNlZ9o4Q4A6/7GwE1dOC24B04BT+TM+Z4Yd3YpXvmQZuxqvKKzeckG7lmKr+v9Vv4ppHMg6
wprh8XCmzyfZR7vQ0Wo43IgYkLEWwOR+hFxo11VZsdSvY2Bz/b0ZkkZ+ue9uErmH8g+rT+KSw616
o1drwN0EHjcqbN8LEvwTXPLCNl68flBKCm5mKmq1A5mDJ/HJDvVSTZhaBE02qtzCbzUKFwbIZ5jy
lgKmk0036+6SrUykXY+1Z3/w3t0LxHTviIM8Qw/VFjKZEyOWnE+MdzW6RnPHfMnTbPPJUYIngHX4
lhH/LzHwtuHj0OeEcldPRZGZsa9wiX147FZTdkxm6/dCkUCwLvyFs391YA0L7HGi8dTP9ip/o0ct
ot3qQY0xEPwB0xyh4HJ6PtSI3KKWkLCcoEPErpBeSLgwAfXeemo9whf0boxcjES68s1gLnY7HbqD
zH52i14ScmXZIHTQFp+RKODVJQBgR35Ycey9qpAlamHtML8XNV7lQb6tMOXLK9NuxRhbBNqbyU4D
JGN2wlGlNwI6RSNRBQ37Sy3KZ0ER+K2gS8Gcwfsmzq7bC/4mKHLfnUDWDdFaDnJO/0xkq/WX6RRs
e0dzGYNeCBWP1dRws/xScvhHZU1A5lozNFOK1Ahvxs3uHPPcqNhZdkaPieEKlWsHsvBEEBy2JkLS
Q6p3/p6GOFv5zvrwV9liKx/+ezHFhpnGWUkxdf8BtuOwmSjtu1zpS06J/rgscW5W2xYxGbWXtVWi
UjfPbyHURMi6AzzbJukBXHXiPniH2gI7XR5lJT1HYoP4A19xIu0eJTz6/rgbqdnNz4mYVVhk+KGM
PJEuD5EJug3NITb0mvndLH8sa7rv20Z3LvYSlRe87Eu57QJbMVFcWwipbQm4pVmbBtrCbONgCi7C
10s1B2ugFQ4E9nJs5eEUrA2Ugt4ZrGpkxYrXo1GGcoXNQjcGb3PtqcKhCGbA2LFUOJwBTMyHpViD
V/kZk9cWNS3KyqkaQuVg3F5ejuBbO+gDQBUak4sLcuGqgU2jFubEgSGgQ5y5tWqUvgul09dhi72D
Z9QcR4JludB+WU9KTgOeEswYI4eXRE+CTqJzmtfs+PRGxHnegoFlpYJlBxRKam99sgJ2V4bOzdFU
Suh6RMUOHUJ7HXp2aKuvGjDUHRid9WxNMidFi4N5AE1RINhtO6lLZ7ttjDBEk17Tj0lQwIFZsu1y
QSr1nL+YNjr54qF6AyhuTjWwZASYSONXuwYhHjKKLBwgwdxWSYweIfOhfX9VUJ3Ql7Zrk6scE4do
z0MZ7rFibzYDuKCpKsSkXPU023G0Ud1dvgwj/WyHDyAXlpbsXjWLM8LEbnA2421cIdl688e4RPIq
cb38uACWm0vxLfIqbdZGkp0KWpz+AUxbpl1veWss6m9jR4s6Jz65IjFrggxjX/U+KMsW35BsbkZX
C+H26HKSxDJY13pl38nKI5V16jMtUHDMIebXzWK76FZuJDZ9qWYYGe7wUvIg03wIl0nQsZJMJcPo
uSp704kz2DiQM/JglFvmfifCNpd+qlFUznBqcV0bNQMdJumi5fhkM0ygUSOc0fhLBffvleTYFT1M
nJ/+mBx6fSM+dFKWoPHUoA9La/5hmQOSdH6ElwiBZoVButdkXEQkXEnZGPDn3nrCMJEm11wxLNfd
noqCJB6Z3Y57GRm+aPscB/6EOESdflz3FRSTujJBNmMFgFTrkdnIwCNzFwlG6Muy8V4ckd7lOQJX
F3dtLgUMGr+tn0BorwFTBJckJ9r8FImPOEuo9+d965B7pIGtRVFSl2NQDZvKj2vbY1D6B+gowhJ2
ztW6WQ6XDneICqYGf4BD3oK5l1yr/cUg8aKW68zuiL4cILzJfIOe02jdX1Y2cegYm8X7b3kFsR8t
l9mn7O65ftYYd2Zp3Wjo0RWNJrhbe7js3Eun3bQravWSxGvdMpMFiPP0zIeOeel4bRt0sbqL4AV3
SSvPbOloV/A49drWh5nuC+OIx3zowF1wSHqar+7tbX4MXOSe06JAXxicfBUuyNEx8tBFgqeI8TwT
+OaKBNsJ4xpmYX3c1U7WfqmvBYa93mRCiwMcbeL+xSPJ7we4gGD4Uj6Lci45YYG8gzYvTXhMbvjf
8T8sCaY31bKgJ42SMY5OMW4WJdOGTqSPuM2k7jMsMYnDuqsqP95llfLP/vWf/Q03jtxgr4n6Gi2K
MBEZMdiadO+DR2NcE5dCVNwqVTfX5r5+jND5212eUw9kiCxStOK9eI/apQWIGHtcWbDIcf1XeosJ
EtSwSb9yOXIkHvodvyOMGeCw4Op7UUd/Wp/+ZCZy+DVFIQ2ciXajjOjYGwssRdr4HpMWe909riaB
O6Xv9m/DLX6Irc5ai0iK7TxOPRqYEWBth4g3F6mk/+tQToX8Hp5hnCBl7mKGhKcTHX7iOv7yEf5e
ITrDdyQY86lLapVPAFmSq1f6UTk6vMPPohp/Pq+55he/JEFKnf0hntUQ4ZeSjqSKr7yZSwCZXcSw
Li9IIFdGctdUDPpzlaQooeX/SENZfvf+wqqD7C40p2ltUTfueFjr7xOLmBK4dpy67aO/ykwmhUBU
xKKgXzT/VEMNFGtPX1HjcDDT4LOcqQk41gBxjrxFfC5fwIiWJdzE+YWs8SXNmQsUf8b4fEZ8tP1N
e3pl4HLanfAn49ZexLXmkN/SoME/ygIy/mCt2K9C1TzhWaPfumqv7DfExNH6HkXVDJkqp5sNBh+o
wd4p8jRm7vGEf+gMq2juJQAwgPzXLhWUxyyVjjxTbZLjWAV9+RMOEShGoNs91FxhVF0xXCSEBRTJ
a8aDYp+PtFidHEB+rPrMYELoLNQA8bhGJ+mdwLOksK19HnJFJ1pQ0txjTXnkpnLWfTpLm7MVFnyp
37ujWUEFVcFrF9lEvEtjf/IF3rNYbRylYmB2oNBM6cmhL3z9C+WlJQNtxx49FxRzqqtHc83G2Oc+
Jsr4P0IjaJMNhS2C31imTUeCQUl+edqkMsNaTZOKS4fds6imWBPwomHS2hlAQJ5eFY64AYcpyuTs
cjYzAX/hj6dPpUQDT1VQtKmHsBp2O8LuFS0baULIaTMCnk8V9vbsGSB5UQnipS/wPEYfUxt/sW2d
GkE3f0d9pd6AYDoxXxxISnBS8vLypFwSQsFsxvPlnbqOELqMVyugqkh28FAMh5J9wHH25oz3Vf8Q
29DdYCAWbr95Hl7gOaRPQyZ3FTfI8phnxL/5ouAbx+ja9JUwAoYSHzWUJAq1RNWh7ZXWhaZWfQYJ
M5JzxVzF9vwrn9+jMuh2jRbMF4Pg0A31a4wQQwi2/kqdyH0GckxdI6BYPx8G3/EQCHvv9xYXD+xt
5NBP+PyO9I438a7u/kOw8a4HqMBSj65FxQARAkl/8Q0ftxDe2/DyeIz1jnr6rjPZtLLOHP1sKIjK
nT0EJlz/1qfQ2pcAExkGYLzmODVEmD+NcUDB4/bXu5+B6PjliCbdi6ycUbDtbECCnXRRKzEden86
8H94g2qdYE41QjCjMBiYg16CSr/4q5ECPulcz0LFMrv+O3uvac/ULIWK+8ULzE4FGjKa3WS6OOox
iNVbtlU0te82gte+ilOa8atluhC8qke7W4Ls4YJIq79MupLZbQ2Rh3EhdbBA4f3uTQO1W58g6gVE
j8aFo2I8L2Ot2xQ52SilEY/zGhnmnQ0e57LMMBGrL+qV6UwM+Sl0OKnOkcd0m8OYdFBkogMmAhCA
Smbn48CvOyX87dBET1ViHhFLy4+PPkH8ogN7VmrGSTcACoRQJaYmU8OlcG2owPXAuQoZde8u2nLY
sUHDLdD8l8HvpIOGfUsM0cs5d5X7UGazcTPo1s18IYr/9tR7TmIORqLFwrTveWkjPQid9aUD4LTz
rwmGrIgRHUBsYfbQc8ZnFxqyzbJA/B7gPFHg0jKvUP2jAsupF+N/6f9JECNHcCOevoiEh9Phv/1j
CEhESt1ZvhlROI+U2aYE1L6erE3e5+QPq8QpW0Xl+nJj62eHFq7s6FNJ8trTK0JcVTmdrQW/7wpb
UYGu9Z4rltkTyp0G0NSRYQ9NnANVn326uzE8LFUCynXGtskPqEohNTzhxZwiEYKULdjzGCUnZkIr
AUGU2dKc2ZMxTpVgZiSZWf4FgD8Cot4n11TfFaGmYiQdZfzhUEFdezBIOaSGHlZvi1BfMwMvPtHi
KuK087Bzgpw5ZYKHDv35sbT23NrJ6ivx0nnlAzqc9TGhatJg9r7RFRxzBphD8uYf5F+adM7j9oF7
vcMgrTNli3qZlpv1L5KGyOxfEG0tQPfAjvha4nY1xIhqQd1gDEvEVCpzb3LcXJ0WldZQx9IF8jXU
6TIc9ogiAltTzM6ouG46SHK/77e7ivRlyVvmYvOdE1gH2SlIGt/2jDqSyQVPlRG5Dhjum0m0WsDK
0NeIbHZozjH4AdAWC8VLzEUE0+w/XgymxpyIEgU2fQkY3m7ezGQ8IneDF1UuKR3RDfE1XR3Q12Es
7bad86pwa+DStx5jSK0mDIX7K47PuMT/6YTKyQOQPkjdQ83e3buQPtkUnB6s7h/aFQFvCHHIT7N6
CxtnWTJbRPwmaxGKU9YNhED+bu3QYmuJ8IUzmP8jCvqU5QUl6CU2tgRUiu4wlmEYMaz/2VCHqYs0
QaBKXfaZRyAUNpR/aK1X6aI1kTHV6V3KxN8ibEeosEIeIzmZPlrCyP3qzhjbhaUfDYr+q4gKHYPw
Kof2Ct9wq3z+gMpqs5CRkI0geNFyKY01mUPtpMbv6IHO1cWIz05rRo6p0nSbrRhz3cOeDetvbfGm
cGr1gIQ463bxCKClRGAdHf+2FA7bU/E3P2rQomomBBlKebuG+Lr4B3yLP/gw4pAjme6/GfEoWMze
VlNjoGhR4TppgfWR/IlgsTFpumKgFRqqSvlxDOXzg0MnOD3EeJcXB0CZRG/imBPH6OrN+JATe/zZ
5hWxQY1/osUfks38e7geatnzIRPjk/7RKcZ3d14L8XtExmmhf7Wqgj/mjiApDoModlzzbx+QoJXe
SkL8OFGXpP83taw4fcaDceGzb+CpTU5YH41/iNFDUDx6Z+8osexw4cmu/0NM1sPipuMBSzXV2ny9
9lVYLcq7lJDj9UWJKADXqYnS/XS9CqtCo1IrqPZmMIk2jNtykIhZuf+LcvHVPGoiHddjN4tlyqW1
XmUemaroXC3WWmb/wbQg/s507GQd7p6Wu2fuV5U2tUdtEY/PW4RbAyjfOQLilfIYxhBCNoU6QLNg
7yYQ7MKUgW+vCPW53DkRbntxkzk3ABE1n5AOyXgp7AhoqP0I/1mmiWy+l/ToJ3WJjXiLYRKfZCdd
cXqscDe6inO2MsTQF6RTtMSnisVW9+wxQz8C8GCm2iDBK0ONjZOO/2dfV/DA1GVAfw+59Go706ob
TqOk9179Wmd0TOBS0bziIK8MdDXSGpDnMLimm3a2rRI0CJ2bo0E8N/ZNtGgqpoEkytqhLO//YQeu
wCj11LpJzxz8Pb/JFfseERpEmtBaZudukfWtQShWX0qeKMqTCtfGIoLhDVLWMgYWpOT3wv+XykLf
Qq2f6kc/VaI+LKabLBIeHiTrCRdvgUp8Vu1OoTEOVZO5yduFFmwZlMEHbXvBNMKE5fKJ9M4rf9QM
+yeJutTRzwsul8uHxplxSsXoPdRXAfk0wpVibec6t0bADxak2BXfHkveI1Sr7clITr/WULPgSZxp
iV1E5KXn+3q+XA5Czsr4KI/VC9vMXN4N7ntWFbVoOn4c6ebATEqZSO+olpSFHWTqpzDPOnkySM68
MB3lXIMbUoLGvcEcPe6Ws48/9X2YMNPvSf6RmDA3dO0mEXi+TgL7gy78G/3XDgQYCDFfofLz8Nsi
6Cfkgyd5AEb6jFnQi25ygfc1FTTvlHPrBDtC8neVn9CLD82A5UaGgMEqa+YMM5pJkdrXL7hyCWp7
GYcE6mtAQRhMzjucQxmjZAcP874HDGvdGSye5MrL8HKi1Ddw1ZUCarNbf0ImsDB78baUJO0J5VIb
R4q4E/Xml2/ucP0Ch4p0zWhulC6qb9gevJqTLCy/X6AipmNhwrvoEjD55MWPF9O71b79gwBv2cKA
/Hm/stA/iGnxeMJpKtCfw9wAMXMQ9t4kWofADhe1HMsvXDPbXg5LFDkbAq2bEGpkLeLX0CFEK9C+
0pPo4omc6iSt16OIZHzuMM/gvAriA3MW7e4655ggE3zd4wOLbw9ZhY6GgnHAwz1vCh6KlBp32Lz+
5wI8ec10PKzOSruHax6hoQCNfnv15jRFoFCylRThZkPf9hWTbVgzKro0Cp7G4KBgTvdHnS1inSZA
X7yDQfFkQ/dZzbYMy5XKNuQ8l+jsCyvIl1lGOnxLaNc3wLChT+EPFrwoYKGYZRZy8m9/55+oQ5FJ
hDb9zii1o0VxTaLcnOhqxITsKtwZ9EfwNrtMZspVzY0QQJ6Q5g0o7SwoqxEAa2onTnDjLTPgNutu
IArNgCUHQf3fYGRINU7kcFNwo9+8+TABllj96jkZVN+XLe6CtmNY9Xdewe5yVWz4w21UAhgJp43s
pG6s8/gHRXmLGwTBJQraq7GiT0tqOL6UqKsYcyQ+TceW/yZxHBkVHdt2xzR5Lf0HNC3prfzT1KHt
YPRy+AAomo1R1qCVUE7HTiF1/hwD7CRmP/z207oMrmkSc8OE9jC5Q5755ir0UnLwRKVOl/J1O0AU
LnqCwlyzJrEozBLHX9der8Uf42eOu5UR8VungV2RAoWGVFBbQAri4TTbXXsqmw/B1/70ODcarIFE
Vc7hZ42Tm0LKcGMWGRfFC/0ipNcPJz19zTvl1+1pkcSyhsEmMdvrYGYqAxYoLKL5TdTdKnjjtElP
SJCnrxc0et9KQE8IokD4Pg6wVXoEM3YN7TCLMgLBX3I6pflz0dZLijgFI4llRwveiSXm6kuxLjvO
RnfpEypKzjHmK9Gq3YlDQoxGERau5BAVbzRL/+Dk+MFGmL8QrLco9nJXx/22VpgdC2cUcxtrk5ZJ
OM2t7lMZtKA9UFQ+hbd1R1cC4UNlmXVtoUpzBAoJ+WXFCibWyq3D6n7ih50y/PGppcmLBV2lLMEt
2knL2JJ1GFCRjQHk3FyR4D90T2yxCMfjELSH3CnrfwkCEkhb67KxsJ0f9LZSU4/LSzKZgJqJSrE2
BXMRT1zvTXb1JXUTJwaN6aQzygZ5gQjf/hjK0TSFH3TW9bYR+zZCaBhw1rHCddv3CAn5q2yafFJj
aFPcK1Wvl1qoN+mtjRW1nUqGr9bacyrf1UmgwfZQDOJ0+v8bylXktFMwve8G9ZLk/j3n1ezTXe2k
ejeBdKpDgOBSwyvG8zsdLQo48kjNIreGl6GG1igOi0KwWM55D9bD4wllpywn3IjHsZeCBdoI29ig
CR3q3hVyKsWvlM33DtGBKZ+yhEBUWTf1R/thTm28vxtWiKD4/5u6+c0G2TRQSSdM6sLPqWYYW9tZ
8QIQ8Lx3hpUOIgIphgMr2+PYXpD6y7dguf2prTlRLc3Iy4RQyL+GGDQvJSPC0/mr/RCGRsIQ/w7D
QBdNWa7czloEkC0jM+eUncPVDzK6VNs0IVUtihFXWddz95grBwTaAyJOQ7iCAVEnmaFFNbxtHuSV
B9by9vgmLo+uLRUfOx10vv7wgwRp0U8qtu6ibIsdcAWuU8Pjhsly+cvLCJKt8ZDY+ExoLsWghKaI
URXjLnmrlqjpCPgv43I59t9NYcwfEN6/OqUwERqF5N1txn7NxTVnP+L3oPKjJlXtqg50aabI9Pel
Uo6WqmK1fSvm0ujWpaoBr6lR1qUFNUdeVdiEZdhPT9CBelYX68w13OSwvvPueDenl6ubCJsXMbOI
HKCmqxSDzqOpkZTuelV7h9J84IphitRUDPo0wa2RvfF+Zi3LeonV1ew6tW/R6BykcdYZ6KDlmCm8
RwLjPi6fYigZPPU04VOTnY6urCNfcXxbRtUe0I7OtA6ZK5eVHxUSXM6kSPfTjb81ZA4UtCKG62UK
lG9SwADZoEwMxY6jbWqitElAQqQuooGPgOPuEUpr4gJiLTzCpS+jiHttErqrc6maaP+on5MFRaxJ
VOP5d8mebc8grec9/UIPM4o3/qv/mKOZjPop+YgnRHRd8Lvqg3rRNXhPHS+1hJWkskoppaKoudAE
1hq3NWy9JkNPvQ2vQ4aIbZ2jygL468G+3slUMqE3DOozyyZxiXp82XX6WpVJFVshrnq3GGcXBQad
fw5LKt219MBYW8w8qQxCHcUrbYvcWsamoqELj3jHLOvak5QhY54cr01AZFGnQoI2LICX7pWc+gK2
Urj/NWGz5PWu81nTzspEPzOqIp+7z1+hB8cYgwQ3c9lH6NF4J6i/g97+EOZ3RcOmFr/NecG6vIAb
ai284ERkyhPJoRgFlgtno1IBaeeWiBOdv3w2j+1v45p5S44d5j/I//4hjKRsEipHUepeZYrOZBMK
P7d/38G8AhIdhS7/nVcIZYOjsUQJgVKv1cruZJMeYioe+odZINpZ5zAwEnvN+d4I9MlkO66Cf/yC
SdvHLlv9I2K+kr/AAG7dBBzCv7mgdTf8/0PSF+moET8utUSwsNnvDcWn3PSwytGJCdDKR1kQ9xqS
Vrvyt+rx0H0kYYI2PJGTo7HX2S6svjrfd47OOtyFktOfwFtoxdvH6I3P2Z7kYOYgNBhNzYICPgLY
gmSMJ8LfM/apBLrfGPKnHcoB1RtzB6F+dOd5goMyzEvLKI7UkyFUAtgiCSisCBIU6tYzaZ6UFZX1
nkvjHJykxCGjCbVPj6KJF7fdaVVTD2RjGWTvSs1fciMSRskoosc0nzxCDAc0mf9JzSLThXa7VBXl
I4cCW+acjd7dJVO3jyDPBaAfvfEGU1xaboQ5rT8bA4o6Qrl7ql9FHAsugluNeicO6GQSIMkwZaZR
6SScLnGVX+dX5UD49osqiuQTYrgD1DfaGMJo1RCtXVYOKp9LtfcLjzJvXbqEr9oWoEv6QuaYWM91
blQz/P4YQkm/GrSOAGFCZWjmBfEMryMo+nvCcYZT5GSzebA+sCK+eqEviAfCEJ4BP8OjmO2qPUSR
08We7DwmvYP4JZNm1jb6cJfbce8guKqJ/9YdX9T/vru5knZx38Lh7S1fpkQze/UdK1ZGHiLSip1E
zBsQtir8ZOxS8eP3Lr967/e/D5l+hq+kgQfyu/ivNsql78X2BoD/spdQUzxt6QXPvxQZWF3obUf2
fLvv+Qzl1Dd1WIS6CQ6icVdIEq8wqBoOiL0Iuz8lYyd8yLo7Mev2PXLdySI/mVf37jM3nSys4p9V
b+CP1IcnXg9yofZOSIPDJdWVzksNlmThcC8jxFyCr17KV3Ezsqxku59YG6n8opx7qWPrdTB4K0DJ
cWfPoegZnxTiUTJWXuQ9cveZzIND7v3Q2dS49ANRrhs5ay1upwP/5ywxq10j2RSdSxv8cKcEgIax
OmMyHcVR4iyoR3cDqi6cXKZIhXc/1/sVc1bwYK2F2ocrpmRDEykWy3U0P6poGg+KgLi//2+RahxL
Vrc8GDA2hQO/+NT5zbGQbtHvur4uqQmY8ZQdOYBPhMpKHkXrUe1/HAaiWoVJBo2AY87veksFeMrG
E+P9AGreBIvOrBdQnMUP9B5xOAEe55/ZkfvsE3jrLM5EJmk9mhmm4vtcbEymZHLt1xRVvBnUSrqv
HUoAy7Jl2Bzc82JstxqBlM9NlMcCQdHvQh4owM6y5Atw1wEKMbGe5VF8OW7Rj/CTbVWBWOyTzYlW
Xvff+9bywVbr3YBqYDDZ/VGjpBYT7bKEuBlyQb+icxziyJATbcA2Kz7V7+JnstKSMkXjyvKQWEwY
W9npxq264aRUKrxdO4W4AqkL+yqDpoL7d76ci5rdu0YXtsZtTFQCKHRM7Oc96Nl7zIjNGWBCG01d
WFW/DY3iJYUnlo4HKMgyQJwkKnBHwRRfeOexo3ONmmGF5H60E0M4VBYSvO4T0Hk7Y0gYfwvMB2sI
qq6lUZvpbuPBLn0OjNkzTsbfu8mgdUIJIeCg89K1lcxFE0l/Hq2NEJhzcgVn+zD2kQdcyGt7e7WP
Gc2D5UufHoPgOd0for2p0kwKZMRzui5i5a9D/dXZq5D9X3Xm01DCVFvT/nIGsV50Lic/5Ylwlht4
bA5mXJEstNLNARbDrs2nSRFznGbH+q/rNn8HSz6S/R0Zh5HtLUUxyK8FnwrfXcXJVbDVN12R8pup
y9FOmpP8WYjKYQJhfKl/R6OSmG3xzFHiisG/x9JdsrciKiLornOovpCJxpzFP0XZKcb/pPYYB5jo
WbMyJVKTxVxaJpN9fWj6tGTzVL9t/Hzxl6D0YBv3snvgwsI22xAdzi2kAN4lOg20aPGXIATwvEUk
BTXbccgXbIYg/YXPO0cMyMZTo8vFZJK8s/5CVKnxlzAkaYxl0Ct/V1RbxbdRu1OpbEd2asYE9ZEr
U3xdJrOEgUsAmeIpirS7kFx9cHejQ5c2Z4R+9eLVPseNU8CG5DrK30EOpE1fy8FPLCU7hwjiXsko
nOmztrJsIP2Vo/o6OkPvnm+HygrUq38EKoJO3pst/f8+1/yUX+r/1CmJHVHABgwdqqnweqYHPRx8
cGWWwwh/z5C9vurAoJpGwYwTYriWGxcumWo/+ahkS5Iy42KPaecXw8CCw8nSApTGV6eI63rVkqcE
T5BBoRjEGlZ/asnvnh5Oo7/OdzAC0GmjDC8uLC/8vKyk1DecqY7wMd7rmLJojeed4O92wI6gxbGJ
vMzkEhq7GR5fp3AbBQoQjMdDC4Q8NzKl7wRRnIbcnLp9z6a+8t7YvMIywRiCQ1sszJ7z7KbRmZ4H
XHAV/v2HsZ8MeQE71JtTCAClbjRmo6eij/zPIriAUS4RJaAeBBukSzQA3McGvsWNCz3vInGjM/b2
q4ZCYeUGCQzGFza2aiI5GFecLkid5TgXikYuAXUBw26b5XZwgPvdO311AY0sKQhCZRIFENFCzjqZ
yYpmvXeIIfRPL63zimbpGYK1yFTw+zzUgtXwEmZ618b6AzkOxYuJen9sGgMRVwvLytAlN2FI1GWD
6+ryDssyNnoxC4Hwx0RBtnxHGT0IvD6gv/iiJjnM2XAzSc0ghd+k1zDsgGJuToABeLZ5CHSAUg3u
kYg4e0k5HfMmcyFFTGb8XWRzwNLfrlzrvVoDWRgiCqoBUMFSbllMih1EfALHL4atfIEermFSqRLx
LnqsUabv3/2v9Ipkk1q/h2GY/Ha37ba3CJJrpJFGjKSVP2wWXDzLPPvzWc2DTj7oZ6fwMZFv7HTC
MsycnOjfp6bYDN67UXr+Pu+5pFIWBbQxqInZ95YqRZpeeAhXrI8nwf5tK+l/rqbaMeJLOTgROSJg
SIyKmqSLNpPAgHH58nXhJIk524QJHY3HDdcupNugHgSoRWj4Bfol7at5iNVpcLUlYr5ll8jfJn91
oX9u3zAGKxhQkPt8hsjKwQQtglUjXZa/LZz7TgxlE2pYFqyIHgeFr5T/cmjruIoUQWMvjbnuPw1I
ga78vY9OCB0DCiJVO7tA927AYS7w5mmgtL1IwuQKCx+DV44bxMuow4B5BQrQ6clGgxWCY56M7Y51
Nq5TIXSW4EqZUP+4U1AZ4+NAo3Ha7L03BtT+z9+IFT8+i1hACOcpzwYZd/WGIUdOHfHYsiIAqS9j
JIkme7C+QOztT+zxCvy5i1TIhENDQzDLBYE3dY1cvlz0p8+Um5bds7ytdo8dNu4VdzdmPzwDqp18
an2W4krddVFLp9rv++jBVjMrHKugwFb5YS2o6jZ95YJiplOpH5tecom1F7/ah+JaNjtRDO56O7Jx
+ZO5vni+EssD6b0ENiA5jgS+Tu8bnx1VqYm3RGRpay6klZ/9JRNL5OsgdN/AP2WQ0HXLgvrzsJIN
zWPosH3HID8RTr6OfntCuMXUA331fH9OE/dYUsHDegWg2rDjDyvi21S1oI4LuINQIPM3PtFKLEyt
GGNAgxGnJKKB1W9Vq1whzBiHF24tKvYYLHROz63uBgkvUi7bc/CTybQNIu2o5jzBgzyXg2mLrUwV
swGOXG9b6kUCjvUQhuQi311IwHVXn8O5uDWcAvcVbDLRAQ6VHRyVOkHTYtPIXjoCuE4ylWlZgznp
eQlfuxKX8tyGWy1ik7hZi+FuTAsbtFzQC1ioQaSA5w0xfStNbmM6aY6BjcG2gAjnoq0mmPAYVqZ6
JpVSxlGpz/NIg2w6bLLyxlaJi1kKMhasRMqFft3taOt1R9fYWlFtcRWcpzErCcaYNzPT/RbLYJ1E
xBFMAZIzc7UixEWEiBywTk/dR/SkE1IYVYEStzozRr6PEk2vdq5YqH/rM/No7j9T2sDbIQQzNB4c
JDWctirR+JRztP+9lE2PGGWR2EXJmuKLaoQlZawAcir8ztUWMQLNj7EXyVYoU416KjqKXla8UbZ4
BCuyqWKhiK/U2IJo/5NEuNa3930a2PwAbqLMouX0oj2fQxYAI6lxdD8UE6SCddLHc2YyqytiXjwa
IOVb0apkk02w3ZGH8gmivYcCD5RjLxv5rjFsX/liA4MaSqsCXuZ0IKBFXaGLIrQOjzXijkQo21wm
qiXwlUsLtdH88KE1t0kWTZ9W6JKzdjAsNDbz+xdSKoLwKdymyr0yOzL72/+8tzBuhTAHd0KA7p6p
9VkxovHqkPzXCnOTTmAqa9QhClmycKv/GPX6v25McI3WneZkUeg9SM5awgSAr0lK0pA3swmgHRrB
/hIlto5iixxncDeq2xykPh1wIAKjZulgZr1wln7EuCckaI8UBaKesXNt3lJvobBTSiy5L5OYxPAx
GKJ131aYcxXSjaRowvRxRD+TwEgatafrT1mpBgyHarjx56ZkNCvyaOSkXNzeTA+HRl+UfCY22b/W
ANAqG7JQZPMT/kXRq7yALTHvda3va2B0UItmlxGD+JU0g2yI3dhctK/bkog5oBAWveik8UcrH2p7
k7dJ0z4WdfESZbLQuajb13C1JjJ1RJfG50ZCAdO3lkLj6+x2SRFVF+vRHLG9GzulYPqkpFR4/2fn
m6gmP0xEq409J+MyXlAdyner7Wetu9sOyAWYsT5m+3G9ncg3G4BOwhxzw80QO7jQ1sEI5IT5BA2o
3eNRuAc8kcRzLtX9I8n7X0xfH/eFYjnMU9bOJdmttDbv2WqC4Obj95ne1RClJ1vaXMDZd1jayHU2
UGaIh9NvjJBGX6q/0K4FYtVNIdi9dkmzqvEgXKZqqDeNprTUWy1LptgBSaTpAWRdfcIci5FrHjBk
UNTEo1/BB+sPf8y9v9XU2Awna2zNwahd8OntteHHPMxhPsasSKRpd8eSjzfV7r5u2pjOAbu3d4kS
GfHK/KQH6FG8cXQEmzKlGKXVLnPaXW5GfmZ4bMJ6zCWAI5RbTI6F5nEz2wHv8YPeviwowIZcobHm
jFEI4sW4jotseklch+to9/+1nGwmXryiesSsLYD1Tjc3HEWyywZD5CpnqLmnO3Zmv2ipV0ynQYlR
aDU5Zts6ID7tcav0S5yvonSReBcKbVhFTr7Is2ASY1Roj2j9FAT2QwH1WpDHx35VDO9ePOeku9iB
wsiM/V8osl/KbEFp9gOvRh9Jvfg+iNaqJae4+YDcTsxlln72ScozoMDNk092Wszjq4PAkn0h3+GX
CnfDi+5yVR8XWyLmSSrk3LbQyCqka1NZrXGbxtJ3BUFzKQVzz45nehWqr3kfWUOeUp/jbQlXDEGW
g8ZwksZFjCCR774c+Boag2zm6eNaydSQHlsUCz2/OyFyfLhiCEr+bwI4geS07/1UODuc82ZnGLcj
EJtctq/uUQ1zeo0VTpd0v9c/87oe8dHOw6kk1Rz0v1QK8PauWXF8+KKYBq7j2SXmxQruIuhtlUbo
+A+LnQc1SHUzTtSVuYctnHAOAYfEFVzabuNROAEz+sEhWJQHYJfXDfllv+pW62Wjq//sBjLiVCX9
zoTRRIcCfdXtIG1pcyVI4JuKAbil6OVIl5oby2dH4oX2A+inyxZkkw1dmw+z8+ErPxchc58tsum8
fEknl7qP+Qo0UCsQUOCVrub8J+bdRhqC0N1BhA6VtOUXyXFslAfkTsgaHEFSVMOJpVBOOViuBL/Z
K5fO4Vz8k75Q3TPWyI/3flVltK/g9k/q493FZV+3dy4Rtpya3axXpTe50iYlbYAKOMqWeJ8496ga
nxaE9rpf5o4ZMIkZr14Iu0HUWE7bB5GvYRdJt0eKPc3xN1Uy2XQTCIgbqlcD0uS4qxf2A0gfQ2Rs
lM/TzZdkGVkSrPMZ4oTrWnS8qXg/gbmomEbr+9/jBU3Qrp1vj/crIELU7GBxOvAc887agcZhgt24
PntcIXK0etLCuQ4xcE4m5hUJDU6DPnrIVdXdUypcS6h81w0wPkK2PhllkeUndguzTw0gLzxTGOuO
lehTugX28lgPJ+ROw7r+7Gdg8QGJXxZEh8LbIbHkpcD2J8EL+RFkKN14yY4NkTdN1YVohgF+JWlH
CALHm0SKEyUfqvSifP1VZ5IHVvYAxxpqx3ZPSFYTNq7VUi40hgXELjqsQK9ephVkQurzZ0CmHZHN
yUln3jjKTbH80i9iDBQiWMYa12FInjlnYNM9nIO9kIeLYruY7x/A2YhmagZtFBx8u8XVABA9HyVm
ojVDUgC3JDXEj67lSqPCIGtQ40iBijh57ej/e8YcLAsI06BT08EKj/b1vu3N+fNrEE+7z5zBTvOZ
0daMQuwpxRoPmFwJ5w7pzTr7oDx5myvajMKU9pdSeh2h3KPJPQWTF3aUzr61JRjQQWdw+blRaWYk
yFL+Om/m78ay55zImFcum7AKdBGZpa4Md844nog6MR+LNUDm/eJF2bwNAFIUZ5sUezB1Ml8Mgn+z
dnN4EYdUX+VzM7GirPqVIhtm2xQoPjXmm+CGm86frqSg3WVMv1QyrGEWDAQkZpFzZLAwLHGLXrw8
pyNWM+YzsQFlcflvnbPyGzF759M6/os0dc7+AUpPzGHje8KQ17l+G7hxvc/etmsRfoaf/vy+ROPB
Im4jwM7EGS5/BRplB3mfF7khQlE69GT+63xPoFvNLeiph/r+4TUygckqkx1PcR577Zm8D05VUWxo
voGVcj3ND9aFP4tzWQL7xaHPvRXpjNnSRu0SbIlixEUa064fCw07ZMZS0oOneE73EXCzd+XBbdGT
A4z5xiTwTYuiWB8l9IqSF+YHTtET2OG7CU01Kqe+rumOw3/3eds9Hm5qAHoyygZ97Dot++hreFV+
L6vs27KAXuWPXhwjapIAXBpnibpW
`pragma protect end_protected
