��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_�z�
�Ã�	w�YQ�ǁ��t���70p(+c�g�'9k.�H�6B(�)�d�y�{�3z�o�(����s�	>R�i�%h�[�>(��ٰ2��{W��M���xO��}&�6}SS��t��Ā�r8Ľ�A��JlB��7RvH]�7=��S[��)=�fm .ȴc�(b_q�m��;��2ʫ�]���)c����׏e�F�,J�BMc�ߙP�덳�
Q��AW�� :5�;��u1��+#��H��	�?���8��	�x���o ������f��6@�۠�V�SS�؝��a��vy�7��ݱ*X�#I{�6�O��uTY�#%0}�v�u�vC�t��!�DH���)�TEf|�n�Z��'[.�D"
dkz�A�	�4��*S{_���� qE�j�S|�pL��
�J��,���Se#��M*��2I�#�ۇr�"r�N D�. O��(�ҫ��F��|����rQD� ��aS/|�c>��Krr�i5_��� �h��p� ���%����,��@���v�y��'ݼ� ���g
q���De�x8C9��J����^���A<�0���ZT�8�S�L��@������7mt��G=ꠎ��_�e/L`	A�C�DT�@���>F??��t�4�'�q�m�;��L]���+��d'�f��5�a�
{=W��(w�S�"��tmA��ҦA{IYj��8�Ff�:)pe��i�����ȓr?wQx���6��l�r,��3�WNNW�����Ώ���I
<���@w�ގךy�4����R'�E�b�y�Nԛ���h#�?ڡ댷=��yK���_��	A(\���*[�.}�g��#e�j������P��y~L�$v{i����#ǟt_߶��^<Z�T�����ǔ��������U�)�@E`�P�9��uy�S���L>�� ����?q�<�b�GZ������;�L��l̐N��D���9�z︺��
�<�������N+MiCi���8�v3!��5�%�I#�W���-�Γ���IZ�H�;�x�Hq�MS��Zg�R�w��橽��%���Q��i�}Y���L^6�z�]�gU���a���Q�9ɑ�?��=�H.��?uj&����6v�ۅ��^
�R��f"ھ8)Ǝ����ӭ���� �xZy��h>�8��	Ͳ��m�s�l5���I������P��1Q�6�<�E�dϋ���:7"[�ͦ�~:@�,��n�y *Lm���}���˪U�d����3�q�������B/��kyt>��&g�/(�N�J3
W�a����K�fU��#���š��UZ�8<ڭ��hwJ�9�I�~P���������ԝ����$T��4Ȭ>���`��s�c�\���PK"c&+��4�;�	Z�)W��mD��1 ���X�=�TS`�qS���oЈ7��t�sPkm�e� ���Oy�dQZ���`jo��V����p�r!0ΌQKY�U偀" [4�c�oA��m�L��/�S}7o5�S��<�,n��W-�X��Jj|�01�5� ����s�xjj�-��cX�4�H�>��y�
��͑ӧ�֑qO@�`'��a�%.��h3�P]��HT�Y��*X<E��V�E�vi-�|���t���:�S<S���D�Gg�s�x��.�\fc#2a�ÊY-4c*m5z�R��B:��`Ǟ�X�*�W��H�ڥ,�<���Nuy��Ij�y�<w�҃�"z[��~.
U|`E?�r�� ��6[������~�dIm���p�^.�O51��k+n�Հ�Dw�Hs��WV	��HИV��0Id���p&��y�7C�h��e�*�C�E'��v���ZsUm���g>DJ�P���#������#��;�pHV�O���Q�X�C�kWe�����2��a����DE���ƶ�r�zO�g��~O���i�ҭ4��G�m��H>���LY`�9��ӣ�9>�����<���W��o��Yw��u�!��g!��{G3#�N�nBKR^>v�Ҋ�*)��R�c��e8O!�ǰ��m��X�j��4�f�˵�JU��8c�I�^��yU�DA��ɸ�l=����Z���@�G���[����crjJ���s�}
OA@m:V�%an��@Pϕ�_�l����Fʣ}a�y~a���Y���ުX�L���7�7��Ӏv��i2:���	�h<Si���F�L{¿�b�c&�\���ѓW��<(��k�
�4/	��^o:���w�ޝ<L�+���*�Ifk:���3Q.��]���q+�(Y��f�I`�}p��L��;��m�)菉�-�w;�=/
Hz���]�y3���JW�#+�μ��gAѨd~�j&��P�/�����/g�/�U���u����Vr:�`��#+�:k�w��j���,X�������0��'`�[K�	�7X��[���4�Y���z��,(������@[�O�{�]�x�4F��ìs��������v"�s:$�,��V���=	w�Q��ů��.�LDx�ع�Z'�S�cJ�����1v*����Ǚ���*e�tZa��-R��᷁|X~�c�:e<��\��s�P����H�]
l��Λ�2	i*���rtz!��37��-x�!��6�Fg��/$��1�e-�e��S�M����ww2��T����3��W�ER(�׬t���a�a���M�ç�/�e~T�]2���	z����3��٪��~�
�05�U}Y��1w��TYЁ�5�/�_���_��`�{���+k��o����u.jl�Ǳ�t��K�T.ۙ<����bx�7&��I���:��->J-lh��x.x���;X�%T��eQJ���?��)��<2ڈ	t��H�90=��	up��X��j�D_� �k��Ż_��`�'h>[��u�f�A�:��3�q�#�)�T��s�E�,`��Y������!߱-�V�A�=�Q��/lI�#���F �c��^��"�(�жn\�R,)�$�Yσ�ɇ�����@��Hy�4�@�TJJ۠�@���
e��R��f�|��.�i��̤��,��˷�F��:C��Hb-c/�@�ӧ:�[0困�1������|��bV�4̱�����T5���x���l���61~�{[��W�E�&&�a���H/g�3T"\���;�6�p��ğ����?&�@���qV����₢N��R����!�~A�<��K��$�}I�����2�p�f����%!>���:�$�Qꇢ�ZZ�v
���p{���U}czT�k�{�c���+�ש�7�D���|[�H��^�.m�f�6��RHZ$�S��z���=�̅�`�x\��/b�"��s��wgD�H	�ќ����d�nE��?zqe�T���ڒ�"^f�^��ly�,�Q�����B��T���@�:���G�R��|�I>�0��5�,��<�2�J4EXߔ���a(ꮐ�:{6�.Z��j���ƫ�H�os���M����w�� 	���Flt.Eu��d������ƴu��Ǟ�x�B�'�L��{��C��-�����AE���^@){�=�F-	�A�!a�{��@P��V�����к���B*R5(lF��Dt��y��m�E���^M�w�A!��t�� N�m�|�Rq<^���Gn~fb�JA������|�A�|��@f�uW��
�~a�#����wKkOX#��M.Uݝ.��ṉ@��������v!N;Sۼ���D�b.�|�CR�����S_�'�(0Ԏ��5nSc"��~P�
�Κ�&W��n��2l��=j�B,����E&B��Z�IJ	�&�;�BC
�Xm��5��^���HX�d1�����l�TY����U����81©��ĸ5{�X�ة�v`7��D�V��@p�>��l"}�J"�pP�6����o��WC�����9�V�Jģ���T�]XJ�c�n��ߵ$:0�˹��<5�S o�B|v�_�"x**!�������_X3� E�p�r����D��qQY=:�g�יy���>zƾ{� �8�z�iHN4��8a�WƏl�:���6�?Z��eL��.|���|�( �-9�?.��y|������˺���I�3.��\B4V�O�q��ᵱ����Apq_FB+	Ne�\���$r� А�ҵv�,PRh@oҥ�4WApp��x7=�!��l�1�vIp�I3�y��u=�	�t���3��xQ��-��\���u�3�ǧ�:�`�SP�ٰ�K��ן(�Y/��AW�Z�h�]?D��@���f�+Wj���p�3�cE�=���X�h���+�}�.��a��I��i8�H���;���(46��3!�!j}��VH�����'��Ry��H\�&�0���߅n�_�v��/@dx�S][RӴ�������Ђ(��) ZҺ�ژ����'Ƚ��!6P�z��#��(�������Gܑ�����}���J�S,lh�Ps���V�"��P��{��ڕ����g ���̫N�j�%��T�/�{��J�_�	�:�a�/U�G`�n�I���Q���LC7�y��0�$r�ыtڛ��g�aLc�]<tOQ���P�6���<�e���s�4�Ⱥ��8��Ͽ�����1���N�X�����:�Ԝs���ç�v�'���E���a��+�x�L����q<��6r�j�;c�n�v=6Mg`&�RޥL��Ga\��'/����0q��t��'����2���bT�o�f#I����2�`���lK�T4�dh�<��ߛ�j��#��7q���J��R9Ԗ+��4�_���'9.�*������K���m5���HV*]�x�\ 1>D��i����4uh G��>��XE,�������ܲ:�0}(-h=���\��_��d]Ԡ�e�3��3=�:��7�cA'	���A���������;c��2V/����4+R0����j�/���!��c�e�8��-��zv]�[���"����%e��<�#�Q��M[i��v���������8W�by���^��e�2'P�I,a
e�K��R =bx��~�x�T��o��ˢuhJnǯ��=�*�zc3�H{���c�.]M-�B��!��@��5 �3�w�n�!~��d��Ku������10�A� [Ɖ���lvjǥȲ
+yl9"��ba�����K��D�c���(s#O(���9=�����P���Y=)�h�?�j?��TE�K�\�!4)�8�a��q]��D�	�ل$�2�k�;Yf�����G���#�r�g(�}��$�m���;�qHI��鈑�%K���������2$R/�_6��,�c	$�6;���v�,��T����Ro�xI���#ma�IC�@� &�j5�����޲<�}C7�g\�9?�8ˠ��)��.���*W����{u31wf�i%��!OT�K��j#��3�Sh�0����/���i׊ܺї�����=2NV��壌T�1� ��j�a�t�8�+NW��@^�J.�m*J�e�zf�e(�0f>�$�`�tutǠ��b��� �<�}"�	Ȣx�P�Óc�U���o��Ja��k������q-�/I���'��FB||��o�ڱE� ��5C��5�p}��~�T��XC�B]��zlγ<� �?�k��@�X��-?֧�G=��4�ZƊ�iQd�g5@��K
��$ǒ��b)��SY�5��+"*�*�E��Z�,�p���ND��Ew1�a�K��=�h� ;�{��1������7�6m��߮p]#��z�Z&08T/�z�P��s�O�xI�+B�B��`+ά �0XܘE_Gv��3�8�vtO�	���t��3�Jt��_\�w��a��395�(r_ɫڡn�nO<�g��\&y�����;�/�(��q�u���J�!+��	g�y�k�ڊ�`S�