// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
QTud5cf5stYtOb6pZRaRS0HMdHE14Hn9XIk/lYR6mLTOP9kd8VjYeSazSgm70thD
MY9gNEexpsBbpmSblTtOIkRfy/Llz5STD3jQdq6fU8qF0gYizyWevJfqcFyNynEB
Br23fK2cjMWRVsSCbP7cnTL69dUd8fnL58njft60PU/C7zPMMEQlhA==
//pragma protect end_key_block
//pragma protect digest_block
qxW3CIQFL6Nci7UbAyTfylDXR0M=
//pragma protect end_digest_block
//pragma protect data_block
m42xeGYGcMswUUqd5i6k4qiawGIzvoFsb3OBtSEmiqKpREztHugqDxHK6xJq4Y75
krsLLSpYfYhk0jjkMIiFsp6h1TEHv9ZjUYNaAsXaX9tU3jg0fRmUGTtAx1M4SG7g
7I5Gronpi2NbPmkpNrKtVb94ijovaC0o0xXdTr7pVKzj86MaaIxUJq4Q5X8N5svo
GXRNu+Ew0nUvQMr86XGkQ9pwiuvgNeGirUEuObEnPm4KPaDz268GmLLpcTJxML2s
bdXcMRaJ6TsDSWwL1sAGKq4TlOKEVBDjmhGOuZJkGYyIwTr7LY8od+FZq/pAobRh
/DtuHCLo0hr2bzmJoEbC1345dSjXu+MAoOZF2/0yWvGuOgw4J0/JvL+bG6LiL+yb
uUt/DhsDNUk3WDlcaRA1ECUREGEJwuGZTpBTddwauuKQCHJrpOVmORchufVBwck3
1/wvKZjWsoXPtbgRyI9XFaw+BMW2K9ZeGWqk4KpuBFdDNw5HBxcEgTNJDSXmDJIW
e2CMGw2igGpCBP4GoOOowGeFqAvaGMtuhM3sv1wjHtCwyRBG5evckW+YILfdQl4N
4pQJoRwY0XzPCaWOJ/wO0Buvxb5P73qTg46ZfhQdNuA4BxteYcgmKu4saLAx8NBm
tRJ5n/8ZT8S3L0ebwrhFFycGxJbSYKEeP0NleKIJ0NG31swHuH7h3s5XJtyYnKPs
vJuA2kV3wVA6ccxToj8oVY4FWUlTgXbC0VHReiRuTBSrVezEYtYWZYR8+bS1Wx2w
94euw4UEIsqtJLXFTZuwii26CcqhUibEBfCFNDTyEQxJbutjW6/30yeYkFycGrY9
M3B66Z+Ah26GnQF0Tx6YcQxAdPGHwBfTEEoyCsbSaYnjIAU8gXDXW04rEJwDd80z
tF/W1nMzV8yc9gvKob0arI+B4FOyFIfprwKDse9aAZuLbNGHGw7QreSxLUXthXU4
L3dWzI9GluTsK9AZjvHDbK0tQVKDYhBhRmmWL02rp2Clsu2tPC7VibrbToP/03zH
3Y2m7IiD0Sg3TyWh6rSytcdg1Ti1AurRW0xfrUCQxOVkNz1cbiTQzemuJOe3T5q0
2wRqiHHmJRsNE2X/UVn3870toxFFhZNHw4Q355qJBESDjdby6TmOVgHgqaFTcpt2
Uieupbf6TJTgGEhFssHXqk329wjIpCb/jf3WOinqOyY+bNvNiwXX7JRMPT8aMOgZ
BMPU3/rpgv6H0m/b/ZhLwnjrUQBytJIuu/tEefqHlXpdSqBAes8DMOWw+lpRSbnU
G3DoYP+dJpk6lWcr65G8XdLDfBKhlf+j66nrL5aPf1wsi/ydlxII0sTOQ8ptroUG
No9XdZtqM3LyWkkFqhVFMEIAzzLpkDJHLYpwVRSvNUsYEQpUB8oSOwpLs8N4pah0
rv7mmSzcm1whlB5Gl6LM3k7bZ7TRqsBMoq5LxYrIroLPdmlPXCFrCRLfkBwzzWaT
VHtHg1kUf8zhwcPK6k3fLoTkBNbwDOSkTImPRu+24LIVC7/L5cWjetM8TDOMHmfe
axPVpe6TsmSZl3rLUxkwR2tgsTMljXPemrWpFaC276w/JUMa1peX5yqo+snoBFPJ
pKm5GjMhda3+5W5BdCGszIaoEQqjrI9NZULEXcvBaTJ4ACLUz4aO33Gh40P8qovx
OGHLZ/erYevTr0FmMAbQjoenOQo4BydJwHX4wGsbzGts8JqCOAOwJHwEdaBUpHDY
upSTEcHJ4hzAF2fbyNIek5iZskLJKqzsfjZCuZe5d5xKeyO8x5X1wD0HlLHGJd0U
8krf20pb5f6q6WMqW3EmDZxH9bSDWaGHRupmmM6hdSrd/uJxWrSyQ8CT+7QIfYBW
e4oydlo4LAQfaik/3XkR5F01QBGvQGY2CcESpHtsrPKglEhsEtOkvgyqQZ1xgzPb
wxIvavLI+4/bR0AN5NinUmDRZDXBxUqcOvmVJiwmb+Ff+89I3MfRSs5ErMwInw8M
I0QV55BWTh76bLcnpaoljNNEUUdbAfTbVexrHTO6QnqCCx/fEIXkd9OfhKMDf2iH
ePeJ/rCkqWHw6oTwtRMISCfxSQQSBwgEhHCD125KRItszVkzs8QttRt13Rmng2vt
lFIzjPWuNVYgqXiyl8kMixIRIfQNKimYalbynNTwf8JkzecFhltAGx4PmgF0/lMd
23J0Dbx/i8Q0a9d7RgiTtzIkkaS5gR2C05lNkIYcsUBq9c8uE6bYljmkjTJFXjvL
YLkANO3AOFHzAdWnyXi6OgXB7O7bsoFJWJjLPi7z20453TSQPeQUEUZUe6WTllI4
A93upD8YwdgN72U7auRje2nvfm4Io5PuEy47aPdp9xL+6jhEt/2TumazhMcG1VO+
+BcEXqv6LDyk29O8/Z5C6QAKJOOijajvktjy5ZGtTN14F/XG/yqbvBv5cTiBTfSe
b1YSNSQQ91Mc6PZfcwv1ElE/upOjt3eIeV6v/hOVJX1bYbPPQGpUiLzLd0y6zoeB
PI1Hyk3h3rfkeDyTpIgNBaRj54oCkDrhGYNbbfioajJc3O7QzLp9zvJKuxbblkUh
WJoXVpy4PsyqhYD3Lg7sUFtbHZo2CLcYRlzcDBvt4hnB0PXAn3iEYchNxe4NeKuf
4KCyFVo4aCgiCCaRNc6xn0PXxA3f6qsTneHLuO9djy+xMUSiTshVGtV1SF7RJWYf
08qgQNjFuJCYO9bjhNbuG12BqgYe1kj+kUGY9DGrDEfZo+FT7Hoj0QTv3mr6UzsH
1QpEmnToDp/8bXL2uPB7jTVEgQ8cl/FLuPfrlz6twHLNunZTiQPfonDnUX9z6SXk
mvjW26p2Op8gO/Rf1OaGHSW3yt4rqj8H/VVrNePmB9ZXti5ATqEyynUoOK1L9dW+
XGLbThDAeIV81AdBWs6EL0746htQ6E/gXSRKvWJ9Ch3IDh6kQCivPaat4Q4nqJ0Z
VtkJAgnPAB48vi4yp0i62ROOOqp8I87RHxEj6Ccuj7HY/CeVv6w0TXCMNgFAKftr
D5v9quRIBLYitX2KtJHYDoUfFzLOPtXNvcLF8BhJ/Qd9lwaSe694WPVRzDmSPbQd
jG9QGjxiSRncw5OzbupzP4seCAeY/04GVNRrxNDlnWQ5O2oMF0/PYPm0HHX80axl
DmY3k1ocP3g3rhyj70Pi5r8/aM0+GPvPsQCzY9Z21G0oK7/AdA2pSGxr6P64rNRJ
7sBJ8Bkw22gTkrgZ921yHob3mJi6vK286kzCLYh7O+U6VNbii+JmAdLEDZZrNKGV
EKlwtatrDIckhnP797Ixjr1Tjrlb8o4G9+ENGs0tHlPkp6AMUcKWgD7Dldlm8cYt
vHJBvCzXgHTLA7IDee2RsZ9K1OEigSu2JJPw/30UMM8DfVRYa634ad/IJtotZCoi
QMr0b+PRtzSeCI5uf85q8Fx6UV3jh7IxI9N32sYOc1NuA8VgN04P9VCKSe8xSbPD
AErstTwfV/6dFnHx8ylsS8yIqA667eUvEEpNdKvgt0cpT1GlG5tICv4P2XtyMVUG
pf4vykcAgj4YO+Y38Pw9HgXyv6BawaaUSpEKuRYzkTLnrUaU9EU4WRn6yWLjb1Ig
Q8S00bwqNe1eh8TWXdoq2SzltCrQm0VVHMSQDfcqMFEXt9h9047iKW9OyAyCPETK
Hty2OAZt4ZR5U9TOjIfT9glQ6cJV0sc81/9qWK6BURCNkSG62AjDDDXKutB4Fyj6
L5227SsOXcaMKqWCxxDrr93z1HGttGYS21lQM8boqhoWew1SLupcqwaVB8J8wYIe
mQnaUKLc4ElMtZKEAa0bnPkLWTmBHKPuHZoeXQM8xKbXkOUH7aeQLzhphjjS+lel
h//sGS5aVZRC0lDxLsUnKX42XWbm+rJWxK68yDuw5kY2CciGweO09KFSBm260sUT
aK9pLAPa1xT9W8Z4Fj1l6I47rexMuPXmrPbjY2xbOKWCRCdtY03/2LAsnQim0Io1
x+JHSnudGrRz7X4WXOv7bG8GsLlIFg0CHiuPN1BSkSuqJRvmjlij+uurJq0gBQ7U
0l052o81M5OdtAXftr/thUg0jaYvsxaUPPaFyzpF13Q3msIWEY/tWI41yeOOeCLs
/7lNpF55TNFqdxo/kMUAKbQNs/hhmt3fO4NMlCK3kSH6iy7TgGWkagagQ2tTdXy/
z3yXCNCtrDJcEh7UHyk2LG6f/S91BI54tOTGkXFdnL0pSzF1CD4xG4Lgbwg9axCe
AfVRWTWVHzp0lQRbRCUu2tkc3DXRXgvGURA7IIaBjHzqAz5GBn2pWCuNA1CvyoR7
0VAzV1TLKUCXeeW3aB0WBtxQ+bg739EFdiyZe4TxsfpbHTxuypz4uNKiJ72pQxOv
N2difz/L5WfboMMBgraqmhXKoH4qGOtFm/FYG2W//IyMiBGkHTYfdKYpzmnoMglv
uRmsYs+7+K8SL2Bcl95jx4ruT0G5ZC9pi/OuyW/NaLEonEj7vv+JfyH5Ps7GgkxC
YDJriQMAy6zCXt7hISJ+7zc2BygOfnAu5sVfOjn0g80UHDpv1Q103eg0NaZiNf69
Uz+ekAi0feYx4mk/IHsCbcS6wQWpaOSm3apcfIEhTVurcE2n4WFi86c445fUpL1J
BzZnYFtBrHIU5Wax8k52+NINH+lBdoU1dQxCe5SCUyrcrsZ0Gxzy69OTeOh+Lq2y
wSdAou6EjoLRk7j/8gerBFcrJtC6/uB5SNsUx01e1lxtrYOOh5nKc8lGPP8iDEEx
p3uH5XzyOTJ9suufBTzF1e7oIddlI0S/PbOY3jG0vV2LiHJAeb3eSUP0n4i6s6U2
3ZiOnVt+pWlSKJpwIpVGWLihf3UNqjgOzgc6YR4gj8ix1qzdBPptDtXyn7YsO2Eu
aYHLB9ozbXWMShULyXQmX/TlJk1d09kJEuQIRqXikJJwpi4lL12pOSI7R13MP3ya
Z6pCptbUcPN/GZvdElun+Hmf4kj9/KC96LaI9apzQNYsGu54gsQJzP1fvy+dP45B
6qKB3xAD/YGDCSkcLBugSrXf6jA1XWBEq5SH1v5+yOwvD92sF7OT02KfLZtf0ORd
x+WPEBjhoYTNjkSeSFpaURZcOUC6TFGV+z9mQl/Ke3NhwB2fAYpOze7Th84/6mmu
fhjponE3U0P4IuOgd6IDLAFPeoTib2lSH7BeCQlxFqF9cvq5Gwg13FFuAgp02MRS
mmvP6whxQWkOwQkNuvdclAz2KAT5eutXMZYSfcZMCbL9rOiZm0X39C4SDxmCWdG9
wwLFuWkyaaKWaIQh4HDRRAD4r5/kImzWrLtBs8WYCHbk1XrgBtLbSjdJz8waaajQ
GV/9hfR1+AsWJ0L1n7+U19oe40hwPdqH9z6wyKErQacZQ26c0nOlSt1eguQ2Ft/e
KQLqa1z9gk4mrnj/IQPIg7G4vma1YcsNwewW7YvViGZ2h9+vFldc6tfai826tZgT
10KljQ/2maBTXmrj+fMLQKOfU0QMjC9JyCQ9RliDnjQIowFkhzhmsN9Wwrh1Wa1Y
NN1dzjS1WTVKFjXbQS/nlvk7Kumz4Y7FLIWdzdBk7IUYAIz0fOVBAIJbzJx/8n11
D6k2Zsz5Vp3QwF7bO8W/DUvIxIHtfT/dqrwxB+UNsQGDS8usWwjFrgF53xsWikcE
2GOYJeehsduz6evie8vCUw1oSLM6Qq1cboCaKq2JOr2ZlVwx+/e25IMtDZPKdeNl
LXwm8sLWIrpSSYUsvPgv8qShDN5W59TJK0/T4tSMjID1N8XsRT45ddQaf/MNGJrG
Pxvt4CPk/FlenBYYWw9f93QJdbI7aHP/JdwZzw3xSbn3j83GLE5H0vE6LUoGWahQ
6rkuxKM7OAM89kUTcNuEeydKDlgDyLVPx+F3mxIptjFzMbsAWaDFkQ/8yqzXhmUr
Y/9m+Zk+HEKz6dKSS6/c3O34EC/AY+g15aP6H3tU5H8xKadNCazS2lBRKARb56H1
N9lFYt+bexlmCX9/+1Gxw/m16jnaqZu9giLcFNkweAI9ISH6Yl82GaiX2WZ1llR3
ZUS6SU7DCVQy724hv0QOMqC8V4/jqNTtBhnFZDqpFavOooe8VVEPcs/A3M5TK8HX
54vnW8lidpYHrjTRjMTdzpP4K/3f5pXYLlne6H/riaBak8jD5KWt4MrLy9a2JSef
H9rnX/9XxKJ/bO8Cwownu5LQm3u/hEELoEMw4HuOlBBNrxUnpoqYUcVLhtHjEHDW
VjKn7FSbtjArjCdicTKgWz9Ey8JVngdPHzwj604BU4z4W0p3S+EP9rZfT4DqSIPR
HOjoS8QkgT70L4qBrKWwDoFV+rCYg3OZqoXGv1xlFAH7x9mXQI4XHbDfS0Ts4ADv
JvAoM+SoA2FG84g3LAekCPWapQBKRb8Ua7/L3uZ/bMvMXUoXFABOaeHFgVJN0JZE
1ysQh+kobR0V92xsGEBCyfWNmCXWcGg0avPj5a7rSs8jpCNLWQa5W5dhSxl335MD
v8y7nvmEdRP6OTF0cMzPOBAF5ObLMwZ5cE0Fcrx7aB1/iO7jFyPuLqB2G8ayB2qp
4wjy3LSA2K3GVefXOHxKfy0jJUylqtfIoSjFcrN4OIxHQJv/lij3TSXfyG2Nkie9
UeYvyTnHPMfaz/3uid1cDvEtnudAEQnxesuTQvtG2IsKlnpNgds2QTtCapA0a4Sz
HBhObuHKASqGhiGGJzhXn6zOhoUMUVwXCg4ZYiadCmeXjKJM5cSYof7lYJNT3IPC
2Ui5bqvi5sNpDIvIlz5lE5XMMqKWXxrIhjwjp+4Ep26wqVuJkrWQ/2KMS4fXpDLf
Kp1Y9ZRNhmVVDHKPk9wZIh5QhA1zWh9sYlKGpjCO6w135+QAXEEpqDDJvYLNwXiX
Cz3Hk0Ulf0iJZ0tLPRc7kca98rjLZtQSTXDx0/3ousS8z65ir12JiR2YGHhSwfHn
FYUPR4YKzVGof45QjI5oSM+2cVYfcr1YXL0I6j9GPz1ySaL9N4C+lJ7YxUE2TCom
LSsxPF8oxZpcPE/QRULHRQvo/GPsQPxP4RxIM1E0erQ/qLzl6fJsWLwkOpmzJ5vF
zoNJlBCmUbcZtta1HqL8/3pmFRVOgFBpClodryWJjSnOlY3kJusUZbNJhO5VIlzc
VTiGp37J23gzok20MLrg2uMZ0BsF9gllWarXwskzm2NcwKSzgOxfX8cl+z8W77PK
3WPqUgeItvYiIGQuKoXJ57aFcLc+7KRqTIMXH5x6dad97SA9mbrahzrrclDw0MZN
OfETD6MtckRU4zV+WSgLTEjb4Jo/HUdszj/U7xP5N8FC0VjvdWq7X1YcHHopcEuD
dXGCvy+BFhVlRfgh9t06D7ssAM7x3Nn6s86Zq8nDxTUraAyBG8hmHu2oyPz4oTX9
0RN1k8AvNC0mSG+dczBb+dGLAN6urf5qjF36vETCVrB9Fm8JO8bH+iSbCq2CdnkL
JdP8PpydJkmMigqN/4za60N+otWoUePnCgBNm3sR+VCMnSDiWiiBixXjHJyawLj+
RJCNi/YBL1u2c+yOsxd3ZuLVrXl7ueDY+QKqyAthBF0N8UbupmJunykSg2MP9pFZ
wMRHZ6g6EDuMpmrzpC/RCTRDgim3uvStH6NyxS6NqV1ubbyG/iVd0zCqvXUzFRIj
74Ig7RlFxhVsTJDcZAhIMyU2iRabTT9n7IlHOegUfnCiPziW7ZcbKHsfBWR+k1l6
QTLOpj7EDfmquzjl5wPxAPX6TkfJ4IO8smrFV7mHg6n7UfFYEmNDDucq/XdMMSGe
hMD2VH3kg0SoLKKAQBp9p1HFjoee6lCu2X3Il6/khuLCCMMHPA1QFLQv2q8hqJsE
9w057E9sr6R4XVIQro24oHObtvjh35a/L1FIXziwehPxD53/f4ZrvaIK6PQR4QIe
ng782pHonj1FHW+BJ+PJ1Wt2EBUw5UUkGeMqaQJ4mhpFD3JmmYz0UCP4HtMwloh8
p0QZEd2+4e4q/ns9O+VVjH5rcfTgszwAVQv+Y18+sgVWf9FQkvDWgFzIn6/H1bzO
qNUnv4Acc3EPb0LbtO6Ctf1ZRC61hWhn9U4J0B7Q6fVpsom6ltUl/N/anV93Qcg6
4QQKqeFAmeaoVh/zgaTXKDu4w1qe4a3TOF60F753N3AqEAp1D8riFMys0dMwB3LE
i+XopNlxHjfw7V+/UFwArVwCrmBoeQq9LyAmCbxaGBDpxYtv/nXAF7w1n4TRuEUx
eG8g4oTNmTFhj4XPgMgFqRbVxYxvMBgxzsgpA19mA0DT7jnXfJUw32lr2tK14cmt
Uij8Ei7WQiqBMJ63YRvPls9TBd3ZZ0Dog1KQfHp0kQpT4DdFXgY5NYDSS+nil8Qt
G4jKe38JUmRmkzkm0Ke8PZy2/Sq7jLOU5mHzGnr38jLYM4r7XSN5EqdCrqnealHg
kcjStZFNRxVvuCwiJ11zI8R9l2FN5pgacRq6dP8OJVOwYdVCOuqurh9hcDmRi+Vc
oMrYVP7fMcCkq8G7AEMzWSNPN3RC1yCJisaZWGbGt11U09/b96BWMBRPoexk5ejJ
aoNsw0BSnB7zwN3nCfH9+rC1dMuZc983nejIVPCyqjvYaH4RvNZyLjfqCPRIFYQT
OZn2xia9EYYWwyh8LJFbX6jXD9Fa9L+0cothDrxlXlhpZu/89vgxw+w3Iqyl/jXg
v1I7p6EhBWNM/Q9u94N6DOAX3Na1k0K83fiJHCQot6al3QtZ8epAnHvFBCa61N/+
jBhSYbphoDEqSzTnaJcl9J6HmiLc5NbM03TJ26NZheeLUc6KUlKljF83VdYV+P8m
pYyIYOKm1gGek5tgm/Dp6YOspkSEM+1fHgITXOywAXW23zd1D/l671b3m/jt2Yoy
qPrpX2lQSgZGrSdzUQF+VC5bzWbVxKv7haceNXHu+8Tf0GYSZFeAkVIbmt/j55gI
1IjIfB4PJAxTDJ4BKEE9kKiJzwXkK9+DoigFmkX8eFOU8bhVDgni3+XwfufAtGcc
42YCZLl2XyWYhr4gnsKckPYa+/jHigUwZlBWFtWkZvuePWJQrAM9tMWx2Ha65ka8
/61IctGtSwNLTEeUkGawVzSsDC3WgOZ4YbKDukzNxM7rtGJ6I0qcbz98wB6TGTTB
uwk18/x5OWJWm7fnUco6mXgSmYaXkq+ojuI4mOuadra6XHDTjgePZhfHLvt6z57U
DMNW+2J/pn/GGqX1XLtbSDvsNf7qi9WgGdiQ2fGBIKt7kDRLvJqlt4JZZCYLGy38
0LNye4qQAuMvRi2prpZdGgnlfdzbjqI0HhOvCC4mBDj6uL4LI5CuV+tKUcPta2qi
MYvzYlGfZZ6tpLZYJbBn17IhYYAxQxu0XyD8L11I77I/5KTdXVzkCksxhRn+nZGL
wyFbbv5kXgV8jmlgVe2gZPECEd02Ma4HNApEF0n2rbzb2ezO2jBzdXsYN4zX7S+R
oIIPlOv50dxVy4mBljbl5YkUJMpn9YrtxoAZfZQmLS69fxOdz0ifGiMttHK9on6H
ofdiINksXoIEW9QWCGAyP7X+3YGZRJ9M9G7wa9DbsOy7URASCLUj/eiQoYlhszaH
vQPhONVEX87MNwTBez1tI/gxF7s+ZjrIf3D5aqS9gmsA76xS5zk9wM6VvFfxpDf0
VqEqumwMD7V4R8Jf7uObsjOsyT5MnXF7IVgAYMYJWvScxDFwhzTFmcVSB6PWE0Dn
fMlYiGqUEdkeMAgaOvx54CwTbKH8R70I1Hk1w/pI7qB+KD9RHMA6FU5ZTbWpMnBu
Ku/Hw43loN6VsczWHrS8P5Q+GQ40RG4vD0LK4v26e/p9YtYgYCO68lISu35Km+qR
GmgRsvnDvD/rk+wAnAnFEFzfZlR22bVOTdv6+VRjLJASjvrZV48VgqUTZX2VV1xX
TD+jpofdUNKqB1zTum5NK99pu7yHhil+2WeyTer4HRFTguUYHNLxXo+7iqO8f3Ig
qZbwYMozhwHRIQECfRNLEnoc4KmUZ4bJZ5JMbIyjEV/SwREReXGKu0eMNPpFFczn
ToZfP64EuSDD4ABItsFxUftWESdKCdeKG46PAJJzYzS7wD7/nY9qAUwCu4OpVCgK
FpRcf6fhQmE2xP4b4ZIYsZzTut0z9zknPIpkyvDjP9LYTEiQ6KPFlBb5OUB9sMJ1
Cp04G8EkBqEL5l1qlPhnVL/bAy+s7qxfXMgA4Cj70oYKJYmhrpzDBJ7jjegOUoiU
QRNl/x7oMz41fh7soARFz/Th2dA3gjETIu/KcEdeBYm0fD36XCj99b1/Rg3wg2NV
kB6kEYds4PGXRkGoHxrNm0S7tFySK7kyS5XgGXW85s4CC/B5SaOsOgehTnowlv2f
apL2ImhrZSm5rvHN0xAdf2QUC6SkYSNUyWo2Q84sLw+usPdy0c8C9L/r95iOVZlc
joSyjF7NY123z0j8LUF3RE9JSTYZA/vdkCaNYk+bqz/8un1477A5tVZHyXfJy6bC
jf5lzmRC7tyuxfV3Kd2ozAmF9rlfIB9tJH7cFzZbpc8s3/xHvwtifgZIvmkvHKlr
lb8aNm578F7ziJhba6UhSBLwy8MZTpSf2xNCxUW8zYxJeOWndM12v1CWAvzKNGV2
bKy5iV1Omv7mc4bUKEfI4OImveej9afJXR585DHdd56kJFMIlVub9N1oMwlnC5Xn
uh5G7vRAFVuIXkbfKaILIrYD016XE3I/ppGSrs9RcZ5TyHlkYsxkam8i2MeBO5eq
IXxSSV0SlIRrGr85T8j31UA7PvYyE93PsM3hx0OxznnAo0X7TKewzlpuhl5KjjkY
1xinpZrPjFI/PCVWQ3NgaQrxzyUDtqmhl3PYUcjkY7eNdE/B6Jjyj0qteCpBftrj
/1gHadHFrqvyiHWLzemEI8u9qCYIv5EjyD1/xScBaz93o9L8vmjXbND/YDD/+Til
wZ2MWHhIuP25hukxx+tD4BFhfCMUvE8PxHvJc7Tt2XQQ2PPLVBN9KSAkNDalRy4Q
F+aE7XhiVetGB7CHqctvjDSd9hAsLhgTv6W+0bF+BK/OqeP38/PWyp3QxnCewgzQ
Xcz131mWblZm9a863HxTLLyqjkg6qHK81RQy0fnUeHsLqZIvkBxW4dimKGWTUWGI
w0OmnN4we3Ccw2BERY2jmJveQaY0XNc3GImo8DJ866FdK7r1vdPplU7/Dlrx+5Dg
3twebIhMB+pI2ERCl9dArEq6V0vM3J6xW0kA9HZ7WC4O/0+T2VFN4BRnfVEP1KpX
blB4N67AuOFBc/rw44dAWZbbWBNfW3KV0TZbGrzN9WplIYdb0Ua8ZR505itcOwsa
3hIH/SHk1VqRwpHoAwHMpzyEu6nizEroQi4xwluMbnaT0JChQGd0NORaqdG3QeY+
cAjIAXi2rTEEMOS+oAFGX/iD8IoU/Kky8miDWYKuZxvkFmM2DGKDACjZKTi1E/+h

//pragma protect end_data_block
//pragma protect digest_block
r7bFMv8sbYGglpj6l0xJyMxmWcU=
//pragma protect end_digest_block
//pragma protect end_protected
