// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Yi03ZrALCyOrqmE0BAYg4mWOtnUmUXH2WVPAEBjLfSYatnX+q608TRQbqLJ617XZ
bFDrgIph1RBS8uA0R6qGhUOLOmpuODYGzn2uilhtoGs5hWsROmRJYE4SB2mtonmC
EFvucWe+hWimFchuPJisd0uFDtexGKweWCDkbfkAYbm3UGBZss9IEg==
//pragma protect end_key_block
//pragma protect digest_block
WMjeD3uhyCUAvZFO08/vUTjWq84=
//pragma protect end_digest_block
//pragma protect data_block
vDP+XMHQt4e3LMEJyI+dD8YnG19s+9mkLKk0j9q3g8OuLQNKc50fGItLAtgUDfVp
1te7TidMM13D64u76VJB6vqI5SNqAawxp+EjBL0pA1Vd7ET4fDTSiYOSxd9HaVAm
FDgrZWMUDVdd9G9TrUtxVAvb8+2/8pbXcJX7Oss4P/JQ1sL5rmoqHOs1g4hExBX9
6WW02IhvRz/mAIZICgrgenHgFpn77KtZi9PdgQhzPI4RFh4iaJNb8VNGP9CUCFVZ
YZUGW6gmuSAIofUjohVScmkyZVOAb4cvQAqhb3mzcmfIaRzHtYz9Bh7TX7vRbUvc
JEFAtJPayr1Xuv3dWTqPOH0wOqkFR8pbFkJeqImkEunX5i2E4zvIikmEd0VjTxD3
o3y0FesBXZhETJAEOwP1yn+elQX/ucC5i9AoNuQKKA7cA4wGFlaMpDewmUs9fXk2
057eCiXbQRLDNXDlrzPMaMvkxj0Mej22YzdOzX/4n0PwoDBpR6EYm7NZCvRqNnz9
x/y/FpiYIy3jlLf461Ehcf63Yjm7wt8uQxeyDhIz5d3HWgocNSyUdVlo9LFesBWt
R6FxLgf2bgpoJj6RnKEd5VSZ0SM0vDk8YIOMFQThJ3UdMVTKxU+SOz8U/BirLq16
w/2mulQ5DX+cMk2AB89u+F7a1ZxkjIdjVdvqrs9kaLvtovI9movUPMXsE7JVKhRx
u2pfInFDAZUqsORE3p7Y+T8eGkLJbzINyFVo/pE2f+Y1tbfdVxQ8S//hlRf4U/dJ
/5+pQWWDvokJecwJdHAD3TfvmCJ6b0X7ut2SlrO4/EmQOgt9iX56gPrC7g5KJRW2
/xi542RR3tudkP5X6Yaz0nOIkzG3XC+xe8mxjz2I8u7x1pWRBUtuBf3lo8kh/Q41
f+kG03v6oWFJxfaOFFF4dxHsMzC5eWW3NrV8MKc0DTeUW7HlV7/RC/nttV0pCqnt
CYK3OZT0HXH2wRgcrKSJvzLS42i6qPvPEuB++aDRvzFzVnCilXjLz8HA/VEz66zu
cmxAOx1O66OICrG3slpMNlGrS0f8u4RzaABiViHetK/T/HEqsDs1f7x8YJUzDnhV
73LeNWCSa91xF5rBKuQ2+77GpAqMQGBQu9a0F0sQ2Z21Lfb0SIrWJoZ0eahz5Zx8
Di2eWKrHxFeIpirpsgKx7HG59Wztk5yNIuuHe2MB2xlgxutjv9BmAzBcRItUxSYn
zJV7BHFsnebqoEWWWlIhzLAX+bVf/LZ+QRg9iKnedbDVvaUcwjVxkmJ763I09UoY
LJD+N19budgXXtqMTa+eb8GzW0MH8T+B65UzjcgFkn15mvrn9b8/lOB3SXxg/61k
BUmoLmPOMib45WIgmCJnhwRL80wBAvlnm27+eo9akX+YmjCUekhRygonzZYC5LrB
5Z7tBqrOU68ec+SvdKh3CnTSrBDzkgwz5OMa7faxKV3HSvp/JZuOpuIJRswUPTt5
tuQ3DlIlCYllJ5b+qUXGxDdMTdzqm2hONJqDSO+T0EvHo7YMK/1CdqOFeVARoDdL
r576n4REwXdszttSvMyL7HIiVavUfc6zsch/4MxJBTO0lVLkdbAl8ofGgUq26y4M
Vzq1x9ZLHl41onmvw/KJoMTIbRTWO7HYprSV29ywtf3rB8fP8iRhCFc6ZsnxUIV+
wjXMqPy7Bh7Q9EUpYwsozuE4rLA4Mlwynpz8eGLCC4B8ZPT8h/YlVI4pqXTNJfEu
nvUCB9N+z3QmMfSJmGbI5mc9k8d0DZNN0NYz/ic88CDnemIR2SLMY0qzPvrqSY9L
6YtfmBOLPDeDMW/j2KfpoJi6tkmRshFu6Cdz9Y0MAuBaNgT1oPaKVTid4NGbnftl
jnC9MuQlEsU7tAIs1KkmCcZDRN1TF5Wz4N3N8gXAQ7paeKjDXGpvUYgjF8sguHou
dio9/V7ua7+3x5W31R0XUS0s5PNlxfjnTMPNt49/5boqiI1puC60EjoOfgpeZTrr
lZaJIlVqUKtZqeISbNl8gnyAVp31jCQqv/kdsJMwPClrwlTiloEW8V09VQaOYd5s
19EZJgcXXe+O8FyECaPMFfG2N18YSQQW46BCINcpirmuytcnjpPlMNGGeLBDcDCr
R+sRdv1QGBXUikm/CXvS58ZKCnRCgLex+Xqa6oS1jB8Rf54DldvKjb6gnzDTzpYY
RGtaTIDoyh+1r/iHmM5OcdgEpiMamJuctaP/iR+b8UeVbg2Q/GX9dyMS1apsmYUI
/alqDQANbAvrGmqRCv95yKe6TsM2f6fV54+UxnieYDMnsHBWPjjKnVwo2jroREEk
6czG06yVP+F8prIY8xRjoUZ2kWjc2M9r6YUYD5hJhY32rMNrtx3B5HkJHCg+yjpD
0p9CeJYt4C3BnoifftKwP+OQkkiM0h2UnaYuCWScln19ZTngBWN4kfwuxm8BeGBI
zI3FSc0AfVa1n/iW9FU5FXgw60zU1IaAE+C5ZgjnuidiyhsYdEjPIsoM07sU/LB7
+1VFHZW0U/cL6jBdI6CB7gLP8pcyGmOXYjK0zunMxDdYxxK7BOeEyv2TIeu+Dpil
ApgI59yhBIIQmVMv0IwBXcln1TiKUhI7BN0vFVd8tRwnoiIQh0wY6INwCsso1lHQ
NUz6RadxO/ftPtgTcNzJAQJH1wly50/PrQQZpJ+FsTa2U7Lwu2J4hgrj11jinyBp
4cdTDhpKb4dQIIes4oMC7slg1i8XOZBc2YVpl5097YQXsyuJcntBKsjKsnWig4Ou
t8XRemn6r++UY8u3Ea99GmSzQAtRstCVgMX9vEUU8wp2q3xChbmGniZjPzkVaXkY
VRNIzoeSFIDN6kbgQo1ujJ29qQi0mW2+KjmCkc/B70ItlKemXOT4eG0UizGAVPox
DALkn3WrXUWOWVCr24xgW7J2/R4IP33olNutWGtggbiprna7G6eGoj2L6bu7bnwC
VoahWo3xBXjCJT/ZaSNB6soXzf+nJqZSKyzaX6rcJE+JbrEBrWhAYn11cin16oRF
6epOnKe1IaIvnqaOH4xAydywOmdk5q/O9eLkGM3KbPGrcatFNOH8Btx+zA4uLjSb
allKmE7l/MJ7YY1R5hynPZvY1NN5xblWCagqgEkS8q3y6lzfDlHzBTsx2FspXKZ0
5r58CDcfwvFQ7TEoBzXCQGuroxZTNluvbt0cczMntDz9qbsGLodV9usqsP7Kzbs1
eAquuJVXxyMVyqgfbnMXHfSCsiJrz/g8Bd9mP94gXDHC01/eJOnTR40xoy6h9Fid
3N2qUyPWrbXDnPAY1nh1GPaGDx1K2SnUGNCfzFm03P1lTEzq4XJepfmBSja/OQai
XyIcePzklJImhNtOJaQIs0zpxjN6+Tn/U210y9ixetIcqoH4ZUK3kMcZ+3d2HrdW
X4whqs83iN9OWt3vEqMJ8ovQJRX070Ln8sCoW0z5rrSAY4iqSqj4fqMQDIrltiRY
E3XUtG4zugBsAGNVSJruhx5fMPfOZrrzZ6qEsjgWKx/dZqgh3RsZh1H5XH5OEmi/
Pq2Fb6yOjoBcxginx/IA4d5uVMEuhI2aiuCePh5kA8kkhKjqoctFNtuIwrkMpnPc
AmnUoMww1/BrrEPfl7YyYMuVymDi/JY7xNoJ2NaFKkL6D9+9z8HTEB/xEhElC8CL
VY3s7c6eJvsLTLSR6PqjPf9V7Ah/+Z1x/AQO3uwxxMwDjIg/byNqbIAag2/nK95x
2+hj8dWIYDRFFeBc/y2x1dwIlRaizmvrxCdHXZL2aixfwVAo8mt2mLeoLsX9yJaW
dBECZzH/9ATTcG+PXTz8gLpTBEsobt1vV5DVKcU1VrgA22ueu0LTgaPtHN1fY2I4
lOcYJ175U9sN8OpwxZ0RlgEhm4CECTLXUx0wE2+SckTWbhgdAO8VIl9FFoZY2Yhv
bE0mqTSHseq3+RuQeKz3f2Tx8vavBZ3w7z4usMEvFz7oQGfspwdk1cJwFwIhQefp
i7i/kYjogJSHa/OTph9sTejM6GqOVnVKOmSxSebvD8YfXmFfQQGrJ+4D9LGA596h
YYiYz5MKpAcCTiTTkY6ty5CWrcfk23tRq63Kjq/qNpagv9kvLRevg7zUEjkw5l2r
gJCghIO2cMadWSiXkyI519I2y484e/qWrtNfK5qfU4hzhRLbRDpiPOJljppStsJY
GglEJjfGfIEpcb29d8YwJnl+sZtZ/OKq7+Fis+DE1AnfK4pqbZJWX0UBACAwtE7A
JEVLCescBZFHTfPwkPDUqxRXwc7oXB+PoK651WcWp0fa4b9mvboTopIIChott9Dy
Gy+vb4Nb9i7HpGdGFYptw3JspZyF4B9SY28MMKNozmqmD1uftIuYj3y35iCysVIj

//pragma protect end_data_block
//pragma protect digest_block
5buk2s//ASzip3finp6TAzInB20=
//pragma protect end_digest_block
//pragma protect end_protected
