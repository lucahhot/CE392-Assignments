��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{j�X.;߅ţ3n�c[�w��o�z�����_&�,}0�F{mQ���L��ҩ��2X	#�,4�����k�2elL��������?�W��٦>�����|��F�}�c��c��Ǣ��Ѐ�[dTf��䛤���a�{>��G��4z.���~�����֤�D�^6�_��T4%��y�:�}�����2xN�x����u���a�IV�j[1D��	\b�8j*��Mlg&%��jO`H�8xm
��=vB#ͪQ [�-�s�����Xl� D{s�*.!��D�{Y�A�2��(�fǩ�w�R�hY�Kl������3��'ixC� %�o���Y�b��J�����=�o��\�M��%����2`x�{By����.��J����^eR�x��t�1��6�!�1~
O�8�	U����5��� Z��^��j6�er������wȑ�㋌��ÓkcIB���eƿ����;�Q��<�阛�2���xM�t�C
'[,f�����&	��ؽԯ�����_�g�/��4���M��;L!�=UpDd�yqCm������^���l�p�����]zw	rFR���M*j�e-��ԑ��f��d�۲^�9�Lcn�'�����jL�8��'�e�֑^�c	؊�������|t�b��Z�[��(��Dz�ʦ�b��^��ʥ�<��.Z��F ��[�S��м>�ȄX��O/��Ɉ���H�X�PEN>����;�\]�gN�>�,���������@~8����3v}��#򶇚PB� +�y4��U���=�f.�!?�����5���vՏ�G/�.|�1�����ۑ��������f�b{�cMU�Ju�*�?��4�����
��|"W�hq1�Ē��q�O�e��t�3_W^Q�9*�4&�wB�P�`f&�c19ϟz��P��b�O	��]]��'���b,-Oi�Ax���kՀ������ђ|Ѓ[Ef:�Z� ��;%I�`d !���ֲ݉�PټC�� Xj�,a��_�i�k��0/NN�F?��TPZ��Q+P�P:|S�>^f]*�@�e�\r#��t���|Q�iX_Dj���g��$�Z�8$�^�i¼�sN�n32ܢ�l!�;"��t�j�� 闷�V��q.XZT֘]�(�0��)D�M��>���W3KQ�#���-��s���>w�"D?��z뢶4E�]����<п�{�R�l��6-~�e�&��N]��@<�Z9ћ�Gkg��%sO5X�v�G5�� ȹR�J8���'������<q��!`�*2X|��H�����;9Y�+�2X� Ew���ڹ`1n��^�0��-�ؕ�+��n����18WnH��7Q���5%�a2�|<��M6�E�� SRG�^�T�6�	��Ji;��׆�G& ���tZ_.fm���gspcu~�J2�w��������Ah�.�p�����4����4��8M��oLn���� v�Fj�s���9�-?4p<����)�J��{�&Ó&�e���]�V����0̩Y�PT��l��\_���#�>tV���4�ӷ�=O��r[w�J�ޓPLh��P �K�D\����3�!t
D��L�Y��n�?J8����h�`E.O�i���G���@�`	����ո����ŋ�"+s�vj�M�;T��6��S�����˲�T>_ک,
��׹���ɛ[�邕rd|X����m�Q��ˢ�"��z]2Ag�Zg�0���}�=;�r�)v$¥�r� jg+4�hnV�벐��[ ,H�89s�H�8Q	3��X�2�9#�/�vf#.IS�}��Q=xw`S�@Rh�B�e�ŗ]���'����N-�J��;C=(ȑ��N֔K	0ג-N+\�c���?��;E�q%R�)rb��UqaS'�@��6P�f�Y`^��k�I��1�����pGOBN�܁�5d� �LgN��{ɽ�ߝP)�Ov&r��ϹO��)f�;�B�'
��"0'cd��_���sx<;��(�r!�������.���K���xA��YP���b$����&ϱ�ȫ�)�A�iV$�[$O�a�B��F���Qx|�?-��|T�o��G��#v�'�~�L;���0�MXA	��$�m֗�L.W���p��Z�C+��f�?O3�!Yx�}x8�\�� g�� r6jb}M�������fڊ˅DN"<tۆ��!@��(㎺t�l�{ky
�V�I�Y>#�8)9���D�Ь�r!@Vi�cT� ��C@�u��m��͙���tQo:�	��PT��&���]մ�d�1�4��|:���]k*�Ֆ�X穗�t��E� ҙ����;Ѵ��ۇ��IL,��1 $��"ٱ����.vV�;�5�MKY�U������1����k��
 �V�|��b��]�ژ?�	Fn��nh�%d���UkI�mg��:�x �yŐ)�D���O)p�����۶JBMy���x�3E4u�h3"E�ST	��䎺!v���?5�&���C��o< ����ջX1��!L[������/�_Z~��r�z������<�/"��w4��Z7�)E���P��h��ɠ5��g�8���7�"���˜����CK�m�{�q(��β�tDbP����q�7��{Uޅ�W��׽[bG�����&�ĸ�)�@�Ή��g�w�uO�ȇs�����\������^T��&�Y�DЍSAdt ����'e��7�5���G ��u܄����Q�-x��^�M��.q�쭁ƌ�S��Z�6Ɏ��L���o*�^�/����͙�A�}%A��I�Y��JBx��_b���4���-�̀"BV'��ҍ��r�|��M�!�a�?^?Z>�9���l�j0�o�&��YlXB}B���J��Hd���u�����KIZ,��
��C�Ϗ����#}�������q[������Lqin( ��5���8�%?B��0;����<�7�����Co*�!�%\v�>/��`��Z�{?TP�o�w��;�����ǚY��-9
5�DkU��*H��S���R�95o��F��]W]Gt%���	�q�����蓶йi����N�����:4I�� -X���5������};����eQy���N��*�#�$�)*Z)|��08>[�~�=)?%�E���c���PqC����Y�#!��OMP�u0[q����k/���1�3��(�5Jr�ߋPY�?��u�{ۦ�Ȍ�_�?������4��MQ{�6ҹZO�ɛY��/��K˝�wU�A�*��˼%���\�7��/LrH��M�L��߈��<��㦿˖�;��FO�gL��-����S�im(�95}�u���ױ¬���m����d��z=��GN�� #"�Vӷ����3�NNE?�c�RI����ە��|����}8��/�
.��#��0	�;�ߵx�n��ʾ[������xs/u�����3�c��g����K�!����Z�L� �,{��g�d�*&��	���\�H�T�����Y��L�Cp(0�Sr��m���ڠ)s�ͻbx��\�XK��˼�($u~�|%!�^t�Y�+�2�\Z�pӇ��Fҙ�	�e�4"'h2�A��S��`J�]J7��fwq����LVL�o��W��AB/:G1��g��R���j���2���y)0��D�-��5$�~@�F�dҔq����8��	v!��A��:��rV �+����� G+#>��uM���ȑ;�ӫ׉*7���7�D8�6�>�]�銻U�v�����䡫+�,�i��;	k����Ln߾�dWjMGG�h$�%�`h��R�F�����҅�}���b�&:��V��1�m����;>�t.�t�R���iQ������`7���i���g���'*�8���@���[$虍�^��:�j��z�����~�ɔ��v��E��-�C���cG ��s��p]�3�P�H�Ф��wDa]J��N?�G�t�;��GUϞ��F9��;	�ti�<�����F�H[�$
��=HxM�g	���:/���R�� �<���.���D��$F-F�ގ����'G*������i�V����AJv|��-���'����Qg�g-_=ԧ�jB�.Y��8D�>դ3*?��'s�DH�{B甕6�2��صW̠���^쉖�QV]��#�qe��dic�g�f.��e�y1$�T��N�A]��g��O���HF�H�w���z���β�D8���Z���.'�$���~{�1_KB��E������}ʥ�:bZwee�z�zG��:B��؍vJ9*������5�ЊOC{i�p+����*���:����FN\ 3H�u������X�SلrY�R��iA��D>���Z��zܥC� ���e�b	m�.�����͕�\�2!�V6��"��C�k.�j�Oы����TvZ:���58w�E =Q$6�hqw�Ҹ�mX�a���:(C��p���B��]�­Ji��/}
�5yڧ
`���K��ݧL�jp���>�S5�Ct�ҿ��9[)BI��@%V]�:�q���@�Pɴ�f��j1z��/�x�f���$\�DS=�xƓ]}��E�am�ºL�>�����;�����6�Cj�o��o�&1�J��_0#�k��+p�u)nMǲ�52Z�n߹�Iq2ǣ����lSb;+���(���}��������A�9u8g#{h�/ݝ�T����Y�z����Q�Gҽ�p9�dsn����G��c(�
2�N*B �P�G�$��q����}#�j�������fTq��5����@#�K��Fw��r���<!������o�گB��imJcnZd(E��å/ˮ���Uӏ��#[H<Q�����L�? ��d�F�;�])*��7����$c�����\�;�Y;�굆̶g�B,��S�٧���w�4MR����Rc��`��U�s��"c���܎3�[M���� ,Tm���r'���^&��(���C˥�G���l�mGg�2�1��O[e����Mx���+�ߐ��70�����f�$C4�԰�.��ecV3yE������觷X��ڝt�Ĳ���K�N�KxGs�����^��o��v�
֧=N��Ct'��~���lQ��a5�xO-,� �h�� 'ɀ�^bx����_Qgu���u	{�A��SwW����Ƹ�_������˟b��K�r��� �@m׆H�j�Ҥ�(d������}�����lG��v��a���P:��R��W�JΔ����)/5^4�x�#M��du�� u�L��f^�{����F�.���v�t�J��)P�U���<.���kB�ؐ���ñI��<�Ӳ�( 9��5ύr|T={�.�fő���,9�_�;�^��������x��EP-��*[��T}��;+G�X������h+��e�l�z�TׇO��'��<���6���me���c���4�R�J#��4>q2��1I
R]A 1|�PA6q��[v���t�@ʼ xЕ2i����)���>�N�F�oB�k��T��i�����塽�E|R�'n���-;���'�
���@�z�cE�b�EQ�R'<��3"+�C�[�n�\7?�P>�
*���]����,+G	d�#��s3�����U{�5�kQ�4���i��h|"!q�߈<�Xw.s�]D�[2�!��w�fa;s�'��.X$D/���OzҒx=;О	>����M�N�:�v�'Gww��U[4�MC3�ʲ��x�f�""8�J��N���I�̗OǺ��D~��k-������D�=f]�O��x7ѕ��>~,x�ĝ%~*�nLKڸ�Q��	��vӪ\�,�����!��2�C3~�0N;�W�m�R}�}er�郪�T+v��-�F�3�B�����Rɢ�j1�M����}� du0��A������Ó7�z�#��?��.j��x�~�8�EO5���7����p	�Tu�S~�`b�BI���1���@��=�{�#��/�8'��V��_���[���X�1�Y1~L��\����4g���KH�a�"���8�X��Ϧ��t��BMO�MH�eX���Xנ<�b����μ��	ˋ^Z�ӱXK�d�((�z��K�P{n��&eD�B���/��24����%��(4��y��I�<�M���*V%�l+��{|�j��o9�kU6kh�ٳ��m�.]�C.4��^�WŃ��8�RY��'���r��)�p����K�U��Еx���Z�lʎ��2��,,W\S�Q�T�W����Ow(b~�)Faϒ�>�W�9y��s��P���h��N���W��������$&�����)��.��z8t�^�����@t�lj0ǈ�\&��
�Lݣ��o%Ҝ�Ѷ�P^��W�I��2է7��*U�&�&��1	��2��%0�D'*C�r�/u�pP���h��4��<-��]�]n3���\���h�@0x��˩DݐHCO#0y�R���]��-����>��N��G;�u�37����
(@T�%c����~N�1��}��4�N.��CF3A����&�Q�j�&5���E3�d��;t����IԪ���3��<Xf�wtN���JUऩ{����Nёi:ɪz'6�%��+�=],�� �nTCN{m�8rh�\Y���ļ�D�A\Ǔ��d�ƶiK4ܾZ1%u��`�����D@&�����^�mD����Zt�y����+3����s�:�Ӵ��HY�Vk��m2yv2�ݚ���dW���=��v���"t��VA캃�O���&�0�����N�,:T�9 ��B�=Dt�b&�cop�*��b�w"F-p�X`��z�����>�槾Ж��S��a�T	�v�n���ph�W	�
�20�]�wi�JNLx��N���b�1#3>���
�f��b��� 6l
��k�*"�����׳�V���(�7�2X�e4tK�݋��!į�x�*�Wf�=)M|� %��*�3��Z�aunxŴ�w���T�n�>��VR�׵��u��8��4�_��{���IEO�-�ϸ�j�����hp]�y[C<P�&����[)�>������yl�K��F���������G�3Jݽ�,4�0�?��j�ۖ���/:y�w�͞�S�8�"�� ���!�D�j+3.���H���	Qu;�U�+65�"x�����1	�¦��x�Ȥ�
	�I8�lo�*qa�?�M���Zb~��7��|�0�\�x�Ue�����*�,�eb�k�^i�ji��_���@WS! �F*�_E	D��B"��� A�L��q���l�r��ha{]�E$fd&y,�a;]�����C�+g?�ˇ,�@�q�|@Q��8\��^l��.����
~�r������.��߅g@BH�p���'X��y�V���%��Zhv��̕��Vj�@XЊ#���M/��#�x$S� ��M��n ���h�|p�)���5\M?E�>�=E"a�^TA�ŐY�^/�O��0��}�`	�@�\���#��O�$d\�vl�#<���2�ʽ�G�=���u��%���D9�P�L˕R��
����>[_����;��XXwPd�.���V��n�M�A���	��ux�_�s�HV�����lu��]C�	5�/PC΅N��/��&n\�tYw3Y0���)��U��
���A6�pA:�����(�Yg���2��a�#A�%�U6xN�'�	g�B��qP�yY�@�`�O�Y�W%��yp���M����(��^���FĉA�C-�D7�H`+�n���d�<<~�_U�����::I��P���{�x2B8r�$��vI�ug�o�b�}%��պ���\/U@P:]��n�ʂK��F	]%� U���g�^�uY�V��W�Z�W9� O�i���\���sx���vSwK��E�>J�$���q<qg��uŝ��U\��KujKh��P�Kv��^���D
1�4DA�8ח���re��}_��o�h���]}�;���O�,����w:KoRp"����l/�IX�`%Q�=(հB�y�=m����2u�f�,�3ǹ'��$M�,���pt0w,0�}�f�=�Hy���S>�q*�YVw$r4g-��q�;.L_�qo�`E�5Ed��)[/�%��S���n����2OW�����ziX��#v��LgF�Rx�L�����M@_!�71)9/�D��xOH��}�8��r�L�;a�	�E~-ǹz�W'�>���*V�-��DG�q��U���d]�3p�J�e��{[�	���WƉ��R����g�i���d%�z>���ܐ&��h��c{>w�- ri @������=ևo��G^}\�m�`}��ƒ��hԞ^��:M%��2.'O���o.xH9���Æ$�����pd蟟��[~�J7�����}�b
RÅ���U��<n��zxUV�4mߑd���k2L�-�$:��ޑ�����
�(mc��n2�"\\n��na�wJ{NV��aM�I����.o��B-���"�g��(��nd����Ȩ���0���Kؠ����:4���i��UHm�)���˼IWL�����mF�~ڒ� ��D^r�����oy����U������~�X��F ^i���1 �?N6��o~�°���*x꼑�4��ig}1�f\�#��ל�����I(�G|�RhԤ&������_�A�������,_OT;�=tL�(@+��
b˙����?�a{���Oȗ#S�A�h�~�m�٨-�{U�T��r��]�+��Fg����wjg�r�oc�iK��l2.�(δ����=#7Re�c-u���(R*෍+�
�o��di�5�<-�é�i�c@-����u�T~1P�7PJ� 6$#����y�����3�%�����;$W�rH����)��o�����>�����!���M�%[O�Z�ScQ-���mF�#P/q[���.���K�u%]S��� U�2��/�ᚡv���{~�~��XE֣pw��C}R�'�}���v�Vsch&K�Sg˜k��WLEֿ�o��M3�A��^0H6�vV���� 81�+���x�A�M0~Q�9�{b��^D�#!/�F
S�A����AU'H0���\�ߺ9%�e�����3l8-����w�9�I�ֲ�׾߰+�;�hK���e��C&��g&5�t�9N��v���l�*ZE�Ṁ.�@=)P�jw-a�*�?����=�=��9n���ڦ�N�݇d�l���׃s/��:�Y�ýjk��T���h��K� ~���5�k��j�!+=�����ob�����lMW��0��7P�]7!NZ("ôl�%Mفڙ���q^�壐�WMWY�g�B���\��8�:��[���S�+!�v�|-rWC�m����H�_�>�,�X��3*�Q����6�>DY�V���gܠ�e�/��%��5#rJ~��"��I���zʭ�`V�r���`�N�G��Yw�4˕��Ȥ`W$�U�eg�		�uⲎ��`(
��ޕ�N�����T���
�\��v��-��(5N��,)a��U�ͼjuY93&)"9.�~�/2K[ou\�d��i�ڗ�sk���'��������~����K̇�S�ac��r�/	�I��X@Db�q��!����Z�V=��y����F]W�ϡ蕫�KTgD��	-~�0hA�}����գ{��L�d��u�8V�Nf����Tgq���N�����-x��bAM�+pתp�JöO�G��Atu�V�Mt�Ï�WNZ�&6-.�,6rt���������/i�zn�>�=��� ��)�� BT���/�68�o�`5�i?�j]^o��氲z}1g���tGz��7�ef~aH��fOX*JAQ�-~��|��Mjb�t;�U���G��ƛ��1��[̓>4���N���=W����3�	н�V}�I	����e��I�w�h3�1P������-$�h�e��q�Mt�I3$z{8�X"OIRC��)�d.���H����"�`"{D��h=�1ê8����3�]��,���%����=��l��n��<���Re�T�>���p{��!�K�CAցZn����a�䶮-�\2B�1���U��5<�h�3�Rpi��X�$���3�ɽ�)��:E�m ��.q��X���d3)��R��=�Z�e��a\�c��4B�9&��=j�o�� ��L�w���l����貆��J!�~~ۡ�Ȯ�
<[���	`��|&z�Rm�FK2I��׆$7�L�6A^��؂	�T�s��{f�H��%���ʗ6_Ð��^��4$�����:�c�0���-����(o�qp��1T��m\>r��M���\oS��V�
��3
��#��q�W���N�=����%��#
�L��f:@ ?\I�~�Z=������u��_~*!{�ț����cP�4�8�<s>t5�1����}F�>7ɎK�s��)����'��Q��X�ܾ�S�X�!{�T�u� ���s��h��(����r yEb�Y��w�0\��g�ppIf�q��|b_�3��ѷ���X�0
��RY�#���_&d���@
3V���P�$�z�E	����qɑ��v���Z� ����ѕu��ty}���=��F����]\��-|��Q�20z��X�e�G���WX]���(�opF�w���R�ɸ�� �Y��̈f_0�
K�3w��@�T��*"�Oڿ�5��\��h�&��F13��a8����Jx�M���JD�)�75pڰ]������E grW{��"��;�/�.������0{�Gg�D�ZÅl����qS���xO
3�P��q|{���&q(n��.zF�P�+?r(^@�a�j�6���l���}��[��}�VN���a&���A�%�)?�}�{����{�1:�ȣ�"��K��b[�b�^]�2�����FVj��4�.+6:\2THgQP�c��`pU�	҂h�����?P������?T� ����� U��R�	NRK#�O�q���ڱ`�>���cP�1�~��Kr:+�:*�R�Gf�5�0Vh"��k�#�=��ɾ�ʋ�-�]���wEزD�M��.�Q�h�I��`���yA��n��*R�vhh�����+���Ǥ�^`J�>��-_Xt����n!x֎X�Qp#)�
���u�^ͥ�������x'�I�}\�d�N�}����D���h�����;?�+�r�L���<���>��mh��\���?&��/W�:��)�䕨Ǽ����A}F��Ƶcx�2�p�h�@w���J�w@��kp@k`�����NB���?��&RU�v��u#{N^��M�O�?f;�.kã?П�j�?Ő%X1e�?�܈f�A�9�@x�}�����Be��0I��b��xr��=K��wA�ek#��Y���s���y(F����)�Bc����6ُX���>��pel?��� �S�W:�[�^�{��;ձ�@I��t��:�3)���Wj۵�$;����߱5��^�Ĺ��\е�� {,�B��;B_W"EA
W�?�Y���a.��i���\��P!.�`�ۅ�$��۹�����{�������:1]�q�YX�+�e��ۑDR:4T뗬tB�oJ�y��v��!3�����rs�%�4�4I�g,���T����M�ϔ�AX|�Y+�5 �[��������N{s�R�Y1�NY� ��x��\k�ь�|���g�W���/��l٘�f����D�}`�-F��#f����=΃�(u�z8\&�
'd�:>�I��N��W[|%&��5.�^t �>]a�sS�L��J�r������Y�zW�:�ʍ���u^�~xk�a��z�^���T�}��L;�E Aw}z�c����$k�4�KإF��d�����V�T��(�����mëG����ψ�n��؆���g�Lo��p��p�lVj������Io���Q[��G�[�!{�3��툩�c�C���{��A>��۾Ha`��}�X��1���T��m���Sr%h8��[m���كؕ.\`�U��ѭ�A�	��I51E�R��X{�}���]��ߒ�<csA�7.�|iel{���8r)gM,�Õ�g~�}�\o�)����� "�Mb㭎(r���'��^��#X� ��P�K3bK�"�5.��?B~| @�2��*�����nյ��_&�b��@�OV�|�]R`��yw�h�n�U4˽��q���=�7�玔ej�t��-�-^���hR����'(��
�����������S�ϗ��&(�CV�o)��\نs��Vý�^�\C!�O�^�C�)��
�BO�Mr�T�]1,,��u��`F��8o���L�$NȻhE���S'`�K��Z�K�/jmvx*����ɢ����TWr�Țc�+_�"����6��%C[N_�%5޷���{%�k\�	>}�l�٣�䳉
}���I�%yеݔ�vʃo��0����KH	�'D4�ze1sE��Z5��ӵ��#�w)�U����=2(w`b�w��MZ_ɮ�(�c�?$j���Р13O����I���:=�����
�P����-?��Ր�G� ������3�#�w��4~��l�[���K��cZ�]��\ XU��/F��T�C�ė-ܟ��D�YZ����ZfC6m	(9X�x��L�+Ś�%,�k� �G�����T�QAP.�rvp\���SU����������'F�8�Q�9x�X?�҂�Ӡ�۳QQ�t���T�h}�K�a���v�<�`�o<3����Ә����
��0��]�ג5�\�*T�x�ۦ�U�RW��1X�!�X���z �\RM�zl��0�]���-����������W�2���A�8�t>�>���P��ڏ�|�G��&�Y�%�R�ԅ�w�yN�HXB����w]	�A���rY��>ݲ�ٸ�`�PG�쪋��-��}/���/�����['@�b�c��Կt�L���5�͖{�Ry�(��Ėl�Mx�+p�XrX�ꑩ�r���k0X��{D�صC+�*>����E?p�g`��	P�K��le&<:g���h&cBDo�J(�0���#r�,ᣴ�9Lvy�[^��Om�����;�(�"�]d����d�\���~�ը1(��O�2��K?�H�U��p-Wc�ƕ��CM��?31�����E�!h�0\�s�B�9�]�y7W^<�v:S��K ��%�$.���(L!��� ��$z�T�D�"
���ow��:z�A����ш�|	8��E���'G�q�,� tG���d���/
n�)&��r� C�y�e��P}�}����Nn��R҄:\6/ŜP�u{y 1C�����*Z�� ��ZޑQ�����rT�fۆ�@B�\��Ļ�ZA#g@�H&�3�D\(�wU�ҍ��}L8ǃ�gZK
"�l2��wh��~�J� �6D�Cˊ"���,�ǽ���^�m!p��֒̿X�3�QX�����i���j� ��X,��y�3&4�u�a2;��gÚ:i�}L�m?�`x��A�֋��[Wew����R��{�����_�����}n��xg)������@��r'����G�[�E)��o��y�lJ����l��cjI� �lk�
-����̮v��0�2��F~$ H���$���}P��G  ���3����h�֚g�=օ����9��Aګ��Q�U?�8�v�?FK��(Um@`��ΗC��ek���U��,��!i�S���MEZV���T{O�,�ji��G��U'9�$�Oy���~�񅅵L)���Β��w���[��BL���� �S��嵅��fj���$Ȣ������K�+F\K$o�j��A�UO��|s1�_���f�Ǜ��rUu�!em'౑����Y�N%�P��B�x�p�|z �.�����CG�uzX�En�G��)�c���?U�sΏF֌,PN��*�P��ʻq���w_��H����\GC�j��X��~�!ؼ�C�8|R��58��� e���FX�������\��Q�?֭�
_{I\��_4$�k���������C�g߹��}��'���C��Z���!�Ἁsn�(�����ug�&����O7�M�S����^cO�yO&C˛��	��l"��,�cG��[�5�5�b'j ń
�K�&G,��b�RQ*�F'D��O+��:�}�d����L�������+����m�#&�����8
Z�)��`&gV ��W��c	F�����ߙ�&R!�t7�۱|_'��⾨�UAׄ���c�tk/De=e-�"�q)ߚ#�$f-B�"̯�;���.lCQ���'�/(�g�f�	z ��34`6]�~Q�\�Bۂ��1L�v�W�_���lv�N�!û��XA	��4�/9z���)��S���2��+***Ǔ��ӫ�n��l�(��{�"�<�O�&:3F��4����ѧ��	|���I�?&ϩ���_e�[����hr��c����h���[�Xb���<���E!���;t>�eh+��)�\D
�k-|�2%6��:�����Wq��t2j��K�j!d���`���0�s��
l��J%dz1�o���ݎ
�I�Q4��w6�d�b"�����O��1���a�]Y�C�l	C�B�|�u�S���x���E"�@L�s����.oA;6�_R����L(�Zv/�ڐ>��#�6
E��<#�:��VҊ].���"Z�#AC��t���Х�2 ��5��f�>��h���Y�N�}�n]}�LŌ�K�����M:-G�ui�%���������#�"��q����A��+b"���6�g$w�⧉JY��&b$3E�]�Rq�c�]e��l�(�_3~Ԅ=-2a��<��@ ���s�;��iX���-A:��ɟ������䴂־i#�4DU
�����)��]ѳ�0i���L��R7�>�*��Y�� �P�m"�#���(_-��6c%˝\��F��y�ϣ�~�.@���Igي� ���/�� �VZ
�dy�b 84�k{V�.g-h�P���L�2p��`��m���pw��5i��Sx�m�L�Br �ۥk�E}Z�Ϧ��,w��E0ze���H(%Zq:/c�D���M��E� ��~Ҙ��x��]wF��Q!Z�p]���}-?6�S�"AT^�)y���r��u��į���PL5|��v0�bN0���:B���o\���oŜx�3�Tj�(U@A���S��!���r�T��ݾ ;�GE�x����t ���'(C���3���k��U��\��MvTֲ�˂���S�W{rwr""?�/�����2YRh��PB��LZ���`A���H��hA�/�S��:<���e��a��U�>"��xj�[s���Pd����͈��R BZr�i��5M�g�C>� �Rz6�
@f�ć�OI���Շ��y:�f��#F �����3��8Z.Nt4[xDHצ�g
m}��3��y���V�	m�=��"����W�PqnFB!�˶Y������d���/Ն��[] ;��Rx��Ԙ�z��Jˢ36��M�#|G�8 �'��[V�z��,]�3���ELD��
EZ�Ase�i�@����yo���D1���12uC����� �/"�n���9.W4uyiь�Q�E�a����t�V�Е`^7P�����H���0�[���	U/���(�� Q�8�針�Տ1�~��]���;O��AX,UGa��(Kl���	<�:��n��-[xz�F	6��/���qcF#&u	<l�Nϴ}��LO/3���t��i7~�N�g��u~E;Ď=������E.76)��g��ck��M�7�W�}]j&�� ǉ��UWZ�-/�Kg�d��H'U���-\d�!��O����[�����O�D���yuˬ�42��j@���"�24��J�����]���W���U4������8S�=�| �Tv�:S�[J=3�:ff�S���#I,x�G?��h)�'��|�."F1ܳV��;&2j�A�0�#��%/&b�`���,�J�1��mXtQ�,�݆es>�q�5��_�7��OE��T��o;hS��>�8sj��C?��-Brt"PtT+^y�^��hnә
^�*�w��on;��	�3Þ�6�3j5J�U8hD��i�,��Et�h�rQ�l�l���~'i�z�SV�^����0N�D�h6m� �r�;��)��/�SoX��j)��:X�{��$LJo�����3���-�����}�q�pIx�����w�ߋ�H�G��
|����歺���|���c���[#;3T��WCy,=�W���mH`��W��hޘ�<�^a���9�%�-R�&�Ƀ�.���f�����fٲ ���9l}S+�r7��]����@t�{�{��a���(��i x�e����}ŰlI�Ye18�v�p>���(4C��f>i��� {��p��14<�j��2� �0�Y�]��Oޙs6������w�������o�A����$-!�հ�E!2�Z�&��t�+*�������(��LZ����H_�?w?l�y��c2�
���U�-~w:~��`�O�'A��p��)���a��@dq?8��V�Hb-.�kˠD|�%��j�r���%sP���U�Zb���,��R4>�,�R�����-l'(]���EpT��s�y�煁�J9�~`��nz�����zT_��|4=���J(��� ���),	D��.|h)�e��|�kP��g�<�l��*�Å�(� |�
�SO�i�'�.�kVT��*�	q��j��u�����>
*�cl�>'����F5���(�{��@��[,9�8��Z�m�|�¡�i�t@�U�� 9
[f;nh� .A�NGo�e��ޗ1�+���zߤL���.N�Z�b�J��;W�Om;u���}�$+Q��i��m:
�G��[�%�0���ƕ�垇�G��?��<<\�vJ��DK\�.��� Ⰻk�� ��2���Z;�g�ܳ6�&���-R;fq����.I�*����!e=�b� �fH�ʴg�;w�\��0NO(T��)�a-	�ΛK;�%ٶ��_z@�F����A�h<a�9��e�?�D:�Y8����]Ѷ )�d�7��)r���c�i}]��J��	�q�N�E����1zͪ���p/'����j�Dޕ�Ķ��w0"��G+�3����Z��@A�{��K���_�Q�{��,���{p&W��Ղ�N��ŠS�~�o�c<��Q����w������4�:U�8�}7����Єm�{c�����Z�W�N�2z7^Z�V�:N)��X�Lr�c���{��KH��k�PJ���xgȠ�U}���#<������7��o��c���YD��,�'�~��Ս{����Hw�V55��t����_��M�N�YyCn�\A�D/"�v�\�T#���M=5l�c�5����M��v�����.	�F>[�]spP�(A���uwz�G�R[lBy�vb����&�`ƞ��Ãl��F�X�L��Nwp���_�l'@ �+�]���������j����E(�G�y J! �qƟM��eݏk����i�#Fz�:;�V���Ҡц�!o`Z�c���4��3j���H��4�ҚU.�œz��-,;�@�*�щG�$nR�Y��S�o�*#!t��/��D��t�A�_�>5{ћ�b�nu��x\�̈́���;��[P"���F��x�^ �p�?�e~���%Y�#k�sv}n_=��g��(=��{�/l����{,�&e�2}��m���_��Wn��u�@8�P�� �ǳ7��i���v 6"gn9
��n��"��&�f�=�Pe�Y����~l����8���{}��"ad�?��ي���7�J�KE�+�R?�<�(bB����*~/�!�� 9A�gǐF��*�SK�U�=���}�^��u���b�{oXC���k��@gEzjɕE�w}�r`OJ3y���#�ٶ$�kpB�r�e���T*�?�n�w/:$]FO���mt[�Vx�3��"&����o.<ی�a[�.	�}L��v�܃��4����� �R�jnRтZ���z���I����g�%
���.�(!/�����.�~k���yA�p�Cd��!�@�E�G"��Q9fp<��ԫm-ak����c}�.��Mw1�M�Hy�c�X\��[���m�4%�u5l�;tS;ˡ����m��!,�)���5$�rz�֡�4V���"w�������&˹��aFe��������Ӆ�b@$[� ĩs�(F�0Y�t�e�;iP��j �ӀUT+u塨zH�*�t{�Xz��X�q�q%��
���E9Vg����d����ߨz��^i�bF���G���,��0@��P1��G��#heg��z���M������4ݼ��(��T����a�9�RڋD&��f�O,/�/a�l��e�0��]	@���ƋY[��mds}?�"��KY���G:�wi��w�W�*O�XGI�e����;�і�������jT$|�&R�� �;�>ّ�S��мU;��o��09$&4��=F�.ԆE��Zީ��+�`�WI�7�;c�,]j�e��.�+$�m���iה�b�<�,f��۰0�.��������rI;w�\:�DL(��ʐ�ME��W��oW�ˣ�%��-�Zn�q{/���z�W`�����8��k�\��0�gOU>� �X��!���a3DÑ���u#�I]" ����Vޤ� p��Z_�4��"dHmJn�@ͿU�b-��:�?H��+#�����T���k4�L��©J̔�3�����V��xu��ŏ��1 W��<'��I����%�{���e��*�J�0s�\?�m�������Q(@>5�k"V;�5S�� @����0��HO6q��k��A��56*.�����>f�]$
fR(�#E`q� 1�E~�0=�[v����T�E$�p��Q�DZ�|�|)��%^A󝘢ɹ4��_���)v,Ӕ�۠��ӑP�ٻ���
fg������'�_��IU��Ȋ���{չ}�lX^J��<�_�8�������?g��������g�g��ㄪ�Q9�yj�q.�f�r��G����WR��:}H��f׈$b�dg	��l8,L�$L8>8DE�KzϋA"�Q-��o�A�ccx��[�+���-�v�Q,��b���hRs�ޖfK���z
�\�8�b�oN�Ҹ	�����ڑ��_"�PS��
�,:�
�=2巢B�鬌YJ���c�u�c�kR
��~�:S,��۠��?����m���dL,7~[��_�ll߄��dF	W���짼zLTy���¹�8k�P��wj;h�%�ݱj�a�����q��P6�!P@��2~���1	�۵���!]`͵V�k�\h�采�d�y�}�t��T�PT��ϒ��_i��#eD.6�#!��@l�dc���ϲ�gL.<�<�VrvR�SfU�'H�#�'�k���t��	|0�11�n�0	��x1�_��L5�Xи�gg��E�#M�R����5�0���S=a��x��ۦ���;��4����%�Y�6������N��tJ�d�K����F��X"���D�� m�d��9W�/a\W�;J߷)�����K�E�T�k��¿O����9���ͼY�ʈrj>#[�i�:�ݶ4ĉބ`�sBi��?*W�	k6����SiM�M�7\���$p�M��!K��w��pu��������1�b�;�W�: �^.Ӏ��HJ7��D��:F�6Ȳ\|���[?�3�j ��Ȭ�[F��}��@�I�5@D�.6��f�P~ݦH��)���Y�:��m��$��+�kPJ|%������Uc�'5HIA�I�i�6���s�L���&�r+�i�aor�_��8�ym�rT�	h�1esd�A3�UX����a��)��a� ��Ǩ�\;>v���t�"��l|�����3q��X�E�!���bpv'���9L2 7���Q�fH@����y��jZWeӄX�i�n{�k80�t��4�
�����6��g�i!�5���Fw��
���p�N+�v=z,n�^��N����0s�,�����b�$f�P=����֢�[��^i饹pe���Ĳ��I]�G%��N���zA�:�T���t����g	�<�f}�OoG��!�s�UNY���&FQ�_�o�JIc��E|{PU�^�_��^������<��?G�z\�=`�b�~;���2���� �`�2ȳ1B��(ӹ�
{5��5���r��3&�"">�'�|MoW�ՙ
c���K��L��u}/B�D�Hp>R����i?�k)�x�4i7Z�p_�j����!<���k�$���2;�����8��",��v!q�ep9�8S�S�vt��]����U�v\Cߝ�y^���طv�V.�T���s���.�8�'���[����IO��t��Z�f"6��n�����%i��*}p욚��Ax��3�~�ww���f۞��a�n2�x��eU������P���z��K4�w���������Q��zaK�Q��ԕ�cܤ�&n��ry
R\팙A��c��9���`������S�<D5�?�B�ƕ��v��p�m|	vWw����tP+��Ǝ�S`�"ͷv�<���4�ğ��Qn��P�/27����Z�bx����H��/��T�	W೔VT�B�m�l��OH�Q���l�&��m+V�r�Z����L�y���e��VWϟ�JŃ���N�#iL[5&�`��t��ԖEt���T�'I<~��9��l8�o��=j��2�M�p��8b��=��o�c���pXܶw4Z8/ޜd_�HC:��b��柉P���qSq5��]�%��y"kp�2�7�6k�
�����Ժ��?�3��F )5��BR�	G�D������������"�|E��D�n�Yr�J-�魣<Ӊ(~+�a�y�������ӹ��d���Fu�Г��y�K	g�<��GX����B<��?��9��V&T������M�QVB�q�ɑ�s _��6m��Y�ML7o9?n����B�Z��}(z.V}�:�c�W�*b7��X�����uՓ�T/L�F+_&�׊fKu7�`����W$����yP�����%H��Ŋ�N��K.�Zؽ0��.�J޻fŮR�yh�6��ȿkF��X�s't����w�$U��c0��d���Ԣn������O?H�׷��y#�7���2�Gsmo")m�M�h��l�a�I����$GPJJ��κfd�{	C�: I��E�g�T�jPb_u�z*��O��ps);���ÂV���G�NIZ V$��J1.0��mV"=	i�Ҵ�_�R} � J��f��jb���Ɂf�n}�4E0$�Ã��+�gh:��5�o(����(�%D炔<����{�"M3Zt��ך�n���Y�ƀhu�5F�+C��ar�P�d;|��r�1�m`�l�G+�u�7B�4w�\3A@�M�?�8? �U��
�<QRr5������὜��W �2kOג=�I�MMj�q�ށ�#��@�|^z�(�3�(L��S������P)����y�.bs��O)I6D?z1	EL�c�~v�$��); p��$'G�QR�AQw6���A�1����(N[T2X�{��P"	�����~��hS�s��<�=��=hR��R�
0��Y�Op(�/���s�η��aV������xZO��I���ub�fQ{>�_�e~��O�Pڧ�
��o9(P�:��۠�;_��{��読鸌[�5
��O��=#8�K0���ř���N?l����G��e�mB+^��@����U��_S~]+C7��Ś0�s��휴�Փ.�C�g���+�15i��j��Eu<�?�~R#�6�ܞ`�s?�(��r�'R�U9� 
�����T���=[6�)�[_�*%p�A)���_�Lvi52��8�	��a7Ȋ�ғ�M����| ��y �Q��[��[�1�0�K��ߗ��h��q���~�~4�W��Qե����91Y� Ϟ=׋hPr��$~�o�@x�Z!mWX��X����9�,�̶�TF�/綅B7��-_iwTv�i����X�&�����E�'J3�æ��^W��7�W|
�����}b���p��m�g�M�뵎�H�~IWҰTO�q*�!��RZ���>���*���u/OU>h�E(�|{��4�.�U�d9�u}DU>l����P�#D#��W'���:�h$u*/r����GG1`>�x�-PD�ߡBb� b��'�r����((��{��[/�w�{���,�=�n�#�u��sָ��p��K�veT�E8��!-���]�(�� ��1q���c`�G=�io��"�٫�H�D�� �fE"Ѝ
�������\����+��)q�I�ƣD�t_.����#�L����v��I}���Z����g���F^�ћ_ã�^ӭ��)D:�E��� >��r�{s��:¸	����x/zt��0P8�QrZB��>�]5���VK`Il�Qm���^R��q�bq�	7W�_N�,>S�!�D��Ǌ���LB��&k�I��h=MI�m)P7�@E�^�L�%R�Ny�f�21X?�c������4����5�v��h����1�����V��2P�0@'�Y�D��V4�W�J�fhy]�2�-zȂ�H��#dק�9z���;k�l磻��7ZqW�C���5�ʟ��b`,���?b������*pPI�$q3�gn�RE.��.IKT�c���O�["�mN��5u��G��.��|�cf���ld��	j9�!ut{�`� Yц�R"q�WB�����W&7 �q�_�PeT�<������S�u��(�h�XP,���	����Q8=qD.;�K��.�nD�ǹ��퉱W�:��I��>)�G ��qq���O���V��\-��}�V�!�eHND)��d��j��4�f�=��S���o�1F�0��\�vgSu�)A���z�wN��k�	�5Y�2�j�.6����Ď!DXT�}�_��	���:y�y�{����X,��8���'�B�8:Q��$�'�Ү ˟�%X~��к�H�A��G���MWq4ʎ�H2��	u��z?������0f,VJ���L���̠�!2��eqo�y7��ud�u��R�AӴI���ꆋ8��r�υ���F*wxs�gy�(�����7���1��4T�_���G贠)�N��]��?v���F������x��L+~x��\�S���`�c(|��.���ߴp��py��2�ҭ��~�^I��.b&/��R�6�aYf�}�\!�z7�Z^�1�%H��!]䬷3�h����>���C�ݻ�v��e�����h�����r��n� X܃S�w���G��7��C]�>�oڳg@�]�ȪKU�E�~�Uu���W�h76~���� c����x��N��O�v㞾<��,��(Y�>݊g&��EN�|��dUus/^3g�K��0af��7�3�\�;�}�\��rfV�=�>���pb��0���RFDc	�x���\��ϤFb!�9��Y����,�z�|1y��ݳ���Yi+��ę�	�)1�s���x��D��������hQ�xf��D���Yy����|�v٦��^*��s*��~n)L,�Ox�P�eIfv<�k���Ԟ�_�&�hl��K�x�27q�v8��M;�x@<�<IpEz��b���ZýA�Ѕ)=��RU��Y�����C@�+�ҟ�n�N۲4�ё_��XQ��S0v� ����D���5��b/���o�E�%,�_�3�\{a:��ec�NU�(׌��
�DX?uR|����RW��v�����Gh��F�OH����%��^H��!U५�;v�'���>_
lw���&kU��a�$cX��M�E�0��e�l�J�bФ�bV��ϬS�s=W���zG	4��i��.ش��mVQ�c�������|�]�X�4�ȥ�p�|X�Ϩ٤z3T�A��J�`�O�J�63�tV��5,���b3�TYa�[ ��6�,5�P.���r�6K��@������H�!2�����F���V��%y�fk����iD��.����
�!)�jp�&��]�$R��_�q����rR2�؋�I�$�G��1 >��+۲�xT*��=���g.�����6 �MW�C���a��VK�O��+�8h�a�I5"�(� ��
[O��:� 3�])9iL4F�$T�ѯ/��m�B�}1�Rcm�C����õ�e<�e�K��L�=(�R�?� ��f.�(ਁ[m=ж�q�K�����֍��)�-���4�X7�h�%k��wK.Gw9�E"qX����sb�g(�)B}�`�R{ w n׾�*�\��A5�d�����!�񬴬E�(���_7;�f�x"��1���I(�x�b�M�#/����a}�n���ɟ����'o�,,C3��.R��m��Y�rE��?R��\��ᙙ�����/�n�բ�=uz�z��j<�	!�n��z�$�~/=���j�?��[tj/�ͩV��&V���T�ь�n�\��1�pJe�H�*���M8RB��=�#�@��}7�I!�$�'-"��ܱ�O����f|�Ӏ��81��>����A#���`�4�b��X\�\\�D�	-��$��4�S����`jn�K�˭U��o���� �|7J��Pc�}�-��%�)x,�a�씷���ߗ��}uv����1���V�ML+g{�D���D3�H�D1��ʆ/���͒p�[���N�W46$Щ���]1�F�>�<��&F���6l�P��U��N?0��UJ�4!�6)����oE�zI�`М���6	��pJ�$��w@�{d�Q�w~�챒J��7���0���E�`��rbsb"�D]Q��3��a�Q�a2"�d��#����Ka�$�5�O�<����4��Y>�d�~G5�\`@M��/��w�C^���f�.���
a-3J�����������9�b �?��Y_H-oI���L` e[c�UZ��+�}�֏�A>)U�-����%�j��$�c���\���bD�n���U(,R�g;x�� Z��0��֛�ZԚ �R�Q���.DԐ��<�a�@ʔ�����@�X2� ��0�.̟����^[;�@��KF��B�\� �y��Pf',��+v��'�6�"D��v��vb�w������?���n���X��dn��J�3N�y�bb�?�ܥ���0O��ax����5��Iԉ謧��ߤ��^.ӷܧ�J%����f�ho�Q�TL��3��eK!@�E�˥r��i?]<�����&PLq�R�Z\1w�-0�p~�F�S9ep%V���:�:6]뛏�|���	O�����ꮋ��šz�)P�nR��c1�q�C��Ϙ����
"_��_�� Ϊ�!g�4�Ϗ�g��&�'C)o�!���5re�I��\�b,N�GJ��?;�[S���+ˍ�d���m��9�_�1��2o(�{ti����}"��ڟ��Q1�zX�ƂG��Ԃ�D�Nh`Ǟ�RP�[�HZh��+�n� �2rRj�F��"~�}�v�R�-� ̉�A�/J���}�Ƌ%$�^�m�v<x���	�n��ױT��@-����և��֏FC�p�Dc.�/�H~���+T�!].�����k4SS0S� #!��r�dr�cʙ�կY��Ӓ���,F'�X�ʭ�G����i��;q�,�0�r%���B��$1sq,W��B�ׁ���,_��K��#a��Q�GE&�1c�rNW=r[qǻ��W�Aiv�X�$.��)E�dR���f�r!��Y����^%��ʥ)�Ӏ�b��>�	��v���ɺ��D�QQCY!�,�v�1��ލ�t�vE�:ã*� u�UJ4k�����֜����e���Be�a4���Ra��:qV1>� 䎤vl�V��A�C�v�}��i��y0�p�����e�q%IR��V<�[�Y
E�<�K�\ʵ�%��a�<�6�a#�HJ�A$��z�_�uw�D���
6�#����aI�ݐb��t�q��#EX]�<�r1��WL�I��l�Ixaik���v<J!X$N_+W��D�j�M}�X��W,ھ��sK��*X�"�)�)��N��cB}Ύ=�Xc�;�>��s;��U{?)�SIT�@�
���NK�ji5bAt�I���E�yK��(��.���|]q���r�E1�����o��h3B��4pSٓ�����$���f�sy;�+��aẳd��u�aՈ@�$�H���I?րZ���wž1`0�__ՊB�׮�hvIs\�a J�	����tEܕ�{W�������`z<4-Q��ƻ�P�ı�i���B����r����چ���ɨ^2�sp��6A()8^�v�7����o���r��������g�Č<�KCڌϏv�+OÝ��L��U@. �mE������H�f���ՎU'V�]�Cޑ6��7��}r�gmSd�)I��!%K|�t�0zw���z��1��5Ф��n��ܩ��)�H��Y1�)�-:�	@l)��l�� #��y�{���q��a�|Ѷ�M�'T���ɒ�m!Қ�2��"r\����֥��,f��[��H;f�
�L�Ҟ%.(:�alfh~[ g���j�*��C����W���,��.(r�F3z_�(�Ir%م�����o��	d���,O��]��ԖI�vt�?^J	ܫ�Ln� ��B8��N^١.e���(���_A��O�ek'7�B�����U�[
�3	��&Y��9���4�ş��xGI1e�;�y~S�p�S��;Y����i׉>IF]Φ�����s����LUִ_�I(�\���yI��D
���o���0x�,�1�.\"������V���^����&�M����<���2��ىp�Q�E�yr?_J�׫���y��#ޗ%�lV.���S��)�v���{+` �k!��$�o<}.����(�k͌��6����R����C!��H�J�4y�-F���as3b�c��nj^���a�6����oG�s�wcՕZ/gޢ���Bt��L��=H�bFQ�"<f�9ܔł�Ar��ey2s�4�e�1�(^S׺�a��7��m�2JDm���S�>�T��A���S��A#0+�
�"�����	\�w�Ү$��r����"��f�g�n O�HF���-E�	�v��nP&`���~��T�fo%p��_Jg�Q4�[���ǝ����b
/z�+M�'xc�Mw���Nt�R�8@��+�lq�M;�<�q%M����S����l\}c��Q�[k��mK)k���il��}�	���c,��"��s4N
�ht���-�#.h{�⣤�-�i��f����\�!��Z*�5�5lf٩���a�<���H��?1�N�y�C($�?��!�c���W�B�Ϧ�h_eK�������D�Hǽ�q�����2�O��K��2s,ϥ�'���IG_�C��[�MB`YW����VN��W�=��و��&?���zZ�V�~��rd�yЬ�w�jq�_�k���M,n��"�#tc�~5�#l� ~���G�Ůof'|,�<#�E��!�؁)��&������&˹L���V�v3
S�	�r��p�BdͿ?į��d���փT�) *�,�����[�Fy�(Ge�y�����\�^s�Ni�F*�s��*�	I��QWPA��V���-K����R�U�}�ث�{)��nA��t�_� �H�T��C�8D��e�OD���c�����<hQ�Wg�-b�ݡ�S���(M+�S��ܱ`/m���l6b`Rw�V-D,�ꗁx���Bi�r=�ŧ�e~j�]�#쐃������F
���s��q��keC�!;�+!���P����O�LC�F�F�����+Q�
����h�?�v~�]����,��x�w�!�a<��,��� �_?=��/�G�w��|��&���[$�$�ϕ�y�P��������_�72�k��Ѽ�+�0�#�3�tY@P}�!�-)P���Tn<WA~�V�6���0H���ckɳqW)cǏ�D��?7fy��X��5�=����V噸7����̲s �q RL|X�j��K!�([��I�0$��4���}�x����0���գ����&!\�F�"