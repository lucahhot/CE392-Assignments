// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
VWtJ/pABBbwY+HAxL4r++1uExib5oXeH8aHTcMeycI4BWxeu+/CWV+e5x1MJlI4Q
TtsNMvsWdfjKLXYBXEGLW/lZx78Rl6nt6mY7LcqStF+nJLaW6PkEycq0isSZ/1A0
7NHANDfaATu1bsK/gh4U+2CLaye4viJE63OvW+HS4XitPtiU1/IokA==
//pragma protect end_key_block
//pragma protect digest_block
yLR8EApjV339G+Lk2iUugxl9WwM=
//pragma protect end_digest_block
//pragma protect data_block
zFJqfnGO4I7mi2mHUE0B1hfhdqX3WEyJxlxLyZpK7O6dGZJPeIBPRxaTRos6yOC7
AO7Tx/i5o3239Xpuady35R9+GtSNw/10jS5ZQE2GNerIb4y5hmwXqCWgpw8MYesh
D5rM3JwAqlHf9H7/6pphO5EX+K8YT9PBfj5z/krXgyFnyLFS7FVIQ22PNFAPJlDi
FcU1d6RvWIp2B6dWr32Cmugh5ENXzn6Vbnrchofol40Y2no+86qU0R0YHYJo+fwq
fbyTYm/NObuyipQ/dLfbpRfmYvWq3J2a/B+N+4JNJ9t3m7gJU8vd7chWBd0Q7vY9
NERGDFzHjdWxXNbKaVAiSfljfwtEWWcCPNVmOwjjlMXiV39IhXaeMT26+FdUxFOK
6v9B/Ws4YcEGwl+hKZ2Nq6eDMW+VY6KwAsDpTPb89JggwbaiSfWZO6r2gTfNCXc9
lQgen5hacLtlURvw6owdP86k+VMl9MLa9gZQHvZA3GZXLvA1LIzHRtFREFwVMYef
SyozZJw9QJ6TnD5Fb+RAqRVH7Gd259LfDiuNIvEjZqfZfrA6F6nkeAPUHb4FNZ/n
fOk1SHPV5yKf7ugvCdmPepVYGVcyD+lhPVX6VPUUaxpehCusV0dbRa6dITVZP/pf
U+L8mSqer3DX5drS5EMYV0+nQKHVkgCjRLx4LMYaDbB5l3bQOScTvmlJyNqVEglF
2V9Mwc4FhwcuFGyRaTvRmJ7H41Q0NSUiWvIsX5/NRFiwxYrpSUolG68IxxYUnwBV
AtdtaO2QgnmpidjbKhX8QlSQd9qXCrIUpFONMkCb0eNR43rMuGxGXX+ZnBwWspQU
MneyrlYeDjTWdKOrWqmhwh3R6NBl43+2oEBrQqSdNbOkHjtHgRl5/wEiLgdj+4+o
ytXo7cnNnO7orFpUlwq2Gu73K8ogHby4RWNUxSmlOhqY00sbdn8vSUEbUT9I88Hw
zwI/Z+7BCXQTYfWkckfKwwhxWzXm9Mifu7HuJzrTKbHRkE/NpcPL9wFnDLYOX2QT
wbx8W55l3h+obbgYQ17rj4TMPcB5xDZEg9QSGxabdIlgNpxXqxBP9D0Ra78bXEko
/4UMQrkouW6LqWnyBiJNLLD2kJo1v68w1Jx3c5gB47Zm7g7TDD+XU70MOVAapJa8
3UFzfK8cjFE6KDS/DCol/O4bPMIxEopeRmmNQlgdGW2IOB7Wi3v36k8T/pI8iYiP
YWKQnST7Gc1fgCEIG+RRlB2aVtJ6Rszwg79FfWaQ/UHmhjf1sf5aYtr9H63aekug
HJQkviYe7IT58xAN1SQnCopi0BVJqPR6UscK53u+RwdK77FCtXxKXJo9lnHOCBpB
flVuG4mGS8iKYsPNu5ILsALJ1bi0swdnyIbXHjMheBPo9Eq/poZK0ejS0DDI7LgJ
7Js7fE5IQ178lpyuj5PW3m0ZZzRF+IeilV6z96+9WIdgXprx1Mh30YwilLAGubnd
c491k//gm55N749BMe2qUVU2jBjBvZb3iQ+5sswmuwCI46JZPd6bPYDARAdj7Ak4
nPxqTpA7iNHqHDeHCqvTxW5Mg8BDZ2cDsmj3z6AjOtlATRCGTLzGqiU/7NUAMhYI
2CY7JJ1FbJIejTty6v6XJ0o8qqb0E4XdFAt8TlLczXboi7Vo4vAz2835uWgpFZQy
LlRNUA4PJgERNLhsqsT4ya/q39lAvoShZ63yLwJ0i+4clda6kiXgyLar1XZKhnCt
VPRANHYWfojbHN66SpyvLRcCPEO7Y8xTT3sx+fvQiWuONe9QEuE4j6XgSCFsp/Fn
n7yMCmZfBpGvQ3dPKRw+jpFR90k/V2BUzHvIlvZKaWzx/2kI3jkZnor+6o7D+3NO
WIsvYPC4jhpRwwvcEZ1HG1HfCWI0e7DyeMNRBC1MtBmBTBzpLBovn003HI7deACN
fwLAHYaapbcASOdaGsD5HcheTQsxUmrFL1dCK+JTOm263ImkU/HBgBZocSHYjUYc
rVHi/HD2ozKxq/LDwjpLJBfrfOV25yU+6SZbJCDVOjNk4S6M3qvmQr5SAmTAVm+G
GNWK7qwT1piI/xex5rU/fq/aPVvUCLdamTFu/xsaacG0wbELA8WG0MxjXTXg/09q
BhWX1j5THoD/HF+vZwrpVgiZ4elIMXFg/fJpyZ/4EL7nJDxbo4LZ57i6srhMi92y
NDbN19ycXkj2Wq51YyDxPrFQLOmKqT6XmvEqQ+roOazpT5Qiq6d4nbZUm0IdmN5s
G9BuCDe6ZdDF23tdLqniS+Pu+XPUd8Sjnoo0GJBUYCFpzsflIqfRxuul3Pmt8ZM+
v2lJnJfqXwfOz/PQ3svsLwUCvQUt88v/aagq2aQZhWGiy8vyYIR0gGdVKdVJ7pBp
zVwBW9yJslBFDcZjQXdc8NNoTnwarlEzPPPpp+7yPcZxkB3BpyNGh6fcyt7wNtFP
H7T89tSoJV4n1pQtiSXom3MQVxTLFJES2kKx1D0DvOz3wk8cC0DjmAVrMUC1dU+b
Vv2SJtT3BGz20d7Aws3z3x3O/nGsprNMBmEkTbPDjQtICOn5j6JPNasQqaHFROWx
ReGPN2pDUw9TlvEOn5unRmk53lBG1t4QjFlvriH5/ZmkuKvKoT5L/bsmNlpD7qZe
n+YgUaBG5V6QKGiewsX4vMcMlZ3SV1AST+6SIZnGbABinABvyaujMiGlClstouE7
R7iMB+9ehpEdCadTJovNHGMMbtlZtujQMG6UX1wpLBicnTOmjbIg8mgJz9Ha4Pyv
3YNmAsGLJbtc6zgca/tJyFQ6RcjGDZ4rR1QJuGKgx4g1VyVig3fkccl8upn8KRBj
zVUQHayaGCzX+nbT4ba33LN7C/gpmrSN/2BqRFFZBGCDJcrYj+LF+JRBr7DVe7PI
F1vu9/dIHTZPFukqZMObFfEHVqKO6RvBEk6+KRpFxTWt8qZ46RrzJzwJb0kUjycd
PBtJ3REdQ0Ji/h15eMzcwh+kqv74Sl/aToHEvba6KMI5MMLRI34/oVKPOUEIx7TB
NXAVE7gGQzgGBlkMR4xKVBxG3FzstVLKwZDwoOiy3pwjA+tfnAp5433ICZSpbAKW
jIwTNxBmaI2Ao65A1fzeVBsKMblghEOPlbyNnyzIEQCllJIMFy2FiYpSuB8ED/85
LQqUMQXiWIRQFSVWkPgQvf58i9Kj+GdQup2s0aF5tl8W6LxXRn5AAotVD3IgEQMJ
ThfPPOJxYDqo7juyFh7O+TJTksamqg0SD4pyeTXiacCjlkFIAtRkLxQuExP69+wb
qIv9Mbrp4OIK0Zd7DJDibh3leZ8LsxdFYIADNGgvivcWjC9+aKPiKqoomIApVk9r
OmmyWlJo0iSWI0r+UdOlNqeGu3mdS64hfMdQMxRIYdR6Syg96kkmtDAY8cgddBLe
ub89wlfrsbjiXJvKwMN419qQhnH+/LVC5cUJ66qYRKcfHBxQ42BcNHmskqE5FpgR
wu/OxRic8Fypb+iWKihk3L+RM+mds1uCPnbl/omy6nz7ct5d5bFqWr9xvHBktf0f
qzgYKUGEIAqCoIlCGdJdE5i4inqCJQsa4u/1SlvDGCH0XCreT0MV9rVEOEQ7G4g4
bfDjIQOe5KU/83SVS9ZipRGvS0sewxK3mGYZRO8G7uFhPKVc7FeLTJg5HC56vwWu
3yvL2gmJieL7xJpRBHlCjKhjNWJuyjrNzfPBbAcs/rt60aS7lg0zgnI8rLVUSzBT
DsuKTXV1AIWb5J/ASLX6mHuBvfL1Rq2ROt5CaGTDHcnI+ZHLxEiDtOe+bbiIuXdD
8Gzco8ZtPNfRimJ+q7kcFGBT+J4dgogeBt/S3MVNbuOwB5S3kIO4mC5rYZWnxFbg
6Yem0ZwuSan5E+tdMrtOrhw3M/NRJ+O+/+hner2/cH8PiMSiqd4hc/we1FS8sGPS
DA1QYlpXtW7sqbx3Kju4ge1aRHRA3JIA7LQWu3KdIU7+txxnMtc+t3GRHZn090Am
tY01EJ9nGRF/+yC/2rInz5hUtgLPcSiQ0ZjzOyIFk4mhAjTJZkAJP7WBqk4T5fW6
nvO1pW0SGXm2guBgQQfqh1MOjFeEgA4VI+R9uqFnRp26XvE5V/b7edHwXkzbVEFp
3oKR7I7B0b/rNfxTF0HA7zAa4DDo4coNq1VgopyD75CvSZWF/y/Jish+JN7Osw8W
XHG4FR/De63Dmw8EwR2kutlvaqQqTiD5RN4Uwrl6WXpQp5PRu6KnA2Xs9BJKuSk5
/2XqFXcUIRSGlAacskEAYjKoUXcrgIxMnBd92HN2tWpdmOBZ22mgm0WVGd7g9wpb
+69djeQHLIf/wAl4Rjiaps+ePRr881EAR3GBra1mrqpIWKRj1ugmVmo6EQJM3Pvx
PxFgP9s9FmvyGfbbPj6dtV5qRE7ANF2itqkrMiLoSxp/X0kPFJxgmARmgxDjrm4G
lDV51fUXyJcKkuJ5VNMpYvU9Etrsnq3KMcq272OwnGwDaDz3Lm6yG1Qsc9rImVlk
uzK1bLfIgnvLJIU1dBe+V/zoOHwbt+gBx+ReZgS/2qautRLSP9SoTlqVA3Sj3CIT
nnkiSCaJwNuiSMkfLVJkvui10WvJKQ52Q4E+NPmTa6X4ouLAHlxAUsE2JJgnxnox
kRTINIw2un26lf2s07LBHmYi+yZ8eX16YNgevL4aE9v4jYgn5hJU4jPblNkjL54N
fXy9o8P1qoeUKKc6E51x3yzhqIHfEF1hoTpCEBwEKZONfi2yfrDbJc3fvzx65rGa
ZSsjpVcgKwKSoIqj6op+ww7LBArB1HJpbvWPPUBSD7R00U+RRkeoLBwRQOJab2oD
3dbG8wamEYyY22h3rd9cAZ4Oy4xRuOWh8PuLAIbeM+PccXiT7m5DLUW0O0Q3vSum
wAmvnQ+NKrZAUmARTt8ZJu8Fjulw1FbT/Dlu5/Wi+K/vbPvMALvP7FXaveTkhiBv
3FWb1e1ttHoDwG5zT4ckVCWWMrS7yiY6jdpqvti7kLpEzwI8MJmjHXoRdjBNtT8C
hFGebB20ZJlMUTUgTNdcwKtEF/W7I39kKXbJLop2t97vewfCqIb7Nk4+kyTlOS/m
DRzEZsLZR0QcuUyLDVXfOm2vg6fi7C+dqahbSRRy5MiUyExQ2TA+mcQkgg48SsNP
RCVID5Q82pCJAu9RuPH7gmylkGWLPDg5ktESYSFwaPNj32H4nV06YOBLpQmh1QRj
6x/IEcs7lgZFVKfVoVyix43FWpphbxDrZo5VPIYSUA5pVOGdF2jdN0aUmGjP3IGA
v/U4c92lQ/GAXi7dfA6xohq9EwesUuiOTBGZT2PgArj9vL1ZwUlvN/FKhWHg27Kb
AtiUCIEQtQ/BS7DfGsyzylxGycQZSMGGWRBp3lOJrSDgiX3VKF79SnS/CsGmiFim
j4Hagku5QwlQfzZe3jxg12Oyg4r3uS5uXt3UXuDZjqXxkaMPw4TeBydX79nW5xT4
ztViImdtQad7Wm6HFrWE/TCbOlo802hv69qcgy/MlSf+inn7dLsCXJve7RWQfuf8
nKKi5TIot9aNiYvbczIJ0hY5wNC3S39YkGJz4ZRqxeWlWuI+bXODF11vWZKDB2Eq
E9wwaZs0BbLTZOZ9RRFVd8WK5ctv5NaAKs1LSmV24ms4CtfXFqCawICqZYE0Ok+W
RK0YuYdkSVe/M0jRXQGFlXcRtZ4Vt/loKEGsujn8YwAk+bvW+A7LCVvKPf0mQRjb
OD0Sg1XegOGl3EK5Edbbkz6eTxlOucRTWMlkxDPbY56mJPTBqBRSrafAEQ9TgdiC
ykqFh2hAZkaMeikDxVW2sZMZ+lmkT0vQyCSdHL+g+z2H5X84haz5SGVUuB7mXqkZ
vKtlMnbVR38Vu81g0bjm/QCeqYrJDHy+RYndkpZ0vu2hfL1hs7TpnhOfmVG5sByd
Sfr3ihV8Ea9JUK6af80H+PLrCPYxJbbMWI00+0+wtm7u3dzXMZYXq2SSqv7Txwrm
fkZyARBIePUoL0hEOVtulSdmEpM8gVYNi+3FAz0zp1H7AgfOHWHsh/i4s0oq6PBl
tDVagaUj7IlWx74Jc7YmWHTr43i+mkiHJpuWnHw7T2NA8Cypal1OVlVs/YHrZrw2
Yb8X/pzvbe07pgOM4j0XrcAbrJFy4SvNf0z6539H/XdJDnSqWKoReDsF9pruSPbi
JQ0d1URZ5BKV2Tup2uPHciH6E6O06XdJV49ZeqNUToQXdYXUdlHuR+cMONHdqWY0
vx1K71Z1wjsmppyUe7YrIzxKYgS8B00KApjYjWs7PZ211/FIDoDXBHXDexe12E1g
ZL4e70Dt86wP/vH++hHb7uU58mJGZA4ZjWpJXtrenHT9zxQ1XhBeN8ST9DnEN5A4
HQFW+61qkOfL1wNqIkrawDTbAsHgtB5LslJybbK9EtrzJszIqTDjh7iyEdG2Nx/x
5CUPZo3HrGBmHVqGnQkt2rdZKVEslSQlKbPESzV3irZrk7kid2TItn3HRpNG0FXg
Qgteb/WsR2U/cuJSAmG/Y030KsCaH74bf1M6HqsI6iHymUdZ1Aq3Dv9Qtkoniwcg
2WyQnzFO68Qh2bQl+NL9AW2MSDuhhPLo9sAkw6mtAvu76/zgcEWPnHldKFnC15X5
Jtt6rvAH81uJNtGXN5VCqQIuZUKi986lkqiLztREvv5Yree9yMEliJcO0uqrX4V2
LRjZLxdaJTrKlBpDHNUTMnwC4cujqJizFFfNBnuO4U55LomgBKVTZ1u71vSWxdWJ
juyJvpkqDp8raf0FjF798uicb5w+1JHQGpHBNC7YKkl7ZW+eTlCOYofmR8lMUV4N
SS+SAwnesjarEZoHX7RTSSBLyHmjPWy+wKEmJWJsKFpnb5NwPXabbLGtrs7bqSaK
yKdOrl+hvi3VhuV934UYCXitRF+8KaoWyTjyd7R04LujCtoKt9y00UjEXmamyyPq
n4I+Fx0SCUh7axy3R8YS95KVHlExd4xIL7TB/q6QUPNLCgPCo9ihVPnssB2uw9dQ
Y5EMlLWEmut/8CORRtB0uPVaKsuoOCSu9KvaiO4D2a0ohzAomCencGoywdm7kQAP
1GGTPh8LTf/3hvriPusu+1Z9LThoJp1s4EcSqGOfycAHGy0d8pOmIF/7ZnRZAu9r
IrJMhCNiu1wxhBC/mCDuHTQBHtEWpsB/qHGvMyV54eOhh3a9pvaHndce5hMN7sPF
LQ4b2L93zdlGISJQE0vEmltQRWvXxyHXgVVU/yDr+Qf0mxpxs/K62VbWP0ibhCnH
jni9eCrK0f2l5PxXIBE8SzLGXLuspvEQvHTgupY3lfsPr6whrjFnl+ahQFKfF34B
L/A/a3OsY89zAsbmHjJDhqLNKAiOQ219DgCWcXqIuxmdnzg4Tao0wKnGFAyNDivD
FzCYQr9NDKKvjXcI0uRSRHD6L/6iLJsO22Pl6DsFIEo6MPyTmtOV82dYwh3BSSuj
vWpsSflkaIqhhXKNUDPGuT+Ts2IgrXkIJP6IjzKAVgPPonO9obmjwM7Gf2O5SRHG
7b/2CnJpIQBRQgYsmXwbTCl/Ac+Tj2SmRNECJlmAHSbIDTcwhngd8XDyko/4tHCw
4IpWD6ohRiALcrRSJ13OC/QracbuOh+sHZUD+OzgaljAvHOy8nj93H72MEqm5b2H
p5C+hxZjhZvAm/+Hs+hZWZO7r1bjXSCZKlSpnIxNbO4WoROkELvNwTEC5Mykxsej
P1PjHk4MZVeVeNMTKYAkhZ/iN6ZABRNpvZQWJ1YihCKCeK/wOYVSgpiwDmbjv+sq
wUQnM+iTAwyfAxx5M5BdpDLOd6oeS9LvPwTg5eTwf4I1Q/rwpcqq+ertI1psniKh
iXiVysdIBC+LFb/05y6gom8njQ5jQ05nZ9yw6l10MxkHz9kpQvHnoGS7d73Q6MgF
U3FZxfwgO/eMBv72TaV4H81R4M+Hv6NN+R/kIXo10AsQSMcXzwSSxCkGNZMSCrfU
42HF15XCBP4wnyOLCX7CbL3e5Js5B3PUGblVGsI72QcLhPqc83ZToqdIvY+D5QIi
P1kD3OMQ/TEf67stXwRrEDUIWJCd77FvB2ewwbAgGwdHRzrsjj6FjO3/XxPU1O4T
pGoac22FNY8THb4gWdnCBddlZGGNFYELSgUcIqV5vE0Hfmm1YXZupggCvVEOODqm
chgvqevIeZp4Fdf1KiUj5ywk82HIb4m4xERzoSqEj1MXyzUVOk7sj0oDh+BmDs2L
PK5L2prkx/Pu6ED6vDx3s24K71FkWxjqVYyUBQ7rgLSs98I9a0a6TRiR9Fy+ehMl
n/hu92vjzkPeEWjeXSj4fv3G5LKZNFk0FkHHm5y+xJ+55ljnOFTGud45ARvECz3p
CYW3XwIGFZSbBcBMx6q5mezJk6UCatxruISTwd+lOg0hH+aZpvQN+INRClD7dc0v
rvrcZYzM+MwjxxjykTosparTUjPahkgXcArusGsdWlp45GIZk25UIp+2BOLjdCKw
yLn5mgXGurbouB1QCSJRJw41lgE8eMLdI3U8c+hpAm+9f7yW1MCBAvh1gSpJVHNH
EZZXY2XmY4Ze9Kx6vmrMT4lSPFB6tU4WCzSeUBglTFOL6917RAuwDrFXv9T1k0LK
NWlXjWuzy5HmTPelyMCW8hXNh24pSbk6Cd365EPIAakOFfigZlIt5y0xajSzvLhH
6KxG6FE+hyrBnbNtKl/dEpj+29uSRxeKOFXkyCr/tpOvZOx1ZFzZdFKc8F8dki7d
wlnwg40iZk4014DqmY2/Y0uFVq8FwDrJB27/trxiDFkhclZeUQGc0bhJKsIfZmfO
upAemWlIU8bxAKsfoISMd1Qpc9tUD4tXtIkfNP0HZOOkcngdiDAbqABlqFmaMp1D
P0CEfHT9bzfWTypeVFq+OREryo71mtVkeZFrWNqZdUwYsXS++cu0/vu5ldTtDYVg
XRUaKEy0bLH83wztdY9Hsw2meLKhWD40a8EPInnp3ffZ93faxVjsBfK0ApaUX5s2
1nyixHeI3wnOFgFI1BSv/XdcNjdYD60upyCK1+C3ky1STX2JoDM5vngcwbpnpQrb
NV9Ba2oIOR+NQMK+29qPZ8bE1vxnPI5wyppv7cIxRJ7J/06fCFIVjmAN+H98UV3m
190c8xg7V2lFfrz8R/8DNLrvKsPcDJM9tr6Eu/X/vTftrVCk53qKTYKfUYkU2qY7
2riBErKLb9ib6HfgMoea2T+tEo1jUQbHto0nftageif8lf2kN+gUwYbQDWLTv+Y5
7FTAtvN6c+d68TLsL/521qLm47FrNozBQ6vwOErDdXj1FnS9MG+taEjVuYzFayt5
H5Wr9tL5DY9stUbdY8UgvrVs2CBNmVUwR/fsclTTn99K5TlrOZv96/ERwMBYMFYm
UJlkZR1+LnYZzpQY7xUX/mu5UAhXVkGQ5FPLBjo0BUrCcskNUGOkz2R/wGq7ZhIJ
aEgbLWzF44wMATA/yHJ3Xk+ouuTb0mbuJX+2vrHkHbLS1/Q1AzYOnmsNSid7Rj9i
4d3H9iub3glt4MjOxKgpBORYyomKwUHbg24stF9/hKDLdCXTARM6bKZ3k8N60DIC
DwD7TN76rns9tm/2BExGkKn8C/pdVxwXeo71LF0I1/GvLXeJfI7XaGQacqqA3NZW
ma5O2mBpskBSRhDFsti4bZzqCkn6nMG9u+YIgMzbNI8J1XjcSIE6qZGIxiBUaz18
UmP5eMPlpwTvqt/GEdPBmdIeMu4h/zcQNHbKkT/T+eZaQDezpWgF2YAsdJ++CXrr
xZSGWX2xf5gC5Zn+6o4Ni05oYEC6tY20U4oJdSi+fdSwRdagJQokKgQpDVZ+27nT
DUAfAnvP6VbnRXWyhWTRfpHYyA31T9QNgzbT6xpx1ApKv+DXfwFu62suxfqPddPZ
IqoTR3TLG7jqkfiCGh3EleubVVPQeC4aA1Sg1StCvJYwokd5JKhiKlp2SLHmxNiS
sYu+b7e5IV2/eS6WnuzBwe7NPRUNW+q1pQKMn+6TV0PCj7zpAaL8r1fUMnjHHT4t
B6T1LvUM48W019oqVWMQVfZ1j/QCzQ8DRF8HTt9v3tYF8iV50BmnjJ/wcAqL01Ub
Uc+8zEUIy6tyPuerXo6Rhmd8ihABUczp/gD1Y7TAiBV6iXVPza72PZ2d9Ly4QJyA
sSTpl2XLg+CS9jCx+x4S65dJIqkM3G75LxKdjz5If35eigkk55IbiPCRwbZqPwnb
/1o9YrkOCk/YFfpZeiNkH0g1sflcyhzgU9H5DzxcBVtGpPJjJq20KIwCfwcEQkjh
gUUTSS035ZFg6GyHmJeLVzkUIXZm/ry2wQG9uztPEPds67m80HGjaQPXw/VU+ZcZ
x/NrEjtq3L63uy3Ua4cZrCUAtHXccaQSdpMy46TzfJ0M3PJzQuP+SBdy/ZFPdTdB
VQteeqUDRSiCRPNn34NrD0sqHfN3wOh0X1kb4N/Njv83Zfg6wqKUfRmayQlmpKC/
1013sghznOb6Qg2mNmiAN0uCAoH9OoZ35Cvxz9Kk7EWnQrS+Q1VA+28ZBlvmzbI2
/MV7LpfFYEXdTP7QXI5b1oT4iSfkZ6NEH3/GEEjNoO/MEAGkiAKnI9nQX4DQyBm5
LZLMXx3NVaboR2v5KNZXuHG0IeI8Bxat2V3WrcEMvYxV3qlqOSUEznTkQKjzzLCL
uJOuXSOoSJTkq6Uke0TY8HbI5nanf1ld+mZoIRffWJHk6a8+B1372b4k8AQo7Xqs
l1R/fkWuLgxustdetCi0iQ1cV9TXJtaRJAVw/JcZiFJRTxSpMIP4uYqXC46p7UVv
3fTyrTyjRs839r6GBc0RT9KKBSQ0xeiHFyjgruQlnvaNqIL0R+9CsXTuYJjt3gG/
1ji0FlW3WjksPAWvDWTLCsvEPc1ChMGGSTc0DSRuD+PqXj8u0KMZ3C/Tc+KnOM7c
3cSxTllkAXBRIZJbmQxjzv5laDyycSxrXQeQgfdry1nA/pgRAO6n8bMjRe3dN8uL
5MbasDlA46I3KIu+8b0zhzjGc56FXvXq/R6S2eEti27mk1f1a1DvrGYFS2tY4te0
nXQs9pIPcBWOKHJDpQip6bSRz5nTBbrto/yrtCeas1oJhDnKzXMLUrKvjqP8am3T
tuuNEsLwnIlqSLrKER72tW6a99icLBViYwyEZOLGmvNbzkvBc0eptCRxdYp/7L2b
qjracCZAScQ1c0sOOqGjDKcjeXegM9nIESiENqIIjszeZo1fke+IkUw/q3ptvP31
TvodL2vyFdT6RFM9iZd+ShHYK7Tc867SdPFNJNosAO/BGZtblhLwgpB0/S2cdWnm
GfSgWXMRHArNPcda6MclNw1DYOQ5nL+qjWx6it7zmBPdw8DcbGQOX1VBqMYVuEgm
yy6ylZvQcWJHlVlNItavEb9TWrd21bPDkWfbWtNwN3i2LHaamTg7yy9OPx4eoWYZ
k9zzGANiFoijtCAmKur5YKxkjHgLy9M8pFxwkDACphawXLBsuAmUnZv4kofG/N86
FHOMeQnRlL38iFSckbUagmazkWn7aXdlBoZ2vNAA5ZpOgEruZnfsBPpUOsx8w2+W
a50ZBQYDe/rL3NU6Sg/WpPKDovpVG+60JhOg0V/mq0JUV+txnd7Fc6Ny5SAK47XT
TabUXLNpUfuaQ0OATbRk/yB9BzqjkZvuArlRwtniOk//4qswL8e2epjyaJCRqsS0
Y7CBCE7FfhFjOiLJe746TMT5vW0+TPtT+g4j7QPuVl+PqmmA0vjyhPtTBACIXvE2
SAV3jIewOPnrhevvuqytDBkuWRLcDNFSDrF6HJ4PZ6TNU/kI4G3pbkPLWu6OeT6E
rLRgJqyfTpttCq5267KsnoEKPDI6RLZ+tC2ayCCHFWCL4oM+WM2RC+WyWpwHopC5
NSuRrObS2lKyBxjl+IXT5mw0AE/wG3SaI/xp3f4QzZ22EaBRjL8kHXcM7htZayK+
+dXUeWLIqWhCsDaatyiPY1porgPaZ8RKXbE1ciBwZrbLQ+/OQ5whERLZ/alwfrJD
Nb/KdHPTRI97ymV4cS0I5b2jD2GtcOSJwTwKMQmmmYyehdLVyvSN9r68oqBdFhMY
uD1vt2VqMgmcX0FUqbBDP7nki/ZSu+l8t+Vhn/460n2Et6xdMGI7XcnYQc++Y+Zo
+kU4BcYY3oUZAzfDNSLrb+kJFjNIpKpY+JFb4pchm1KQCVOLQv6d8Ov2hvaleyWB
W3t+8kP4QC5pAetIqSHWjMSm/1Vt135fN4N7yxfri0SPuScrYoLMXj+8bpxUMZbU
aG4533GD4CU/Qk8Qg4cQhsIAEctI/htZsJkG63qiH2F0cR/nO+MCCo1X+EmXtmWa
/mNttaEVMGZtB2sUYfCn+k1PSE7EfzgMjN4KbuH2iClWvKYW0o2oiQnHPjXjV38w
ha2btNSH9+c69OH1HiQzwKbJ33gYFdPOdn9WHJXVxKct8fGTlk3damg/OznVGBD2
Ykx25LMvAQ1S/4YFzZeUNJk7oCQ/wcEOFZ5AZnVo3HJsz8oZaRx5N8j45my3fCa4
5PRoWAV0QWRIwq8iHFNiZqVthE+wySkZo32zOuRUw+AeoYzCadB6IWqbjpaib2R6
quzTcbf2cspRwWB0CZG14fnwsPkUX1w22MuHvZqSr4VXE8QfxJgbCdHcSVI9eObv
ADZqwPfiGhNhNzXrTNC9BXlHouw3T3Q6eZ1k1sw/dyhIkz4iGU+fDiY+hDk+/Sft
N822StfjZT1DGOL0MAT1PqH6bYcVv74bcUEON9p845z0reoGPD9vXbiuCqh/y3hI
mhAnLiwVTgS2kJ1GeD+iJkewilIBtmpn+B1FaYIDF9OaJLUiKqGqCX4LVBvwxShY
C5qqbcAlqV4oahu5bNwUlU7/c9eAeMxM4Fwy2x+ZXPRxMqUw4GJlg4nd9E0O1Fm4
zH4CuQNYnYchgW+QdahgeRzTnMPCRVZrU1L9y5go2uG2B44jOMFEA2JSXY52A1Xg
2i73s2l2XFmcR6O50qFOQwtadQLcS7nJC3uQ+mv69Bp4wdFhrrpQXIdx2h9TLzF9
L7G61SwaTniPfM6NGen4Pd/PQNyVQaHCp5HAYkNhgnmAqTqUSaMCN4aTDnGi9kk6
fXRu0ZMc+2N14pJxx4WEosOHGfEheYhTtHZeyp/jYjK915ZFK+Ar5Gmi1+R5ngDc
U7czHZgyeja9i8xO84ihGXIRxaG3f8LOXmRuA/ByTQZts8P49QhBzc8pTdR2NeVD
wvoQ5W+cKVFV7+74467OgP/4akDQK+P94wjuJiGQxMCaCo6z6iYKKDxCGm/KApKe
bgpD5Bp33MkPG4YDdIj6ZdACJai0XDwZg8DaQX2RrhsGSPkPNhfC5akWfX+KWnL7
ce+bEKBexDlXYZKaQLBFbCNUlgUvzhiZXTYxE0Ib7X2vmR1uXxsEvmaZRz3o76yx
gGfmOoRfAk8GZy3NvWAktVcjEQCbJv98R09/+S1FFxFup34Af2BzCfymaCAEiPd2
uulORBxY8NK/ud7guJn240SjXWpTt9IT4CNC8xcuCbovvBVzsRSD7/H7uGxuxqxx
slYVfG6CZNOFsS+TrcZU9ESiBC8bzH1btWwIak0kdYN0KuRKeFvlw9AiTmjk8/o1
lMOPGr4FBq5evf+2P31hlKqjsFSEoJgM/+P0Z/Na5BmYKJf+U2OWCXKqspZALL0f
Jwdd/8PqGLAZPIWpPONs+6JxEanyqdrRiSTFJ7aMkPOVNkRytbmz0NuzuyQwoAub
cvovba0/gz5A7AUD3/HBfZXSsiusv5PpAJJYzLyuFkJc80wN9wpbL4izt/PlJlw6
ncuDaj6lsS0PAuPriTwwaVaoJsyrsMfd5yN1I2FueWUlxAnOCdtN5HryX9f5gZ7u
IV7RiKPlNTyr9RDQLef9/HHo166XnBopeUuj6x4pTsX+sLKQNp52rK8HTYtC9KbV
ox+fVhH9uOhJZcqRY6Ifrqyuv2KQxMMvGPGakDLRbhuORV/CVqiydjTNaFRedBll
chnVqAfDlnumGFm38IdF1FqdGKVg2KVRSpT4Rkz0VOMPGHeK93HObvy14Cp0U9q6
UXub4iPqHyuR6xs8IgTRb/hGMsAhlV833te3387sVJhZhfbiDkqE/t9BaTy9gRr2
UJ19SDdXsbkxsr29i4sgmBnO3TjHheF1XDGRIo2PdQ6t9FJSG7X6kAjWi9Y+KDM5
T0/EnWS/UCdslE0G5Mt1kY5FnEA02wZq07L6uy/D/ivlhUzVdnFXgPevySUjycdT
9WcQwf+pZddIqK17TgBzlSMgtldwGYPUfOhxt2c6B3F7QHpwMDWyHPppvtOOQtj6
gwvcxKydUrIFK0934dnjBwJzcijuwAT4lq4bd/KcX0AKiq4BrNJx0rMxI3FwtGvP
SvnLYPni1uzitDFjW1vUdjIbIgQOFfmKvKm5MH36Ilbbm8p6XSgEfLiIyCpG6gxA
DlaSx/Ekki33a/uAYsfhTKjQ2uj7MowUhVP2FAGZEUwyD3ZMuS4Z6IFrBvjEuOfL
myAZQ8P7JNQ1/ZYS0gcML928k/BlTo5/x0SwUAK+4UIHJ1WmDFygZFIOLbHil3je
A7gmnaI0rHYY7Mm1HrTUnHUdegnuRCOTDVZF8gjX3cP+SinDrpS0z/5tGeTTOXag
AGScUIjtcw+gcrN6yiZnO0GO7mUyFn4nJWUIdK5PjEgXD3GbHAy+DsczKHiHwVgf
KXhYttcDkel8MoeBL9YLjRKG0sXsClH4FP5sLbM+9e/uFzrAbieUETdJ+UmXjqTF
VfOahOK0y28ZGRDsaSIArC3dRoYJ5KqyKNmd8qWzRPAhU/muk4AshBmlSXAVUA1q
LjHDN9pPMzbhcn5g7ciTvCmQB9MTaT7WTLc+okp5pz7E3rmRL/Qp+yBdDAArQGrc
xkOPUeG+XLHd+J151rjJMMPnUeFhijomLeeSB2hcGphU1luVjFIKqtcZUqIhHRD3
Tzpb5kgt5U48wyuJk+dLGqJQNOmUrFkfYjnOI2fRkKATiVj9o3toqdYeOnr5SXw4
j88gWbXb70OGTrCavkk30jY3AJGj1fpDN2emCDJiAC25fUCBQPQkURkMxittNJVT
SBxMNsagnW9pqXzObE5Mxk7+ZrN41M8RgImLexs7+h+YzYfIqzj51Zy09y2cMDlD
h+Cm58KuH4C2L/G9z0pGKPey4JJYNsSTD23bNbvOrwK8+TyYu40SrKXZ6qvVNAMa
RBl8He+21UVU4eOTR7mxwSaO+mS9tj9tiBKr+9QUES45bTbOppcQDd0yfn0ymWuG
mXaLvX5Ib2hMMvWBcb301mj8dlekpUp3aBRD/IFaJshP6rZTiEoleJGcSOoC34to
eKluePLiquH0SK1zN7AgenntliuE+c7s6GJadMdNfTwJRnzvqlKlVr0hz3W2Ly4v
cgNecZFe02NP9pKqUzKy4WGfyIyDMN7MX5XQyGfv2AJipSX7gZENC0++QkrkG5YG
eJLkgmbUu/CrFpQP6UpNKfy3ObHOCeVs7+TKkFO1pDqcICegyg77lw9dgbjnamPT
NZiCeUxjqaZzaIMCABsdULucXORo8Z/EBjMilKfTtPSui3eBo6lbPPqurTrAEF/Z
5mtXECoarifBOjNPISuHsCbnSp0NLzk8aOnD4M6f6vma7zUO+YSWtjCPgeYiFUMf
EaE+LxBVCReG4XB5WIHqjhqsN3BJEvxPagAdHtnFh2uAefOLWX2gBGEVQNumXLWt
JtGzTk5JDGaMQAMwymNjA+aZdFSxLsxvsi1s/VbCIpnS7Sw8XXfeRiMb3L93wTiX
g+NcQXEfnsMlzX0+ePsron6nS8P9KDVUkid4o2dm2ShSb1bUgNusXDn6saAcygXh
oo6YDZAUq2aa7h8xmoh6JjmN1K9VY96EfaLZW0tlFRvSOMLv/yCliXT1SFCj368p
u6a/8s4bWpJLHZnTZfSfmnjMwQs1Oz2cKVIOzjAhfQTr3WRo7mEev5aK3ttwsSkL
LqY5YxqM0WGAqX8DUSqxP5oWsju6gOt6HVYoim0py4EibnGizxOZPdB1Y2gaAvic
yoAMGIK4uTfy2pygKMd8LAO77PxgK6nf4r5HCIPlLBa1AOqknNCbv/cRc0TNqvYL
D4OhoCUsV+gVhuvcw41YDkgMo3hK4TrJ26pcte8Q9f/VU3k8Gr+C0Cns/+Y689jV
I4QDKxHDg2+zuTGYJq1VKirmjv86iSbmicfeBC9LeW7ScaaGDT3Am0OBnpYfLJOA
S7+5R3f+4scu+S7LOtixjHQrYg8Y+Z2kjS24/f7ducRsb+F+KCYHVJ5hINxJqbDf
bt6S0iCnQM6e/O7M5rBsiU8Txi87SudpmKGsh7NFMa+msDNTIgO8z5G2zJv4fbzh
6mtN23AH303LZPr8ckUv4F9EGoVbUHKT+LMaapEF2UbP4qS3Xsd42U8CHXP4QL3W
AldMRFdNrMKEyMfECOtlAxQVnOSOlQcPvv/Ez04YwW3f/f/w3+WP9LoMtBgTIJry
mpBuA67d636NqDwRWIxdKC0/UmNLegc3iMZGutaPe4wlutJmq4CgWgKNVAeSMOPh
hJNbYR6xBbWidtHHCvj+hzKIwALyI/4BcZE62Tx+MOEK5AjdAL0XiN3ItNZ3+PCg
ouA1KQVQMk85PMuvCCkH9KgrcBV3/W8oGhr1prkDPSQaDJ4f3nhBDl80B/QVcy6H
GGr1Ep0HwD/iP9RjolqMrl90bnW09ueb/qBsshC8NwgAxEtt4sq/d7a7SuQ+Hqc6
mn9133anULJnQGUvpOjQk0FtssxtumvyMTTt0sf+JJBQp2OxbsrjisaUI32T7RFK
trP0ZxaL8sWTOhdZS/gd48aw3u7eje7+TKR57Qhr0Tayaa5cOvR0ziMXDSbslI6T
Zew3xgdHqdl5wdueyqpMqGUmzLhAq6WYQ0lGciAIh/u2pK84qZVCgK7Uth94vrE3
LnyTp6JPLVt2IoK0QDwttvRpk28DClvXEjhQ0ADLxaQwlsivyi+NuVfWTP5XtFIC
Qqgv1QnLvSJPnkuOsr9i5b7epSEjG75pPpCs5P+w0rA/b9ow9UlwPvN+fUinUSXk
dxxYzioJ8eUa54UbTMymuKixpZlV5bdhOUcf/ufACR1aeCZBxX7CBiLAllXjV9Vl
RgWocOJA8otFZsgNg2KW+nwqf0S+uxdR8w9bOR6k1dHVLwlytCpWMojq3rHFwEzT
yvhfx2+A4ago8yuxSVIcZ3m/1ZgVYc47oasfn5TzwFcp1jNgfeilCiFa0jU9sfmY
Vnww6lO3DLe1vKgWEys+/c6Q5vYX2gk6PrZbA5rdIhd/pwJ5tRPZg2tR8H/9O+IR
27yaNAcVhjMwWsJLK3WIgFmC+wmKmvIJ0gLIq0mCMTCgrNgS3VC3TjjqLPxGe7Rd
S4ixn9mT2pCgUolo3QxrS+fU852C6PlMcwv7Yr7Bu/ccvzgfDIKGfQRG+7AZn4xz
Qqj8JD/kfXm8+RJZ3EKze5IMzhryoSEaBCN3xvai8cExRn/tO1NzYgqyatq1m+LE
G0wV3Z7yRIkRoSTOEmJ05oYw6f5NdoZ9FBwNwLIjHyYbJb88bdan6GnL6L6z2ElN
9ObVZ8c143sl0kczUG6U/ZKoseA/hehRbR0xDQF80MWT7L42LUlp26OzLWmJ63j9
qBR4NVOuACL7vhsIZ2ZNBlrb4pP29TnJqmzgF3vPc4ax2ruClTm/ZXxzD106QopJ
3GgLXFiXSROGsIZ/6GH4DluiNoAgUCHRY4uxXvbHXpb3GY08MWPdiuhHPV2chqTK
KxES7Y5y/v2J7nUYp4R9fR6NIkIbJrJIZytxvXjEuH79spHY/rI3dUvH8SoWKjsE
3j28dTMf5nA70McdYG7KbNlB8o0yzrjfERY1OAoQg8r1JzWMDjFYRMAxXsRK+v2r
smMvS0Lucc8QQ2GQ8aq2VhDTKW5lb+nYPLQiFpat+2E8jOdID2cBsbdyLz90flpH
59cn88GgmZT/53xkQfpOtQ9OuquG/c52RXMFVBfGF5LH3A2PjTm2fm24K+MEuIJC
jWkV1ZPv0+03y8HlM6bl9Uwv/3BFcfm9kKrLKUvqfwCufSMeXUueUn1CkXdSAjLR
Ded8uFHQkiW9/ZgviUzOPdbNSGcX2pMbnrvRYMe0ZS0qxTWTXCXWtpfm5Bp6dEs4
Lx9AtNruL7nyOcnSDVFZaFIlEzEvhkILfLlaZtat/QoGO3hECy/DK4bv3pgVauq+
MygqCEH91XM/kW1oQqm+ciPiCnblrT3LjLGqcxpZ88XC8nqIkubqfxDfQaY1Nq1X
OMeYtYz1VLDMs2q8Gnn4rn/pc/SHFRFkp77Vj1kdb33i+z80CU5pJL5JjoRqDGwO
ajJiNgKa+5GK6jIMDr3Fc+JoYpGODFpwztZ28NCQVAIkz86A64Aei/xLV4eYujyx
rC0yLO+O+liqfg6h5/2Q7L0NsNrsgNPpDbVAVWaxqwX8jaKGWBXt10/rxZ27GV77
DTk+0mmvWFeKY587hVigPGf7aCvRnPm4cPWkirOfd+hp4vsJxbcyor2tGo3y7Hoe
8ieyjf1ZnboeG7kPWcSvI63h//bsqqEPudKe6V+VLEFppAvaBO3ngHWPszfCRbW1
tTDvKGaSEAwFbWBDiNiEiPAmTVh0QiHNMoSl7CwHlWPDHgkAU7V5Xew2zvS1Ochk
XTCSy3PstrOsbsFi1QOi0kx6G02YMWEkpxh0b/mLWwTDrqj0WNZ3G3cvkeUzEi0E
r4sZxZ0VVOB3X9uCYKv380Cq0RJ8qLmpqGD/SC2tDJBmBzgcPR5qc5M2H4Pr+pdM
Oc9/uPix7I80Z5wtvH9N2R/lFOSjH9HcGthTy0AzOb65qrUk2NvfCeF65srG8xpE
dTx3M3fKpVLqMwcMmmAIJZWjZPhUrvq59EetIMtMCdVww9QbbwF+yhiYyGc77Zmw
mY96V2IhPTl82pzPEg8la8ihMljT7pO3cVwtHw+h4NWaS9GObrFN+Zq6279wnumz
qZTHCzRdyz1H/bsch90mFcFJj+02G7QBMGQLW/ihnjyoBI0rWldEU1fxy8qvAwZn
8aOApiBiZf6PoOu4/wx8am35McR3oXl1RCq4I3ewDTNcI6NQQPA9NxVXhnc+5kal
0vuCleoCxI3B6JA+ZfcCitjKNTh5wyMKNaEtv0xf6mk2Lgsel5ZEFUXiAU55RDth
vdo1m9aAYYMLhlon7jUtoyih3k0G2VJp8LakQol2Wut0VfFFIZfKNUWU5OH41k0c
vSSuPHkcZdaDc9mOujNMcsATh66nUxn1k8bwdb6e2n/sKdegH4xkfXfIFgv44ViM
d7wyYNxteGlIJdMcDQoifqtDo4hMSauXMX4T8AM9oCH4iKBSLmQCy3KXDJAHf7BJ
W1XPakXWuvGN5J+ze+tnvc6Q6sLQsy8WZEPDdFVGfFzlE2J4hzwmWC1gKJR4h2DP
VZ/ABix3/KiK6JyK1RyVrFEPZ8RymqlPX9FiQLBt2q7NcjzwlGG0med7ABTaRi4Y
zEoHYoqrzbcczUSJGB920BJxZCTCTS9XcXg7PHNURSAr07VYnsAczHUeq6tT39QP
vO4mmM5IVQ05nnjCkhW/8nz0zkQF2LtZHvKO5Wec6pFgOigOcrvL4ebOd4uBgQKk
K5gHMOH7KWxE8ZAm4+VA9qJhK0RpWbFSmCWyQA2y0QJZdkLkHfo6w0M/FWgKumk6
C6uf66VqWdVLuBfkLosTkfW8bwZKrzla2oZXos8m3DrDZ5UfV6Pa/Q1RD5scjCIZ
GdlCBLGythdld34ro+sxI5E2OXILnUMb9vbeYbnMsJbV36j9ziwq8NO3dR3uzG10
KARCjMGC/5klsO87vXVs345EXSbNWbR1J63U0albF1Xz+stZb9+zaZJ8tKdVYJc0
7ALk9M/jDtXz62m2fOl5kwlUSgmL8NZVL49uIc9EnAcuvvKiySKVX22kztFhS/+r
YfD/DXy8fQvnQKSs3pyFLhPIXj7SyoHoBfc/22FZfanPAYC49AmMf5Eg5me4YjNi
XzqgKkfQujWE59POeDjAXHi3UWU74LJr1X8SmuLAO6TjTdchwkCvLME99Cer3Oaw
PJ4iwg53WyAGoE46FE5L93jWSVSznVe679+xfUVEDVT6q+cBvJBoY5dJkLNtJDa4
P3Fvvevmp7Bb2gmWd6sq7bevll+2pHaL+I1aTx4+/GkeZk1/8nPx8xJlEQ1W+x3b
AmP4VtjAEkKyxV8fge3yrB5xYOWiaTxxmKyz4jCmmMg80TEazGZCvfzfoQQnOWM6
9QJqm7R2nIIhYhJsCDGREkQd5pfjhYjBO9xfLQe6p1cyvKW/1C8MJvdao4xkYO0M
MCYdVZX8yHfeSBgLsLsxImd80be3tfew1RVNpJI+vXCg76fnjxHQNO2vJNnrc0H0
vbCkrvCnn8pC1rmYmC93jO0lVyT1RqQmPoZVpAgqzdbmiWyokhRuerDjW2u1Oxkq
sTTjkg6AcCfARm1yy6xp8LkrphYABgHDpt6fUxewG6nd48OZilrn/0CXhBoG0TDm
9tXMFWzyFeapKi+iKptG6Re6NsNFKPd8gw3Dw12SWQteBz2VxwksyyXR+nsDYOlz
ym4qYyiCuROVhN7Fl0uGVCzpcqS3VoULOyt/mYGavA/34/DW0x36YJ/158wp/P0S
AjIJIZq/LbATLRnohEhCyjyQoJX7Z3wR1F6oGOjBP9PDmFO0wtqjw2NgwW1Jz7kY
ry3gNBNrsRR9Y0XOMh4g/J4i0KQI29iRknXTR5PTaydrHDvOhNVh22FbNzrhaKNy
ZNT/M95gP9QY/82ltgGr/IPufmSHFlJ4hthMY0waSezozX2uozfrAga2SP5786sF
Ps2MvyLZYhgqw2utoPbaif+4vfAY5Tq8X0TZEeNVVNXuuM2BoJRsTmJ4T2jjCghA
GRBzrAWKSpOBAPKmQ0XArhhtmZ+VLzPKsGk10bD49q0tMVgQGn7xCp7b/NQ7TPVA
MtkRRerZayNy3zdb9bxzLWJ80VpzDMPisK+4Xza2meSU4BDOF45P9/jVgd1+RrJf
tkrhM6rOJMRcVWa9Db7IIfPwXpa+vxDlchJZ2d80GY5AwmWPX/PHhaHRbRdA+DC6
eCrXqDouja7Tr5SBBZWBv6rMiT/LIglsj0nezUpxep5h6DWUqbc8J21rcRq3ww1O
FGHXmHe2Ik7xPrpD+Gi2f0Op7rZvK9rsTk+zRYCcrX2iVswVVMq8k0VU9Z3GksNy
2/jdZsmpwCX8ley4XBfTo8iS2LdkubhuZ1UtcK8umldGxydBZLok652s0aZ2ztVq
3IlaCypNLehF5H9LAZK6QMSpnAg1tK7+F9/p9dtUvC1VVXQqDnyZd8VY7bammWxZ
YzHsoF2h1z23++eLjB+7MVc/bghwkP+p07SV29BuBAukhVl6t7y+iMdzg9gOnyym
juannVSxHjaqegN1B5zIKbPcI6dYSG8eyUndcnq90NrEZNS43a6kmKS1oI+/Isd0
el6ALHhsAJt2FH53eH+y6OuUr+7WewpWb7C/xhbpJZLSjChyUrhNatZnVatK3RSy
EITQIber5mrSYn6Rz8D9JBAU+ME/s9cIGCW8+64w/Bp2tfzddAaeDlP4sw7HhNMZ
NkolUR+D1OdIwEn3ZFs77V75fqrH1GAduN70YCIGhiPVaqyoQiBZqoYD1MRdb640
LUEmtqE0YhtFAM6Z4Tog7La/PHKJnKKL3nLTuMKLGQZyH29MQpex0esEpYWTtYyE
tD88DhrKMjoMR7sX67p2RQVC88QTgvkPyAb7xu3zw5XOXt/mmcqHTb+1SkOQ9BVY
r+CsJzLAQK6WQMhKmm8pHqVpZf7lsV6/sYelG6JjPba7pXEF2CJ/21fDSBl1gGpW
iZQANBgA6V6B5So3iFb2AgJK1ykWIReSVQlj89BLmaFgAf4QFQnyp4EP7g966L05
c1t0h81rWbVu3e0W8dYmv+MrK7hUMAuoLfxpMKEeroC6Ih+csBNLbkb4ddlry9lV
WsRiswwUiLMw+373MwlC20ycES47BYq7C3Bn3U+7z2WRGiej/xCMev3nSAyVrrqh
pSnxfJNHNBjWEhwQYB75Z1Vwt39C8Q/WsC4DTgWi4/zBu+WPbuIrmZlwIxMVPyVW
CwyfvKs+fJcqPsSDsTbvfcBKhrZAAFeeXNVP9nl01/G2TaN2E1n86njZGiVzf2Ji
nPmo9yNceAy9GorZOfBVEFGBWisNEJ5F+emHVOWL9y0Bzu2jHa31wEouvPEA1Ysn
YUEKyGWFQkj6igEFFjvJT10wpRfkk+qlXLu0vElAIenn/r8oOTesxluSkUWD5A3D
0TMQilTaq5E8SjFUZ9MXE66Lji9AGd6GeN8YFFzttF5G9KEspzmtSgzGLe5bOpbi
6SUulwXt33lgj4g5LKLQkyB2cvM/hhyaAiWkUd/Ta/OUm+xM8Zua2gCiGMTrzBf0
aHe/+w+QLmFBYA72GBJ9uNGU7DOmAa0cVQs11cYCF7ksAqfdF46TH598/Frk0j1z
mPSVrZxsOrZlRfTxXKJSeXEn0dVvqJ/CcDzMj9c+PiZXUkCiIQcA4l6LwTdvdSey
osskPZIGyGwR+oGk0siZtK0ppsx7CsCKD+lObn4oDOZxLpttuQ5JgiTxRkm4FXcm
RAupgvNskD0Uzy206ihQ4eRta1uLsGeYkQ28IlK2NGUdf646FFZ6p7Iot5h0aegq
E6gMzoQce4oKbgpr6O7XYQwzd0SiY5DISfTPX7/GDhKWMN8KbD9k7I3FSkeMCfYU
3UY2ysfptEpbItU8QbJPoPSJIKCYKA2oH6nU8FN3vmzodhq/buIgjZyCo1piepFZ
ERP1VQFyJN0CtReDsl/gvAsvW1BdRWVH+VYwzNqM0KmGn3Qg/BnLz1f9PQ+kFuv6
N+MtBoqaoyRvLLvr0+rP7fW1lV4j1AjlIeqF4Z8kUnaEH57iOk3VN+a8noeAVaXJ
NR78TmoIyGfCheOAfriB2xdq1RDiePqWqhmEbqyISlpj8rzGs4loZefsxac14dT2
Lug+nevbPsdE1JMptDZTxcA0M3EX3gvpt8ujiO9wzY5n6Ieb5gpAz6tcUAJUKZ+o
NL2Bf7I6dTzanqUrvG/r+Hk28yFGTOCm3kTTKiMe+0u9h/+zG5m6s15A+baZMi/a
NSZvzxjujgtKpL6eUHwROQnT5vdt1aN3rKAVNgjT16LmTsHgjnFArZJPy3ef9MJi
OaDKLzDc7ZI+XGTelRfReq/AL4hDvWFL0X1SHvR8BUakTqT9+3PoBdfXuq1aj2kB
BPHi41V+DlHNtiQGaxD/ONyVbtPs4pex9QTuQ4q8nmYh7/tWF0O2SRHn70+/ve0H
nwmc397PHPFCcWEsegWvr44FgQOrhPNRnVkN9JQOU00hv6fRGbVKOmfQyWsLDJIm
buUtberJ01ZuYxUO6fZrCqn7QscfyZpOkJOT6O6iKupKI9hcbA1L1rJ+xFGsn2s0
ezUYJVHM6H5yjZJN36QhZKy/SikxmnKhAQ2DY59Bx4hGIhjLjfm7i77cKoIeNMYL
8soxSEQT/1KzbemXcgGoP/LW0g75ZotivGWpSCkGdVEZ/MhqFG2nEU2PLvts6kE0
vdZUq1cM7dP+bhvqxHFmxR2lcfFGIvNRmX/SZuQI6pRqGhTN3Ls4klFrmEWRGXbX
eDDCylbPOCuLyYVW11yHF8nqa+jk+uwMBM2K6/CrGrts6JqIev6ZXE5xYptdo1q4
+eLC/fy0bUHQSZ/20zJnev9yU9x88f6zK0gfrQTnJHNMsc9vgscipKsZwO84MDK8
qXUQP12rYa1ozLNQrtseUxjz3uQIzoHM6/G7ebSzMEZhF3/BlrU7mjBR54rCFTX3
aNn0vLu99ZHx8r3h0ZnclYWPX3CwImdlvKOe88R0tsyRs+XMHUaIqgSZcsO+2UjG
guBiVRxc7j36hV+Aw/cEq56xGj6SiQm5v82YAhIK3XqjJ3uiN/rUsu/Sp5Rb3twJ
MqNu6XB/+0IhRsFh1Pf0+2OKvLH9JqK3DiLxQfKhoqyNbisRnt0qxTYjmG+H1CLY
UfkO98AZa0iVRRBqZaDFV96WE9a8aQOuRi8SU41l07Uq0BCB7sJhNHDU9SyKIqzm
/e8yIrHVj7c48hwDxwJbABfVKKREkZkJUMhNNLr6d3S3l5UK4nDm1vFqkI1TE7+w
h7b1cb68P2ZvRNIMBSdtR7dcaYQ+V9skp3slxA1qo0cNUUbbFqlMcYh/ydtl0SX/
ti2O963ugGn4Rz3rkxVD8Q5UzxSG1F0J62q/dgKv9wvXsz9bHfHhTuIryDlsZZ8j
2iNaiH6h5urbKWqsOa6c5cQKOcXEsqB/sYa1DV9vUmruaUXMPsewEqXAvVwvR1Vu
XBUPydXqFyuVYR0VH08onVlhVg0EuCSctIQFIRVoLCBCAdr2bopLu2GrqSGyoe7p
bYqPemvKwE0LqeHji7JfpT79D9wqc7mIgRLoUKbr+m6tu5H3Ff30LBl1hyb/9Nfc
6I2eseuEqVObku0FiGPEOxYfWkeDsDbdVBOIJ6+xUvCUs0IAo9DIQnN039h7cS3D
UDf7k/uiK8PAALc9dzdf5SJIA34RBlcLxopmzuMtFEGeAUX2WvuLxULHtjT5ZP22
zBWOq/OQqM6IxCx85/C/oMvuvpW2BCJu2CzIR4dhQa5c9L8MlyWdBX/hJNhhBcLY
OF3nFS3raLldezEmnI7QTLyzJgsG6o0TsR9fd8BonLoiC1C3MMYmVhQ7HX/B3U/J
vLpnQDaglLBcWfVOJsLAJ7fYQhpNwSe4w4b4i2WO5nk9DCpPFvmBGEUs3h22oShO
xltNDWIFrrM49a8/jwSy1cqxnUSwVoxHk8YnCt+jPQQjuXEvWNojtkgvekCJVnzc
0EPrEgcwXwRxDzrXXKUNzthVbTq3rab4OthdLNdGjgBTETMemYOgRcLi+FXBViKX
XBv1mGpBDpwMaCcqlWQVt0b+UyccKAhShdLDxk9DTUUYFxWQrl/Q5VVBP5nDo63S
0xd6nQPCD2CTjOiaurTJC95Tbvy4r51wJhViLWqsV7UMrNlOv0Q/iHyVVXYPCJ2B
/V/NXjQmxfSgovlUGRpctLXMOat8S/7LHSW0kgvn72t6uRlkXZ7LgRIrMRYBjV0N
eWvZqToleBdhy65RsnnFiLRnOaOQIUxoy3New1OGBBo17VzE8kgduQfNwavh0ADK
UkCwFR3Z4cPY5Cr/2jf/ZvKhqjNTVWuFvPJ/t6wL3XCxGSZIYyKUDKAZmK1leFt6
SoLA6ie5pS41W0uOaWfH3KzR+xNIeEyyRwTouOt4Pvi/GTY5DYVAnDms8tKhcCUe
q9cIZeXQMwbgH9gemLsdaR0Y+Ca6DGzz4EfVa82h8IP1NRBeMQmuv9uxvA+wbkFL
gb22Wkx4OtS7LcBtqMv0FlPGQ21ZixRQsT5yegeMo4dyfP9prf2s9NZQAT5zHRfc
qCO0ScQ+6j6X2yizPyKAeY/PWp+VZ8/cqBHBtV+2lUa2+BUfuFRCIKKzu9xGV4GX
QL2zefhqz98EbFk14hqdg/Oj1MobbAnLw1ZICQ4XNzRqZnpxhSEx4Zneueb4oCTn
FI7OgKwjh4hbx5pAfr7q2bHBskmyu7GOKdeqwAgyXjrM5SuyO7Ebk44F0tvfNWIz
py/ZFhYqmYx0DKYOisy0g8GM3bViBJjFZbOduVjs/ZT1x7U+ltuOfV2HaFUrdQ0M
NayerHINpzBFmd/J3J4EMgBCpQXgM+r0ZQgpsp7ZX1zx/qMk5LtdCbzghWfZ+mQC
OM5aYnxGj3HDYNotrhOWmlWimN0YWLBLJPDP0+pVMcH/XsyGFp2VbaPcdvdsT3Pv
/ZQ/k/kAVdO38Gby9zN6Vy/OCNWzwOYPA38c84m6KgqOaogN+y2MKoWuKaPB4qi6
bAdPETD3YjO+orD0fo1fJJUlORwHYDAmmCUWxxttZvY+cr6VXEg4x+O7KobYpNII
5dVAaTeRTmKY/vLgIJCxSrnO0xuYibWI7oDWNQ25isAoYSv/hhNsJaTL4Xg/Z87S
gvHF4Hj7vEIDL2zb2xXonoka18VG22yqp4UztcZhn21vfwRt72uBbx5dszJiBosZ
jJK9Z1hWr/FDG/d+50EiHjz2vlty1BGdrasVmGwHFWJLkRxxtZWC6daQAmW/Ntvi
hS+mBbVaPz1tnqqurR/2KTUOtxFq4xmKoDa8tBgUGCbLS1Pz2/u2NR2TkHFvOUPY
lRdE+jCwso0bJUM0iwi+GBnTTE+qxqxp7TrzppOyl9VVrsVGdyiHD1Rl5RWKtxZh
v94x+Z3lHav+mvujC15Z1+J7uiDL1odaZOqacEgdAP9f8UEPGvvBV8u62Ee+0Db2
pWOE5QOMVH5PKhHEGzCfPTwxKtniOnA6c/SkiKoDIXPRDj9PVdpKF7zoC57OUjxA
iig3Hjy/vEAirbgRvWLRaWQDgvPjm0Zny7FU10SXz6nWopR3gvHHLq743zCjIvGF
GXf/PwJK/7QpI8xsCjOsnWtzIV6mKSVahWvZI1if7P82ssO6vLvq78kq0x1U4e2f
OfrxdqMQAXX4R1/qjyx8ogPL4yHP6KoTw+5LCaSVFrgZ5U9zAdewIIQhrK5OXF3W
cS/gZzOi3hTOdQAdKHnP2VfEg4eVwZUwVH/Rq5jIhVleZeuW8H6gDIwPwzwyBvNb
JzAB7ONhpByz/8sEmKIo9vRDwDLMC95yhO05kK6tWszeMdnTytLbaweqGJVlsN92
NagHSk1N5hq26jeJZVPrtbfRmZkWrAh3UfHSEBdJAYcFR95EaxUeXPrj4v5LlGPA
bJXtS9YAhMDx6NQEO9YiBctWjaJQ3lWVrqJ5ihY7tuJUYGDndRDJdwGGWCUkzROq
RbomM583V6zKjG61864cN+DB9YQZdAqe9nRHWGgeX8Cq1BGBQnFfWc5Pm4Y+co79
E7drCfc1cBNHPRX4ISlUFcb5zP4hR6wYj7bQLwg7aoNynwsB2ivD49mkI74ILluF
VuOGI4Y+ksD+7Da0lkjuTWUDAsHJrasY03ak5poCpnFSs4DVr5CKMa+GzdaA2xuh
UAZu6zu8/LbXvNUzADSEXRmA/ulH1AgkeHbJ46yiaA6O00ekazV85J68P4KOCOd8
91doDaZ5S+5J3AIRLTsYSDlClwNSeSfDhmFXv58SDmRy++9+vIkXfCiZVKYoCt2S
5kTa0gKzdIVjkU/LoQDwTZPHdzp687vEhIZzINCozAHSFglRGa138NqLDt0w4YMr
aY4EX8m0KkAei4+aB0FsBp8MWTvsHfSckeMq0Np+3LxZ+78vcMD12WfPVvq14tlu
xqnsV0KCt8Mm5lV4T98fCzX1sTZefjCh6o/FUiUA2vKa1bYy6YBpo7VMKsWn+JOC
iurO3cmkD9K4S6NnTEr8UhzleptFq9n+dNtCd4tVuvcbJ7krX5UIxMVPG3/tOiyV
1CYUCAqYRT6XZhbskkf83/hkitIrSKMz5Kt9tvcKjqU4nb3+gLNiCu0a7uGA0O2W
+vyLUoFbWIQ2bHhn2qkLAtNUCim8qkuYTk/YHxCghrBtRpZb+feB5URCqLD9yNM8
Etwcub1cGraywd9DIBUyzfmrcbdSCTgSRTr07CP6x221HQSxR5skZo7FCR5ToRKz
u+4pUetAAkb4d74RmK+NjCu2/DD7Efv54eCZrJznhGz8bCCU78sd+bY/rXnbm/6L
e9fDD3iMW6DO/DgIRcQ1ZBaSl10hHv4LC0jihdXpKsPjpkWj/LuCPq/mOZ1qe3A8
xFlHNt81yUsaeAA+5c+AiebIl04UTbwqgnyBopYlI3fxxVI49OrShoy7SB+dbJ2e
4AK7LbBU2gLo51FiVicN2s75KrTu5KNyN3U9FX/3MX5eU3ker4ytd0lEQoi1ZHWH
cu4wBHirQkOMc9VwL7YfCas5CkSJ2difoeCRfPu+cio9d2W7SfTgVMgRRNtfPXHD
6haQtPlhfDmfT9zLggzGPsrRP5qTguP+yiucbCNlR9r3EkeaV74IUvP02hR0l/I3
kbIkLZTVP99b8HCMqVr6Ckkx25qmjgNV8ICPc0VauGgx7m1ugx5x66dIvxuU+eRm
G1OKtHMxikOl0bkEL2KijfcYc+9kNY0pi90hvqYdNQDpVWXjRWlUYKjHMxCf4mJu
De3OalQLtbcz9M1/zVivHRGay3DGynVNWg9XuIRkQKNOJK0fyIdK8iHd5++SOE+0
3WYNsqtd7b9TvfZ/w38eIz7u2Nj+kmJzYmupz7C/YyILJQ9Z+p9j3ge7Ka0tANeF
+Mqs9pvkoDUWgie9/vIzxbAay/6up5omzob//5mM1N2Y79ROhbsub2uPeWXRcXUX
vh92YYYSEvEScQruyIesCDVpKJk0AaU1hSdNCfCEmLg6zSciDBk76k91y6wnlivM
19pI+wLwUBFzqpy0U63PhTQlQdFwWSI/H9G4fWp9CMHZKwBNojncmZRi3KUPn/O7
2b2cR/aiFzb3wK2zoR7KNBTj8tRQ+/3dvjg5i/8xFPZuYUA2QtXzyoaZ5j6O3+cQ
93uYuWqpAruTnuDX7ooJ+TbjBr9GZFMB0ECoEyMgqdlnLCNLf5hzihGWV/pJY/Z0
ehoafR6D+QXGdGI4KK1gy+l6NAuUuo2GNo3JGBdcE+a8aSs2ZjPvDOSPzmI9I1Ug
flM2V+Xb1E1R8Dy5QtZnc3psZ/pp6wPqCAVQJOqITDwUGn6cqBcUF6V6IJm9uYFL
qnZuORorhd4HXBKiJzzoY1/TIs0VnIWCeJLqgAxFNdg7Dom2X84vBOqfC+8+PAyQ
c8Td6oPBI4zbko9euOLHbouxdOOUoifI/RgKFtsoEfCyiL0ZRbanWRptu4FaTyYr
dQTp0oz7I9fe3m45XtYd2U82/wU3VYksBD8MJLbGUP3UDzqGweTe9kveDvCHjWFW
4EqZA3mNQZGXVJ+GJ/diriEBX4LiShAgfXashsL9a7loNNYqaN8fXeJaWLl7Nbk6
W0ElZ4OyjipTAl3WRRAaYo1PdnkIw/HNvNiAFsp0zr+AynsOdvVh2eheI3955IEo
/VsrbAbgbzeUHcaadPpSXPKcKNJ61Z1ByIcpxOPerpALIEo3frXha6yh+wn/AlDw
pT/Gc3a8vatG/nJV5TOokGWaMYtxvHAdmTZwMReTDWkVTbp/lMqUH0petVWkOge2
CVe5NasTnCD5gbrTPFcUV/ibRi21Bh3YckhIkQ6u36KE40Y+Vl5Y8+HKg+0WRiy1
j74QiKbYTDzL62Q4aQjec1qEOzHfe9eJfFY97WtGTu0obZBwHyZZmhhrgO4DUUM3
ALAyjpDEwJOmfUwlnsZgukbAUl34Pq3rPzRYvBO+JpKTZhciwIbB+e3AwXCai1yB
zhwWTA6Oxzn4UbT9PeOZwRd2K98WYJK4nb3sgC++LuuPciZ9CujTm+rJGxiRpJZ5
EAZqHnzBH/49+WoDtpyIZhxEuSXw2q8W0sMWJk5aMsr0kCdrSZRlwCBA9cr01jPK
jVVtRI3XDvlVrzWt7YKEuX4LnBk+ol1kUewJtuqZ1n5PgzKujpot5nLRestrGcqO
l9WIo/6g9ErqvB5k4DfFp2MFtXOEAThKlZZiUcIIEV72B9uTopMFqXH9sm3yd8Kd
K/TgJfBQ3hwX07DvV3Yx60EQOwbdk14D2rcZ9IFaXPSZlaSRZTQTxmqmd+5r7oJi
NG+epRrUjOWF4gH8RPCZo7TXvv21PJnPorP1be3pOsnU47F5ft4obZ+2uNKKZuIy
SBe5BJsSDVVJV3I/aWFMZcu60rlU50RSYvLjgYmcji5AtQJ8X5BSq8Ft29Oi1pfY
Q6ng9FpuXOnjBkHqmowGpyqQsaRFisPe4fNO49Hi1DJv7GVrrKuv+U9nGoRJxNYq
8VGs3VLMUma6UvHxwmgRR5P4rxDRTfSJFdk1DyxBFPZaxOG6PQB5cCIkD2HKKV4W
mVo1mh38O+4hTaBwOP8gpuESN4LT/CzvmJmE5TusfnCAy7yPhmbgFXEtSrPWUuXg
dg+XtAYmVuw+USKb8hjaFRPHYbjUoX/STIkkMRcZvHrsg4nNwrH2ljLiCpcrS66T
LwQNuv98AqXqkvj449YzJACzu+TObmorrTeRaX3USatc3yzFh7WFL46x94VNXsvS
v2y/nc7cCkXYeIUwTiZrnRvK5YAq020LJ3lB9kegFFD3YY25kBjXDJonqHuoAYbb
dUFDvcINGOZOvNzXlrc1A0M7A41XSPsyDaSxBaQs6FnEOWQDiykORyZF8DMALTj7
vPwfgMlLcuPvMZmZ2yARP7LqGsSanX/HEmH26SwyYujkxPQmtGCT9Nni5pLTxNMe
+XRKjErgfvnC+Hn6QbhKs5D+Zt37H2th2pCeMLRbe1lCw2NNS49i10xidAyfgbNv
JkTJRHnQiJjVeIU3ddH/5Yj2q769CNhnJUYNjEc0uDw9IesbZOnSRQEnHp0JdZJq
5nxwXcwLlN+JSZ/glHtHxY4mUgHtZaxEy9WxMUMi4B3wBWfjh6NOrnOSK7ywEO2p
ql4fZrDSA123UNnDpG7Wlz1j7np6L8s4QINbelRI2M9Smcv6qQG2bXk6BEJNeyy9
/QQ6/FijWZ9NSmOlyF2Bc2Cjk5SBol835Tw2BrTYlKG+u+vts9EgcLlG81EukHpZ
l55Fowj5OCjsGAr9YheCph2qMwNf3UygyY/P5VRwri0YVGs+TdUBuadQkacopL8g
IgYi2pvm6PMx65IlcAMxhavKRYJ0HopTKb9qyhFYLd4n+kC3ut6wKf4vpN/NMX8b
BWtGoTaZJlA3fS4eLAQ2H4xTQkCNKCPQ9zM2z8P1vHUnO84E9GvGe2UzFIw18saM
wiaup2V2zI/l/p1DNOgBW5Gbw+FKjFQU7qzONnmp0y/+HsqyVX+799jPNp98R+nq
DnOK7RRjn38koxOCDEF6vt4lAhuWRW+c/etPuBz1O833dSmihawkJYXIxoFXKkay
rbZhaLRSETD0pIsGYcn47AHwmf5z6TBqL87FUF3e44gt+NAQC8WYJXF8dWGhAKd9
TynlQXlQ4SdzoYd57XlP2sYDqdY7z8PX3KpADs2AMVrWoI7R3hMADrENSTlV5QWI
CxXbrDydBP3xrPTzYgo9VIiALa18x+c3JP78LLlUcasC6yPezXjPRLhxgG9Xvvjy
PV5elLL8gtgvNAQFrmpMx4MXJhqrD91wBnavjGz6KVs2V2g5BC2jFKK9Zs+7bwL8
Awl6RqiyCUTvqEn/GxkHKC2XVNtw4M+9S2MdAxhwQTcfPTOqoCnpwlzml/SYKEbT
8oVRXOSX0bfMwSvT0qtsDxTgEI1j3FzwSXXT+jXspO2cs0AEvbSELtY1czI57+Hg
0Kf5evvx0uTPSIH5Sw/sHQMMT3RMWD044loWWn2Ee4J6WROscrvZcSb1pVdHW+JY
kjPzE33oLzJdqcjxps8MwTs6VZ1efS7yo9aPwukJat/R0h6jIQ7wfFaNFUhSjMQm
e/o7IxS6wM3dvQMy8ZJoa34w/rM9IjYNx63c5iuLXicLs53EqDPplbHqPt1D+LoU
RppDQuzdyeUl3rBTKqNp/EOs4eRy0vk9MlD49UpxMb5Y7NR3USCCEAY1qtjCaT4D
/84u9foQfp9jpYtwdPpsSI8+jcFvW34wN0qxt4NOauHX9e/Gu7w2miQgpXIqQo2j
sawZoRjscyJzEUtsgqe2OfyGmaCW4tCldikLwRBxwHSXVBUSQxK5S1oMrm3XnuBR
3xj5UsPZgLdDclkvQ2Gu1YZFODg7/fN+ZvOfUbGZahY4bfUed3alFKx+mVyMRpZX
xJg0RmTI9KliQNdiz9tBrUpWog2MQHF9OUP17geLD0Z89AGVBPzPT8a3qfhngMOg
WVXD/US6QZ0l92UJXMBlKv5SNRby9i7X/fxNQuXF7XK84HeMjkTwdb7J2EtfxdWu
Ym6dgVUg6Uwzgbuij63XrB8xvZYumnGAnR4oi6Y22la5L3R4m4l4JXZLkpO29xcT
v8QrTrXu7Ff5MV1NJ1LNdw6Co4uD6IcJsVYqWKUHAxtuCtjjblmHDKpK7ACXsL8X
CyYnvP8u2fEusTaKB3GoJ5LKhOwdOmPxY0wp609rTmfJKTjnJ2zfeV4qnf2oTVfQ
1gn4sX/ppKJJwMq5NCs4+EmQZF+9mBPJ47hc0p/7xukqTruMAQcaziERx5FJ18sT
D0t0IBJ9j4DAyX54KZ+4fN2tu0+E/R7gWrDMstHGFiDrwAlNXw0VRfufea00ZNxT
23fn+Fj0eG/ZA/LEvcPmc2nELmjq0kYS3GbWHaM0NFcjnQKWO8U6+ZqqhW+ZMcou
Hn+tcaLH6SosQ7Y211F7itgu+xIb6aXBWCltjP4qgfS/MAK38PGUXVgaY6KXHSW8
KoUVTN9hMruXTgjFKMo5q5az7UCVt9bDKJz4bHVjyDKoRny/Team+dp//281pe91
EUz+ZEl4PYhXiKHHQPC3yvqhyb1mwbBdVejEqAkpm+lvabpIY/LVPW+kgNa12zKe
0X1gaA+2rEBnpmxVPy2DN5f2g39tIZym7OM6IdnYs/xm3YoDfmtW61ndn6tCS/go
PN0qT92IjTc5zP71EKK7MLiKeBJ88DeHOOtrlDpzcgOIozzrcJZwgDUkCojT2Ljd
0/trzBskrsLaZJkZK4QN0kHrWgwvlhI5/qZHAkXbzq/wFuEWiVPD3OHFB0V5YNnJ
6tSED9k61z0qBU5ES5iZ7SDvzFG3Xkr9RUEcgD2yB7Vy6a9ns7lFcdc/PYco+KHa
3ufJ6J6GctAK1O2pOa5qCjOITGSini7wykyVxGkDg3LzlQQ7JVNv038r4wqYh4yJ
kDXTJfcw8qmDW4jyte1yEmTTwsk0sNHbX56w7Cd1b7r0zRPMqhE0LWKTqoIMIcRq
oocfAwIChcar9JpFhfGq2+itKkyslquIo0mZhBpZzmvBeoBXI1rXoH3twgsXD9GE
OUVwSev7q8gEBhbQBqYaRNCXbxSQrZlnIEMmT0PRDGMymzkECh+xkmPxs248PMGn
154+V9IFruBdHrou2XHqEQEKhTDa1zBQexj7KjX6fcwHU8UaNqYgRKx0U1/qsOQW
92Hg100oILmqRINOfjfEn4MK8zlgt5gsBjeJ5Yw97+8EbJvXEySquhgw9ntSQsAT
VCDThc6Y1v/PBAyhuewsaMqVbtgieWIzWREF6i233XHcDm8HUiMA/EkQ0elbsSot
FcSAQsAAsTrttL8HAQd5iikU0VHsJa2wuksRmDGBfNWnHzkow5Y2zAYXFq6Noysh
70NaslIHRjKzW537oLPjeQunrbPFj662TR9uq9JQK5INA2NImciBCdzuFt78N8NZ
Cl2BkuFJ4Q38J5N9NcwqkLRLWZ6whmIN7VWnAV7ra6j+qkC58JTq5428L2vfDmEj
wOvhYo8UpW4n3gw/l4xug7VmRjYdDm1E+KG456jeShfk+H/J4M43idIm2T5PwR0C
SL9t85fRg4wsX7Q7pssblwWngkssTWYYAbmu3uTPIxlL2W65CpK5cQNZLSPiFuvJ
khGjN7kaEQkSA0MdJiEENKe7J50Z34CwPuwa36d/K+RAT/C/SJ4Do31rXb4bx3dR
Q+ZG0MsuhSV8UceUsxddzt8JG+liIP9OvGsiwDnNbICt/PmRUaP9ETGMrhVF21Hg
R0lIZOxPbCt8D2CRbXmvmY5wkeZYAYTOpOnAr/4EhICj6hc6IBEgIe9F603HO5kr
3+w2pH3dQQU9VP9/r0qObhSIeS1hQm8FfCNH8zQ5rU2naxKuFy53m8R2FqvUu/09
6d1JCnaGh6q8vNaS0NdofOxCiU8YXl4vu73WF8jVHMaIOphYKXLFP7h4EV5O1EIk
lHYWMAbgYatZBpyP+6H9VBqhZbG2oObJU9vhZYHd2WmNbken4KqwHgY3lUmqO9gn
wdBJGK/vLxdS/GYdLcfeq0XkdlQHHoPbxZTzawfXuEqGCRLNNiipFI1ukPvcjMXM
ZV5GnJsxx4PfA4ryEN9pMZObnfR7rvPXS3qKa3eAa3YG7tMv5d1BAsFmfZ21S6gL
LnPxkmSTz0zZ/ptOYYl9NGlqUz3MBmDihD+XRBQptQaHAbHXW1YeQ0hfjig4sevK
3Y2Z81wLD6JE+gcUe3YZZYJZuPYDM+zTw3nutYdqFQLzI7SWr7KnSYWNFS6fSl4t
rJZZASB8XQpRrFJuGSnuGaaxkrGLItbxcbKfsuyUeeYGmix/reAXiBlCyX9YzANw
EMfF0Wcq/X/o3JeKxTpAYiSvE5SdlrYozb7n3dm0XsfD6gXHuG7kzZHCdDWm0NYd
T/3FCIK3rOFJesIc3jc336eDDjP2jYALhhFFPgNe+n4m24vb5dmbBbEd77YQIStN
CDwmsNDgtbCXaEkr4Y3IAnQKFRrq5/Tu/vMjzNirHoZlRFZV95BAEH/eqGkHbBIo
bUy78QSgVlKocRz4XaSO+BjBs9NuuvIC3cBxIs+eL3v3w+DtKSREYRdNXIqTHjNA
1VuqIEbg0FXmuXvfBmfh6Venk0ndhrAj3M9Irxe9v81NaHTwnw30ft8BLqYNGWd/
slwlsOn/tv/5kOWcn0w4w0o+mC1llT9QLl4V2UW3EOzDzYpO/GtrCvrhz8Qu4P5X
d5EbIOW27miDuhfsCD2L3mC17fvojBKQYIup3BdMzFDJzBV7WU/pWO7cwl2GubU2
JUbyVbuepBXL8Ss7Xs4RPz+kYF7WsTp+bBJn8pf6kno4O2mnAybSYJSA41olgsXA
VCKfxrHNbnwtZrn2alr3kZmoEmn70jQrCd7omupbAhsIQAcUBG3ACo/W80A3VSss
wYAmDUrtfrMf/eFtrpq8Juxj4wSKSgYFihq7vfMd0eBcmWV3HdMmGq+n7m7QoPKh
LPi21OnEwWlzpW2a+f3LlliiyClxHr/0L3XpVeKRg4DV3QOSxuY917GuxMs2ZuFi
k8oL8qFZ+hodF3XbrR+kYsi4D50CVm0bSeMuGamgCcSEXjolaKCmPgTBFhYW8Jfl
m49grr6Te+t30jefR6OJRgAPGK82+BH8ZC34sxCpQBVuJ6hKV/PWpleQjqP0nRpN
4775DTugS/fRpvSCiP7emGoCiRY4HjWy0OosmZdQ8tO/fb5yWqOxHjpjtAs7hgsK
Zgq9dIvwFswU+i/yPA4RrJ2kGxK9t8fWHbqjvU/tERk+VXplaM4rQBcz/b/5ka8F
LTp8P3+IB21t8oXI/kHgh9Pf4WpahWEfgC6T+oMusBArwg1AFcAo6+XGjov6XkB9
jy6MCViUFcPRHDXp1FcZ+4foVi+bhxRiZ43sefv2argtWyvS2ex2aCQZQBZMV5sK
bUYnvquN55pSE/ckfJ3a32IekxVoW7lg98afb5AFb4Y7LCl2FNVWrkp6IBwzUmSx
ybZK/21sOGsfTkpB3RgMSW/5C2mVingedcK6Ln8JJCdSLLwLQGpB/PmYqcfw7HwX
mpS0oTX31euBPoJfdYHvNx6yqNG5tJRbKDiwp+TYJba/AwR0a1VLnjQW42XH/h7t
jcVu+p8kRPMH7sbwXkAssnjgwSsEXN3qNq0+zrpemsxBR8VG7ZorUbKcZjsQNbZP
jCMhPJhpFySl98rd4fQ2gZ4EQKIWgiBqECj9vJ/9Agoj3qrmS8T+cKTNFtfKdNxs
bmu8PwN/C54ZfTb+5zlyLgx8qubLWw3J/z4OdzfMZtldzsvEZcBqFzDOR0RhG1uI
Pa2fU9J0qvRez17MGgI9GsKCxNauM4CqlSnEcT+zxRS9+9jSt1+ueZT/68VRgGwc
gG6F9EUq/t/CV+QzTp9VVuBAo/Z78GeY8Z9tTw2UYiwCQwFJxEyt0fYzkOAzC7HI
AWxs4CXAmunnFYOF9SXnKXu7HL55jetE6x/6Q6BZmTs7cuO9aXmneciDWiuRjS+R
FE0fxWBXDVo7dTo6S0oWBzad0w/PoT+Iatgi1CdAMXFKpoWNlUXnJGakOpxI6x6V
NE0codXEZgOjiqRTiioUVE9+rYVpkLUfFlZJtdR7Am4pmk3TIYZThrsYYZZEI1un
qXtDk7LUOuf6WSsSFOx4M55CYoD6WmOsg8rrv/SZ/OTOMJr6kCxHBG/MiLJTT98D
AN5S1zMFCge79EM7wt6nC2o6pfg0wT/NpZy3dXB1q7uOb5MEw+1ysGiwqNxDgaB9
KU+HyO9+S69ptH28P0jMJyqlfoF4o8WwZfcU2Fwp4MB90kCpZpxPlh9cMx8+T3MG
dtTd4UYlhdpRkqUpOh3PMBWEM7gX7uAtb2dxOK4mM9mI7QJcj3vIk/7tqw7K2wj0
0VW4wV/8XhgvGolhAcA8RcLvu0xoP2wkj1MeDoVcLgavYP+BOQ1p94jOxeL36gLI
jLrg/Ak8MZuDau7WiU3GqeucjZYNsUemPQz9NgI+BhxOgkfZNzYpxwP0fzqcAXeS
Dp3THNRi5wFWBViOhD5uxsZuzPcSdOC5zMbt8RGSMiWsc/k/NBy5Vc8jm4YaReOw
+dPNz7sFGF5uHYaHbrGNZgW/Ji5iflMRaZRBbgqwT6oBiLOcTFXEcYvrsDiE/Twa
InkYp0X7BV05ezAlcWXh5D4sI+BRXbglAoD3apJx+VrYlvztQLv6RIhudXh3Kgjo
b42Dlpcol3lfqoL5JvGkpV3ZFx2QpBNV+c6qIE+5KUz+mzYGn8tr5Z4mFm9GS03+
AvlkWJospajwnnlWQhb0N6aWU7HPZJBxoEcMEQ9TlV0xNN0hsyWoCTgwsWA6TUxC
WZhZO3q7JZdqeNsi5BvygaKZWfCTvlvfMYI2dfpM9Nj+sH+kZ8krLZaCIl8Sw4tZ
pyMyiVZdtie/Y+SVBkUm6IKaJSxlLyIAqaoJr4LZwJ3m39w+2pDuOw74g39ILnZp
32kJZg+1z6x6tlZ9ZZOpFX71wd8Ga1INd6VIkvmvNPyZw3rDP/NCoz+SI+A/rTHX
kgqtNFY59Qep9+LFyEtL9+TBmIdVrka9IoloppSMLLvXcr/3oymTQXYTQdQxJEIy
CA4lkwaekX3fdhK5HwRBytbDxdvVO63nsFlbxRt/87S3/GwRUvo67YyPEfFyWA0w
NKKxSu9mx0Q2L60AfoP6ChpjBy1/bLPw5O8xvGm5lERK/IlNPvfRFiJ/iWMYUc5M
oeYZIYSOkBN+diaBxBJAQyMU5Ja0fxP+ssWSf/4z5n46jc2fFrtcITiMFvA6PMCp
6cvy9v92p46iKKO0+zsEKrLAcxGOqJ1e6Sli4BofAFq4qn8tlc+AShgLHQQAApee
PYe1mXbzcku6ZqHuOpHbA04amLo3hnyZ3tXMvhO5ue1qjetsG1riuaC43+OD5cO8
ZYXzXGjk95GishDLnidHafDMRNWDNJ3WPUtGuymdb9JXneOmUUwwzoUhmz+XiAQS
RNwJKKJfBIw6xsztphXcvbnnYVqWgksB8bFnHzPsc2Cy1BPvmEC/WZrKvfDsvG3R
4046i4sW5jHsYGhqcLd7JSW7GoEUl9ZGM+M9kqQm5bfZeflgphkcXFk8zxUbGUqy
kwhIB6I16sjK+rKTBam054NUh/ug2CnI61Th3asLavoPXWx6uf8ejiRwZl1cBZNP
QhBo8GndRwM8jb/QjDcLG+kwOxdCRN/3vQTFTZ8mSeDkxZKpPUwmFSVRFFHmcCAb
mPv+R4jif/NCVQ18s0Tvu/tQojW+9DdlcU8oxedHoGbivLRFPTSihzjqvYRa2JeH
AhZAltSg7dh2BB6wYd3hP8wJvcdhsY7z06bux0+kw3Z9wPFCuldRDXES3mOf2Q5s
j4c/JKHVRxjqN1zaNY2Bovx0vNTngXNphzlm02Y95WsrM97as41d0l9KHzSfR/8W
UR/doAR5IjPHybeo8+dKjMSTEozBAa9jsJTlgck71EW3wMecCn40sxo9pwQlmMDq
W5L366Sz6gXIfAn/meQj3BBVmq4R0tFS4yNloYfU3FygRc3qsoFzP123Nn5usEAc
P5kpLFr26P/+fjiybdb5y+BcqSyweVzgK4u/1ntypgdNji32ZW26oWWfLawo7VJu
xilXs0PYn8UChSGcnFv+GIQRRf148rV67MjvHzGn8s4RDz1WB/DFJqNRq0zOQxV5
tJraHNWa+w2g7p33m1VrP8791b/7UewMVXGEKZTHR4gCmsAeWZSd9twLoLRsayOs
r3nhu6O3qv2acZphMuAATBT+pR9dxcpgwymIGtaqMgD+WF2Ljhf9lqceq0zq01JJ
tgLWNKNjf27JiBZMCr/HwDc8JLTRevxn1VIlyshspw8H2GCGDyIpDc1opLkuDwMO
bjRXSFyvl8PqFC3sm6kEGYpnQEFb1mg4janLLiu/53eIDORx9IAieFX2s3ikBG5y
v7TfLsfN4PNm4XYopjgyLeB7J/CsZI1o5Nw6Zc4PbuJcG+qPrZgwPkntnaJzSZ1W
nFVEFu66UBTa4utiyWwcRuHxRtk0h3N1P6EwBQaeEMMtohIVkFMuhQOKVXZNPqXW
3jYqBOH2wHH+R5AjbpTpjB6NZrh7F6Z5qQz+/FUfvxONeN5q5j+6p7sScRfUr2Wf
am/A6ImZ4V7/JU8zSxtkOAWx6L2LDFWuZbI87f3jo53sU1TZ8jprw1rQ7Oyj9mUO
lhBdULGmcXivZd3LuOUMHGyStDdqXBkVH+sV9+jwfn4FoMvNXEWQukLAt/YY+T58
qWb3tdWhXsjjPrFtcuCx3c9SFHrc5Zp60+3sazuF9U6+F5+T6uTHX+8w3KPSjcTv
V8TE7SPOdxPCUU1ysRwU4DqEAwp3lQ1G4lhr7PXks4c4u9SVJjj0q44sYXFYDidA
442SP+ZeNbNHg6O4EzaX5oN0Hpw4w0F1BBHstMQJ/1V5hlWeR9wlhNdAi0cpUBS2
+0TdXFrBWXBwjXDvtNCZTHdTeh8E66rG5y/ofSX/kioGrcj43Yty7n76NuConlhA
boGJac9D6DPwHHH3Cv8kjxR6HcwBVz+X2coR6JSHd6JEgFEJGp2PZYffJnubFJE/
aNLPbvxTI/B3uqdNeHpSJ94o52kaAgoK9orBaaartCFwzyL9tDv91djGrehYZicA
YYG4BxR0LtgH5QoShrxnPHaj0Vt03S3xMgOmSV0TXCmvtbBLZlUn62JmF+xoT5fx
JTzdT70lwYros1OidlxiJjysJ7dPcEUkucDfZXGv4Vv28Jve2zQVunrIGsBZiDmz
V5NpPjN27tyLE/lUbi8JRbUpaGLvzzkoiuPMqAtWmvKBgVdFka4OAWkosYaIbuLq
WIV0RWe047HYrbPJsh3Mef1eSAZYHAmrGOYrnJnotO9RTq6joqrjTpFFjPNYLG/8
OnpnlCNIKUiTJBlixw4yQB8NLxH8uq7PjaCffT2DiwvQHaZMDZareMeP3pT4b4ON
Ma0Jx+5CLVxggUp3NfShu+B2TsT3Gl9P9+HTAl4NFEDIgMC8ioDJCAXdKSw2+J5S
NLVWTWsg7faBbCDA2P8PBQZlgyHbPVFM8HEq1R/GhljNzYp/A5AK7A1sW52DxgJz
8Tjmdu36D8yCqyEKowVH3KeRaE5AQ8ZtlJS5n4T3HkytJHrZtunx7ZzCUZzRKaWx
ArlrbSN4CkWyj3fwQSrkdAmpozOSFp9yrFcHUBL40eipZUDx1HBsvwEN/lXNZZbe
dh35lO3/5N4iSMcaUSO4em/QBFlqPMHWZpFEAnOJ5fTHgVioCVJSWt4Lmrzbs4Kw
TxSkrrMdAwz3VH4PEz8j45GSJCIGA1GLbcsWzlnVdq8lrOmPnbiu4+7j6DogqLUn
RBTrSNCJy+aiN9UKsvXsVSR0r0DXnnNEmXZWu5bfkSa8h+gMM3hGsqhW+BTX63qf
EF3+RBZV2nC7Pdd8pQjIm8+hRZqHlixAgSEFJXPyGF3cXhqcO8+2u3GdzLhWNFPF
Purzq+Df2fpohuTxjPmJ7Vhf5EnfyNtBVJoN6ace5y9wpO7mC7Fps2/npu5sC/M0
zhYf3VkH7gyHksSgRrQeBYboDXaXvzcLfVnKxRTA/xWkuMxEXDUsH6Y37igJHHVg
AKVohQbALxLkxaM15M4fjq64KHjgCWqcgdVx6Fjmt5B4xJrevTr+LKW22PwedMfv

//pragma protect end_data_block
//pragma protect digest_block
sXJuM9su1dVGCLYveEHltU07vXM=
//pragma protect end_digest_block
//pragma protect end_protected
