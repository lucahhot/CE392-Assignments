`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZwEvShC5IlYF/nUm4lmROMDO++SSUW6QKp+rSsI906q59IZX7A24vRmEevuP/xH3
b9NudxmWYlTl/MJmaQLZpPUSSBxVFwcw265KoCvNzZjDwFkRTptc46mlOIG7mV72
Rz5W7+J/v1OvyhSQu5LMvleQ+bSzvsEY+EAKcWGkH6s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 121584)
1/LlGZCfpTmb/o36U9wajMMYhCbM2dxpT0472fs7qCwIdw9J0r2WdkWIVgKZu/zi
fOuhFaGYCTnmrjZP5fsH8m452AoWvlFu8K7fwv1/KrRHQqZWcFM3rLkYZxYAu/TK
4H4j2rcI7fgXjziLeaUVwAsio7NtHWMgr1itQdl3gCxebydoRYSL5LEpwwuYRVlD
JD353lDzubVs9tLUb0kQihFsZmfSXA9rMzhjJc9pO9korZTRISCPY8ylz3s07DKP
FRycKluOYm2SaVXhszUxcLDrJTBxhiOCh/lrZe0tBGTzIAEo2/oLG5Hyz81neDmp
oGAklkSoZLZDQEulVmuAM29Gtagv2A8VsnXcyEJzuZYnDF9e40F2Qr18egb2MP1M
0JdbNYRBMVIwpIV+TAKlfvtCG3W9D54OJMQe8Dr83DJR6qDBLgUz6KW0LQuBCVGj
c9XtXTEoXNLpF7yVheY2++69rBPnyXj9hG5B/3dY218eMf3ROd7jAqD3I0yTe2LJ
7PJiz3b1LuGNecJUuIH2ES0V1O0q4+Fowrg7NcyBjFw0Vu+QSh1pjq75rgRN5slT
G8a8pQx/kjeBYccx/Huk7xhz8o+NxB4N/SUdXJ1Ad1d4ajxXxaeBO7sX90iA3tm8
8Z1lwz0RSvmhaH+mlqyMt/QZjH5SzyzABgeDG2Ys4bn9QeMFe5DQYPsNEgGcXgjb
fdTS9ReO+haRebX8AtfornY8x1ED/Akhzd0KhYCnzF/TOcRKXIS1jMVbmhHRPk+0
HEXdVeBHqeg6rIrl7aLfyVE9PDYEokDK14in0PlopHcU1aW3HeJHs4H9X/uRy603
Q/ls5/FgNZxHYDeapx0aqC+B5+ldGvLZoYUOHS4HEe1l/XxYS53BnCEehpXe6qsO
PrAdNhPWT8kgNhKxlZSmJs2X+wxTDGHvEQSoiChSsf9WeQbENduKpfqTo7kHfBZl
VF+CIdr35HHOwbVXx1+PtVnL0Giq6cdhvsYD/XOtmCRUrc3/5bVlQxyKY16o4Fk+
3sTDqmcw1IIf+RJznWxemkEMuun6amju322xGrfzXZ8NH62/UzzDHqtI9ml0mGY6
86+Sd//kOo+GJj92fmktGdtsjhb0LvyhpsAXd+InVdKGpUCJSA7HdzToq7EopE3K
o8Q93hu5qqUO4rYau1btYSIIpoFFh8Q4OUHjyils7BMfI6gqRoJPBXCyfn3b327D
e+obHrfs+Cq6G0jvWaJcvo8KqKoNCnHEUFe3SGJfaxlnbFvLAkejIfj++5pIv0RM
UGT1pnctsS8V5MEA11dK3FIc+bVPnV97bkxVlT+H4LbEjE5gmeORljCSYdTjbX7Z
jdmNoUvlLaDR7rWXHaKfdQ4hrzJgEP7dVb7TAE5wOSO9S6VTnOQt1UsOkAMcKRiZ
EDCHaZ/4MqO5M7BMvvOuFDV1pRmjbdmP73qL1fxCbwTMJq1dMvEeZS+OgX76Gbos
Qbp1PXBsi4LxaMKgCanTNl3RHC61i1JVuQWQelsn1zFH/707iLEPpj16kHnT/75m
j+3TCtAxgME7ker9qPjiwxMVO8dtOcrxLFvEMhQWuXZyXLsR6Pg5FL0RbUX905wr
vIiqCHZ/MnpBeLOXjP7dnrE6WrWzIRmWmNSQPtxHo69AEIAXCRdWGQqOccr2KKZN
77PBc6lUmcIaDkFj5NLgrD20imzQr4Urte9clpNT+Z+qIFcIOeg/wcUlnzsVPpmG
Kva3cDmJbMIUQ5qTsA+3SJTrW5zhLDfo6oM5EDjdT3a4SxoEnDWAwf214ieNflth
Lkjc0J0MWBwmIotNvDY4j+Rg+fwxVY5pGqV8ksruOclPne0a76j81c5V3VXhXRwU
M7NOuGbUjMVlaf5eV0+FTV13U2dvqMq1XGh2pnZskg+6N2EvMWvroZCEYx8UlL4s
9xvuyoQmP6AVNi3u844k2dJMPK/NZ97i8nR023bRpiqMTFNPbDrDoFInIBzf9J7c
/vAZQT0WyBXfVzobysP7zPok1h3bU8risjJsX5p49QnA/DLfDP9sVmQ+1LDt1MZR
9LlMw2KIhYPz36EmsAiZ4PIH6ICiAo2pp9+H6MzPJLl+xsuYgp1Ld0Eu60lubCde
Eujwj1SYp0VCaj7TNrH7Z934uXwagVWMxg88I8Ly25JevXPf7iOeQ8Q+ctLv8U2O
BMq6G+iCnDCVBDOJsdA0OlWxeAH+p79t8yEF1w21EzMaNspaig6lYYcyP8irwMmP
SSQwKnz5KPfTmnU3A5HMts9aX/yzWIF1iU0Z/JS+P+U5UmtcZqShPvz6oiLC+OvZ
46+yg47/zA1wCztD5hx9v3nzKB4achI0Dof0DgRIL3QSMB2eszqkbsXNAHGeKhls
xomD4KANis+UHfWbME6bp4YoEdv74xZrQIZqfFXNNSu/S/1poIKpZeOS9/M0S7FA
NKdS2onwE9hGVXXv+9uo24BW0mmBibHaarPAYmzhYknUHFwPYd9rXl0WKq8O4Dm2
QAhzNyCa8+BHy7TcWO0oD6VhLBGzZXU098u+opedfks/bSU0NduS+1GE8U0iy263
yobtBmKfMgea0ouCFYjgUqocCtoEHKOLOCK0UMcrKc9tBFpVwgyK981vNSJVZOx6
VUr5bWaUGc5iUmLAntxviooYgs2B08F/1vQRARfdFRxGzM8lNMpim6OtHgMAzfK1
tQ9i4TdLOlS2UUshlZwWmvMXGNcPoIb2T4x1Wy1MQFefeLEhc8KJjus/6PIKW9hp
GhMJ8B2VfSkFXOYSQaek9JTasWzGjsWAI13Hli4BD+v1bWYbn1XftPVtrN8jF0Uo
8r1fVKbX4A0mbepqtzW0Tj0xF4KZvYPisVxFp62sEDkeePaiFSi2RyxAm5DkLfji
ZHf3eb7RQtjJAyV/EE47B27BmHXlH0oKdBakZZ2e3hKl397k7S3ZrZes1+xgVHMV
9c37rccSWynRbUFZLpxKuvBx/ONd7rfQf82ylIPq+rzv6LtXueHcJIRmlAioy/4d
KaFxZC1kqN7ay/WOCzT+QwARHsVf9r4N+pbzduVvlKtt9SWgUJ5rulEdaWWarWTf
qRPyKPiQEy4rXIQ8e5YETlTQ4aNSg6JldwEJSsW4OpkWcMJULyL7NmG/DlDJFlrG
ySjwgWITDY4mlzSFDvjxqS54Gya7/88DzN+WHTlXRkaE10HGebwEhnNGABtp2clm
50vHHRGm2TqmYEFQdDH85ayPQ9FgS4SL2XY2z9wj2HDMcT+x06dyZcQN62m5y4Wp
wVMRz6ZvFMkN7xfMe5Ganq8nv4sHs9qYGb8qo5C1NmCJUsbYqAAjKKBsSa8uEWoV
E8DByCTDqdz+18PbR0Moj9mKg3QsbjYVC/vrbNtxBhjsLQg7APzXpN1Y3+yoSm5p
eGGKDSSZywPrQKhBsDe9xIveDzJLEAFTGO5IrWz53lDQFN8ngxg+mbe1e27IaNvL
KqA6b5BWpUAjaoL86K0D7MUAxJJ2efDsAxIOZCiGN5LUmKonlByJxLqvsCkQ1+v/
UYGEfieWDoHV3e7ZdjRuP4ALwpxL/jS7/kmQIFCq48tBvNnUS2QMfGN4l/lKHBGs
diA0q7jy1o+IYof/2IhSHM3xCzu9gXnobuMyAHhgxD3KIX6HuPHwpV5p7u1bZqjv
JnG7+oJok8ZlHQ/0LuemBmpRV1dXIYvjnoO3WJV3HgsZf2FLzBEoCJJnawTox5HV
ZwuyOCrDH1TTJuif3WMQd60rDvwISK8k/sdPjIvByTJbS9ulLTaIPh1B80sLeQtF
jEOHwzZGjDtqbsdv/rfe14NpmtVOODHdkCWImFRPgNSzerYSX2fYXf6BAohIhqu6
rLtZj3RvtSeE4Ai5husEJmCt2R/9Ynpkxzl+sBINOEXr7m/Z6uh52z+lUj0cuDtB
WSW9jtdo4X4LVLP3TEMC7+pTw/Os3CconP1c6qyULKnHdq4AZWWfR1vO4G9WLYMW
AdRWbGjq2kqOUdTBKfYBPjV/xg4TqvMA39g0qYgZethcyUpVizx0mUROpj15Q99+
H6B0aEjomiWpvzAtdi3VORYHvKVm1dERJAoA5Y/fY0Annt4s+Jji8VlHIxguadtM
TOEZ6Jg6BF5NEWT7Iij6ZAVnw3rsCT+W22Nva4ny450kDY4F0lgWFp6nW8x1dBuT
GPMuKhAV7KKLqx2KGIVM/E0Z24Oe6Jo0gUo+ZFHi/Qi6nxqAHFofPbMVZZeCX7fm
IFAFFsmom5MxNMSxXqaQsBsHxBJdZU64NpYnO6BUtSX1sf21ZrKBjv536eXvpTgf
tXFVIYzXorf1VelHvqPsoAI2K75HVFMd9i1KyYPbtOWCQckXJl6T9gjNyrSr/1Zq
av+GE02Khq17KhxnImltXGmIxvNWANR/qYZaY0wlGEiM7qgrGmX7qjV3BZp9r1Ha
NytdPLD8THVU0T+W1RH/c8eVNU3vGP2t+PUMM8x9DsG5amgZMWGdQUY0D87LxMF2
PIo8i5U/vPE4Vi/wgx8lS6+efH6nWXrN5Vuz4kAVziMHMi7zVWruWyoG0ZkLfC6i
myv5Fv/WHnkDV4uySGQgOKrBQ86YLoxAa8L+17J+gpenaB3U9kJJB+WIaaCPMZL9
NjdZNx+D8+gYxsOyEEdvV/TzfhM5YyxR2Y+Ofw2PoSBxHu7bkb30eGTL2CC5xZTj
kj3E5wLP//rqE6bCc7BW1VlmtnMWZGlNiAV2/wgmuiiWcy95sDH7mOCTP6pCyGhH
YhJxDDRkX4MXxN+x7iZgJdsLxsrVSSZ/1Pnzs/hopKp1lV7IHLpS5o+NhXdL7UGU
7FFLfv0At7ARwowKT6bJcleULXk+jdE1CdTtPiE10Ut9arkTqJOdT4bO6LFizXGu
Y9hiT4L7uXCYYEKwivh+ZaqX3jPFuoAF5zh/giLGZSmHcmip2IxhIzY1QvSLidWo
MZd+XrSuvNZ7LUw+TlsHwkNf3yZiR33RWFT0ltXKbL4F5UxcuwviAF+gBpua3hNZ
knDC6xFmxETEyY4Ljp8N6GpS3seDnBrqAItjLvydUmlfsyQy75FQVj+l9/j6QJk5
SMtI6Fa5l+Xb5j3REqQPaPX6LF28TBv3zilX2Y+Vf9yuviac2hyBNs9Jcc6G5EiL
BIJ4U+kaBR6DLMR7iaWj2mrA7qYya13gpJg+UUKTQHcyA26v9gGBOAB/Uf+9lQpC
VRDcGN0DxRiGNudpSgwcH23SAYYaW3GS+BUwlbMZycmaw7m042m8GWsdhslxQgKe
aTj8B0EWzAeMBge59gT0eKSNHEMLZdoZ2GFis/npKivirwlbF5wuqSIS16yqp2ax
fNLZQ6UOGCKJtffz7MRVRrJWdkIzXQ7YmXfQLtKxw3JlveBJw8gmWS2b3ZpzX83r
y0pybE7CG9dECrlN0t//q2hbyKyf52ZNdVLXGc0CheM3PLyTNF26pxEYEU1/Yu/J
UVIlhaifJeHg/sPjf6s/j68pbRneZRMmdi7p1MHzPfXc0dLqG48qQAsS98zoULp7
j0+be66hwRurER1gcNa/bq0+sncqpgShujN+82AKvlIPITj59VIaojIL0dM2UyUB
t74HXfvd9znGUPpxknhJdqXItx5dWWpqn83IsOuzYBpdQPMwF5VugxtZHtF5JkrR
9qeovVPQOBjqwqKLy5bT55CWv9A/k1k2dkIJ66mk3etCgiKp6CZ7HFS+fdDGRbWh
nEqXcvESaujtDRiqzN/YTrANy5wfjUguoSIShGlginGmQHkUW5ABswBDHX9Duivb
xR1BZf3+17+DgXcR8cQu8b2bijOivHPPHxIpUKUjPLskP71zi4NHtkMaNdGyzkwH
4kpPeTHdnxVI/EGjywVzGC5fHC343qItq9Nth4wrH/JDc/POfze1ctiTw3q4a7ip
JjNLIOTKjIuhJNze9bLNs9XMX49G34St4Kv7UYFRw6UtydcNBb1ZADzO53QBSIoT
ZW1rdlfo8/jtifZKWUf/UZHhIG1NQEoMwfsZeCt+xNFy3nCKSACook4huEgnxsv9
v9EozJeQhT9vZRsXO0lcwOQgP588QBCxxJadFeXhQNrkVrIRHylsZR0XF7KK4epP
RwWQJ7qRkB0XhbIATxg05S6G3Rls1yasy52gjWWvyjBOku+26d0Ov6oQoqFFEiiY
A50nLWRdrlkrj4MZGm3kRgCCZsF7oratY533BdR/mDr5SGYcOkNrQ7bqAPXHCafV
bOc02NlGgJEjZFTHWWXh+K+wghiRHd+WuqcHLf/3lq6LYQ7cJpeDPgnpnCh9cdg4
CBmOl6PZrFb9pjJbv1OR7SXvi8UmEE8t/vgbJLRPOJ0iDZ4YW2qx7P8ZIMs2HYmm
CqgitWQTxVcdnmQT0cCGiktXpDX0tB9tskeU9nItKtWV0yH1McXBUPzOPT6PGSmX
/lzHxeSPglLubLf3DkBDKFivEzDWFOrJpQffn4Bj4poraaBQIzx4SjR6oOknk/Yg
/Iu+/iGtu0Hbkm4spq/8YIS3Xr1Xge9o/Qxvi4Hr9eFR2P3wCi+iiGotnhdpssJL
q0kTEdvE1dKZEmVMLgIxQiUKTerkHIBnssTl/jkCOshE/34KE0eCgrXJVpDtwPtK
V7R8ZvAZRx7/VtZ+WPAzAWGW9Ijo4NBo1h+IBGW+e2TvBZI9K9ZqDir24pUqI2rQ
1Cs4XaTZexMVv5uEonproE6TyVGMzPjPBjqNOktsxD223maHoWDJQIiBAolaH0xB
Y/YuKq8bmmTynepjS1V6CQt0CK7JN72VelXSKhmTRhYCPE2ueqC4l2wlI93qzK+r
0jRrB3vqcHBtJebbHgsNHa0Fwo6QR+EsUCUgfYouv09IZ612FGQuiYtuV074efAq
VaJoZkpxcI7WZa/xGvYOHKmd8ZMaC+FeNMh55f6VqWDxEen26Tgj6HYcE1DIyYXD
5EwkzbF65b+TG/gKuAPa+xkf8VZzwRPsAXMctks/pwONxomPp3HrIuKofNAaDSUc
QRz1A7KuoSodt9bfpv3x/MHyHllfi4vfXy2ATeJb3iZ/MPKKRmer0ej8WgDi05ku
umNB6814n+485hebmcK1Me91SVak/UZB1rNvDnNC04EXJ2W5tZXNaXV47WgbMJTd
pyzu11CkM2C9evEB/vrGe13uIZ8bGIr910vvlLjH7aTCISQG0os2bW9Csadyj8Z0
IS+hV2eTIPaRinaU9e2Tjks3wnt6bFUsLqCV5RkAvZB9xc8Izh+2vyVjWxGcQYzF
vKqMXF8OOHrO7b/P9WZRCU0DZA+8JBm9DIsQDnNVN3ayw+2LJ2xgjJRH3PfFm7BE
3TgCWgkVLvUBEI5D0bE4EPFTHcFJnJUPBFOgmGwIAqEfp4IuBrwzYZHmZIe4pohh
M6pBsZ12qOqkZVNthz0qmmzWfIjBEkuq3vM4tWFLDpbn9L8BjwZkvnpU9RBLLLSa
WEIjUJgW2hERkEEDRRK+t4ynwG4e8RzDIeOnXIqDCFV8lQAL3aVw3OPdJSlEwhsy
4gvhWHg4DZDmiZzxqIobTTXr+1WqxMcFzGf8AVFPTTtYh2BXsyJ6X681EH2/sRNX
m/Q5amPHkLF7nEtcCYFAyJ3qpT1Hc6L7igRnofvXtJVBO4mwtU85Fkpfu0dWnP75
1noEP6I1yZmWBewbROEqmEJjNiE5gDnqA6ZSYd3CvDL/bF0/5BQBP/v82srx+cgl
UoRUY/phcbgiRrkA5vpsaDTvb3ZIA7wDFtZiOUUVB7f2IbsAwm8TX1QY84slUnnK
RW/FrQNwREADeYjwBGlrdv/r1f5Vwx58MWFQIzZT0tGJ+vJYCJBQBoR3as6BNdgN
/CpaMT7QH4BP8HyZyFnbC8n9nsEd8mCkbn+fxEIX3OP3Rtlycaa7rlHYcSYmvjkV
kKsvc+XSzFuuFsXC7tL0zD6okF94c1xZqolPxEiVgia18YIJZv600r/RGmparB4+
szXCEkqUPazqxK/1e2q0W52lc710kuhKTGpepmiHfod6ohBuIHw4uYctPJJh3f5n
BTLswYU1hHXgTfiZc+BUvSL5OKoouwb0NTFBB3fLnas8h1duDg3yXMI8+rDpl+fz
PIDcxHVvUk5vUamWGtpKjkxWw0Jl7Tjvp1boHRGpiDrB9oKPsYWGz2hTOtGaBH/a
4ODjxIQihx9hWzVOv3WK7LzlbSGjV0S//vTIcv7nqQtkyY/nME4p297nq+q5ymYZ
O9i67iCxF353MveQKiGz3gOcr/Rq/YoY9gHj/FV5Pmfinc29BxG2BB7odHfrd2Qb
vqKx/KH5WEeLaqctIHLJFSlmX/1hRYRA/NCTTdDUg3CYZqDFBibdg02HIaVjIzvj
RBb4TEN76hAjotrQHMOqW9YIkx7s3bxJ79Oxs/AlxUIWKgJ6OswVkBi5WujR2mQ8
aGCQPbJSLckjrRJWOvskbSMdK4k6/3dK9E8AUAN1490TyTNVXyGQ1iTPqFF9UskO
TOmv7rv4MTebZdRiDuOyrE2uEtHvCGyEGFvYoxxOKr2dA3ReYAxVk+jC17egH7ri
CtYkTQT5wgXYmH2s7qM28JbtmOnOUzgpUaaNBbbTyyfNuUHwWUgO8FDe+0bC/tgg
nZBEoIgkgFJSJjeS/xOjskbVNUptUbzHNLQtg4IPq65m8G+vECVMQDFfy/+H4x6V
/2uMrtthhLkHCAKIf6y+cH/vbJuDG3HRUuQ2RMvp1JO15mQU5k5yjEuZy/ffubUr
W3Jzc6ZF8TTJQDDhseHPEejplXGvKNUv81bDjZDBspPLSQoXJQTaB+1fgy+weQTr
j3So19Uz8TJf6/tGQ1b5G9RL7niYzsFCqxAs7IKi6z84l633fcXPQQSFnQh3KHil
qGe9ThUVkLzYHCMamrFKwGvILnWEyO+efzQlPh72r40V7bpovA2zGVUOUGsaZc9i
lJ60oFaaJ91HSWg1KthaBdvI+szXKpZ8TcHGwVkihu7GAhGvgNqrGK9YIL2P9ESK
3QsFt2upADS/QvkX6/aDkb89KT3efIG4nMX9LCDmHLUMtizqd/99z+M0Xr7dqlw8
zftMalu/7cHzrS/3kiAPd3K5KJM+mzBIUZxTt3terjVmMZTAK8wdK8akfV7WGk9s
QoivuyNDvS48ChOAAgSUf2cMqyr0AKsp91j0e9O6JoVv58ogrj0PLAGZkjRuTN1i
zfxuxsIeSqAeFvVi2RR0eujUBpuoqGZ6rAkm91w06ROTwdNsHjGeM5GLESjS5FRH
I3vu7k3RiQ2qdPK/cYA6RY4ThGFhQqOCkbh4mGoho5rI4AS61r2Pa/dOjkkdE7KV
N5IKa4wlemMo6c6KWH/8piqk/cPWbNDIxJ9MCbTTAkVfUHxm2wORsZ58nQdGG+Ir
TZAWNGm+jfpXv2oyQ96H0k5qC3f78lsiKcuKR7+sFfa7yho2XVdICcUgLnbO/dDU
tNPzl0k23GDIWHcJMyNzzJK/Iv1uyFI7tEpXKX6mkAgXpqYt9iR/mMXschCY7AcJ
AmwUG0VuZc4Gj/7q2eltCWB5ByXq5IYK7sMdVP8KXJA9zXEePfFdTnUybsAAngfK
uuEJwxgWM+KH5fyijw7X3hhGdJddYhpaPIxU6AoZhKcZs1insuCKdBzSSriPWTh8
paO7nW6z0REHvS82M0Ghw56HoFBle38LCz0NUa13U1wb6VqfkKtdtB8cBPBG7mwU
1T+3ZTSqPhDcNhCXlXcT98/JU64/WhAmvZQATJeWthQJimrIEkjZHOCLrWA7vgRa
2S+6ysZaL3/6bRPiVOSY7xAEvLH2FOMNFjnG/z0Fyecy13W292q/8mPDOftSgwSX
FZoFO/cIkurgu3yb3NXPGXL8bju6kIMy8f5YNsXFlXmtnNxWklTUmKPfg4dWJLcV
dq/2EoN5eXuK50PacHW9r4sflqh1OGrS95nAGKIkFTWv1qV7xYBAcXwHg8+qHWgy
G2s5cjXDx/CUraHcYXZ4Ibv5GXldtrhrriHnJJTAROiV0A1AEqjXx1vL9/5pVL9X
pH75j+M8CH1WRpdzuCvuXnYuSAf2zUtY49/NNqDtg+o6VR5am9pWaP6WnEGNEmjr
lYVANq8xl8nBxOn5A5TCSi/c7UI0pTfksuRbC/4K5FKamhgm7NsBuzxlnCrL75zl
ns6JfT3lqfZL0qAS/AcMGbmvgadK5QhYuDwO8W5tJ9/ZKyJdF4VFz+OFmZdzR6F2
AznrTm26G8bO+T7qMp+qVb84mjo6w8czddR1XSTc3UwEYvX9GcL2l/GacfgAbVpx
BKtxruw7ochTDG1IBZBUd30HSUpyvrsZ8QzDG0SO1z9zZrmlY3/z+ym8tPBlM1k5
02z8OXTPsLUO86JL2wZIR7bUILQKJpBsx4+IZJuKsuetZhC0NOibWafi7ezQ0gMj
/rRkjCSPIzoywPq8TDZ+qCJqfbcRMWtOacLsae/Px3g+XbOVOxtRXj+izEcV+lhc
qOYvqa7w3p45NMTVOJJBwPsEQ1okjyxsTgZnVA0X5Zuup4wCEFolGLSbX0qGuBLl
4J06o7000OlMuTFsOeekjiAZxk76XvSPSFXYR22PhaQW7fOIecfldUCMO5dhCvlS
vd+KRsqSHJulhU/x7emNJoyxNr7wDV8uJr8mX4/NSRzfIp4UfxSfxAp6AH+dPOMc
lYkhJBViNRjQQrEDe1eBgYJxVAGJAXuCDh1knatu6nBmx+4r5LGxoWiZWgSgaR1F
rQ4ZlLMQIxZ/knQY7g8WNpwAhuxhzk6qShHanW7lHtX59jPoCOmYBHBNj4ucLyMr
9i/6a433UMG8g/8uhqveeY0C2/EhGLIGoAbNtNwFsEg47BC1Vi/D69lma6dqc1SQ
xQF0uQW/BDFSQDtFD5IwnOEm8UnVxPiSNRtHDF0vFZACj2EecRZR7LiKMAkrljR9
ZcMm4gshf/zI41/rIqDeCLCNPrb5qVT53hl8YWL/S4nGQrbrcZhxelIaw1XblfkX
44KK+e3gWn3sxMlB6auu9PJo0ehocWNdcNff9Hrp/yc+5w+yftXPQYk84ZPL2gyP
g53MFelSxXEcAdIXEOU24DAQ1U2j8nyuxegbFwwngbvEwxZ871n1J1elfTjlQVm/
H6TUeGrt4iWYXu8XpQJOxNv0jl3h8wQa4J8dHUKc20L7vP7kw8Cw6xvv5UAvPfgg
h/tKVGsTLJGvovpJqeIHcq2xRnpK0R6q5SZ0PEWnBXw2B3x5wAY7fNvoByw+TX34
yBDKGWA5rWodSFPMo1cAwhTr0GeDUJIiQWJGyqDfw1i4YvrF4iq6bs10V7SB4YuL
ygaM0vRKki97Pc5Yz2msRflDpIly19Zsxs5wCRECeGGuzFyZ9RgyPHpO3GZDCcEt
i28mT2UW6RcnjxPMi7TX2bCnaYBMgbde8jLvP2aVsbAqgqPfmcWEAlN1HfZvazkL
zpBMnmUkTRocPdNYecQlN1VbfPYAs0SFEsvDWaHgB/dDBy2a9dhaU0oGGnmF9YXz
+D6tc5KGSaJIKZJFhDpQSL033/HgKA/nNYoqqYsN3L1JJ1c7hmf3u/dn/6o4SXY6
1ponFUg+IKYDFAMH7EwXH5gkybABi+i2n4dhY436/EPMAOimNr/O/wtV6B3OKtUK
4zDeZQzi+/KC6qxYcV05x9SjUgMsNrKvZGcpTER2n7f59eNT+MfcUoAt2u9MyWz0
JS2/JAs6nyJe5z2mlRXhBLZcXYYqOXgTrR+IfqrZjX2WEvvt+ZhuDgMre9rd8Pg8
8oEpKik2DVEmNeUTXDQAv533anMmsxr2MXydSiJo83ZrYD5dxB+yO/Z+YnSAjGgU
aLku9COg5E6D+hyTUubiiWQDp0DjOy+Brd1d75sKRTsfF3b4emrVP0TQcJlwTP9u
kX2amsq/dyO1YnOvRMQ5miw4XV6VZTwe7fx9GJM2S5tNj7nyKGR2V+RYq+qe3bJG
ZLwJavU3hNN95CBHsTXA0jeqw/mMyg+kkRnPWXmq6IBFxPBGqzVQqYzs+6Xwc96s
A4tA5smSLi2dxQ1Uulb4gkfP+9ok5cGcC0552iVa6YBqEhOk2vwCiTQLpX72CEqg
6wrH5UwsOPioUBrpYdfJh4bzDCCM1YQJLDJRqOD27iQcmGKn8RXIODaHaBABMUe/
kFCY7iOlBJYkoEn57CuLAZMIpd6BYpBCVuoX1BZ/f5QAy7lZCfZfxRBy7E6Y0IRi
wlk4b3iwJ3hDoYAMp6GV5HohYv//NM0ITmjzUam915E+PioOBHtoQ4kDKTnxQ4Y/
VFR/eDRjPNtdKIoVuVZZE9wW6RVzuqX2snreDZhM1cQaDoQP4KDaSiJqmXhd8hxn
tAtLk3aTsCjCVGzFbgHed4wPMkDZQqoIHvrJRY2kuRX3BmpBr6UwIJ8ZeOlu1F+H
VYWt3U8PjJPSYuUAa6E3u8d1BOolcQQntFNbU13WAoEN5OBshNNt2tdTOXGrJXwY
VIabDw8El3Z4ZyvXtNPD+nw7UJ5EERt1NFPXEnjYo6jrs/L2Z2iTnB5r14UJ5NrH
fhvVixsu2vZGEeDH4psAmWV+kYqPqJBn0YdHyqqVoX+tOMlT14Z8lvJwO9Y/utgw
skZiWbyizjS8UuA8xeIrQhuJNSqSvpayu88zgaBTf8gzTgXZnso9m5b/9tR3Ei2W
dR2GeaF5reMjwLEV3giGcE3SLbe00jXzR4y0+ONDIpXAcKzCa8Wp1ecpOawbjxeA
qlpCvROk51UjuAkHTlPhcoaFG9PbixU+PPi/PkEGFqewF4Rg3nKfEIU9RzaeasXg
wRxVAhz0wGjIv2mGIeL/XJMuRFIvPuKBJM4eKb8gy1x0TT3Sr4V3jzN/EDWEUv86
q0eLx+NrP067NeUdAuDAA5y+lpN+sz+qSmlbNaSBOZXJCb/lgUrx3me5IeWfOegA
FmfUbVAl3XwuHgHjsu5M1HcGJMc4YF4Asv1/LbV7uUTZQj/wz3xrGhQXcvI9uDbw
yBLo/HZAWzGo0KMvssCp1kvo1O7b5aNCuqY2MdU+bWP0KfIUmuVlvoRUHdUU+ENm
Qzvvh2sU1duE9J1+sWWT++nmBOY16eOBQLaiRysyFFtFcF0+ClARJryUt9ITNzaP
H54DTg1E7Yhpwz9Dx+OSHXYzUavF/+2PZNHoaM6ALXvqHANZ1SkGWuXmMev7HxHn
6cdIQ1CDJAdTbBUn9KLlEktPMfVZeGdxbi3l/de/Z3HpV6NzXiM0VdfIUnBY4Lou
LAeyFHmAVw720FQRIUm69IFHlJ+efnEVhALvYgfn3i9pMfYYJx8mt70/yptinZ57
2SmfULAg53Oaj5QMBDCSjbG0E07g0oRfPNrM4RPx5cSecoHaMBRUMZTpq19EAT7c
3o6C5qmvzbnCi6P18h7S48WWj/lS118w+v9tJaS2iZUdRUR/k89zBqMzjKLV7PMA
DdKLAI0CZQUEJGvtDlwHuU1/dqxgJPnLEcpbVmcJ0Qg0SqXKWnE9FJpb9++R7uHR
5faZsLUO3z+sbqe1aE6l4O5LWubH9i+3vgVrGcp/nt5JnDcPE1K49i+ibxCIRqR4
MVck2Adi1Oe2eCQzLsiyKzTEo14vR4RVAkRhokv7MrO9j5yfXwc6qT6LlyE6Im5W
NdL9jLuV8ZzFFmToFbvTHt/MKyj/CE/doHsNWuKEw6GCZHFl8YLDexlYtYbtvJNw
bR23A5Q76DIrC1OIGQ2qT6W5aRT1Tkr983ZDs36dVaZbTCbXzDemUke4tDcba0fD
iqmmOEgpZzvk+IJbBem/m7K+nxXItWUFwh+Jko6eevL9MyXXKMi25sYHDHn/3Rz8
x/JjHP6mc8NBNMSMFPduB3hIGExutjIlOY9PoRtRBh/ENhOIn+ieAVZkd/hW90r0
OhwtXDCPCkKZZzp3aNbJZEP3m+4fiT6nfaWk4HmtdRs+6/+eIaLfHDi4WA4Vl2EM
QrNKc2UFYGnKDx08azFdcrYhFO2h7QOa6j7mbfmb8+HbqhtX3Sh/ZbsDXK4XOrCB
Ohxpc+4c+0sXw4upyyZYb6WfnuKFIGLip96kqJYIONBR88UYZDDM9bnpS1xGoj5L
A7yZZUJKKOJ457Fb3jkdStXXB3GE5fHrje2zsujHkVtlB6lRh84ZynqwvoaqDZ8P
MOgySHtqlyYmWu7afQ4E9YoiIs5y8g8cnXq8WTq4dza9buJy7y9LBrLc8mcP7AQ0
hSRtuabY2cGxfQ6nakqr979Ufo48TvC0yWVHvoLgwiZPhGteiYwMu+x/GQTjiK7/
n6HEq9X+GMEUxWuSs2qZZsRoO+BJ9+/3FRfLjbAUSCn//RbMJK70v7IGQRWdLs/U
obtXQtRhx8yWaRxnFI4J4gWVk/Qo2YvADLcNsqY2XUKd5oc5AYnzzw08qgOo5oYz
QEH8ST1/btIJcAdOETlMS3U+kXHUBK879c9L8bNnsTVqQBlhOLolzwn5Fhiy33+A
k1oCh6GOJjMch32cRFSw/mlbydG9bZWOp86EeqpCOQv5l4GwLZqF6TXp3l6cfZAY
u30EolA/mhrNGeWKBnSO7oyZDEwaWVSLe/4HL185BttZks0SGs+qeZEH48QgSqNi
zjo1vHAwToG32VNjcjx6r/72pHkbctFM9G62fyVYHpQWkv83YXXU/6B7bBcXnhVp
pW9sltE+65Dx4+l8QUCyB7ZxGip1yboFwJNTyxMbbs2hy4BQJl+xMQ5legVoEQrG
KnoxyJ3YeWng8Nu4yaDwBRlVVeTRkBnoIAVd4ms50KB9SwGlLS4/ARNazP1YBJ9/
r0Xd4araFozf2N99DtQ8+j2PS5rcSe4dNxQBQ8UC3i8XQ2W+suvt8OgYgwMae17c
IjsaXk8T9Yv9TVFuLaE8VGmfp7DWYVpBYcZFbXFkbxp4rRCk+IphZ9fzJDtq/9MN
e4MwNSjQjdCb8saQhZu6UvEbsfUVF8q83J7tvut/kLMq+WSr8YLtohpfitK15cTb
XyuupRspofRlY9nk76mokGOSeQ6l1qM/KgYqmLdyx/YjDnBCySlxTON6NeXFMrs2
qKxR23KFlZ/0GqIQ20TRnhtqCbK5UsEe4zEOsWZiFDCi2JHWUWb7bvhqKXUS03Ng
YlcnqNc/XO/psBSctMWHRZ9GCJd2TT7VA8ainZcxIPPuIY4h1J9jDy31xKnts4lw
TtPIPMwZj0CtL1PY9fqaXdfldefIuNG5e/JI90y1O8R5KV/0PGwrFiYT4vXStwxd
JjdIXtY/frmRmXO87mJsLd7DS/7TWvTVG8y+kFxBrtuOOiIp/xZ23Tqo8MPuxwa0
0np3XIewH3FUmz/dgZzXbrYfFuF3aRGfyubsu/XIKtSsWTAWDPmrmBGSNJyPfZJh
BPxGlPjVyx8qEpPTBMHOH5aZOYQR5WCI8JA9enkZ32ULPUOrLWSXoG9+JVIXfsTh
kEzuP0SnmF62BiCejmvrzVe1ZX1QXpwSnkIH+TmHXufhrbW+uL384tqEs5yexYi0
Jn+Zn18WqAPHyWspmny7clz7ElovLdAhw3bwZWZLqZDToa+XXP2zcrLRbhMLgfd9
FG/Ai1I0mpO6cuy1SJ/4yCvA6DbZqSToPLu1ZMI1huuxhJ1hu4w1Hlgwyy9vAdgD
PoWPKJp5bLN1K3m/G3/mnWY8l9ZR7mzjfG/M/zjR7VJkAGMlEGw6RJg9Xj+qQST3
CufpllG4bfGYVDXlmCcRMNqpEm6JlcSE3rqGgTZiCkbZGJ3dZk87MFb+cztwg7xN
vntXfggXvqKiod0t3L/3ZMhFWhLbZ8URLw9mmlPOJo0tA5x0UNLDH5yAaQ9yuDqR
HdGx5NVL0JzXEf9Pc2aigEE26vCH0ZBi8TO6D27qL72rb2uibD7pwgRj0cGKJ2VR
XUYCt+HVsjAIgBiFw0/ltHXDKbKr1j91rHC0KqGwzKvkEll67UkIlgwJuq6uY5Nd
xqtcPjvBuaekakRYidX2iIbJnRRIALcw63JleOHC09pRF438L8tQsHtN6wsDOVGm
n3EjeI3jmGTfe6f94EQGGoX63aco3wt74ZI8sAsuuoSQVhDciCOz3xMe0foYm7dq
34WoQhQh4oj5GzHFeeMz4CE6D7yQtPncMjVj2VIe1efiOj78kQvFkoLL4+Idpt7+
dOeZ6y71UR30OqZCTtJEwGZKboCH26TRJzMDwtVCD5UBiMRjkyG3uuBXgzcXqqSF
0nsQZLvJrDxob7vPsLMDBx/9/IUcQIigzkJyKFJl+5iSjjwsd+nkhmxfEuquP0lo
bz7UZSz92ltkid9IKTo1gft3+0NG8pZ0maVZqNDSWD2/6WFWKacF4WwOzv8sLwoZ
36COHF9m2krWTdowWzjkwweb5WTsLHB7i8nBr7WVZUn7C6RXwKnSpFnfATvKUpvO
vv1f7kUlnMQOaCT8CA7CX6CPkSJbpV/cigFdK/j8Kxs+odtWc8oU+7YJEF0ym46i
BflRKSa/57lsFaUD9qOuRjT/NMGj+1NADOqF41itQnZKKUPOtFLPX+ZZuSXkSrFE
H/0q2S+6Oclk66jN+NnEYrjC4JlTGKRXCmBYQuthM/4rPsotsSH21DvoTCrE/CdO
4mL+bklfPQ9YIDDPqZyNEStYa4B/fdD5vZvf/YTkeKkRfE2E06XPmxGTUTt0v/d4
9hCqH+yZ+xBDcvmFi/7anOXYSXco2kFhZW7WmehT7ol+T+auv6Ze2EtlRiurOtwd
XTrTQIZFVhakPAwlKkIQkFzlTbZdw07mxI6ZBWxiJjUvXbhKxVKMsJaKmxlqnStp
jyioi6kqyBYAJscKfTjBeZZ2KQjiLp9aNMq/xcBDTQazfMBsoyoAwmbEScY+nOcV
wZgpmmhh56QGuGB7gTjytQjpkGSYeDbCJrX7Naw4fq4R+vyr+YwWzSs0V1s8m9Im
vHB4qpa6sy+9tpArx8kXj9cWZO3Ks3xE7/uK5WFN5Tuthnu1sTO7OjsUdHp1CTJK
PABt84FRyecC/iu4Fb/bY18fqj4ONP4lX5TERNXZPV0UQ+V0y/ygt6mpEYhX9ihs
4IjyavUXIZNMJFPjoLQDFQ4JfKaXVxemys+X5RnUbeiYcIdHtGWSjVfhcvYtrX3Y
M6lqgRDV0coaVXa1WlpC8n41WnaM9y8UWEoVm51XYIEtn+wEvU7NYYuEyfAceZU1
ZRqAsRpktGCo9fyQiwjA3zwieC78zmeI1i+2qxwLzoIQr/33qeDpGcsyQcBn2cTn
d+Lrw0WoEBYJN1rY9MbQAHYmMYf5II2My0gbuDoycPk9+GPeJxILWS5og/BOpqI0
ScHASVOUbEQpP8wnzSS0OOYbKLzaFtgPF0M4f0f2rYYV8VsRZ0ELo+poZIgZ7vo4
Eg/hxdttR+78TaBJqQDpuB8BzLgRhcJjbKH3sTR/gNTfe88QeGsinnrx1PDpj2Y2
+2YjyQ4KoAEjIQZJktD4fqd1OAVKLBamxwkFP10OVgoK1JiTuASqRELrzbd2Ii04
kxu8R7AIIQvvBYOAkzuLTOYbRTtU/rgkfZcW42xTPu53kSDCR/4IdcqwCtYZd39U
w5DKCyfOMImeHIUVZwQEKxepYap+4/KawZqSvOOn31kG74xgxZ0YCA2hvvO6CBEc
AQEp3C+MMRURlRsx4bqAW8Xo42qPWtl0jQKHeviEcPLml+H0WPNYrSQsJ7gCfjIT
reBS1ZyJBN1xaRkmqpKvVw0ye5eRpC7IZeSEabPWwJWOaOFFKq6N4ubaPBEESj+7
aJdBiGa/hbL3SWE1ibOQe33ZZqa1P6TW3fIFAmjFqROIyij6IQmtuptqs52/i3TE
0KCqBkCX1K1XYXUtu7UrwqQhGFD5RgKRpCwGcpJP2squrVLOBkBdWB3FsaNenJv7
ZooLhUyIJeVZEK/E6A2rW1z2VEGPlsXE+FXS3BYlFJo5YqwORkOp7GqOIlyoOvGu
URrmgEeWpQG/WNgtOqYjUG2R5YJAWiym+h0hys69DRN1jBs7xh8eUT/vUs6vLitw
IOjigyExrvIYpCn1Uh2ZLvhgSg6qI2yiA+2TwxopUsSkILVn3c7IkwUh65PPS8TP
wwptKbyu6fa8a4gErtfbR1TnN7qqtYoexLtZddCljBGpu9TbvzNkwli/DDTPCHsO
JOM1Bz23tR6fA1As9dj68d0QU/ctzlp7+aZ1YaOcpmJBFON6mHy//XrT+2rH6DbK
xrrw+ZDWHCT1XjrISeiwL+Osi8qcNlB+Yk9rw8Ud1bfDM6m4PnxKcmPzwG5+jBUm
R2TaHup46qDYR35pigHxSiss9NxG6cQ9v4kne8ACmPcvYI4NKEs29Qjq6m4QuwRo
iaM4sfmZwMh72bmaKj5BWKA+otq8Mtp9/qUwB1R5ri9kaCjvGPYVZ3ELGnUHloMG
2lw2XgWqkygW7ZTjyjZz/Wtn9tUwAd4yox5+g4Sk0ixQ6klRhxnuuw0aybn0LL8Z
qIvB25c/FEjxsUUnbt28uj6cXP3Cs5uUC/zuRLDwdEcwHdgR8UqLmfOfMjswCuDG
CK3cSHQR8MP45KkhHgdozM00j+k6XRYHMa8TC3cYT9eSntmnLZsiK48TRv4VEL85
e1nfIffbzMlOLD6ydZNQRFZ/AfPZS1ykXUDivVoZoFab3E3mH5XlcK76n0mf2phz
yShgh8FsYA71EezvxgladOedXMqy9UxhmD9s7mIuonpVvKODIP/2TVsIXxmFJrq/
m8W/q3i9niC02buRZHrOpMFvgFeX6SoMVD05VkVsh0atgYz0CYYbvXzN8Y2nPXld
T6LTNJ+JtT3K8wB4YXN6aYQsKvTZ37Qtt/kttTLtel1BAKfRWGHw78fKV2dwHv1K
0383Rj9tHcwuGv7sa8myebBeTFmjNj+tZX+Q9Q7w+F49TBANnxwCQT+lnIdeNfcU
nzcmUFpwhW6FQE7448IjDIhBEeNv9aypQpuoMoHqfUeZqRMbtf3Myb/cs5W4V/wT
xKk7SXS91cncCH8TgFkHQWzgHQUFK+U1VciqgSEwGhN6m/XW0ya8gz+393QYcKJz
PoFugNfT9zRdXGfQhTcQYQ4eTL1iHpfLTk7TFmWm3TDAGlk+sCgn2kxEzbj2LVs2
MK1w+281QhrUfCMlUrGmDBlRZRFCwkdLh9swJZFx+OrkW4YIDGCe3t0XXAf0ec+N
klYDJ1LlOXcj9O2BhCuGx3NcAa3Mpi0QgGqrh4IY2uBo+7lecgz3AgHtUx9IqkYN
JTxgK3F/AjtRB7uuZprSTGXftqxM4hJz9V+FkYBIKFkPRPQRcDzKvaaGkN3SJE1E
mpWrQ6vUsqvZB6pL9PkBIFxlfkM/qcAa2IhATzJwlJ4euKu9aJyNfT0b4smBVMns
ocqrEdztnERJLRHtNORR6TalVof05ZFiwp2NrHDG+zLAa3UtY5pVqys/HmUpqXdJ
PlS3PTCsD2/kSyW/U1p5P7GLbeK5bs5mhJiCvLKh+7DgyaZoFHVYUmy1cwQVcZ3Q
AXkY3FAkCzpkoMJ4U1suqjUPavVhyfYRycvJAQ8C80M6DgSSYSia03aJ6YEtezkn
F53N1egk2SF2gYW/+Gu4GRJRfHNfO3gpuMXy0oHx8OoRDWx/k9Bz+Wd5RdkVLIx+
ArYRVQ8qpprF577fmu2pLTw4xB0+fjUMAAymo4jfxGnKaROzuA60em/pWxS6BmjI
vCYDU8u+Pruscy4SzrOj680L9UKdg4YTy69CZl87JEdw0FxTgMhdVGjFf2+Xm+TF
J56abyrlFrJB+HJUyM34Uzq3xa9N6Tl0hydq2B+jQ3rk2X1zVNUx6S8x6EOmIsSZ
8Pc6LSF1EODnEiSyhC8FKml2w7TlAmFqggC4pZqMmRPzp3TKe6mcLHJa+BYUCNul
c26pCZu9sQmjm4/aryC4s4a/SsZAZ8l80ovvRweUOn2RtV1qZCBhza6bt6WSW35s
SxksJZhxebrtZRHKd2dssKIXyt2RSzj3/YvoO51wVxQiJUd4fM8k/ZYYgPO7vU5/
JMULweAv9jI3vdUVJqo+L7oJK8kt+7GvYvaTLR0KjtYOkhJLzeZrVfIabk9nmddv
4cKfSepwZJhH30R7GuV45O66IjnSZtp9K1SQZIxaz2Y4uKP8L2qSqR4/jQPzgD6r
oYEW0ev8HW5P4NNwKAihKCosTZfwSg3e74meyUfJSiVJlsQ8ei4Gnyb38OZF7sVX
5GauHB9ryQAl7xGpSU5Y2lbAE7/R7wic90kntfGZaaCXikPFKTOln3FjKo881vrh
0kZeblKkSwPRvqhFBUerZKGTMAmFDhk6IQNJ7bOTBFxFTeAD2M9K1Uot3+EPtOCg
tkCjnP5WavFgmuf2d9vjahrsNtNlKVGpV/iHW9sGr/FS4+vNOFjaIiyOhmg8lX0f
J0Exj6U+27jKJM1KDlI7plfurldE6ofqyzi6dQ0xA527ElBT61HUMsmUkjNwb8d8
tB3ABnMoWa+pV8JCm6Qv0omw7opkeR7BLZMvZhj6Ru+OKQ+n8CL1OEg4yHKJ4Ft5
b4dUsyPcKfApqtmo4xdwcCWX0HFw2d3wA1DUbTZClJXBUb+8mVEG1kDTR0M8Gjm1
jdhrCA49hwEkTlf14xquz2ONWlDh3cU1E4HeGxwAERirQ3wRXpheNwmDc/s2+6x4
i482hM1FflKR44wzYkuRb4QLVVdYkObUZIMuF0axWyp88jYvEjV0qZnOEFKYGZGa
iNyYyAbPjOjk2otfMT9KUhB12cMgFuSC7Z2hoebg8iqrUel9zDpD2XFi0ZFOylee
nTvcd8513pIzddSCpPKDVenWh+77M2AuWsN8m5gRC8fLL0OKbcbXsBgCFWBHZkCx
a7BMVrIoMTeVqFw8b0PHXqXmHXwLRVbxPDDe8MSGgo7vnRyWwHcW8bruD0rB65lD
ozJUG77Jm2Rpgu1g7gd4Vn6wLe4CTDy7P4JxqqXj6E/+aChHW7te98wLPnPGcmDQ
LpZ4z5M+SXNJgZiGRDSH4fE0SmmUTYWiMfXiUKWeiXiOuc1ycSSdiAF+vyd94okT
Rfz0jX58o9vMePF+g+RSLZ6YcjMgxf+zS2vQuN1UQzFlSQkm/imDFsvCDnpfrPud
NXH72WBh12971JfSIvVpti3zGClHaKwSAU0U63NqvSriX7vPEwZaLZWzwEV9V+Wx
NtY4pVK1bCvO1SbDuWRNt5PYEQ98AYpEWpQ/sdDMFxmkhvroZ4h4qJDtrKatTa+7
nHNzduNVSS7wuATGkWntN5Uz626vj3YoEjlVDa0G/qWnKbH6kzpM31q/PNz58Xj0
CLQvZREa/Bc3TLdBQ2NpafoWJ2JN+ntufwaoR5mWLBqa/W+7pdidQpHz/f+LAmXh
9i1rDciM+L9xTmJDSO/MRZQZP39uhAqV4ytX/d+/J6mVVXSTmeSxU4+ECBvTMHg2
JG7yTkUoSpiXOH1JCnPWX+G8pqi/ycht+gzrw87PR8nXWAF++0TPK1eGacv2QGVq
8SYzIH3b5zdV8LjlsCuOAj0/8MMW2p6okYy4QHr1+qwLGwTQ3NliXjhj+Razs9YY
/+EGK2VUd8oG5rgfhtxPIfr108Mne5uuA1S13DTIzyhzpRvs6yYf7gbAh9MSOSFN
/eWsJzb/Wbk3rENqh/EW013QJmN5MLew6hI/peGn3ibs9xqFnkKfOtcwxKCV2wiE
kaocb+ALPgsn/HKasTwblZtz/VMEqv4HFdrIdqhFRjc6SJ4cH2SWDLjvFjrXyUIc
7xd5EQdWahkW+OloPX5ct4ajWcouTYyT3sGRBYjZvyU2+u7pRvdqU7tZejo0A907
H+h4gwbzigDk1zFnFrxw9ZxF9hpxNV11sdEnT/5Du6aG/vZzeuP5ib9GKoTQrLBx
Jwu3Aosj3esfwgrkPyQfzNYpdXddXD0igNBq/Poyq/NHXutqlQgd5tm+cv4B6O3M
ObhFOzGE+9K3uGvVsFZU58ekmznGzsxazTJenvlYmjEqMJpgN/4IzxO6dFgAojS7
3BOPsmNug0cfYuFUG4zM+oLxZGq79xOMR6cNeqbCWryMO7G4i69JKZFMo3o7FyGO
PemToDDLkBCdH6mcI0bwmn/6wESgotekI5VW+FEF1K0v1OWuhdJut7WteLbW/WHH
KmfOYccTJHs+HzJDi7NrSk/5PXatb1ldc3Ubnl3B9y/45MIi1CupE1RJWhIQ/kPH
2C35pYWN5QZfXhYJ48B1dJFaLKojjVRpa1lIbIElOqhKOeB70QuMYhfpMgoc5z52
/41KVTPmQBgHjXuZOWQoJacPQdr1fVMg3x1lZi1P3/qoEDj1BFjZ4iUrYp/we68t
2lJ39hxq40+jPGgRAgfldqQOP+ucnn6fYQJVgx40pTQovmYpKt7YJWIe6S/LnePq
cUKsKbC6SKpAmruOe46jXn00/f8uqDurqT0S4Q5e0nilr4MUr+SGPv+eCuJPWv90
rwIEH3bsNW01BS7KyDQyG0f2tNIpAdcyZ2pG/x/S+jkCXu5rwTV8KYGAkL4NO0Zx
HWgWM0JXgGPEKXdaX4nAdg3kDyIb3HoaRj/gxDo6kLSoCOYaQmsfsVEJdwYA8uTA
UwzRtJVUV/+u322Q1fGoC1FwLslSlcLoBuV9bHPmtGI9LNJ2v12UlBXsmmFku+/0
mXQO3/P19eHHQRxPazEESc6kS+a486YFGsuCIDq9iQMiYV86Sp/IG5wWDTTXXECs
pJR6KcyAq1j4r11pGKd8u0DcmQZ++IcOHv3+VEQ1IaVZS3cNeE5JO1EYuNWd9LEX
FbKhEpOEzjZ95e8F8ZQZ4NhrimvcitoUaEDhFoW8tCb48RV5gzy75NRiGNMuSvk2
j3CFhvRKEM+XG7E7yoLezy2tFTooQmN4N5PwDkIk+QWUI3eqFyQ7Pk74NES3Z0Yu
hVcQF840MjxdIdL2MINOZ3fTLXyiAjaiXFYhKLk5NEXvM3eXOGRk5aPUaPFpTB16
OYftIXRttvAUoAiRwEJZfvMUVTplbpMGMEoUPnzEILQv5NgcMYkfC35QbOkuB6z4
IDPRv/hMNMG/Lt4Zwh8qZ2NpXF1Figniy/DwBti2qvAaxqKsLqvy/JzO0UkiUpNp
BqjyK0LZo5wSs/aXS5YRIQF1U6gzkePIxQTWLm3cddmBhDroeuhTd1NBrHzT8vzw
tkOiQX+OFxWF+RiQyFe0mdNuzlCX09Zi15SeyGm8UENI2BboqiUPCY9R7JebdSMe
trW/XESLGHjVu3DyzJEp0T+6Bp0TDxMwc4zDoP5QF/hobmd5HAu9pt/Nk7yQq+XA
Q2MDBUvam1rDpwI1q2Pl5Rq5qXRyEPHrafywdNoXLoD0MVlMPzvELYCC0vNfBpQo
rhrmoSnH6A4SKY015+WZ1+Ft00WNkt5FvqmkmQzPm06lq83CDMhvS38hMzv1bJrs
GeIB2eqWVokf7JyFQStF4l1U9Zik1V096OYvFj9x9Cj1KYnWFIIt3FL13WdMwwsk
yIyIBpAfkTdKsjvlnRGZcbEaMyB2GdoTOowyeg/3/1S5foaVFsLDSLkzqEOxDWbX
TZAc2fxkXcqT/r7J4OkVwZb1KkzHCH77xElyCmQega1jkmpya223X7JAPZHMrQ6k
pBp6vreZg48bDAw7cs54/8SnnkleSv/AKAzmSWxzdRbfBVKxuRTEqRpmPr9EAzRM
JD9cvK/7Y9SbM4cG3SYOXIWvcvjeDmNylD/PRO7BcBkFDOR99NzDTATTFfux1GOK
bx3hMUDFxs6AsyOl7oUHGRBb94cN4wqx0PLIEY7MxRLseC3OES/e1IjTZAaAKYAY
izdRP5E0qkv3+WfuIDdljj+mwW79aBT0dpjgSddzRBsqJSiVV2YWho1PtRPttfT3
5l4xTBQW4rUYv/HOIhpnL0OAB3MVyTkRl/00NaDMl+H5YXT+WPwC9ytAW4kKrYsk
Awvk9t9orrTtbfE7FUcid07lztPCi8PoYA0h7UG7Oq5F1k8A2FMnmpzaerR20Qtu
UP7LI6kpt11p8LHjuqyxbmWaoFZhwWoPYzgNqygzAGgHzdjilnGybdMxFWQGx7nC
jUj5N9BMOh3VL+/mVJq8BbBMM79JskSapYMm9zLWuXLbkF6txfcAJFNiON8Lacfs
x+WzaWKOvy8flLpT+gd8ukuSGBrFFdMRy70vQLHmfg2j1T+Gc9Jo2DDgxZ1C6/a9
m1iSCNRotIYMAGm4tPenDbPK+uNX6Li4iL9ZaJujBzvMri+Z6E2ZpRgtu+oJd81M
NizKqPrnEcZJHYWAtNOPa7QGLTGN+Pg3jA7X77k/Ir1JB4pUJDJoO/DniqwdSIKX
WIp6Eua3sPvAWfoeW1EK0pgOwYiRA4b5c7TL0CI1fA4t2cyMGmUt6/eFJj24CP+I
0XLxJwZRyc350hptOUUetBvzdXKf+/uLIZigf3S2o6uFCJ7ppFkppuP354FKVrCB
BHM22+sS28iw/vRJJKP4lUJzMMZiAOLnNqPovyPJHvaFaz0d6IaYwU+tMJdPlXyN
NLSRuSyWK8frFgtsqWU4/HFR9gOLTI2vN1jgBzMwsk4067kQ45VAHVK5n+qa0r7o
RWh+WUWgalc9BlAGerlq7fT0mSftAlPIjO/wBFx7I8tCeSVN2FwFAauK9KhhA+x+
qqw9F/08IDeJMXZq9BQzNVIFlFfTIkfjEyfBtQCB2FRanbrajoMyw8PqFEoUqOZM
JSJvpPFlG3/5t2ijexv7ZrKWRp8bMqxXRcWjux/s8jxyXIQlw5de+D594ZaH1twy
yqTh6ddaZ7YCza2HX54x0w6vX/nBNjJd6vvPyZXEOZMn8qO8oZiVNQc77HH4U7Kx
3r8M6TyB1E0YPWxUfeZ6Qq9auZuJUtlSAK0ZUCfLx69/UohO4v7SAvP9KteaeiLx
+3ppkZ1knfJF4jEMXzE4NtsBEj/tyPS9KWRLfwykSoUeR3svK7mrddPpA2ylUA5+
Nd/hjPvZYzASCrnu9w5o1TDhUdILmiHmx80x4U7rA3fAf2fCYxuDvt7cQkat+FHX
AaaqbFZ1M7BXMkuyALUNZkTH5/RkCnqSshsO2tJ4t5mWeAMBUhliUMSIdboL8t/A
hXoCOLfNbbiSUZX/7sYv3qUa8OdxMV2ez6r1RN+IR9bvWwvlrkFcX4kZ2RR0pAZq
mE6YIAEIde7zJxXx0v+G1m4ZKV1DNSRoc8Kk1h9XPlXt0ptSDzT+LSCeJZf2kHxW
+EUD2Vsn+QTG0ihAUYbN0nsqwLTlaS2Ee8gysZhutrZRW4VToFAi8natSmK1+ek3
racftn/PQabwJy1EQVX8agFU/wMnp3eLl8nL199u+r/PTtj5RIMuBcQUBtTfxCyU
Og8WVB2TMwHecqD5Tx7meBPqDFsxwi5FNePREE/a2HvtvSn/0kyIV66EiWVVDuLZ
NQBETGPnFHUyWGXWogaB3Jg3woup5w1fIVCaJbsl9Iyj3iry2SyZfiJufSqeCYOx
j2ZEIfr4iMBL05ziT38/rleLSjDCgp7AzUaS+PAnYseUYGsMJVgY+fkdVMRIUhIk
leqRn9nOJroD7tEoxkHXKlbxyzxArvNdo5cHFBKAt+BiHgNZZAbTOyF9+k2UgMnq
lVx37KVSf2lIbwVTmmufOq2q7i/KKiySAz6CGc2uHA8dKm+QRyqHdFI6V9WBnkQJ
feafZbs68kAua/15Z6aC/R9XjPOBz5m9ZntYHiiF0Ftlmo3VX1iZixH4Kd4xbGw9
72nTbi6wyXAW9WbDzaUtJzftbRRO2SBrCYnm37dNKKQO7HHN7tCh92lJ8IRHAjWE
I/oyHMjDZC3Y1gv2DYvE2durBPUQtBU/7byLBu+1SdjtghCSsk1l1ku5+qrbCRC/
2aGbGOW604KI3BwGH1kCKq2u8orAudwYQoDlqv66KSsqe013LtM0aNe/8lFjFD30
QyuriM3wSzpCgHV03WpOdjs9CtLZ+dRgj+0/mOAXuyibjeSd51ULJ42l+rDr5aku
nny6+nj4uJEzmfWtgcCurNDW9tgJJWMJ9F2mOEzdWPdS1LuGAQyJytSgTEdZtLDw
RBTEHwFaRSUGPyn7Cw6QcorgnZXEajR+ruKhKAkXpvmGhWU2nemd+hijadtaQalV
jK2jCXmBjKf9+Zo95TOk4rmf5AJBKg9PaKNVlYOcMbUUs++7ITstulc2/8PcCq5I
cm9iuQLqTUaXG1y4mI5gmOKTXjx0ods8zV1yrL7GKJ7edjcvTG0b297Zakxt2dNX
ERU5Fppitpp/nFNKfdtdhq30hwjDSTPIQB23fcW4acO5mhgrldsezLsZpl1aJTAL
xWeJmC9fbI4YjMYVoyWBW1wIK7/WerlTqLKncBMoUaKYfpoSdzJ3CxMG7CMgCsuw
6SarQNnqfp1JOQTe5BMoo6CpuJJXSdrS7ZWLG2TgeseqEwyIMm2rnF6VBefn84ZH
KWzJZOgznqz2VmuW/642aoIsU+Qyt/H5XezqCQpuKkFx5vGPJQBhBLMJtZg/0W3D
5bm9HO/UP5A1WrfNPApNdDEXn2+gaY4LaGK45g12Z3fNJ8qLJ7cfuYleoJfa4B/V
OySAJGM7m3Mf5hXp2Y+qOOa9XNCd4uU+LXTwzS26WRDq8azIold5fOLSVhSZPAZT
GfSGxG0KMM2XTiTR7lgUbKNCAVqym4FMV8JMtH97swkOHP40jBoA8qM6h1NTzJ/B
SrLYQNyyWQV13W2jJgAYGZM/KsuBF6Bt6/QoD4cuIQZxiqsRwU7o6WkX/aJBX8Rj
vSOjFTxQyACW0s3roteQqxEsfe82/+L85Zsok22kE9YG1OomsS/JIqqrYwDEycDB
k3g4koe1/zzmrelMlgs0ercv/AA2Fxctep7AzWkLZOaYqyy1g7AGG8RDHXPNN8AV
A5nFMt5B3fHq1in3YsFgX1wTczvyJkWgkDBAyb+ZWXyNqqj0r8du9sf7+g+35paZ
Y/1MOORQcEZ9Qf6KFw+FBQm2Y0i3aIrxCPVTWbXbfp8cbpyAzwSzZMpj+pVjw7tI
QLawmC995vnS9FCQMCUAALCKNmsaBAg/BWU2/pP5UyBsHkZENjuOxC9T6ecrlIZP
n4UddCt3dnQ1lRGBfKaH5YJ3EqMUpnhbgh1chV3wbi9w5YmBQ5JjwS1hDtAQhusU
KTKfg/4Gxw4jjQiZI0GbYUkgoC8CuojK5uSx5f+PMw8ODGL7lG2ZcCiiixAFkIRf
4aW4qGa0ILiwAMc2BRSjE/H1JvE7wP4IiShF95z26FMz4FSKkusNwN8nxi8jtiRO
lvp9xvOBL+YGfmMSe2iTASgmeLMHEM2yzT0KdUqsh2dUiN6kuWxWh0w0Rfl5fMaI
qOEj4eIekBDyY+ARg9jrVRcJJhg1rGuy4oyHmLxkQGUDjB7/xkgwwAgRA/p45IxY
nbtSQegvQnDYYg2EUSyx7vQpjSp001PXfYGR6A1mhXpytBXzJMemQAXPuc8LM2Sk
gTWEROq3vOfDAKajwa5eqpBrOkEae3YcKl0uTrD/UZe2CxfhqcZymbFw6JDczARf
sWJT8Bl8zsUGwsEUPrq1D/Fat6L1bcRzsFa8vp0CZVisUNt/FfJJnyoAKsrhTTqh
COc3iKPsNQBy1hDnNSS2sXNvBoYEOLC6qUhGGP3DkLCMubZxUwn3iL7nHjJJ27wL
YDz0aXSIglCWgmSkgfPc5nfhpSA3YMAKE45aSC9KYhecL5nglPjf/tFvWSElLamP
PPri7E03UquCndVApBky8kRIHKNstHc7xc3W47xovGuAZxWa1pe2obRs/MIevwRK
HkXBbQfUvF351oDwQudoZwDQJ2li8ZVegyrAcUJuXeo0JuxwIu/aZdgZPCOYQVHv
3WTfHa0RXxkaC+EGyPJ70yGJMRKb6sbkbgTx0Dvzg2XE0oors3bUJNbqzYxsRkVk
di3YWPT8lzaxHgUc/gtYJ+p30LBGlmPf1jlBdgSpg18m1f0VT1c0kLFHA1r1TqKk
9Q9xxuws5bpv/wSkqeIAuTWlyRdcsqCPvqX+miqe/jgw75V9Czf0pnQSTLVyGjZm
+vt7GS/9pYrVGG8zzVBsjLdZMWmq6Kt9vAkTFFdvNHPYCAwLSlpukQ5BfQ2lish5
g87RhasG8FgA/6Jg+1aKvN1Uxw1pN/y9gJevbhKG3o+zrXTpP1m+WzQ7RGzCy3Hw
89DoBlhx1BzDQ/UwAUK+nXsqUG8OE4GdYCEAEYSmjEw4ZJ4PlcFobQ1FE4oI8sdY
KKC8U7+PzE5ETbNGZe+fKIUYrxE6biDLzn0NggGNCDhfLqb3f0nSQJrp9r0friB7
3kGtuDXHp/wPOGVDt7FX1CHm8KovmLTjqEP9qUcKUYRmdMhRzOfrqlHsrlD4FDG8
g6RAbC1jwRFTZyl673NPQVy1OSgxJwNZs2X3KIv/Oav39KsdgwYTXx0+RTH0q8rZ
z6xYneI4k7LgWnZbjgRLRRF33ONl2ZIoiZOYkZFTxaJ6pyi07SvgNYVxdtQ07Mtd
FsQlqjFeldglV2vYqWU5ozeo8N+8JuxmWlewWcR6DsTZe8y/IC3pnZHDJGebTdmi
uyWz4UnA8OF2OuoY7Zmbx2ary4FN2IWoCIqLuRYLnyNAOsZKhbJBI94sZ3nkA2UR
O5lOsEp55/SBhxxCna8FC7HJRxqdqprsuPxbpYAYUFN/OFF5F92LyL5Xc1wNlJO3
a93tFabIoCbA4EkgIjWSYEjuoL8vsijmf/Qtg39mFsW0P/mZYD8TiW18arEyzS12
74ZnhqVm8J/e/o9DB6aPwUgnsWmTyhVrwhGEefG56IeHUqdtry9dFLZNPoFfBdUG
cYWYx01IeACnDpgtMeP7/smtecJ2F2UqK23mh/mvAfYXbZXA2cVEFKDwxmPoXUda
bYHpJLdiEd0u6lGt/zBqsN4mhc4+fUWGAd656sG4o9BwqbYXrO1LnDkBVRxtz2+U
JuAou3HpK8Ed9NszaBAzJCGxKTj/ir62t+NHYwm20PntXgkQUdC2VGgaIOM/O3uZ
y9Vve6fAEtOqN+AeHTyWrHzaHzUBwoDu8QHelE2t6OuPgfyXFkyf15l587fAhlnl
bokHjFEdQD6y3TkhypNaLUzgyFrTQPUJxg2Rfr7XbetXXvLqlba+GDPqTY9MqIZe
/f+s5joAPG0LrfYlj1r/Z3owLMC/6YAMQZ7ZyBrv/06prbnNMfn1RSkV55vltriZ
FqlDgtcWmtfTlFuFXfuRJIpheXuwAlSwGep87gg0T0IrpF5cl9Fqu9F0VI76FdfA
bQMOVoZjV6pwtI/pN6Mkf1OnI/5YOm9oQGB8Cm9Aap++O4vJNvcXbmnOF4FNLKVl
9GJuTorLpR7leA6xna6n1Fi0GviRPFmW+XSK9kSh9C5gb8nPNkeKowlXt+HOmPE8
4WMAU83VWPRXljOBA5m93J10heQUz6TT2Iy40tehp7vkF5VJdPiygubm+R3wPfgV
//CIpveHXx6nIB9XTeBNDix7gUBRugOFaDexKTAnsnobGvraEnK9Fm1An+RW2PeJ
2gFIJ8hwOYxaxCnHdvhLiEnUQqSsNUjIJHCfCWrRjDZkgzo6+SIJhIDvWX1WLbYH
jnaeRQSEYv4sQL4Dl6zfwnIKyZ4x5e8zveFgjIV1e028lV4d/bsamH2DlSqWSE4e
DOO6uyNsK2tgRzvA/AxaxtQP04DPv1vyFFi4/8NT6E6HpOM/BmXcRP2VYtAhYCyS
EXkHxW+RQ6HojgDuHCU63NmLMVcAcpaJu2FJ5NoZnTXWWYebfgMizwYPRv4GjA7T
u22jCRWVUbKE8NY511B8P1v0DnDEwn26oxq9kIeMazgegmimPo7oJxidRcLhvM7R
hS6DymquNzFuOwq+rJN0pyPL3WJS6Xml9Wqpc39U5x7HBcWBevYJW4xsxFoJ1zvC
yHmvwUVNFD+LLkbH24E4mzRaNsCVgcu2lZgdMC5KHK6SQ/JCMBAmUDxeRL2CSxPb
+mN4IJ7dVx76dQNzsSYTfqDGPRU8MzASdsn4yAemen6es+/2R1V+fGo7zARdEQ0c
3tuKG6vdjQrVzLjmrHywEBOPaYZRA+cPgbgZtUNfIeoNXYbc95/dNMOvDvQfMXq2
mYuMg3mU92vYeEXwIz3Xr6XEdLMA5gBxFdVifS0Q5eoRof2O7uOdNPgwbu9ywHOv
60sHph+odRWQVvjGEB5i1ZSZeLCVjQbLsX/3MLwS94EI3IFn+QcGGcpjJ84e61od
Y4RJxTXp2QTUk56RKmDSUwsy78qAUHko6BGyGQJDS/KJ+34jNFiuH2rQ88oYPJov
ro7/1o0uSDb2wgoz56LRyOwKWhvYZCq6kO4hKrg8eOwZfRPM7OQMm2oKUqnMD0kz
d1hHExJ5wRXN8v+5GNjXGDpPMtdvooIcCivwXrS2o+RSVDg2MWfVGZkd+c10sj+z
D8S9IaohWpn2wZd4ewcm5/QV7DLBtl8ujUJIokjZ02OBUsxWe02MODJx8acqwfce
QT1N/fQttR5bDMkR2uoGU4UwJJn6987WV3Kx4R9Sx1ZfRdxvqz52GvD6wu7W4Xwv
98Ir0Gk0IX5JJLEgJAldGtqF2lfKQY7GFbZCo/Kzhneklhox4OxIlLqwrWOfg3I0
/5MJ79zeheVUMKxjw5ZywxsiOIsnzgcNaRhgG7XCmxegJ57zbPEN42ud7RdB+k44
HGVXcnH5B8KnCmGiNBfzDTlt67GVYAff8TS6cIHSx7FUHBm4ZzNxFTgGjb8ximHG
VxRJzxmTMdsEeneDoV7hgimjgizQLh6GaxgP+AWzfBhiSObOojADk6cgSt+TKmJi
Wzm9k0HoLDjJIbDOXyHHm1zxRq4G8028GKZkde6RUFdytpT6ACvtZDJwxscwygUa
wknz+QApuKKUzbc+OC1he/ayqMfIoVGAvm/I4N9PycsAkyvLXYoFOY/7bIus1ShP
pbJFz9ufxZ4wi5hS3FIoc3mggE1g0aXv0WVIMUTfCQ3rCTAZr4FVPwvB23wG/SRM
atWSvazZ7/gcbA/tpqUyP4TAwCsAshKCZLh4/PSV75WmREtfN4xpE91J1LvrvdWn
QHRiY/2oicjTCDAWkXbP3DSSuwkJx0MucGREc1lYqT3jfBiAKLEC8z4qZhwLBF4F
yQfOl64iewi0InBuo81+sUnB2uYHG1HBFw2CRRCtNFHZGIXODDmM3S2BbKm9Fvpy
G+bHAAuntnPaPPeYr/fPMWjqtrwXaqgTlEs5TZE4dWf0Yumgsggoatmew97N/fo4
paFgfMU0Zt3VspN0LXv7Havls4TTFToH5fI4N5gMu7ah3PWW+7c4AY14KFKMYxcl
3giQkOozvvhZfM50UWN36kfFOhRlcjzLyEh2FGcdjWVzHH2cYEkbAFTgBIPBArfF
5PvrRYp43QRKUETn1k/u7xRBhnyIrWDcpgobHEUtfw3bJnZu1ZVbtskai98RbcYj
i8LQavVQ+NCv/hKAMyS3cIeD0U0pNHUHilhJxZZASJGZEHv0CRXN6K6mpjv7Nn6X
7GpMRSUY8niMA2mtGaFc9UL8xqA/Y1veV14CPefpXEwkrGjM0BE47Aahgldc4Ney
q1tJDDUkhdP0vwJtSGerO0DWcVCNXAFJsruiFHDp3lNpD7vZ7DnCxKjpSHXm/GSz
hbMZujYsAbXsucaP8jrF1lnsPA/TI860t5ex4ws+kf08QI3DcEwmk/1pzJB9F0eG
FilqueTLvQfz38h581nKzPtiCkiNL+rMMvmE26tjdTRk3UcGN9fKzQRH3M7Lo6A0
g3sh9O/o4fnyrLkNax1mHszZNRMgaDtoBaJqOqnlgrnwWQ48Mah1/4yg+xzse6sw
9t2RuoTfPe50H4Fw3sKwed83C+kPb6s7wy0T/+HJSHDm889RombXwsQw9J/pDPJX
zj1c3l6h8LdNf1NUqNMC9mStm35LPuEKpxJbeABbGw9J5qzY6IM7NgnbJrtpeNxD
M0udbW0dzZp6/9sbYSegofEGqwuyCIePVV17A1ONRNWjWGVjAOW2Eru7Rlo1Fheq
EQ5GDLd7YXthqK2qAcrxpXgGbjDLpraKb64+ihDBs6FTFuQhd1AJANEQCUUp/pgC
IWv5PcxSjrsHBVu5sSP4eCv7NAPXQkZp51nORe37QBZV801U8/OJA7V/D1kmkJDN
9Fa4vrLB9R6ZLBxdJrm6yuFrjRSMD18+t6Ho6R4lgr5xotiMvnMMG07nDqXaiYqS
N59qTLAAHLvKmXxfak20vyfy9OWMu7FA98nocOM9RrjGdl0t34VRbQWW7nf1HCHI
ymlGhCmKpWFGL6JSdBCHCyVDjQY5QMSnzRhV2+aLmZRd2YBFAmJXro3LtvyzkED9
b4jNKoZ2b1UPZHdj+4b5E1hFHGgS4c0tBGr7b2mIXN2voqGexFYTRbmaL5AhpbL8
wNhja3RWShPsoApGCRkmz0d6CeLbnEjODR+2NBLvjEZ8UWIxtTymCpKudry1jQqd
0svQy9XyYhp3a12Odebrlw5gy2oGqtfUeSj3Ie0U+ldYwIg/TSXA/pMF7bn+wnTq
HncbEHAdnCr4Mk+B6xlyb2CLqL27cuUYTUGOYi8bxm3qGYp2BjDUdTQmFKn4fBqT
Xn67iLyJIPz8qiJ8JrfYhSl4Tw6PXn94IuVswUFwgv6xGWjC9P5lliHGHGbaE8KN
gQlvK25edyfExOMUL2eYZWFcFC37mL6WEsSv8FF578MgNUMhlDyg3vYcmTmmaaoR
VN2L+npbMYxuGhhCe8UfLfqJUqXzFqvvojn7p/+Kg0fiQzm2ZG/T8IrpHgdulbjj
CAUod7esarqK+UmVJbhyrxEVkbHm2+Rs6/UOaaGpR/PxOf4UfNjkiLCUfDkpAyAN
rLxfHawk5+3PZotjXKHO9aMKJbhCAVlGKC9AOad2w+0x2XZxFlraHdv+B/+nELl5
Yd7/1ZknqGgqrt/b9sNucOjA5SZ4Dl5xCR2xejPa8FeMBjv3knxBQN/Fz9lJApMy
P/e8CS690URWsICcSgFW7d69I+wE37OlA7jX192qyZoS4zzx/DW1xgQflV2tc59/
gYiLTa0wQzeRC/8nqjSMjlGaDsB9UkW/GpyvmPBeD3Cm+0stSa5SfCgiK9nIFnn7
QGnFNqSoD5bFsYhR+mJWCB9sJw4Ir8uqUXXYApBDJLsZbBVtB1Ie0PTT5gZKjiXh
EI30yHGHhGv0h0gaaw5xiGamuplH7tfn/MfC/roXZh713R+K8WwZ/RX+Fpz0QZ+9
+ykg/CrYRFNyOiQ3Gw3brHz2MM2eGwUWJFID8LaR/Mvgk83SNopyyfro7g7zZd2n
A0mHjzW/mUGPhy0negoo/giEzeH5Iz1CQd9eu1jCuKa6d5puwUpJBqAj/J7HwPLb
76qeX0O9jePWPLrpSISpnzo7UAaIxLjwtEockg+UJZ2SLxcPipJ7mfUuI0VGebII
vJ4+Qi/rC9Jug9wO2WN33NDFZkgjfG9oy9XpUGsF3RLgArzt1XEn/2m2CnNpfiNC
WNtx4iHqNgaGaxK6sAp4oCTqqkbqCi/DoaKOQImjNCCDYC96col9xxNdnmaJILvH
ZnK2V0FirVq0K+3BTzokaMAigmJyWv95t9DxR5SN1YwOECCQQ452wP1j05IREBCk
r4Gg7tuky/ny87/00t7InZlQhiagyPXA9ANhiI+CfCHThElIgBYOAgaQ5YKWMLAg
tNTbsfTAfc9xj8p9cEgptRiOZU59+h324siPqAaS0fRKJxt2pwgoKa35pfFzLt/o
WQo0mkLtsUJNrAFklMbm1Vjv03dbEPDi1Pi2Rwdi4f2MP0iXE/DfZjmYLdhrCGe6
Lb7U73NvMZLafKOVW+IBjEGJUb6x8J/zA4+lfH4NLSpFMkw5sw+F+4xJGcQ9Niix
YxGSXI4YWrcMS0kUPRgBNi8V3fGe5vD53tEqzNexEXdGfNTG7FHN3bIwN6wFe5xI
ByA+rmJ3Vrnsknu5NailCo7/UQJ3TyZarkKZGqHvlBIfoCrw1mvS7gvWbKve3OtY
L8JzkM3cUDk5XxnB/bRJESiOj5Eq2+xgGN3EqkbgcPrKzqrlDhwxyYgBsTchs7h3
xFy8jm4SWhN54Zj6TaiQb8F8WudQBhVe7v9Moa1801B/9B7/7N5hBz3tSGPJsGbj
HgOucLyafkHXMexXLgKhlS7uutIi6UkKmijkBHnta54KoXtWDThhs2jiOJS6oeBY
GU+FK4Cjvd00zbhPOMKeihz6rEfKlpDpcHsJpQpUSsF5qpoNbScf1iXOjEFb+/ui
TpXQsoL7MOYFl4uw5Kz/7w0GWJcu4UXbsxc9HpHuCOfHBbhcNFE4nCl/jJx4Xtco
lL+Idjfz5bFdGIV0Um0Enz/yQRJdhYd3t5XO6Hps8CF/S4ttKj01G7ZjuoFSZXGk
3JWAMWMlnP35Hpq7WGlUGhMYgrfiIcdgd28TlBW98w503jrEGI/9F2j2rydrHPND
z0OTP5GFbgLbDC2IJqfgMjX98YHaKaPl6eIebqpZgLp76/gfHWfdbRQgEb6M8bcF
krbauZDDHmuIOMSX4SNmtRK6JkBeOlEONXbQAzYR+uJxSismNxtfd91f5xH+4Rbf
NRKpIM7XLL4T12P6wjB31skmAUlHyeJ+IrQUlgKloi1A/7iUTZinGO37Jla9lFJe
woSOaE25NWzmBNtZ/DrzFMSrL/C0NpmuQMG06j9mEtlMcRSHOykg5QD8hNqTbynq
zC5ezYW/JMWu8nOYQ7rErTTjDNFtixYL2jJ4qeKZXV8hGFTbgmnkVX5NRWpJcj5J
TleTKsrf5xdW12qksyYn/AcBZ76ahW6SnOkM8f7tEwWsRnG+TKXtMolPi9QR5uN4
34wWvLFH1qOFUUDjC9XgGvBP+oZDxqtst2yJ59r0b3wnYvGD+xihD4OpifMPS005
osUW2Mim1je5al+r82+icv7A34WRL4k5KX8T0J8Xp5cxKNpYm43D9hNiAzBCc5WN
tSLpzLW/CuYhP+YCVbEUbFq8FkPXqHZvtuE4sguV9ax2/CsHDpZjwC161gQAI3Zz
8wUNDWo+gG9FU0JmH+GGntzG6UhLBY6muYiPwL3U1NsafQ9ul2Cum2PsO/rxXaHo
HhMtq0VR4AZ2Wp4zUpu3gKODu04nKYc4H8NmB8lgDyk8503SG9Y7KJprUDsoKkik
CIzmklajMBwEdMFuPQx9L75dCefHwYOkMKEh0an7QaKeK61KX87pVNTNLuPqgw7L
osAy/6KJTSCJgHAwyz2o3gzzMloaXfNrh1zwEzdHBG2gOJBbKyp+rjSRopTjRrR8
HSCYDkUErl7Zk6ynnJdbw8JiEqt6deL+OYUFQMUbWERb9UqojFenJw6LVHr8flC+
s3Ml1ARKFCs9jh5c53RFNeoUFRkCqHytUKt+dVZhMX5rtOBV8Y2kOZKnBM3IIIzm
FlApq6qxR3AKcUJfuUfkH+GaVunpI3vTFTuNT/Z6FGePwsmynUl0AVuK0C2PK2Zw
B/M3mwgqc9W6DfozJRd8UQcizE4tVMBdSHZYNwGfpwwBIKTzrbofldvGefp5mvK3
t2FcBiyEkm8wXOpR9LzppNy3hhyXWUKXQjnk6eCulODPs1oxoO9Xos/7GHGT5F4C
rqRZm13jTJrf36RsWWiQBW/wXWdoXhXIYkkHmRynoOU7mCfn7rTGVO0AMZ9wyArT
oXkyImavdD1QK2DGb+01L27xSS+wbR7jAPLvi2Nw5EJsBhiDYVHBtWzLQaOd+qXs
FaZWOb7GHE3/Z2bLLwQhC62KhdhSO8YLuIYHmuFIg7rclukoVWBWiwNvDr+uONp6
AgadQ4NjnoqYUwp5G7x8Wk3uDlEq0QqlaU/yAofXH4v1yN0/ihhNSKxbPxQYTA1K
yGIoNPA2CH6TbVAaRBETwbwiviQvU1qOHakGxn2fX3TL1NIXfDt5lY5OjL0QpveT
VrBOydQYPl+ggAPPCb9n6nR4X+Ern6L0gb/R/r6hQKpgzEhtq8RxG8ndcbLj5sAk
nJwokYK2ji56xhaDYZH5xWvFxC2tT0VSQ1PlF3ef8V9k/QoXcIEv9pSmYRhjNLRq
UJ+g11hpVcrqy/TcdMH8vz2KFi3O4dTWzbNHWx5lN1XLVu5i4Oqo9HqCLYjP0sGz
9oQuIFYVuwHFY1ssSBMNGnN7ee6I74IbwRt11xMbQYeK4fh2wnLB70WJiWTMaj1m
aNE1Qp/+vE2CCTnASkNaqjKHou+5BHIrVIOKE3NG/J2FHxeFqxDO4PVk38mtZt9j
wWQ4cBMDGCZvQMKGy2XKezzCv+16G1mIxghMyLF59P7keHSQx7Z48QealROJCiNR
Wag0InysgRc6jvKeMlNdVGBLYdzKn06TT173h/5pygImn1i71pK8EFqiSXczUrBc
CEvOof3LQIKIu0xxPrwDyyvp2rCBAmEfsINCBqYNUttqBx5SijLYljkFIELIPLba
MhFRCbQiPRVsNwKj4cpeFm2lWfZcySoQEdqAiqwebG59OS7eK/B9CZK8zXyETQwv
wrEcEQCrudRpuNkv1reuc4RQ6jmwXHG2kZPP4kYza+E+Es/HGV7wPbqT/TRsEbiA
+jEtYdEA/bPYZier6VU4BfthnLpvXl7g7uZ7glMFowQ8qLVCF6wHIl/rKhR2mVOw
xMThmohdwy0m2t+STfRa3ln/VFryxoLsBFoyWvrxbfZhMV4L1RbTyAg6V56URyrt
IS5rwu4xKQD7XZoz0unet92kczKTGzmtQgu8AN7TlZEvElv+TlZFk5FJGlukFAEC
AYWyfR2bv5L4rK0fi7cINCDhjYCccc/IOTZ9H6AKaAKKaDWWwpTsSjbJbFtUhaMb
anexR8AnOoyFi9Wcb5fhShJrbZjpRhIYzXr36f4hyMcXeSSFVHoE4DeQibzZxLfP
UhJ95ta4XNrprvsXOtrd+cyB258T69GnNoEnO36GgnJb3SJ5IW63zeRI+GDlgqIJ
TJYjN4IUCOQMKCso+3J1LVcuxGz8bGy498s0nOiF+9VLtPQ1bi+0yNwMoRIHuztM
rtnmh6WoxtHHuVaCvmkYbxgagYS2gk4qKbCr+1bCaulT4vkEX9NpnIytRXwn4kIF
NqBcZbyhuvij0HJixoQNQuglvhpIPl/nOl5DF7i0mJtXejIudlX5SQRV7HXpUxhy
iNBy8YWRBpsg3GN1nAArLioZ7TsumJW5HmTD9QrvpWECunfUS+EwIlnU1PaY9aor
/DJqrKE4X0mw/waa53EWlQxNp8IkaQau11r/hG/ThlHAXnDiEVJRwAruDM3mcwN3
7kq2EnmrB8dHL4/akuoBinG2jib0a7QDp9kobRJ0YNZXY8Zc3vfAtKf/6E53o8LR
och4eWAtXb+S8G8GDXYJ/zJHgb/rbONtz3V/NNDMCL6qtJhObFTuKd1y2pEIdVQb
nX/QZ2XzpQ2JaWx74obGHqLsZsCO47hj0JOV5zq7ZeyTQkD4GWe8eThSMMC8Jh+7
BkiIseEyK7JcGk+bihP7X4XG9qaFkgLPI8Dqn2wXmHMPQbpxwhhuuwFQSQis64im
2XuthoFnf1uBddZTOlLcYHU/8O0HF3VmWGxbnsXfb0IGdpqZ8izAUoGantxjdSLt
E9vxOwkCpb2xPv5MKk8hO5k6lnAfHe17JOhL8342vOEkwLZgsrBWX1ywkj/xbcN0
L3z1kfNJ6N1gprlFSnWmit0wCC1YHYtdh4agbhNc/7GZO6o4/gLq2+gVtARFzjCo
BKcsSvT6JvbopV5sDeHkTZF4CCvNwa6N/50FYUmKAkfVi2v2h4XYc6L1OgQnuLQ9
+ZgTLJj+BTZ62mhR/JipxXvTUGTkQ5RO+z/+9Jtwr3omSYRvvDT0l2sk7d3a5usS
6izpbXKSsl/qZhMZx5GFBMmzd9ZGXRCyPh+d9p4ivk4Q+bovNGDcU3THw1RZREC8
cstKC1+E+5PQ23s8KxprMN3xObMHeAdwy9VOwxX2Gjr1tK/wDV2j61PFr0QBihGx
wNHyyR9Kz5W1/DY0tzj1PiSO6q31Vr+g9skYduLYbQztCjr1eBVpvPzrTQauuvcy
0O4I92XqI8jyBkgOAaw88KR/Y9l8YSzD5jLBYOKshM4N0wa0tmqspmU1wUYKmmIm
LJm/7++JJkLItb5cNhiFwPecud0Fi4rgKCaw4wBzJJ6jLbAMzmHdUJPjmJW1hhwG
XxNYcnihiMgYDY4FMPs1o+yk9Q6F0s03bDDoB7vCujs5O8MRTYV5xtuaqRc2FvlS
xm6bkZ0pbFQYRrfXNN0yK0AwcKiH0elJD0h+6PbJ5Bo81qgyQjnuZ+j5vB8G8cYY
CqIjKr4d6MZvZNPAJzmHb1l6tXBfQmIHrApHbOjLV2hrEwJzE4FKODvcr3YvY4jC
zWWGBKk9s7LWJBJKE5ZKyg595Otytpgp4j0MPO0DpldKsf7RZMSecID9pFFSwQ3b
CNqE40v4m1owQpikrwYn52DmQes2eDAZ21vT9BvMp3Ji/Axbqh4HAW5u+9J8cClv
SSQlQIcq2175lwJZsKdFcHZh8rtr1H5Ihn9XvE4/ZOfpJtHeAclvE9RSklHr7EkE
jDNQf9RngbvFTSV5f3BPviZNQ+lkZUtSnoeq2VIAiZfSvz2hruPb06oO6H7PzdJD
VSFlexrgpMrvJf/pRwCu5V4hkIIDNyCjSqpQlU+b21G9EMtn/K+WBotC43it9g2T
ycCfqNzdZahPjRhRCVF0rue5meOZ5f42JVak8xNh13DVCo1YnwWK63i01Rd6PK1s
KzUQIdwUPEy/rCsqizFggckoybmWTsel2/n6UXwrhU8B1IOW9IevaOSRvzdjixvp
IwaPo7bscy4KQKpZRPAa3JVX1f1e1egpvEz5wms0jWNVgtMrET6g3GQD0g2e5QNJ
yODPER8arCSFaXsRe2C3eiv+FFb9fkcchEwiGfL0GcqLJKLZfuZNnRl64KjnDFid
NhzdbyDo/8BG0MP5MZwzug/g2SYxO8Kx5z4xTxDHdbs/FL6cjpWvm6kLwP0/HuLC
Bqv5fkZN0CoD3qUCQ3+s5zVYtstz9fPT8CZF1MmuQSZzLoMVdP+daoosX/XZSzK0
Z98A6evM8N7/aZ59v5T3cJthoCJHnjWMGkqWwlSlrDMO2P5kHUlcTBMK6dN2zQLs
UdiLXEYgCxIo23UKd3fOUVU3b2ruGkalwk++Cy1m0cUTAUiuGsl39HXAFh7HU76G
9lfStxm6odRm8TR/8FCCSKlnXNi0FdqY7xWM8LdMYsHwTYNtlOsO5le+JJh1qA/P
F71iqqNPNQbxn7G0kOp4M01aBI5Hc70CzONgGqAwnICKY+LwiRtcy/vPBKpcEwce
ezt6VSul8ZQumLrJ4syuXnus7VLqk4yB9CLo9mr4QG3+1vBrm3ZQshTsCbV2bluh
qbogO5Uv+gB1UNWCs/telJO3cwqEYoS0WIhPXDs/smoFxqdO44BnS7P9ob2V7pxd
KLbbsJpDM1BKoZjEqRVH+c9lQQ8j4YWm6TBJOHKopyKX42UNFlgNQoy86opfWDsB
gpaARRkiQQvRJUXLepa57R8XHpNymOU86a6dr+57b3EPc684syOqcaNc8r7farjW
O/LkTBrLtYQ4B6smPBvJuYWQe2CTfmmGLRjGalLCyYkaEZusPuYBLHiAhBXsWEdu
v8uPEqEAjfHI1kA278eefII7yUE1OtWLiVNFt1Nt6+TU3lKGtH/+cDDn/m9qkq/8
SitsLeEvANuu8ttTQ38/BZttsxCMv0JYY9/Q5Z9tiLaBy+nO+3M/xlY1NMX50Xpn
fugrBCu8FpWkUYzBKfc1nmrULmJtwFrNkmEj0eWIw5qRvqgMfEVbEjaww1eS/FIT
KNdNxT3DUbj+YoQetgfPJJvYs7QX9MFsE1upYVFjPG8uQPU23vncNiiiQGvw09PU
S0zHNMI3lLDEqTSqdeenHZLlmTZ1U70PI3Vf5+2FF2jnyzi7VCIaN6GL1zhJg5I7
387Ep8JENBfc0egkQF68FbbOW5Zkt38XBPx+DAV977a054aD2y5YPR1kBMKvAbNr
fzTYH+AIkDN+n0ZBlPxp56p1GEsQbVIpRu0WM38kb6xPRDRiUqQ6fB9dHUXjGPje
xQZ6lsxJ7FAFca0anjiv9Y+eZHH4dB/rq0UIEhOLLSDaLzukE9V8lQ3nD9jNK4cp
6Ogm2IER5GGccSXaaprtTG+bhY1gnI6wG/sBup21fFVxdVy47tNplv/J+xO81lkO
6qtGokjsp/FLCM5fwmbX5xiUjJfSMu04R81Qu0oXkx4dfQYuwPqFI97l0DmRwFMu
wvcPZx+e1lMiskZ1ANpYGTG7MB+saIjgXeCJ9bR7YWyYcfU/MjwWKH0kMrz/HyPW
xwUXjIm2LSst0bdwOopUOPlo1100LdgUXrNMaLp4DliApIj5i7blrKhrQIeRelEC
e/iItsG94bTFc8FB1zbCoo0RaMO+8eq1/p2FgTnXaGCByxSCQ02bLsQRoltNkQg+
pdd6BI7UzmFZX/YT5S/CB9EZfdsIu8MhkMe7kpArx4a8rTDLLG4Hdi7u8sx9+FV0
2sM8gsHKnIgO8Y2t94vuyeLq1tbTLSLrANxDLPxt4mjY9mfkRLP7V7d1Ss/czt93
b/SzWOiztbiwTwp2Jg6mzKYC8rtumFbFqs60AmD840BdK/xaeIWRHzYJrzVuWNM5
d6vtJcn+DXRCSQEGNNVa6dHicmZD6SVOXh1AxWq2I164Nei8hOLp9GiJCHt0MsNX
sD6Y34ibXmnoHqQSc4PtMk7CRebt5vIYY6sH4S/Jbhr5+Jj6m0XaLg5A3GQSSORE
SobfLmeSAdD3c0pf4uSU3A3TUx+rmNAjt8iD/SH2eECYCgzPW/WySw2FVUJZvWGg
GIhgANhAz+f4jVHuyhRYLxnXXB9QLTVPp5CDdZ13WLPsLFZaLcAj7jBs5Fy6mUSd
4AkFAtTfzJuvD5EUoX5ZvhQdxAL9bs+1YQpmdPxf97lpEswRsqDxwBFMUiqJz2UH
jul6+yNYttzWQpRoHHmfMUAcBXkYX4YKlacPCmcW493KKH/xHUOUTYy0kyD6Z1pB
VH+LLGowq8hmj57u05VfXtB7YrVWk2XG17LFBoW73EOGkkpo92PjcDNEZfrCldM+
8qXpVlHH0+MgFg9wf+RNhyzoRODEkDrwhkpzfQfwolsX+BZSaaus8DNRdN+Zhfit
ihD0i0pWiUWgl0jB+Tbh6T1Is7eo0zvaSbvco5DeeWGWWZ0Zf/ADB/k7vnOy/8OT
QjHKwglrSWcVogYz5zXjYFxDuD8fg8mBHdH0S2dP9u6IpC8drao9dNfFKw6k3Oub
w3LtGj0jijhQhW3yc7rDMogv0bCrq9f2y19/0CixUnEK4i9tEq4f/WlhO28IuXuy
9yCdkALrVxOuuzYqZ9dQplYVbw4IogxlHdnwyEkH7ErygPDXL290AT1oJqq4Fnqa
fPbPSz5Cke4y7v+WneiuXGKYraL3er3TfmBwnjjQgCHSKZvTWIyJzD8GFpRLVRXn
RvytOIKE//VtW3DzgIVfg7oHBU9B/edQSJPcfKrU6WklyZU3A/Fokfv5ROJduovW
LHu/Vus/7+0lM7vvXZXF+1dTlguMa2JFw47IUrLsnqR+odWSHz09xgTgaDP8uRyU
wmbcD6s/vAURJFC1qoerDyP81rSeaVwwaZpkjsnx4THKb+RiHWXn5hL0pt1kDwVG
fi1kIeXlDySuZczRYa6Hm0XIsnSCsT2XOgX+IgcXA/j911Q53fPg9i45OVo+lSWF
KfHWAYH1Mpsc747Mp8+7kJ6/Ql/Am514VxXiqXTzXVTF/wPVmWm/OCNi0ujw3utZ
CMISTaY88MSUkjO+WediJuxshQiGvP+3pWnmefH0o3bgWY9q5SVC/K7MHnMF4xRS
XFQhup0ehMmBsQeMRSxeuL8RRADVnHlKSsPnSRM7+dkbdpuwgToCFbl8wpkumxzP
0pdYNTzkcfT+ZDohar193v43vNr9FdsS99egF3Pau5Jy0IOotNGNnyScMbUPzldM
m0+xM+B/OZHK4165GN0wn5PQXuf9XFciuwwFtiXllQxacWLMPMwYbJ3leVSWANQ5
9zCMwUDFu7qpP/6Hs/tKsnoHqQ4uETrY1qZlT6Pam0VUIDdV0EAZDrHWipf5b7zn
zWKSffQZHZHm2O9eB8aimknXljAjx1C6fN09f6JH+DTEK5wMlbsq3482KXwKcaB9
Hc+IzFbF++qvs20F6ppS/+/Ggy8tbXEOp/5G377Qg0L/Hv9Lr+NyzAs/S3dfxELy
XYCA+1SnHGSkHSpru78YHQihoC7WNAXKC7KGvc3l/8WveHPs2lrVqB9dArwcS8ck
33F4HT7UJFZ6oroCKJsVzfU2ETaJbY+3hkTxF7MDWfyqhG1CzLAS9Vq2+4lps2qV
mFPLajWXS/LD5zgawJs54ET0Y+14owT5rIMaOwbCvDOtt692cCcqa0ldQQvZuG8O
PUJNOE8am3Pnm9CXQC47/ey9j/HW6QNsIrZdFeaYrXNlaS9rscVBVI/4/Gif93tH
1ivZrKejkTUBU+1Mv4GWp7RGCdenHsLP2hYsr9s0P1/+VHYvLCHZX5rX2Jikssi+
tTHBxGccRoVT0z8fmf17feX2lMtjgTbHQCCjYfV/1IsC4ETiU9G94KEr7aQdTSZU
Rjw5tzNXzhS0tnrYEwg7P+FBp3rDKaNFbxx3l1gB7LmSrwCZ6zDQIX6vkmfsWwBG
nxfZk3I51szG0Hac8A9CkD2vX+M+FxBeb44fVfLYiu5prpQiHbcgA7sUzdng1OdY
3qRH3k8XGmhTTGbJFkhCH2av4n8B3vnP1iui/oLYMdMnFUZQhPCI0qCuZxnkg8LN
hw+NqOduf70yzqmRTqtEfAON1+RTKVMjXYtEY9s85qYJ74aPyUfsLGB72eIO1sNy
lxxmdPo1jAc/tjMMdH5L0iDRPiTRCozd5oORzHm4t/A+F2S5Sjpbwb8svHyY0hLZ
GdXKRckvIGgxv9zKCZ3By+kiEUEPCWi0NG5Rx6xgGdpSVMzF+rataiypTAx2lbWS
zyKYNNqU/9hdsbY7eOde2JHSIwQYY/Ah865ObVSzC9PKkvmaik8J0Y78Y50ct4Y4
asR9A2JHh+otthhiymu6k3o88zmbqipoZtiumJ7UFldsqi0uiJsDR9Lm5VrKCQKV
G30aM4LKqPfA8iswZLYvAcggJo0sKecjLteyI7CQnEOR6NIjwtzf4F74GgTaJ0F+
c+OMhYwDAT8nxDYp1yXI3mu7NEPpWRpsk1dMBgd3mG+OW3iwyeraO9p9B//dyxvM
PkjOEwrp1WGhHF+aW39lQieCnYXOEw43BsgM0Rpn37Dnm+2jOnLm3hmLJ5Ht52+Z
sdksNuJ9Oxg2GKzhunMkfvN6GlQuTjPwKz935zlSEcuteylTFka9WAt/l8Z0l1al
L5baUfuQVl2B8HoXhfy6hGnjKwoV5vTIncVhZEaMjakUr8v5cbolhxlHnW3A+VXY
d2ewHW6+HTM3/VX1i1MKENmPG/spyk9LxivCKDW66+V5sDVh7Q6DsMFIQDoBlrpm
h13ESb6tRvKqEyMJdHd0M1cLc92e4YdsfA511DY5zEKyyZb+KSEV+rBZu1amD0Uq
DoeicbFtVPwaC8nt3QMLHoOruNEci38EUJ+x441ulOaEwuZofdapQKXNLzoNSmc+
hqQdcVejb/UqgVJOPDbZL/AeVIeACnIaT6YljpnqjmebhP4o3z1aN2HPu9cXQliL
ImiAXjwJ08KaPm04DQtk9LBv2tHxTVUspwVt3QrV+zKqtq++0n6KLWPgjvufj1bi
BjDtzh4PuV4aGQ0g/EdOuyBHoLOMtXPOzXQqeHsV5SUUOLPS6TZ23ZFvJc7X+kXf
0tFX4PTjNX+rsBMTECNlMPEKd0rG38L+oicof+P5TCZL1NISRefvuC7bh5Q0V8AM
kpIj78oW3Vo2lsAkgaR5bxUI62bVPHPYaLnaAqddrJJxsF30CUKr3Yn2/cCc2+Ln
hDQcQDaUGMBt5fQDgPsJoPgh2qYQbqexXrEV89s/xFZ5gw1CmGE/iViGduzH7coz
DE5uOaeiTQi5QqgS0UcAa0jpn0o3zYP2whPlB9udFWJ/pK6Z0KTJtuPBPf/R5hvY
xGIB05TaKyk4adYoq6CGhgHS/gAmlEzsFl0xP0tM8L9ThYM4Kf8iCFH00FP+5ZJ8
jCc2x/cCQTdZu2L9RgPWrLavRTNA3GSuT2Ap9vDZxPhmU2xosk9zY1WQIUKKrXbl
SDNBg9Wr2YU+dyaadDSa073cbk27yS7jd/iluk2GQYcaOzQWlLWGGb+PzBXu/Zqq
4NLl3X4XIZklgO2vCxwwOm62erEsr8OuB+PeuFzAHqKG3zhmdQ0P/yRtxi+VzEi6
nUmJDiHheudKnQi9vhl4Qi4WDRH/5B3+jox1fkK9PEhvSmw7XToJmaU3xHwTCjPf
4Mr06XqmAU1Tr1njfeCEC/HiCm2lDQa+cg2j+Xh+wKUsYb4KEOz8RPfKBrajPieu
vegh1eU7LZiPHcisXw57Nkep7Shp1ZoZD75IQwTQAiiz/mFdYKesWmiriDfq9ObJ
76CkEuQmg2NpF4hKKqK45MrBD5GRjnwauRfVtOBWjB1cfWFCxhvx7/apDVTDfi3H
BiBmZebeNb+CM1FfrTukBlOEfckS3RnzcbdHsWq2P4uQ20YCO4p1vpwoQU5YHM+i
gnpUbH/xSlvGX8Wc+VeVHjE1yyuBhosgZhLefutoOjiympXNEPozbfjqd1PpsXCt
H2Wc1Yigl6DjThM7OabFcEEkksBHONVYYdonr/XIuNnBecwO93ydM9WUhQEwb5+k
wXd41eIdUrmA/1FVlQ98twX1hHxudtHjxcvNMyxLSz+cJBsNoujWMSdOmXZvCsmd
c/V+2ZJcJacWLSErmm8v/OCXTBa7SubakE/WqrQdfzXRFHVNqmZW4G1W7gErI9wP
hR8yRxUvVzn+ehjW1mP4QYC3ZdFytKxdQGWaTdOMkeqRg29Bf0XttrrhxFh/psRr
ADBeguSlAePt5Cn5y7qB/LHjC4SrX3ikGjDdwi0P+AdGoCQSxGFaBlY2735oCM38
coxSjHNVTuYuoZ6sJP1M9FUH8j/o3W5ITqsilKOFmPIyyLLtE17t3nQiPZhcK0Ki
LNx0v89b8q60EesyPzn2VsssPcnXMdN5rfnLmJU6WZ9W98tYe7pavb8ihk305Tlx
agwwxUsGUtcoSMJYTZNaS1yu1fgZMXpJ8J7zjPTYTlFfGtr+8cTVmrcrCCYiTb8o
9jabcImA++LjrC9EgH/X3seA3x4y4B+XFU2RGt7r//gjHsn9GlPH3dfSuqi7Y30j
vONT2us7q0INRovMFEJXgjxmIamrrdtxv0mIDUqNO8QVjFUak0buoGQuWJBd7l5C
3Vbvh629ZM+UaCIW2EPnv02aOiT5OWgV3AERrxO9wkxzibumpI5GGwhLEP+UjoPw
2uRmSOn7tPgD0FolR6vT4a8SkuPaaFkciv7nkM1dOvpN8Q0Wce0FVW0vvFtn8qL9
IquM6uFkPfBwCLNve2ZONjd/NcCWKCVZ5gGgV5IBGHEC8wJWEUxKXghJrP40BOOk
28gEDD8LN2gvbV69j/IYIfdNG6/myS+kd8ly6I6fOD+TRpV3OA9LvJ1pWA4tvcia
BgL3IL8/TjJy23mri1q1d3DCzKKzVkukZL0l5t6uFcdpPvdqiFndOawSCvGHxjX9
bGiFm9AiG360rZH+UjmP8S9PtXhoFtHw00hIr2tUX4jQAfX2U8zyKf29ISotgUjM
Br1cMGz4fKugzYXXHQcChfbPdE1IemsxX40x35Sm8fTIDUvU+layYBC8JE7vnCFl
Ws1EgzH47aw+pUZMG90KrmNvMRhXU3hKyrhHSClid0E7harYSQOKMMK0Znp+y3t6
q9eovfMpRbMO/ckLmO+oqq9R+/jzleys5Zun9Cqm9d2GDqV7rMfTNerMX5I6fA4L
0a4tyxTSiuhRpOlhytBmA38YHRGDiVLLR/Gb9hJK94wHVZAqfUT6WESAuWu/i0G8
rupJWfN/vL5KoRND0DuKKjtzqUYl0L221/4mF9gaom7LSke1jZFgHhV6FAbV5nJY
x8w18kZoxD6nYwExtKVKbW9tjOizjq1TTDda2xEhidQP+e1ewU3ofTeF2lc/QzqI
dCJhYj9V1vT1mAi6h0IPfLVACnz6WdIEedEMqGfOxREMc58iAXaTnZYH3woZiY8I
H9186WsEbvAHF58wPhFAKgvvCJTZv/POzdxiDhjd05Dfn3+TuyOsmwpMnqcPLmRg
qsjAMSrWetFuyZtCsP+a7qVsxUIlLACrrhOIAaKCptk6f3AQXhXVrMp2JHSiZXGo
cPQOUV1ckxjfUuS6kmKqqoLpunBPUQPbCoxbDVJpWw+sy5+BLnh8KF+W8TXk6Rv8
cbINLhrRagcJWNPICIiA++EZQh+dq04W3IzM+vWw3PcDpvHx+k6sJCUQo8tcaFNX
DcxBEjuiWOyslASZaOs5CcS9EQSLKbYKrPhw1vc+wRNxTzXALv7TIy7/kYUq+Vlv
iUmIVmE7OoNYSUO0Ojc8eXbFsPMBdGNvuzMJOl5CLiU0u+tM2CwXRTzWEAKiBvlT
aMERHEUY1p/q9hSAywsvw77hrgdptIVrf3hsXPwT0h5YW1C5wubc76e4YV22VS6V
lHihPCBQTIA2yljKZjn4JID+8UX3hHfi2M9DZJrri3jQVm/uFQBeNA4zf0y9W9TC
Re4TK2a1FYxFPmAlS0estyBZ+5yOiSoFm9GrwadsFhLFF4l+rD3y6JUiD+aFlt4/
kIx3cuXZNWh5k3KmvowVMi7wUh25lT5l2Xd2mv/M02VtyM11lEbnfnImjoPAKOKc
b6j9jeG36P4hZAqATowAmUE9q1qOUJLUdoJLO5VoiPyth88AF+DAWbEw60mDaC8I
Wla4Jc2b3YSRDZVg+A/CWSvCOmbWuy8XRenDq579AtIyBnuQAVM+43dA+Wr/CDKT
8SFk4qIz00mHpx0geuieB4zGCyjxcvw9medWvXFgKI0ivSqHlBvB//y9NGEqXAVb
nuyj/AB8kdJZDv4wu/Iotff8ZXmnPC5A2g6Em5qNcEwQQEQzUk8v3UXB6ArgNNgV
hlvctpj56GnWcgYT653TLrmEC25e7/soP34RNggZ4qdRuNEldLhZwcvYqj1FwyeU
0ENcKz8M1JAnD38OaSrkW+KSRYFhbnWzZM6NJiFZsbb8w/aZJH92tnzdOh7cm0db
F/LdDfQAUoft3Wl/WJVOQbyQTOVbOmNoMiV0kAuyuA0OwO1C8fzaAMTfTf9XKQGF
lht7pex8mY+Rw29NJ3UT5GgY1K/ge0UFeQKmjuGZ6tOkGvA5BGno9l2LVTvevVAI
Xr6lcByKIthlAEcZ7y+1SjC2QG8j95JWrzo9frY6ArptRbRb2gmj+Mf6qIFvIqB1
FTmrSo3vrw45ATCsuubp8UYVeHotje9OSuha5Z4i9lCg/q65Vur4izaCsa4vdta1
K3f8hMT+Z4bAAiUc1cZakux5U53YkGUDPV2aLXzuRVjnNJgVRLJSqRTdB8p08/Jt
jUlWk+bgqfQPHmm0F/NgoZwrTFIUfmb7SnMcLnzTC/VQq1hKBUaRiVg4FSyDhwXN
AG3SC/mhHb5qyf44DzLM0N59F4lVloKDNICplB8MaH5tV07SrJMu4oZSyqe0RY6K
QLn//GImLJXzRQSGgxq15RdHyb2JBiybBxZbzv+h7i+mVCtMwVPqETN6bAx3IS4p
62dSIqFLITPibBi49L+46e4LnZzzT8dJyrt9+0QLeOjJUfklBZ7YoJ0XZsNluR5r
erpI/Ue8wvhjcr9fiLMz3Ru7JK0Knr3CbdOmgosemR92VXDXtMYILDdx+dgdel75
RnmjlPl2pqSG4uUlHwnv4CX98/r6XTFPVT6kZSAHOk9X66eEba4HDVTJxkr/gSjr
LinLyObyCAi1sk/BgP66UsayZf4zVNAlyIdUkyb/wBuTt/B7OELANoOe51I+LMuL
o58Cj0DhMZ8i/rn/b0aOZTHYkBGwYw+COwxTPuiDaxLhdq3QNNk65gVVtZYkrSd2
hFK+54QiyMDY1kz48K0b/BxkHj62vOeWaT1Yx0DkG5bksNU5cY4l494GDR4UQjp4
g98eclDXbGDzrm4SF0a5R4D/u4S3Ciy4AY13xaj1UK0bLdWOuScP9g+WglNK+lEm
6THYTUc1UUFHnkf9Wqh+JuXtl0amGspRL806l5IwGb6mjnRq3U5yOMIivykikn1G
mRtZdK4sK0+anVY2vfVQPFsfM8kS/HXSOay67aY8CT6ZHalDvV44K+225Fa46dgq
B+rbe1ENNjbQDz0cQWf5idyPQRpNmaKou71W6SN4jEXgCbJCNcQxPs+qxIs3tuW7
cB5wNkw6W9eQp3LkjQ17ftYg/LWyk8uH4vqYm77TWwf5NW1UMozjqD/Sq27m9hWe
o1a22ZU1jXfHn6NWxhztjKVz5kQ7hJ7slyYAXhe5ZV6NGKQ4ufV8KZ7l742EpgLd
E7C2Pm6fLhbrx1nHZoiJLu1UndEdNxiUDeDS0a2xU/lM+5571Dh/RqNkCnjEefKn
lujj5fc26oRt9ug+a5+gpF3Hpmis1UXazn25rNvUU3lR2VLWA35loL4uOOxsIwi/
tt2+e9z3uE1BzYw7Fd8nXBOtQt1zaFYibxYTHWn/Z64c1j+21KJ4BIjIKx8pXsGx
zX0hLKk3Zz0Uf4DPEvPU1+gKxvRddXtjVydqjFtdYMxpw1agMi1UT5d4kJP7F5lt
ApB6ZLCM/afuIItVOx3Mz5k1GzU9caEWxPGzXj1GTDJC+cQ2NHfFQMoCWBjZHx7R
4GKkUBwi7QPjrkkL3Uo2z++MsR0rEXDruCirvpt5ef9+4q0f7AMUDFEPpmnOP1y+
h/RY9o2GaWsb4UnHkBQke3PJ5H+xnuDu3SbQMB1YId/ohnksG+/4CKT4H9nAFI03
ZfpPmDldoJf4bDsiZetlvencEMSGAo32avYd0iZ22aEXxO9uJQHySdki8xMpwZU7
s2bt36jt7k/RgyasBOv8X9yLIeg0Xd1VHiqxFP5fngZLunf0HkKwmNeTO0C7P+D6
xRVezAgUa4oiNA/4uXHQLjiVculZ0ybe7cKWJCgeGOeYRo272a4729EMUobpcdkC
rDxB1UTG51DaxkMmxYvU6oKXA+XTrW/xK0wI6wBUyHSN+sXOgYVK3LYHrojQtu/J
3tmhlxYeGGbSOK4uvlEsOP1Y5wjx8CKY5owSJXpL8cxjJ1j4DvYlLjsG8DPpsxsu
HZuCpukefvVonyO3dm8g2d30FeIh/G8+r1MHIefFZmoVeumPuIPE5bEkSMHM5clD
e4AKSKoj13MonOqeMSWl3+rgJTnzbD7BAAB7n4kLQE++4+n9RmtQi13szX8rRkxJ
faNV6xf0QuYU0chKEyZBKMk3KwgGO1bc+CPk9Qfpq6Gb/1uxu5Q5eu+KgZUqNtiB
Vlx1MHKoYbUqXuKK+MBh9pm2zeLfZbH7uyEAZNoPNN6QTsGhTngCOFJHWL0s0GJC
JlSFzHZoyr/6ICaYBBizApQULBGIeVjtvJuaJOE4MFnVtgNAbhSBhWCqzDwnlfR5
JLlWpRUtPCuRogPgdGPLQSarFiTx3DC3LZo8e0bKkwltEavQrSehWpBcojTGh8sR
NP3MxKlj+Ky5cEnVO+cY2A/8XODimlILKM0cUdUt/chjb+nrLTdSWvwng2Qwqscc
tKwzos8ZksESEkEWD8TUZ6qav0w3qWscW0jUnksanPc1/hXsJFZElKrB86Gup+4N
ey/hv1noiDSjCtsdxCUkC3vZb9KcosIXEyvabX2QQnWMxeUE1sgLYW49YHt6saHY
n1NFerl2sKtZ1FWoKeTFBDxBpB9o2O1vWy4w07BVQS0U/Hs1Rhsgz5zVmw8vceoa
3Fmh/9VnvbTYN91oIpycEZQo7Yw+Rz/RPABoYKr1IQuNeJSoifFX/xSgGgjlRQVT
bZrL/ePxbmiEtt4nulr5dwEcF0ioCULXq+Wg5x78dDfn+SC6lZWddGqncVdwzUCn
7z9pqZV02Y6uTSzhMNTq96+vxDRc2LUNJmnMxsNEoWWoaCNl3dfuYXxASdzujhs+
qEWfzWxHbsp053I1FDN3v87i60VtMNu8Udh+lriWEq7gQuCJZjGFCP+AgmW9ytew
onP/1bPdJEOXI+tVdV/0BRZ7F6UT6/djiOuVhnUZiT++VmfhEdcNWsw41EFv3dxH
x6uccnc0Gs9cXShiZQhdGVFMaw9Y9PxtmajcUzsAUXfmIa2ockuNXm9m+aef5irW
NREI1EG/WB9CfHFQcIlqdjFbzCaWDomHWTOTW7XSRJ4w/FyRzuijgQ1DyvOCdI4R
v6UzXb/mmXi8BvXH7nCS5wvxgYZi9VqP5om40iztQTZtpu04ANrIFEutHFMp8Cq7
mqriXaSRs/zWS7mz+ZbJJ4LldmD9YH11n/XOXMt/bqUKC05X6NO5F9YW+8oWK1Kg
U7eX6ReSJ7y31KyFy1q/Jn/Y4HFynnj5BNlL3N4F8MQ6RvTwT/pGOegyYZ23mq0Q
ywW5KEEl9JK603J3KHZyW4g5iOBwaKbPZEfJyrDSTS5yISiYLprvr/pEG3imqTNv
98WMi8frPIZp9tQL3lopVJ5cGg88ifwP+yzCQo26yZayuiip2OcU4OiLc/FYCEQG
hz4rudgHykxLikdUWArCDZ8F9F3CQuVE5SkHepyaxBWLfI/GpD/7VLxqHSK55VcL
pZtZMNUaiyakRaDNa5C9fcErqZ5KJPmRo76A1GjWm1DcuYLps86kf5uXdR5KNb3S
Eh/s9WlcGOvy6qv8grOlvhRYAaIzXtEuay+vd+OE5BfZDdWOKJwTDhM7bf7aWo/7
XQaHg+lS24Cx1g0e3z7N2x7PyMOEta9WAEewQA+WQrV6fVu9zq6aZlgLsPAROTcY
EWu7/jumxUiGxK5OP0LIFNBC/f4BhZzitt1k9qh0a+NisBhAxnZUap0wnnm/6Iej
Yoh7/DWabVMBQJnNjWk8g+KAfLO/XqaXo9qL4Wa1X5cW5BZMDAUJ6t8KuRQww5+J
fEqvFB2xELt1sQe+yO4zB0UGw0FkSok9FYrZmVkAel99TMLY4Bg5TUgC9R5/9zBn
AW2Hw4F+ISvtGigyDZhoDBHLKo1SCH5LG00Z+TDvujugtCDcq3UKzSvPu/6rYUnI
e9D2/6dl5Idhgr471yPTN+WL5gXKRLlSRsgjRGBIfthWXLO9PmbMiukiJRzUrsbR
PZ9KJHIPF1r1+0s+b+1Iu6b9ISrZ3pbdTPIG6oCzFbb8cF76LafuOADJQa8KfumV
2iJ/+g8pGVbzrtlJcPIW5VXXIU0/oqW6+EM5E3z/tDUudBxcA81rcT862lLUtzUV
Fsbr3LRyBgBODrv0DuVFZDauwWmB7mCNYDIS9AAVq5K8dOoz2Ve41kPjaCt267HW
1lOTnLCnoA4hsFnB0+yIi9e2Qm2ruL3y/1wHhOcIBLVlscokqQAEqqH7f50Pce9O
whL6ShQVVX41PL3KosBErjfHyvw2FlHmtU9xSuU0eDp0JWcIcWgiuEoM+I0TCBD3
PFkeSm2zwzdnlQRRP2hWhPJuWbZpA0jfuTLEHbLTePZAKTMo/ANI27hwznS9COHo
ISqp/i6ZX62kOUDuJtrcUti5R/pYrsYH9V449neWAouL4rjV7v4ztHTAuyfYX7jl
R+Gh7nERYRJVRVuUs4N3KgAskGNc9AaAvO1rw5HJD6NcoS+BGyUPXPERkpYuhEwr
HyS3u4PeGqGJ0ta/o4+sGN0ya0gf0HmVxVHuHvQH7LyP1xR8xPDy0oCwE5Djs9av
CmgV1s4s6ImJ0X+lxPtJdiwSkHSHNK/KBPdXLKvao+Fb58/q1cywY89NGA3KvRYd
kTdNa8XfMpwDqaaFjrHy4BwsNSjcNTwySOt438KnYRUvcqmOgnoIxdIUKyN3YqUu
fSTQWGm0MRXFEvZIOyvRtePhus4/1rfTGUBnxU+YfMATrvdN9sq4WbuhJ0KNkcqg
fwS0Q4GRuL4YVAFKq+YzWFKxOhsBO9fy6vKc9XT4DXz5r16zxR/nmkVv9vGB+93z
nFpIOoC41V3iA9hKU9AKbbFWnG6nGGbn2m0+BXlR++y7scSqGl67iMCAo6C6j4At
IZYHfSrDr3JErdNFbuwR1+QeefMTyHhy4gkIpuj28nRbejbWWjglgiwa6Y4C17WO
0DZa7bLll2q9bJpLJ9VG9AVXiCmIZ0R7wKL2CM/+vBn3qgEyJkbvhriXTydKEXf3
gNs0+KolBoWemevSUddS0pPVwn5etziYqf9TiDzbmayh0fXkhQy5204pg4V/6DPD
5lLKcMT+pvbth7Vw9KDCm8Q3o+QcE2ZszuVLOHFvT0IrZ8+elU6PpuobhI9E3IpO
ZgtEM5nSXYr6/by5v9FJRnHw+iB0GRdA1lqgxA5PTTZf+JzWurdgbBljmwnLy9rg
RVOLHhkFM0ZVuMkTBhnkcx1tMbnMtPjx9MUyac0Oof9gYXoeyWvGBU8/TlrV/Gy7
TqU9zMZNnfO61H/cDeCFAROtk6ARKOO7JOLCRoXr4gDaOoycH6FtPQr/1gsNpE5J
qIKSW/AU0xypc4D9ypAvz1T3/1iT5j4dlzoI23ldwLjH/ATL+JhB9HtUTDmkmdd9
zSRhM4eZn1R6GEeDYXDwkobh1jBoQiPUFh7Ej52uuW5MxvhKHV+FuUdsV+hi9LYF
Lh8s5QUdPF7VxrvDJogyUPbMQwc+k7jT0JcsyGrh/bOlrRpNFo/B2l+WV+gsIkZ8
vgSnA6zpiynI/kTv1boW0/lA5zGjOG6V/43uaitqBJ/4+YekS4dB6jhmNSFpsQ0Q
YsdZGGpQ/3kKj8bteCFALFGfD5HBh0oq9DfGadQvngdVemBLtXToY3ij029WuDAU
QomeKvlvELBbGSVRfP9XPAYEwHX2ZXO7MDTrWV2qNgpb3OsrS3rs8i0i259Nplg9
lZaPoqDmxRgimGIViLRP0M1ii16Cctdl/NzFMpURc8NwGSX0TJN4TeU/gTRUv3RQ
p3fnk594lxoRYlPMLEu4qeeenHBwiO+FUzT6b5W08a7kLXbsDeva5uDy8BKxmkzq
nXBtkQZHcxDYc7Lop2VQtV7vXOEGNMzLrhIZaavFeUBa3fb+fioAKTC5PYgMe1Xr
BQwcLULTqtPphxRgQahUhSCCiInCQK/lUJIkIAmiJp84oq4wJzX+HwyZdRbJV6Na
zYc29Ca583xqqMs4amfnO48EZMdtWYzy4y4A0a5HDZLL1IVPOX+7ZLIUuh4rY5P3
jEwiOkVrr2Bmai13rWwjmu9cOIDrulb+AEMlhj+G3S/ib3UlMt8So4HEZWnGp7qG
oE/ZG+MICjRaP40pjVqohF48FXDBv5TwgI4t6qg4g7Wec9/X/j+2I3Yr3zhqvECK
pWHy8zzM7yB2JpOTzmc2rHbHxBJumBJgin7Jz+XtAmzGB1wfoBluPOwb5VJDBeBv
tZHuBziUatyrraFMrUKSeGh5tU8VuNaGhTt/U4RB9Uqchhca4KgOV/sun/OvVadl
qKAJNN5U/PyXO0D624+lYg/I+wArtVSKe2EkyEy1xnl5Lm9lDe1FDAX9bl9X+Jqf
ea2KLVd56IUiDxKhU1zP/lr/3L9lw2pDkl+3ucSaJdUPv6Eav2n08mYTlo7JpwI0
PGa4XnOyGX1ro50DjbEzcT8bySRgCCu4ljDr1xic18RN5NiVXZ5gtDvH68tjg25M
oiidVRTk6E3WES+UWIWHMXq4YU+khj4bhdV22TUtudKyzc5KwhjasTH6Ph2TJ0SV
6t1rCG/PoaaB0TxKXYJbv0f7oBD7t5Ry2JHwSHD65vL24mEx2mXZpaYq2WW9jpgF
Ew5uQ2JK2EQ6y12czuykRmyxWu/3r3JxRPbLNrPM83h+jwJWUBs1pl8ZzeVlwHaf
scML85puiReGwhrn/KRvNmNl5LWucqamxERcKwFtmGG6xwRIeel0Y9tsFbgm9vHH
AnjUy32uFjhqxiCLe54m8GD0j8Jgqg2FsQRx+4aYJ13yjW316yQCjS+MoW8QFbkh
kxzoGyecryJoWfA5Ys9KPOfs1dcqSJRmFdanatbtapvw3vzB3PyXu1u9XTmc+7Fv
wQEP5WskWNW6ZYG7V6vp8XMret906JFIIlPbMk2on4CKj7PPtokkCujU6wpYpm2G
43L4TeOQVhcom2HvKvapiH/Ra/QKerV8qiVptyj95SVNY7M/v9/CnE8lhhfoLth1
GRy8G/jTPKi/tJD/IRWDlJEWyYA2QXP4Or3sjHyHrMa4KQ8NLXSLSKPsDAQoAyFI
3lCXuUYufU5PjD3BFkgpQsEMy3QZXzwugrlHVzLssTH8Vol666bDROVqRMTDQsKv
fSvkU5K5C95Olvba68+lcqShNwOtp9Mkx/DUO1n2ckZK9Pz9tC7jqBIIN4n4MiaO
IJW0EtVRsxildW6PjGQDHZXIW8jx1J4yABiXTJ8/D8n10oU2wj0XmBSDKomZUcnm
7ZXSLtiOOeXUzLgX86An58TQZ5lPf60NafifXLbJSI/HnKl92d/0JJGmhBc4QSVE
InuE7uLPKVBs8oY1MfEajfbu5UF0a5Y1Sl5GgG2J3cbYs09Bheys3zMMPwZOEiI6
JTj6+QQUlV3BK3BnEWI6UMUS/4IwTwEcFMMq9koEtNFskhwrolPHNeorjCiLLd4h
1cAga8d2NNmVj0zSP5U7rzpK/maq2ELFpoQKtQ9Q05r3m9tq9o+vFfxyA75SCGUG
kFZf2rFNr9PKK5KplWFR025fBhy3rgse0s/qM6c32+aVJbjiS3QrjjAsp4uNGEnO
9lmcqThEK68S61b/xwTePLqmssrpQScEkxjcDI2jlwfhFuUQ7JnED1mJf+l6DNSG
+XY2pu3amvAhz8NbBvaVKdweZjEWsFKdnEXWBp8AwkrIqXnplZ0ZolirfE0zvBWU
4ZsNYNZqNAOn7aIF2IGkrHOgebufRNJ6xop41J49GuUNhI+o+QMurPNRNWl9VcSb
s6OMDchG03XovordxEbiWKBvzXtxWp9PfsUfL/lV5sB2dFzA760mxZN62HsPsl2F
PnqGTUCK31i/7IogoaYOQaCgkwacIejyV/KUh9AwQ/wBAZ/FJ3Z4nx21RTfknAc6
WHD44ew2suME+WF8MUbMYydDGqHBUsWAU+l02nZxUnmqMYAHSaA2qtq4TQ+2OLGf
raDj82ATByGLe5sNju02k2ccr/gsrHssBhKniu69vWDKRlJxp2VxfvbB5j1QC4F5
P1Y7Qi5enFMmuw7WFUKNEAXuPDr1PisMzALyLBktmqP4z/qN4smzGp1fgmnDmpC+
oQux7aNB1wWIHnCKhyqfmPooBLrpUvhdvH+a/E7m+WCnpuV2+V3JStqkQ77W6yjT
xYnw7BJSfSG06RV8t8K+0wmJ4f1Dbh0DJYAnjvO0KRDlXOVJ7SWvHFPsGpqowo/S
p7L5mypJfefpfucSn+3/URiBaQUXYTqYA0IwvWm0ogdndpnoK3xH4eCcalhiNSDm
XMvpEctBIK133fTLoL09a51IB6bDO8rVKKIbSROLOnSbGxBmdR/a+PnZaCCzlHr+
ZUZVCBpphJqX8QKlA/75ZbSQT0lk52CNZ/7g2mDIQaXVDEcxsrhSB8BFo4/Tt+DL
5QjRbvJKsk+ULSyBd/SKfTso3j2STlzMAWBnMoM3xyHqvzmDkTiDEVVvhi0VCpBp
PbqLD6ZcnbFnDCwitaSAuHSRuW0HvaRkTVvbShKiZs1mhECObQWEXFgABLbYKqER
0ekUWjCNiHkAqpZzUkFuYMvB9iyZdFlIxkcR/xn73c6/KE4LF4pB9/qKah6UKqDr
00dU4e2RBscaD369tV1J8Rjds2TEq3nDKpM4sdTXbN6b7S2eWi5J3bMrtaPOe16K
HLteD1ScXWOy7TxzT2++EJn4tDA0AEvKGZwNCjUKO8FZltC3WEi78lZsYKTVowF4
UCGGMZJfb2t4updAxpS4OsAsJWLcaDaUGcqJcCStGcZIkv82W4L1ptimobt7+LTc
PjhTFv/bMXMrVORMRRxlP5rENlM8K/qP8+03ypQ1oojasRYckxyURDUuub0yMC2Z
/xZWyvtVMSFiqQXedmnnLFGp3jfySvah5OtH6HfoNzrnVNdbS1RdoYKolXsghkRB
wCogu1HQyl/cpt+/3sonnnNHbFOil9PcuEPGcpZ5I++Dr9nsp/t1oExzNDfUd1Gp
s99Xzg1XC1jB2LUTvZDXH4+0nbjAEqqLLJc9OJstSzK2cQXkYF7QeexVtZ8yYaJl
Zxj7tYj7OUBYiy6IMl2Ye5yO6i/xMq+xBekmlU/UYd2woNV8pEj1IZgLJ/svM3j1
mlyxcrTV20yasGF1ac9y6CIj/vEkalio4YVtwR7x1KH6VxsfUtunk4CyNMn0VcMH
9ixIhmsmdP0mY9VmFgKbUx1P3aUajoFf2bhuFiFYdwbXVfq4DD65GP/UI5aBHY6N
GNHsgkWUxfjthX0KCUWwjvHQngd7nJs4J4owzaIxgb+64Qe1P/gGIVWHgCrJ9npJ
tHNq5uosO/I8hFud4T2BuSKwdo64GIo47GC5AsLfxQt1Xa35JwpQRv74KmrnzISY
ttl/rid9IEMn++im2XieMzkpo1kgne5Mar8GheiB2LpX1zldOvIHl5cAkwf77C/u
sCzywCv3tC+JjA/icSQyUB+Cd5SBml6raVA5nqLY/a9VlcG3qhRCRUA425uTtsx6
5UwGz11dsitZ/VBmIv1g9WsDIOQnDxumN/eRojLW423fDpMDDLmjBzhq75W2UwKa
2iIABFOyE2mVQ77UyXG0S+fuGl/Al2utcV1JbtwvghIMruRuQDdAg/lUQkafUIPj
Zte5T0M1boHYGWn49U5AoW291dTVP60rFvn8Uo6/WWE49316CpDS0qwLFOrJ0x/s
WuWKRQOZjyYVhdvvc5UmNKXt4gefqOD/tJuobd5QRh2V54y4h3TlxZooWd7b8QGI
HtN4SmfteyKDlSaJK7vKJTe3jOG2qUTskSS6IAqJnvSE5KMk+Kg3CU6XNV+3X0rf
cWn1akYdz1rok/rD0kw9M6RxUtToGcjh39AueRKw2Q3dd8d0nbOT+/956/rlnyW9
+dpwM+3s51a3AKyLQecfQEykS8YVUuq4cl9dWjZAemnALVc8APyCrQp0NieziJVs
mp5jGkEsSN9iKG088K1AYgi6jeWEkkqwFGFBSpHwz5njmoe9+Fnm+0DIeQ0g/A0p
TQAAAn9EUellMPOCKUE8B9Iqo3CgwLmMnI9mq04LMxeJ+Opa/mEFfZa4x5XRNW5y
a0jttS7GkA2HJHjhrMBGz+KAKwaNQ1acqh5fw8Xo3Z23qXzR1zF5OKi2gpZyr/rO
GMVp08/ru6TSwUsYfRb7ZNGtNqNrqB97pu3supkcoR4pJIH3Ic63a6HLneAQUcAL
sTEDc8KnF9tQCtQSN4pVVp5Wybz2VrCLZHL8PCbs4XUD3zWVaJgMULtrlIm3bEUA
+8PssfBYo1TUhXGLL00ELLmHU50ai0p9pTrN586ZRa2h91OKkVH9dioqQoORkORx
ngI5t/7vwp/IWGC0x9zGZZcC19ETLCDNEAWN3Uf848ze2ecIdOulfIxanb/lc0d0
VKCSFbB0sY1AlsVi+/vOdyyRdNEfsMfqhNKkPT3bcx2LKJsMsj+cDvnJpdX1KBvO
nS+Or1JaYZ/+bbucDGoGRl5eDZUEQpZvE834DmlSio9zwui/QDFSh2+pjDH9TntC
h21NCC3o/jJIqU2s9flvLMOGTGVMPUMgUEqPgIQWbr7BsAttZdl4WmdDEpEL4HQs
Hyzsq8Fv9UilZM+dFBVhJEmkX0KTwQ1Dsia5Ep+bfZbfZO7qZyqGCIMwbuzjpbIj
iVqZ9I0+5ejgoOxVoC5ZPAJQii8p2SvF7UncceIkVLFCqNsMSk1vJpImVOuq/0NR
BJiP2e14UR1rZbN0TnQy+MYvdlFtUTw5627fySx58qjaDv2hJrx29pykYT2H4zsA
BetWIln6VN4tDhwIoLVLPdsVn4uVNmx8CJq0lOJLCVFF0XLADAzrykjrVPX8a0Bz
ybK/RRd+3u3mtYtWgYITYTSLid/VNVm3u9tirEDZREWMimZrhKR524eF3GJxqO4m
0jWVhcTQTMVPyLh2w547TY2LKu2kw+RLtGwPSfO0hm166GMsUTUDzSzvlZgN3CfQ
v9Cw+saen2LOXLUg8sbFcQXuETQRJj3DJGartinS3Yz2xVb7/ikwaK1+6xxobSnB
qDFbmfMlUX7KrnbInhOk6eLIo2QENpSpOGHVsj9HekzWOsY5uemMumVdkIt+rLWZ
trvTph8RkHtmuN5vlhzRTiyTKVdfT+WI/G3fQEAjMAPJOoIhF4q52jyhklfd4tHF
8wVED7s+ju5luVN8i+jeyVK9Vr9aQntEzIyqXMosImmmZ3bdINhjCtWiPuTkDnPt
hQYz2g4DPTbkz/Bi9EWBfrvgm4wNm2uu+1yRTEs50Cvc9EGnZKIMhXK10Hc5BkVU
MqjMSqq7lhC+cw5Xf4rRMozKXoMoEUnJ5jSMxxbC85tybioRSC4AGSGFw1mYmSpf
CdzH+6xWflmZltW915MWz/Ck5ArYxrVh5gAW2zkK8hEBOK65NYDQkwNBayKy07EW
AYZ+JvHQUChwtwKIe5sho+XhC+HuYqr2ZQo1iGgWrClJ6ZMkIaNqvAWPx0v5Ao92
ANj94uyZgzMOG/FcOMffnedqj4vGNiwq8nPbStfjAl0dVA95uaSzqUqkaVDOXRCF
sB+BJx2BFIKtXOG8O6rBu/HNovS+/NFVRFFXOrnU7LJPit9l4aCTJacTP65eu0EX
T/do7agus0XVeZLdpItHNmPdIor6mnGEjDXjWnQEtYFauqh8LeQJuCbwCnFLAgoE
LmKuA5ub4EqRV1GAw+SsqxJnKo9o6ENoPsrxLQceF15U/TmgVD4PAO1HdQ57FMeJ
sF8xiGLt2SBhaR9FtIngwX3mYnSBhHakraezThuc6xf1oklT6anp0lYvf1xH0XJW
y1wwEn4fAWMhm3LtzoMsoQqqxRQbMkXnkZQ37KL7pjYfDu4vQlqF1k887+jUzxQv
0nlEQ1yybjpo1FYs90zVUL7hB1cl890/GrJAMIHKHhM2kXxXCoQ37+2CD5ows8Ts
yUvf94TROnuZJgwqxOkWJWDh085MUrHzf6G4yu26yNQKe7uVEv8OWLd1YqSg/kdA
jw29w2Bg7iLaRFNm0YrGmFJtngHMlSbCOSMFnvv14W2K7UDspMhg+uhukksL5ttp
jTkIkB69Vwh0OEU+3rUV4jDcq8veowG9QTSr3yqTJ/kH59yqKwtcCU7JfDXFqgdY
zul6HD1DSl9TZrtJz5J19Rwt6qLunMyohoGljhsocGgBjIkFCWZkdVw5o8YVqRSQ
UXbpcMx3X153dG8D0sxy/LZM5I+eITYKYEuyez3Jsqhc/7ToyAk0hSOqkb+nd+zO
V88G+y2NOti3dlEKoBD/JEhcIi41Qc9LPRuTtZiGR68CRyxwVWo5RV8R44oSevIW
b9C93uKqulpJcZAwY80heHqLKNfNbBsQHfuq0bPlWk1uumisgre4VBiH+2bTaaXY
rQYMdw27trtBxi7LHHpwmFILuN3QAlpYa4V5FGZUGCHLw3IKTqSybnPyPe7exHHi
w9ubTU7chsnfDHt9kbN9YC1zj/AqSM7AMi7U+IDK3/26wdKUbNsS1dffXH67K1Fz
FFP/DzypwCMqUA0SAO2Xoq6LBdLxSFRkykDtUytIfji39eG1ev5WuGxuNG/cJ1IQ
bW3ncQCOT2hMoUZ1gpC14DOFNOTH5aYw1zZiON3tGGXgz6elE5bL8WQ///NcRBwY
5nSIgtAt1MF84AQEzIlO0+mrE4odDAORMoDjm0uu97olPO8nRmXctqSWxc4BT158
wznXe58Wp4LXEr/ErkswIuU7rZlRM71hOmbOeQ/ktU6Pnbjsh/pnnvzunVIfcLfE
qPU6tTlCGPS9tLOYNC9cJrS98vv3RS2VABF+/V+Y92R53caajCYGP23WtEdwZDUZ
avkscglh19apqW/sx5A5Nr3ErlJdq5zJy6xpwEaGq/4Lxk0YPgmTIgt0827UKT+6
KmWE7UdB+rqSeh9ZnDjx8yOx0u9uSzIne459FoqZkuR62EqDnO4TPnwLrq0WWYw1
gq0mWIAHC8sP3fNSXMygOdB1cYTqfIYsj84uobEYP3mjJi3aOz0kU5hubM9d0P2a
6O2wbo7nrUEZw/C0W70xp4VAGNdUZz6EtYYeT3BpzSCBeJxZoO0B9XaDvOMxCRY1
UvXYh5gcbD21Nd0XH/32r9w0Efw/SBlHgXfqnTQkvCuAsMrwQYyVN8fdqcQ0L6PL
auTfnaGcGunLWPm3e2uK5Sd6DqwcX4xAquCCa9uJmYls21HdCimCRHOGTlsoC1ud
qKv4xrQiWGDvCK0Ri9bu5df/pmW9EZSp/3nANnv77k6OVd0t74KAMkqTfudzg7Sl
QWow0unlJwMAxxMiHS8veYoF7sgW4mu0RXzuvI2o9b849JzXgyE/1l7vHnoJAk0D
jPdN4XRSu+PBTxsgYesfr8mUm36zvQRYYS/93BbNpf3xEgShMnPBfsqP7jZfXSDv
Ri2T08I4U64iN5rHocCZYqPJHC63dsCVGY0Ctg9wVlfPX0mAdVaxF01sxnA1E0NF
GI+WRXbY8gLSLvatObx8tBZzAxYmW22NA698C4vtgUdmoW4Xl1dg5OJ/1pX0wUCv
xwZ6SFg9s4eEbCRa0SaO7W3LJaGskpP9QsPfhx3JBvNVZgvJ1nNZzvBPGQPogWDQ
83CLPGdnrJssvihM3rApIlGzgxBRTD6c0NUg/PQXQU9S/LaXoxGGXwyyezJRHcUo
HdYAvEzfD9aGJRuLvlkolep/C4IlxsLjzy8V62A25jO96uU9hHXKzP1vduDVg1ss
lRz7CtIU6Oqy8FywHcAK9R/QsIxse3TS9OjwuPVIJG+lYuNRfnsAZ5bYia0Gy2uU
aiyaXLFRq5EoqXwmBUnoYqedcFhX2jb4CSrGcJxbvt9AVrsTd8MmTzdMid1Oxcbz
zqFJ9oNX/yuhaEaNT8R5XX4/MWLHz10yeqtS4CQnuWU2bnCSbJ5uzFIpqskSNj0Q
YokrmSpMTEB+zxo7ayKOfibH+5rzC/V2117IFo31+Gst60MWfhmoam9EhaztBrM3
sFwfwThBDssxwH4tRnTMFmoQ9WvBgrHXeLPK8OXKLoqHLsos6n4ayTS78R2vORrA
fk3NM15/Ymeqrh8g79QXEEdqy3/R0vk44XJR0bW+9wi9hXHHo9Mn21Absa/cYpsK
JYmCaKS7f/B6wZLqX+mvQDP9A70Lm8KFk5BBhf/QpbkGDCKx+p2myUKba9CvUOSr
HSlI2rochQaeSdNCFFG2eYBgIlIaXqUkbcb0LJKqEMHw2W02hIMhoGhKu2j8SYZj
G4/gnc051l0bBQbc/v7UOsoNxkdRT38AhvC5/ipsAofPqBTo6oI8dwGdwKgjNayT
LlbIu61a8KLNpFbjGUpNjlGSI37HK2P2tyV/a3/dfpI08PrBTkG9bwIKRleGuuEg
KvPkNmJ2HiECqVPRMzVxIaII9PtxzztCD3HUQi2aALzcZiaJA4zDJPUpDDEaCpP0
ePHlI3nRoXiLBFwA6p43TAhu/uta+yMzvGOLORqgzUWZ+/kUbAT2AfyeswC5KvOB
/THhC094fcC9Qg9JiZStjFs9k5Jyyzmvc6HQQfcMyM5PnvTOuslJE1N30fqa+nkL
NcVC4AM3oJN85Jx62XWONdbKsotS9fj7aRMVyyqGQgf4dBxOA4ZNmxkyyKOKLMCB
jaCFjuyCL/iHDTBB9MMbF5772BGmDCZYu71h/h6uox+m2qOjOlgJZ41ucuJpACJx
+B83c4jd6EdWW8vkFAmBIGC2mx5Cb86ndhM9SKpIcKt47JwkB/3740wbUbEbdvh1
0KuYe8taQMTHqkQTxBjg6oVQJKBHs02E57t8gONYNHm7LPRcaU3OkJmfot/837nk
NZQhAmAFDg52C0+T/pq8FJJAnOyNwHLL6WAnouOsYb5qtCZVcHVHo9qtwxmcDIIy
yU8f72YAWqTEhwy5uRGhWFYir+UQzUaTwD5kU2pMKCRQn7iNeRmuMX8/VmyY5Zzu
ZyLjV2gN6tBEEVyw1bPfPY3riWEufdTGhek1stT8y374F9VEjT/d8RSX8eQ44fuO
6R+KGlTt6YRBAG8hnQ7znnhbCdaT1i0NayAUae8tUiC8uJ2qjNxNn4we8a9U1r7V
nTz1YFZkp90gFiUbzWuETHuNOhexntdOBLx7WMmHBCScRGr/tUB//fRkJ7cnldDc
kgPqBx/xpIPZUPowtA3x0yPyrcn4XCj0aLxdBRaHLgI+2O2QoXB6BEmC/ANUzXOI
T5DBSrWLlOUjdS72OhGkg/QjNcyI55DIufA/+YUciIms7aLOHWuvYs6JI+hnoYCn
eVI5paza4sH/q3B7irx9cJvl6X3xV/4zN6nrmrBYx7A6RWkwgH5L3EYgMoR7nLWm
Nup++V0ie0aYLCDBv9nRBfrW8HDamKBGNixvct6xZY5CGyQQWQ4QfTcypyRMP48H
2m8rDszZSM1CUHq5yFpaVTeC8aHq8qp0Zftv/lGbwi8VdXtcAp7tKFnlt8hmCa0j
DtINQshQgthxFPL6Too8daPUhAJkGO+2tfC45rUSzyQPdbFiShJ9RO3aN/8xjK3+
iVjMoHFcFCyXJ+sDo6iM9MFuUCgwpmAymgf+tX8L7e2TD+/OGAHtkICSBycjQjDU
RV77UDsvuCd/q5fTJQZnnFRFg4OTa5GKXAoku1I2Koyv7d8c6SM6hwAMmrFMUQnI
AABMZeTIbTRCPHExknjxMqvmGeQYryXtL7D5kISaq9KafugH7MwsrTOaZaBhfkn1
iefjw7Gguz4Gd6CIV0zKoW7bdNITWGx5Db/gEOC6Z/70bhwv0jnuXoZfD3h18s/t
u8ZGiIeVGOg7ZjXroaxVA7BmeUJTS3QqMTwURjVc/FH/dJe5nsQZ5Led6UP3kxx2
7LwLVuJCkGyVSOTDvKcr3FIf8qNEMQpCPkmqbFhoGUbf/WWnev6FN37T+Oz8/mt0
VvBeWaU+1rQexY6A/9KIbmxaR3i4vt7BTIZR2Ezuu4/OrYPxcHFw1EdBGid4nVuq
YvFIvefp5WNncJ4aJv55LB7EoQTVSTr7IhuB+xq2Tpnw7o/6Hl8t9mSpBWhcDpJy
7ao+lRuMKLLwHlxzf3CIeQDxwezV83+YuiKgzErnZfRDBZB0nf6uOzIpSupcYayx
1AfGoAaPSz86Mu+NMuoJsjP1Y6gwtS0tZGsjja0oaVcAIxmvBPs16bER9fgkzVIS
aajSemAtymRYk3XktH6BOtCUE6qqTaf4RjwjjieNPCzBGttpAaGPfrpMTz6WlJTa
zRYGSlEdgdz1Hx4mnkNcuU+qHgBn5A1VivHw/n+FKnFQOMUclEIyvs4u8jiGCeKU
HGxnUceMz58gmgrh5GZyA8lx3HzftzZ2234/VSgyK3So6iVoKE/VckgLiZ87Nn9a
FLZZfFSLIIxhyr+NAJIGsxonggSbMXvzE1m0w5wzUufeJcx9SXpup6gt9AHd8uvQ
fA3jJJ4dGmJKsjZmEiS2K/JtcR7ajHfV8Eqt6DFVVkrQY+OHbbqUv7eRi97UXTxp
VRBsmOdZAW3L99kmFbHrkE4xFH2LLCr250aYyTi7TSRWVc+rGQBQyzYZ8DBJGjPJ
Lh4AQbPYplKfoZflpeadAsAY1Df/WgIo2Y7TMZMXoofr8dqLs4sK3bSl7zkaSaXF
lNtmy5J0HwKBBJk2vma6ZDNtvay5YS/IHeTHZ+oVNFPpDnk4HORVqhDUnxCh4oNl
WQtJLaj/NkPmSqxHp6OnxC6RW1cptW21QjCXnVtn0ebfIe++gqAxdNstxRTHOcM+
RK8NZcr3+/BVE5eD+Vsjjw2NEGSgc4c+YcEkiWLnkraBmbH/AG3Ic8lZBZDqgOl/
DXDRipOg0p98fXC+RR3Xn5M9fH7+L1UzYHAPVebAxtGDVYUFqspI6foO/6wUYzvb
OKtkr4RP3bu1uT3z+WK7RNHzLt4TKnZldqTy6yW/6tvbywlvTMjjTV1YgQtMFwIh
kDXy6ctcmsWfFynhq7YBPijaH1CiKliExyqMTRMNelKprFIxf25OwUxXQU8xbbK5
7DFJ/zCP0vRPtg2Wn2NQvRmqJwNM7UbCvVaMJpo8JAig7GrYGlC5+eoA7hELKuN7
wgpv+ls0GCXdR/PkjBNPIAYJlvekmniyujPkM4enOuYKU2icmJjqwNzQHaa8yr7d
hDwMCaVbh5rdCHir6gNrUqrqG7JzwY5nCEr7hRMfaNMd1107dQ4BP8PU1IHlvHxt
NwDkNpUJ0K5ZSE/Myqj1VldWE54+YThEpS6+8Cl8GP3S/oQ4BWgTieKhs60m0htd
lZP5llBjcG7UE4KjZZYSyWLfK76kPvbipVanphQRQ6kmvUN/WsC/Mm7w1exLQeQu
5EY6oLxkV1106Kfms1B0wqWvC1OkFQBAUMbgyKDYeN4KN129oZ+r59eFiRi5EgtZ
vihK76qaCKgCHgdRHptxUia0+1jbC8YDCu/SFupfuKfueWyyR92GYP9JlKPn1SM/
OwYG00ZSp0Tz4RNBxmIgjdq4zLVfYv0iE/28aaNHuzK5m3kFpiKr8KIjoA4a9jkX
dqGLALI9vOxePcgOv/OUh/542mT0FwYp3idjF7yXlcZtfL7Jnfkxy4W9PTmwESXj
KkJ3xOVS2qEpeGYQ2jYPRCHpq6IhI8SKeEPJaoaePQTjDKpn7mH9VlTBkcZdb1++
DpfC1y3JjUFirxUy/65USN1QhHPfPAVKkFRJyQ2Sbfqu7pfipigJF+Jp9tch3hkj
A8Fqc5/pIB5cQ3xbmh1UTbFBkohtD8mVMhYYYjDF4fLYom+nT9FAvh8B/jSC7yNF
47+aYoAk3JLRUYppKDOt8PUq539F64UngNOi6bHHvdeh34A0XqS2Ul44tqzYIrNi
JrRjIRBy16Ga7Di7qNJIGu1ak7+oJ+P57rxtVvzD0qX2CI/SDmon60iK3nwUWY8C
o6Xs17YQW1jn0f1hfqShofGnVstvlxR4t70bHBPpRsYULxIw90ZSP9Tx5dCsNLBp
EEo/ZYjAPAoqVokMg2zyKs0gdlQacPD6jkpHWukrYZB03A1/8sgD44U6X6iQzS6l
4PrYiZiwdZnQ+6YQkYM39QYRtj4M7fk4EGMAN1z68GZMMT7TslnKBb4Cm0gymo/T
1nkqs9LxAHCQBvtrTYV0gncl5Vuvs2Bw2W5NVR5CGjL0UKpoHmsyvvYz937Ow9u+
YEARc406+RS0ndZ2zEy9+dullorcJqSBdA6iquqIp9oWa6O+pcAD97/cmQKmB0rJ
B4539pPeaU5D4Sp3Wn47p5QqU+1g8FXjk90/20e4upCXCxJzY3Otd/tvEB6r/rQ0
JkZHFvLirF2TpEEpxZwOxI6U56nMA6zf5CT83Rd2DUca78kPCKBcy5bRiHtmQrZj
x40gQzyVj90i7/tfQTljbv8MAgRwpghDdc6GMgporLeRC8m+gDlIUkA2WTpN6asf
FpIK+Mi5Vh0ENnLk1yTyxGasxZMdgomXpkrjRucDSy9XzaALEVLXZh6NOTAwS2F/
UebdEEQgPD2cIQj65easYMtl13xkIVFo4aD7bMZUJzLA/yWgLv+TxxvPYQsL8ZNd
wnShPVBuB/aj3nVH/fEtf5/bZByXzx8yP5mJ7tVcRTeXEyjTNNhC9hdPV5UFcGUD
hAWlubCyjyXXtjX6A8iprY77Bb0jhpC5JLefgoaUubfjWnuqETAaEIWCQHNkRxAH
RFo/dUmuYRmCNV+gdPk2wAWMz41H+y3ar95kYj6PkqPZoYc5lWC7CAYLF/+xk6Nt
jgaRgvEkQZUyNbuWpFiIf1BfVOiMsbUqmyAturo5oY2XO9I1GNHb0nsmI0oOwwJ3
j7iSO6xU9BquxMveDSgc8SbfmoLezJ4ZHBWOpsEqLkswL+Mo8s1doV63LVWTSQcC
Cb7piHgVUR2SCd+8AvKSHWwbJDb7SMBrul+wI7kEaFxwOoI8wVhWSWeKf5BpSOEU
gvjbCjLbM+0jefMDn68y1llNPPaQ4EIWczzeSUHZ4NGNLB8u/be86ccSts/cUaTC
KW9a6HH8vhJvbVy7sCSFRi4C0I8fn6FZsFbAT0PBLa9jw2ntFD06IvPwgwOj87VJ
cY3TX75Ma5Q2KpIUBv1CfXBYXfMZIY5lwTUvpv4uoQa27M8gE/Ehl1fJEb/rZ80R
RT7d82atNZRJPvQKkDlbDm75SL29b1284zSwH5ytSyNQqk95+1iWl7clvbcIbvRU
/824H8CGj2aQrSvN3m3UFl8Boi3UCpKsF18WmZwjGiu1GE2ndud1INvS6kzUwObS
Ut6lu4OuNzJY9LgMbKVw6c9W4oVGtZ0NOLWCMXM+aQz0b95H676FSM4ZW/dBN5lA
yv+utW6Akp0UuvVkt3hHurdBDulBwcfxoP3b6GOgXlrC5+OfJv9mgakx+ivQdgk9
H4Vbmc2cfpBFb500QQT20L61p5gDsY/XpvXSmq+p1hy6cLR7yXDr5soBboI6NumT
fq+omwE3kqf60YMuqO1HjVP45ffhuAyV2QgSO9A0i/LyoEWebCk4fPnRGvHS1lyh
/hTnxpJodUnxZZpFp+aTS+FQ0LVBs8OGiEdtDsYKJwbHLJ5wFmHq1UCgm60ZLh1S
YDc1hRHu1QBW8ihAf2vS8MQJz0wZL2qtqrwT++oYQ1EP4ErfCenNWx3NN7Wa0mWs
Isfme9LL+uUtH0Mra/0JU4o104BhQdg9nIpAcsDNOmisoblP70sT3dD1X28LpMnV
URfJQSqA5LBUMY5+PqIP6mSconOZ+ML4WT29ph+hEw7AmdeT1lqulsqxdZJaSA8Z
rQ3lovalzbs8kYmGLOwo8Jq7ruISljVlbJI/IR4iixorMd0X/ZidUlB4yxqq13vu
hdeAPnjV8a6IMc0liZlkuXmy3BHb4iMcbyA9h/G9+w6x/ylLyP03OjjJwcnYYRSS
VOdgnJhPZDqE0DQb9PGz7yMrCnmzINER07U496eHb/b34Z9L8ZhLeGSeKD3plwiT
naMtz6AvClhI0jv4Ju2bUsbSvmwh/vP0k9JCXdoBQBnH4EANcPI/ntuk3IQVDxn3
dnJi13qLUw5O3RJqdLasIZKEgUrMoUqVRAnvPOtCjJ4Yhd6FKF8bWqkV0JJKn3KE
P2p/HaLyNiUJnp0X4VJc6rRuJ50v4aRUvpYWTaHm+q1ULqL+Yw8Fue9cAxyDQAYL
vtHschqaZQVUnpw5ft+O490bg47qDT4YRZvEd7ZQe0TzIB4AAHC0iy4/bmMZ2XsJ
YzBJtAzjytPPgLT7sQ2SX2EgkJl6SHNK2H1bVli7TQJN52mnK/eh8eWiZxAxbYWH
fvtMBvZvgZ84z+3VcYbktvuNT/EUtUR9UX3JtVl9pbHS7zDgX6sIFDdBzyhYRgxM
8cLz+bILI0H0Yqf2Vlw8Xj4+/EXActqUyP8rrRKrxuPWmA7pWw67Hr1hE2Zujdl1
LD67CIE1Y2vgSjVOlYXBiBkatojkxYGUtJBwxF3flC9ytijhMl5B8boEFxSj/a/h
ei4mSAHAuBjSxMJT9kIg/GszWxy3mQwhv/oDrHjgPYZugS8t4s4ceIHfz66dquRR
DRAgTqX+QeD2HKjWpKjpa4JWj75WvsUklwWEFZEgf4JOy3helsy3BOP3SCceN7f1
JEJhmSHwrOxJJ2kJLXEYOGDn4IujIG7roc0lpnZzPXOpz3ncE/Q10bvw++5CuTHC
tiBmiiAhyuDSlAqqcDGahnkLAm08/QctdBeSZMtY8OdCEylWKwyMoF9WMryxcHEw
tx7mP1iYJ2Q7uT132oEINTuaLTsIvv6Uhk7Xi+mSKCw5TzxAVCKtwZ3ERWpyDCCC
+EwB29KeAF+Xtqvzzv+/WKNX5iRvQAB+LV2vQ9KHp+lCUVAMD+RGEjn27Jc6ouFr
DQK2Tcgz+gu2sE8eNtTBWqWcyS5jCJcoXhig3oq7NLRJD8IMXdhUibs9mqkuHWvx
kiK3Tvz6Yw7NPczHbmhyeJaQiztL2pF7QPtOXIMeec+JgE/cGaboqav3hgBfpBHr
Q9//x0Q/eJhoYVzFtAYPc0R9pzHp5mw4TKUGyla3x2aoq5FRGNP4MAwbPvn5+1qY
OMQqd8zo+Tt3gEktFmGa4oTZx6SCmCMg750EzzAp7jB70Hqxlaxr/9anyI32lxr0
d6zUq8scJ5H5L8O5RH5oz/t2AkTZoYSkvAZxod7E8X9ERX2kfpV5612KO2Wc3P5v
NrMFczt6oXHE1HICs82OIB5XnXMKjstgHJHrk5uwLuPzwMdJ5mAllV+ercq42DMX
tRyM54NxmMmamfzVp0oqV9PI4HShb/PzSz+gTyhelNbj6kAZRQjjRFLm5SaaAXdX
X7yJt8VOtr7P+WNfN3aHc6OB0Yv4I5dwEqkRt4d30SG9E1lSywGNV2/4AghqNTn7
/TDEx/JjM3e3VPhWaNTBC91DltAAVWjmzU2X72f+sNqIbEdslHlu6J1FWlXWPSjx
gOQhc167pHQ/Q0GHtPI/Xlp2YtFmwQr2kre7iMluRw8BUduwsAl1bD2Q0QrxA/sh
4fKZc6l78Tv+t6OTD5wgvtarzSxNOFO6OlIVFIOS0Vsqxie7Ps4U1M1P9tdAugxy
jNh245lNtvsAIQoF7QkHkFUEPJ4quimPeqUxR2petFdoR9NdlHK9NlmKORvQxzua
c2yWuXRRkW6kZ+I7NBUR3W7GclhluW8nUOB4MoLtM8iJaLYT9i0jCzSs2M5NeawK
8KvC/LP7zMtRubPpqLZMN8daFmn/vA88pCoXHAGaqYkEbHk5f2URQUd+UhI0HRvn
sV6YSwMbYoTUzQ1pfFdtSc9EM4wJFmTbzvTzBF4bTsvC+nq8bBw02wUlh1s85Pmg
fwida4D7Lu5PjGfynpzFHkXCi0s2j7mJzLGYmjQlDrR9DPZFG0HxsI8eE5kH1fFl
VtbRI1/ezyQuXYcqXgDqjlx45OgFaBenh2UEA1GjhDZEl0Th3CtOK07KbdRz2zb+
asrgMEtwhqAXW4W6BMJSJbGNzL6vDBNYPbwvpKdjUXs5Ij0qE3r8b9MI8bRanU1u
OAeMD92TCshXUz/UId0WqXBoXd4RG4ZnLXnzItwsEM9lT0y+xqYU4Th7qMTkgXq0
rHy68Wd90/J4mklr/kpdcd5UqK3u0SoPKLeP5e9qXGhkFk42OVThPT9vNAp71ER+
m2+TokUtwh8LgpUYUMTv1U0LhfDc8IJum+MaXgc05DNCTuygRIGUhdc0LWomaza3
ynAUBZXoNz+TcNrUomrz46LCgv9yzd5QmjwcwreAhtfyaC1RYGDy94NdUCUOKar/
C/FJYy7MIjx27VYcwiqBppV2v2ywv6177FeE+rR7VeLwvz1C/s1o/j3oeaHn0iSa
enC5SusdTXoFxcXWOtfZTCwujKXZNyq6b+38649R5nTOb9/PzE1G02mu9miHBE+O
nCwqFJiZJwfVYaKTJAdFv3qAqeYWq2zXfxbeXSjlJdxLyBiOMPDWVKWKW76FrSYe
sgXS7ce5vhIk0/HDhUodvZVfAG1R4UAHy3C82TEuyr88fo0OlrUXSTbb+te2xphM
n/STbD2TeyLX3wKSLM9nsdaM+/GM1N36or9XIrBKcT6ta51ioH4jLB+ZylyADdPt
QDGgGKSwKezyHwqsalZYb6i52W4tlvCmmua/gjjFb1eAhhXsKvgSB8r0+MXO5P1O
7Us1RkZKZDR7NPcP9qf/DAGI6fPJ6gI+vDYRz6Cw8CUE2y+IjyAayGkZA3+LQHzI
yAq4n46+dVVE3xw25UCVxxaHnd+5A9+8/X1YmbdF7V5RoqavhnmQtAV/F/FXu6WT
bGDgd21NO+k8h1xr4sTYD8e7g4b3GtyZP9npJOZ7POEeEHzvi3YV6l0Wl3+u1EgS
dC656Q0qFq2FbR7ONQXq+QUnrNxjqRvBh0VNhhhczWFtcLhek4nnsWVYEcVjCRnn
Bs7jb6hK/xRVu9iKtapBAgOvJsIfm3dUIKag+55ctP1KZw9oT1Vy73NIMDe3YLli
3WeYaEREKM2lT2czDYDMx8QKwO+f37+bHyPYFfGMdWdmMtk6uzDNSY539SNY2dU3
fH14z3K2ALWzkStJS35BaBjoQxkady6a7QNN+ORye9pmoLBm/lWt2Q7JJdKBbDyX
PLmFIXynjZgzKtdaB314L8Z3MmHg4RKu6EnFSTLqE0xNI4FZu7tXHUaNBZt3aVct
Wh6o0ZPP6pQP/zTof4IN6Dv1Eayy3V9KOhwhM0P+VU/tZLysaBJTkjYJRAsYf5/e
61p5nxW62h9FrZJ2u93VQ7ybHe93YrS2JK5CZo750DjCWUxPSj1a71FsNv4mAsMJ
EevKU+pSh+mwgQpwh2WHbopijz4lw0i5KIO6CXNvKcPCQyDVfogXlM8Rd29+vG4X
HPhanQLHmO1O/I7jATbV6aOu5dUikS/WAhRJ5MGo9IptDyd+eYT9waA40jnCNu6T
TuawF5J0dlYdkjMvfbde3vf3xY82dTf3W5Tx/bDKodb/hgK9HFCTMcUR7jIYO3vj
GdepjpICI68Dqks0FyCTX4Xzp1vqhGKOG/pisJy4eZ/RYLdEPaL7QyNiY+vEQhYJ
4SIkQnTTo7HvIRZJtdipygZLbtV8N/AEyYdfn5vIKHaJ6JcJ2pqOsjW/BmBAmN3z
XuAfbudTFlk2w7hCMzq34LC7qYyGiTwAyO1PAe86vGWVpsmBOwFzJH+w0bp70bf7
O8p0Xx7RvIKGb7ojb/aliprN4SV2Jneplq3P1dSpEFHdda9M3z2a3HS3UnPGU87t
mQAusIN425BgDmsJy1Z1k1PiSYHZfE3GlBsojnzuexeDPy9I13zve35n0+wixR6Q
CP29jekm1dn1boAyQxW7as5lgZ1jDqaoXtuVfxDGNO+CZcCWX6acua0fEwYOtLER
DF4olUhwkOoKveEqGWtLlwp3IEnFR0LcsT8EvbHse6dFl8BdC9wrqElwd8TBb2Ou
gWcp78Ouk7lKAJyo307uIW8OFJu+fpT6gGOXTqVKfrymVMOhtKCM+VaRyYi57Mam
qMRLQP7QSGvOV4LO6nxrSCzoiNXQ8y1/d+T5J45H//nN5FmrZVsTWYxZ26JTAo4P
WJlkvIzvGCesHl/feZd7HToEyBrtj07SWeCLqn25Gfb264Vktrf+noLr+psavX7c
bfoQuxhxC0Dkcu4h7ek0gqb/0RdzQ4HrOSVSqbwqt9WecuQegz3Zj2jsljJtMrNu
UlIw+QKuw5mGPH1lIB6XFN2nBHD4+uJ9Z11JAtk2KEheEG1edJ7aQvIiOhVaMAYC
mednvs/svQRzEcieAEaKSwzROuCpwQXPuEIAqinwE8lut8nBW5AR77x6M0J8lMMD
er9XEjI/bBTX+DWI21rSc9r9qZ5EPnskkLgHJzdR1E+q9jp80Va5KeXUsxJSD6to
5IuTqWlsBdjUFuNFKK4T/QGSZBTDaGZLt8gwbdAUJkUvtddxetZW24loFCr17voB
yfyYdS98KWTjC/AWWsIOMRXwYYFP9TD6QrVHNRel3AyJyRXBn/7MEt768wW2PsQr
drwURwHbTmVD7tWX7BT/6zpg96AqZtoRjQtDDDGlGoiTI/M6FACxjNhCCtMg68Pu
3f1bEX0EoYsM3Hlgw9v+1fqonSpn3JWiyoIpf+GxBFkDcVOMNhEPputDGUtKR0LH
eASmAFr5j3Bs7OSK49HwoYRoEil9+H1ZSwZNZkxaeqDW4xLfv66gKWLSP3IjKyfw
H9CChT3m3ECedD+pGgmTd3CN0RQAzdVmRtxtUKs0wRsVdF0mCqfJhFosq+uho/WS
CBcuMqGiDACZuZuMxZeKGGi0L0Zpp3WMk2xpDggAaGYluRxVOIbkmBxPMf4Yyy7N
h6yexiu5i23lww2NY3neVjUR3fNDmwzWsw6Z8k4XYpADb/lkoGT2omXyYrVmaDPi
wyf8iJSJEdZLgCKEU14GEg8J4eP9h0MurlUoEaxdUtGRce5JHVMKJjo2G5QhpveN
YAVC0MnJ9hBm9B9GwBUEorBn9a8GJG6R8BVTcanY3y8V6vfbZ1jRe+rL3xBHV/gH
UWWXcaxlCL/R3q+aPaLBQhYKwFvC8ju4z0Xg8DhypFWpbl1q0maoZxopOLii639j
yRyyhjfEjocbJLw4y0O5iRoDx3KuUO3gBNew3TyEnrCqeWGoji8LP03KjoUCnSfH
1/CumrQj5vLyVjb1xe5NHfbmnIltKSG99kKr1QKp20qTC15gky/y4m44hz3QIbmC
x7mSuZtU5QKKMNqjp559u/HJIe+Y+1KwS6Fua3TXYRV+N8zOdmxY/11ktX5gqbE1
Tpp+LbBgzkWl1tBaC4CN2pEN0OPCyCn6YrLhP10ZvO6MX194Z+WN+W3tBgEgxTt9
pAfBYcRWjzzXf4QduJAyu82culY3yPDTtMRs4FwJQY0yM2Ylj+A8DVVVEDBWM6aS
r/QSRqP6130yh1Taj5uH8ikzv9q2A9ERwUL4l7R2DZ7Q/H6ooUHZNAazouc7sJhH
EO0ege3OW2v0FA2o4SLBHROPkaLpzJWPQshzE3x37sQGbnW3MOpn0aykauVGFl3U
ircuF1jmmKeoFSyW2MD5BWN3klDHBTFRPg7dMJq0nJ2BLi5nTvX/hoVtWBQGLdDO
rRKR/rmFx7hrahvLtoYxrYEGrof6N/O3X9KzDz+3Cl2yCqLHm+AkBsMJko6dUhZj
IZkGEKgGSwU/j35I+UPZidaDSYBFkBQWbIYILENIye6fEpnGHIsDWRxhMY5e91XT
dtlFMAqBZkSrPnJE4oqEaM3EY5Z6bMiP14wqShvCGohSLBbYbYthVKRZvKCn4pQ2
7YWW5GeKOhnzJqtwyJvBRA7VM+Cxls1pDLVp2zzoRP+agZQtxqlxFa3tOk87kgM6
U4vBgG2V6ywd7FqpI6fQMff8nAlu+JtTAmfc7YVrOZT5N6DTdPoOxb0Nhi4q0yrZ
tqaX64Va0sZPyGCwZb0UceDenjZZs5qcNavQ03mGNQkgtnhaliHaPlxsc1DXsRNO
XjyUsMVLnMMX15fnXJTnqhQ/IZLPF1ym1NaW+skSkmZdzxFB8KtjB1PBw9lRecro
05XzRoDvL487uihdZzM3CS894LeliuuVJyiw2W2cTJtzKqm60dnaoloC6nXG5VS0
zR8r/1EZqEXYcY2zUjkjsajxVIaxKllP49flSMNi97stzrMfoJt1+hRYsVwVrwLt
eSndF6l23YLng4vrJsUoyXWi+Or1v00DEFuzBkhvswbWNrE8uuHSlbLpudCoyb+a
k2sF1FkqBT5jvhBFPlzIgA/fyucFNoGFIrbVeLvZBUFjIhHFTzTcDsICB+Ja7Nmv
SHbFcz/E6O4/bQJwFZlm33hFuxSDoUoPU38BN0j2VIEJ8r8qMMygfeqhZvF8p/UU
EaQUFCZKb3FHt2sEm3I/7ufQwUgf1STuwrx8DSc1G1nfDADcPXICOPpUUx0H/W7C
5CPk85I+B//X7sjP010ggYgay8CZQyUbz4phVWEeEE5teT9nlaHtsjw28cCcqyie
GL34DojW8m6L+V8I3TKSNKtVgbylh79TwSopoS5ZJJ8WhzLMRbMJCjhdY2yAw+a5
ICUYiW7YAQwusIuEBV54GKiAd8+UahI8xlvaRH3v0caDAvwP0Ol+46QnTLgfmcbC
Z76xzehz10L9K/6dU/9Q3Pfb4rUfvtz3PMK7eZxxbn7stsTEqJM7wIB85Uq3BMSX
VGTsRhtggAupHitMsW2+fxNBd+5A8fnx0cEzTwPKde1BEg1qzVNAHmucoA7k/PZ9
QBM1ULcBNDq+HFd8fqrnwUvnWBk8vPkiUvvQIfKYspT7oWUfPEyqJJvwXVORwIQN
snaVHHkXrOHepKEy7AzsE7KtfzK42ovdnWvfwTTLIwtjwG5NlnBQAdN0AXOj8aP9
71+nYh2tGN70X4ki1/epbm7tisWCq+6qU/N4veE0PY1Cdb7edP/eXZJxdNjA70m6
14wRFI94LF+goL3EZKKAKDbJv6FF+c1IWzYBIFhxMGg2H1Rgi7mk1W9dWV0r3otj
ohqeRzjjhu/Q9TovJ2BWOVKVcs4r1YSbJVVDoo+JFAu2btWCuz7nBmAbp9K4B8Rw
IakNqFUGcA5/xmKDBtnkPUviz14/+cc2asez0IGuGMB3ypJdc5jswuOhFCHkJOQo
AqHvMQnrOKaDS8i3ONyErpe6a7NkHUuL0ligiN6oT65e4q4cYKB4Dny623MwRhIJ
Sk0eWs0avJiZv/dGpLSv87F0ymNmDWxr/hkwZ3YG0SGnVa2NOuBIpMKKu/YwMKOV
XrnpUI9JhHHllMqGTYK1p6Kv4/RxSvF07OI+hMijmxkqefTn7+G8n6yzAHyr9fzu
1KlOSrqHGCOk6cBq+0OaFUR7Nx0IT7EKfcgh0/XnhUYP4TELGXOFlolMKc4/6Uk/
Ey+h4y11/eOg908bGt6K9TuwoyTRJIZYEpgFoDnmAyYUMUU9JI3QfvGVE7bjIn2o
2PI0iAS69mOw5Ejb3bQ4NuzonsYQSfP/MHULf23vtlOSUxbMNwSNOCOC9p5CwZA4
Dipm8KUTmTO/zysBC6bnj1bzZCCfrkwI/eOonVNpOD95qOr9vJHoC7GKl7A3FVNm
TI+kThR4jULQfeEWAWePJtxaoll1DjgsrOUQ6c9A4UKkJLPQOICOfXsqpL8IzJjI
8Fx8J1Uus0aHQ5JsbrWOuxBi7quQSUOjtd9+4l/020L+MHDpXZGh3cevH4YSMDj1
SA2cEC3S3z76kzo/ArjQBlr5wScn4Dgr42AaPQVle2Q7XGvWm2rhMwKvzDc4TOlp
jgBYW38Oqz4UUtIJGzE++cVpfdpAV9ugBe/IkeNEPCHhTy5UeveOWrDAhhmR8uOz
I4W8P8LbzfxIkrBXC04tyLwaXS0w9uZ/BluTZ+yIA83sSKKNylPiy/DtJ1uRjNKo
sfTkDtixA+3DWadO1hMVRebrnoq1yseYQZWNYkzKwDxBEuBkTR/vu0ySuS4xVJm5
4w7Zzef+Z16ph3LbnJ98KzoYKoOwlmlQMMgY88wWzPvYmjT2bqokhg/53T0Zd5+d
oJrlK0H0uFdEo7IhOZtuDBIWWOBhC5g7NJizIgfpTCkYBDI2WMCO8v7wJa+XghRe
/VMvIPbfgfhKB4Ch46ykOKNPmD8WaLhuSQ9BRYbeKfJoY+KmcuC4RoxNr6p3hhYV
Vt4504m4cd1cHVZnOeN/l+Me9T62z+eaNYgq1HYEzckY0YGb9D0V5Z2h1DPQZVTa
+FdQZPJo6bFZP9hvw/YgtvDFVdkcxbjEXpzhQi4xfYPvZfcXLcPiNxyWDxsZcsf+
3GWtRFR5OAzegxbKR/i8Th0n569sG+XfOHlZ0u3GtORh879tDur69ppplOo0hTcY
EBsl8pbF380rwIbRwXzhVjDFeIuqamU/jxWgByEXBpTCBd24WMD3Pq0z+Hk+dbSH
CaIixjG9t1K8KBfW1IUMWqPidblA0IyvPrI26UP5r4+uIEsLKbfn9FgQeRE8sy1u
vG8hn7+RSJBKRYZntgSeVmPAto6yiY7D3n7yi9+AakH96+zrPuwVdXZkhjH+2GNr
5BYLKwYyZqMRRunZQUsbTcqrNvgWoEqa8jYWyFHmP1azzN3PkLdG5zNhn2vgXVFU
pwIKIa/VzHbKEJW0N3350SKPsRDj/thu3gJhaV2vLKqQ8um9PHI1h2l0YQA+MpRs
r6xSbSHX9WgXyxCNKfkZO/zutXVJWZnXffKcY1VqCsZdOOLzUboncCECkeuc4Jnn
QumDlD68YIzURwVNETHgka3QGXkaX6mYI873JU+u4A9c2VTzUlT2FVzyne7ENUc9
GjHHQBwUGcKiP7BV6oG87hw4PAtCKDCr5bfIuS6UMP+Kj5Ai4Eaf8Y1FLlY9Bey6
zxFj37ahXehqlV4FQUfXGXjZMn9vnTJ0Hc2bwYurMG1Vm9EMcAVjwc/Kt/XrrvBT
xT7k54IZRHJ6XUVE2bXNIkPB03L1W4yum5fPt3lJkBt7o1dlgzRylbmtTpkgrnUm
fzl+WnJyEO+WSid+i0kZBmQBQymt3gdz0//qbgbpnr7y2x2x87Z+xacHiOdwSIzV
Z+WMGTG3nCHUOOy0vvPjUD8mdIvqaww/W/DCVGBWz5nym4Qn6N+dxMOpa0INNePp
vNxLmTAN6hkI6cIYDT19W6D8RTcXWIQtciYWYlgc5qkWxF8jXnwoLFi4SjoEa4dt
13bj8GkLBH2dDe8XNce6sl5TL81ZWEf5KwUe9Or8yLvwVR3XGCy48pHVFeOnG4K5
aS+/cdpoBNGmqlrLbRE98+rKfNGKvCsKvyXDdkIBcjuVwHA8JomZs439QnXt9XCo
8roh4qMOvOS2c88unPCFt5f3izS/69UfO+xgamurQNCGDay3+LuyQX+LqSkW9F5f
VGC9J00VZcmPeLAmPrHE42yHKFd2LWQ9NHDYCxonYEIZ9Enrhan56CpOqUKn0yZJ
G2BRJOu6URTpjSMIUD+atB+BF9ho12/MmbYPGtIVzBM3Au0udacoFEAEIc8ll0WG
0i64Jzay2Xm8pjHuRH+kOFmu7nNugbZZ982kXZGT12rg0XuV45yKVNSXfXT4JxWb
7R5p/WcoAJpRV/USEK3ua8+PcEfJvGcjceVLfUNl34Vo6N8KebpoBuhJqssigyQ4
t3RsStJCtCi5FvfsyCRij/YCGGfZJ2gDm074cGtNrjS7C/ScfbdNOQODuhj3IYIj
4XsutjUaaRFA1twmJDhZh5WN9Gfc5f7JE/l4JjuW3oKdN1WudVZqHcnZa0zSVRcG
gKjJNiWMpo6bMJKioF7zM3JkxG3v0GptoWnlm7e6H5HBqWyAAekIt1JjfFhSrAYQ
kA1pD2FO+zIaC7TiJisS+zFoIDzQRu75YoSZcGsOJCKgizumGwGb5wyd5DH+h6uL
0ka85KMKC935fEb5alE++R2ubdxLcDtba68a+usR8ZYliDJiY/0zUYX0THi4mmPQ
8fbjzG21tOXzKdIVn8mF0V5Kv90lf2Aaz3R/6Haym7z7+ZHOHzqrtTxBsWa39hPp
Hnqq3KwE03tJRc0GI0ZoMsIM+lVmndhPWnxhbtzOYNbBucWoXH8R1LBAi57/ZsTg
hQgRIUYN6jqvLpHMoOwuDac6zDTSDmwWPFl6Veu39FWk1nZPAeGVVgt/oIyHZJCF
KnpusnhGk4OfwHYJZx20PGvhEdFeaiuqvHWt4kUA+msyrq+dx+rbc5wEmEu0OQh6
7XU3l87z7VOg8oQtfbzFlPvRk1My9OJ+Fb8UQCZTw02XivU7jUqxMfwg6kpVBCF7
Wty1/wmJaG/TEZAMOSApyUdRPqvOK8k5Kj72SXdevRaolbOs6d4YkLExIBUGYVcr
I0Ho/Me/fJo01mBIaPTxX4GqveEPDFALCIwP5RgVgALiUTCHSlI5b4HQgVbV5WaX
Ve0HhCGChSoHjEJTPYEqfrMYVCuDOSZr9bLMSAat+Erx6P5ZrF2/uMeJ9Z4Q1W0g
3p2W2TIbOtbL1LCidUxjZ5KcurX6A/Ok+IRVXxNKPELWgTxOkkzXIn/acM/IokvQ
81EFwjHfNU18PuDrMfRU1Ng8fSqexo9SDJQC/4bDZNYNmNE0rQvu4cw9ulXyNXqN
MmMAWu5c1vcLC0fcwzVfrwfqgwR9OIBsD3DqglaesxUVteX4dVI33GBTvXluoDVG
GotSvrT87YiRjLwX1RnwiFpDEeMDUlMOZPLcQhr/FMkhoTcl3Lkm7DmRjACz3zhm
VMVHRRBtJmSQtDFM/CKq+LDb855BWuP6xkbJVVUZWKivXMZQNLmPBPk3vdT0y00P
xwsbosaYD9eWoY/mmwixG8wPiVTfoUe+oE66VF0Bey8fyPXDxEgEx2uOyr4T/fX8
d2YDduWGOoWmwDT8pqldW42cy5eqdDn0xxNKFNKzYwsLNsMhquJ/stEH7IsYqo8t
iAL+qSQL45ytQtY19sglRSjfCzCryVzxZTuFUZwHZyvejnQjJybzG9xollFl4Vcd
O/PYoDQFgAGCzyu3yDvMuBBuyO37DCfon4gtmhRgCrJzb6PuAUuDOKvPIqiKsM6p
OGOf+vsptt7tDeFinKqdFUI3nrxqrL+9Fkr3RVOhzzwGvPDSVCJ4YPyFHnLwPvTW
iZTAjmRD40+s+uudWzNVDJK2prFsc6mgNQHlFOupK6Oe8AR16qxsISdNORpcvik5
X6E6qNGTL48KQoW+GQjbCtnXpbBe3KJ8RFKja93f6fx7HX6DN+yLSodICdLqGrLf
V/e89ouyHyQRqKpmBBmZsQqMNt8KCBCy9YpcVfTX8/GmblqNIruyLJxQB7urwOpo
tTIAcjazR6AQgYdji1j8QufnInYVF9DviYf+B5I9vG6HJq144FhDModSDkdW90Gq
QsAxLkAkZZpP8VvYzvddNt2/A5zIrMj8CxZSfoR++6gxvBdrl9lfX/W8rsxYARfX
9Wjs8i1VZJeBBl0T4mJRibWT46uJFc8XZyRkwafJrHjyJcx8W+bsFfPtT+dshDKf
BXpom0LPTW4NEWoErgMvYZcEaA/8jLJZS6LKiVsWhnsQY52zU8h1iUIoiMWNl0Hj
jh5vU/lSpDMTfHdfcze2S93X7JzxLI7hl9IXxsNfEASwSXopxiccKvIZXRTmBlwW
SioAIR0fdLrd+WwtIokosZt1LPmmrY6TI5L0ahs9/T6eaq9U8cdHcpUD07tiHgPb
FqAS0IVpCgDSh1EVY5sIKHag1cbkgoyGfdqaeLAaHdyMwu+kTaMpwv8QlgNFnB3J
E3n9iGO6BuG1ipJlPoKWIczMHC80n3d61RD+A7CJ5Cfjrw9m4vECrwQOl87ck+8G
dv0u2PFaDOjvwC6xBZ+IoLdzEF2JPTOnAA4l9j/3e7MroCl6qHbkBz63GXH2OCpW
fzLIkU94iRNN7Qli7HFQ6u1cYzL0tfs1mqYWV0l6z8wc5zMeEm06umzb8Ik++2pk
Y2MxHqKmxiOOFXUkn+b4iw6MPRql8bKv+ccfyIOl9CL/oBS9N5AYB1NZZ/eZd1q3
FyLk8eHxT2BiI6HmXDoXLr2+VsCRnRHIeDTxHBg2nyQ2CBSnZbhNMCe2s1ZbPxE2
SaejoChcoyxNiI6QABnWW+pwrTDXTrn5O735ZoFbAFiuAukMtptW+YDPqQfxmkPX
ps1GBgx7a/kIrcGb9QLb+a8ImJJa83K0cDC9J8QGEOnnZ5DVB2WjLsKW1nlClCxF
vGZ8pbVXo8cNftaNI9O70wa4ipUAGgOU3f30xuqDfj5jg752wIDwmbXUTUIEPWOD
FSTsoUZDM9+ph/UD5NZ/sceMrFGr1f0/UWIgEQN8WeCHQQ2t5LHAydOWvQgWGgb7
OBjOqtYOWCQA0WGnC95FUAlMr9JDEncqHiJmzcQ+g7NUKj84ar1Sq+XnihkFdTYG
oIhrJeNARKo9L4Er7MnrnFi3xH6nuUT35ZbbBArzMT9V21tSW8+9XF1ctVi5ZXUf
qnAcY1HSIaQ6sSbP+wc/gzhfLrJi/oIxe0c7s/x17ASxoACHAJtFWWi2c4PUnfW5
m6dI0IPb2axJpqbgHv3Va6kJ8JMEEWmPyGd0+ouTKDDLalELeIqFW8Hj/KH5pNx5
+HfEGuaZSniS0BxfeQQxBUKSZJg0KKObOgQT1dA8BRFly4dBCx5uOaEwyC9E9vwL
N5ujDtypQiKxH8h3Ji7yBXrTfingj3UK+JCVqlP03n+TPRY30BWIJ1Xl6MBVOsOk
W835BeSF+yeBYEBMf9nSmtcgKCkvdlJOH+ZMaYWqgJ44Ojsm2NNJ1rOLIiZGKGEx
dtJCz7Od1DwpLrLIZz/OWMfxdm4NY3i399a4fbASkHByx94aA9rutbB+DLGutnYq
P43d9o3qKpN1UohtOm1FcNAvAvqn1PAMfXK4jg7Eq+3oXv4WeWZhnPEE4lostXdF
VbQDp+HaYO7NufDiBYC95mCa1W1rXTDKCG2y3U+Xl4BUyMcGXCfsU2854LKQepf8
vuqC49PvK+Vp4x4UsEDSowTN2mJlz8c3J9PcDnRRkvYc2anFbpYhOLFOV/ZXOFnB
orVzdInbSqHXfI3XY+SFx7etuBb70eXkSI5bjzcrWn2h8PQqqgqgR/54DExY6ddX
e3lwJwEHeh5w3PVvj6UmX+si52MJbkI89QbE9ecr8hzexE4EJgV554RuslE/YCJ0
T9PYjIQW1LHw3RLtnfuv1wf5AqDqZACrfEN/G4Nbrt9u9/AqPfHX4eGQ7lyL5vcP
oFl+98De9x2qCP98hnomWuF+Ah1Ri+q71eMFaSUtBmgNr+peGOL5eji8LGd2UIeU
A6P52W/NuTDz19/Wc4Huw+Pb5JIfF5wCnH3Jg4VLHPVKBRMBetXvhEDw46PBSX4c
V2Z672dgHdY7a0fxME6kHcmdl83i2PxMjYuyCDVY0a0YrWNffP2rU7hzSPL1x/cx
x9j4jQXCyytJv0cjXuXfHW2UPYNsjJDUXQsL7IkMjz2QlcCvfWeKl6jB0xxM/A24
wmRz+MO/Bb5tJfRhq1NbLpsgCeT5FVTDC88uqXLB4aDHdxZ6HijlfZjpVzh/oGG+
iiLhHFN3QAc5XV6txfGjBmSyRgoSxyaz9gHyaN8iT/vba1DvBdd+8708u1JXci+l
24/xe8V4ygqUx60IICELGXGNK+KvKwM7JLzhyHBCPIG5W7SzQuC7TW97dO1usXNF
FjoCodD8DLSSXLFSQRTlykXXH8UBV0M2spQVSQltO74yk39ALuCYqO2ra1uBsZh7
BH9AeRyoAcuOUbhnqdv2caXhFAH43zzTVRuboKCbcagPKZUb3SRcZ/DhErMM5Rir
zzDpjX5rRAeFTJXpBmtxUuAh9x1DUPUtkftrlJ0eGH/O/xB1MmnAYi2jXuGz7eK2
nxYE2LceWlcA6SGcvbNAXSXDogN5XzxCmMZ0ZNAqb4SJFt+tBVpfkyFAxd4Q322C
uU3SYaIVo/dvM/Ai/KsQkZlYh/Lj4Ck3R5dOAfbL8+eGMKZietYlsUYHucEir2KY
joQM/VC9Gr4I18GjwRB6TjIuIcxSrVe1suO3OxgX9HiND6gJB7iz+jHEuJUBLy34
dIL+JBmeipSwiB9/eKx1mWfHElvOYqoZ+1UEALga9F0lIqGmxHscQz2WZlrhk506
B64wunSj0ERu74F8Iv1LYcGBlEljkPn9j9jXQCZbaZUmxwqhAsImXCv6hCnuRFeD
SAPYXH5j0uPQNe4ZqSvbf9cjWlkbLkaPcwLB5ywGDk4LQvAbAhLunnVa2NUwz+co
7opH3VB7BB2JzYr7kMef8lVbkRvte9LMJMUwBCgeZRl46qnmfUhC9ZRisjUSz03f
X4E0H3eLKM637dHelhv36CUso7nTsKcgebMlAqKYqg1hTGTEMIFjYqPM3X7641Tj
P+g7hfz9Rxkb9R1Eq5RItcTlJMHGUf9KHb50pcQFw9P10sLP6dzt+Zwu3bZiGII/
zzZA7u3fvS1p6kg13TqBqbq3GS/Y7affPKWPuLSB2OlwR5/IdzujZqzXsTKqKPJP
3MRJjKBTj+0k+Fzg9nD/dQFgiZcGpExVLlNp2h0TA1ddzU2Wg5612o9op1nF4Qin
pGmOViB5RAUMp2iWUY/5ygwdXoJPWPPiTeVlMrUtsBHb5XUoxhDs/ZiZJfmY7dOt
RTanUZxAzZNY/ld4nWmF5iEC9MctQqPoRCy1qpunnbQzlo0kQqk7hBgjww7lewn4
o2R1pIaUNlqWMR7iWqTTbKKkfT/Qm3WCZzqi47D7+ntqQWW5ubzpBJaBTvyKWpzG
LwRQUMoxYdVSzGvVZ7yDehikpFNr0/XjpAltka5gINnxW2S9pYVtf9rn2/5eQ38M
b/14NPIQ8tsPgjjdYFAUYIIWJlFrzm1nP4IXnGXAdoNm4l8CNe0pW1tn53s6LoYD
WTO0Oef0oMxjSmN7PbMAPy0IhKZWyj/CqC8ru6a05llqtUSQaJuR5HMSfusRGtjX
RS36+3m8E6FNI38tiN7BP9Aps1B/elBGlBvKbMlzdVyZvhzfoR7V9PXQJ8AOmeTt
k16GNqY1P11wGOOUCr5MUDPxCKor6D2aNccoXPP6iXCeV144sH1JDV7yqPppO8oq
s/NI2LtV9uZftuieoZZAYT9oQ9imkF4mz7N3phoCKDiNQky03T3zvcZJGAvw4cWb
0iWxM9u+RZLcLgYQMxpGU8P1Y4YJro+/FqCYP4K0cHevXseLXrDQBhbRctpMmm6a
zh5h34jZOnDn9FN1W2Io6o5mAqEp6APIq4OFi/DreqQdmmulhVInR0Lin8NbbhVZ
AUaTujADTZEzTggwnNDKvhoQFXxcYcNIn8SImTVBcBdwBoyBbMQrm2cl0p7vkvx4
jBWsziRJ+Jkthw9HPRxjU0YvCt0c2KaFfUIphfRHnAz4e2zCmlut3ZqYXg3pmFwG
HbauC2rxtx0snM4X000Rf/CoaiKerGMDVGVGSOcTEozInFDcQ0yZ+atd0NAxf35M
uVZHKg6wy2vqZTzPCRI6l5k0LJcbx5AVNygm8oSJaTpszs0uwKIImrywK8mCTEUK
JuR9vFF8v0rNlvXoTwR+GFuAOQ9q2Pj9e+TwEJN2Zm3Fiy+SCCwZQWptzXfsYY0E
/Q5UTkMoMniN6TlJLkH6dhTmow8sJh9xUqHt7fcFzIXQsL8ld/CjWPSYv7WPV0RT
OK+OUp0h+bWCBq/U6Lk5tguDC7ilTWjaNa0bCKzZckHkO2Qp5+gGKt8MYdsS9Vs3
o5lJwPZcJKsDZm8Pd2TaKPwccfLMeknwEg/6tVjsL+E69AlE18t4OKbvETxSfER9
mpFEfoaSnhi+Mp1QU4Zmq71sCmm8Y41HUa2bkvqwANsHGK2WA3a5lrQFLFnhG+CP
Xo3RxDWXSJ9ADJd+TJyPjRy6512JQQ911iCfVfl6CIfhDS5XOoRsukPb8QlH1yKh
WgqFgI6b7tDs40twE1H0mvPCHwG6C88jS8bjtk1fb32GuDFk6DNEqawFMYZXL5HL
htCR8vBVDupGg3PZMkarf+qRtmK8wMI27Am68WL/OhMmB/+FQBHPfoicXAmzphPm
YJ7glXY4MCvIOHY1BlZJt8Dsq+CLNYnmqgRhO6+yTl2YWj0VScUValc/WD61EhFQ
bHSzEplUmqlUjTLFAL51JmUOsrZbyqP6Bql9wMG2WHJMt2PFa4DWwrZ0awB9hVvg
qpLIrT/nWyMsRj3ucP5uwrWqHN6jmq4Coqe8cCL9TWsNZoEcKx3dIexK03CFDPrN
fkpkCiSzKo3nc/1qJNhYQBTo2GFNPamPpIzG7Wt38K1WhA7WyaFlP5gL0kOXFV5h
I7T3Mk68Kbe6mXtdupVQ8Rd6MFg4NxKl9nJUsbiaS5TO9Yv6SLSWYR0oEf1WJUNz
IIbUPOqvTllnmy0L/j+Xq7e9WAt/6gSWwkOBhENECfqfD1Zso5tdkdqgOSaoSHCd
s0Ci5LVxlliVrYFGqc3kWdtStkEow9gs55eLFkboejDrzojydL3B2gnHRlzlaRGl
+1GFpKeLki45OUv+Lmxsvb0dO+9/uuNGW+g2NqXXnDOUuPT7tBjeGsNkSWn8xfnr
FKhqtHyXZOz1RxOBojtU4Q1P76eDaSc205Bv9Q6UE9teZTNbIxiQPczbnCckbuI6
I2YoKqN5ZHDOe+1J9g+WposNIXmFNirg2Z9xqiSFIV8jeq0TNurKNGAjb/Pab65p
WP6wEI3ZYO0s2MlrADfnuiOBn4YnNsriM22aVQINTfy9xT/CDfxWTue7GiYwqaSP
S42YL6ggKxt5wUBBKOtVE6PULDu+iuNEQZQ5HpmL786DrEK8179VwzwOnKPMcxYG
zuA6izIeBh9AsTADtRpbQV8qNGX56EDHthgHEUWXIoQysMlumuUJBpuK2WVPvnfh
y0ASglF/4RSmuLjXd0c7jHTgkrr3zFU1mH88iGijdmNMBdVSiGlIu5rVITV1f8RP
H5GTKire3IzMqW5s844i3jp6hpvoyX9K1OhI//u3f1m7IK/gutfzYOpm8/fQ7vh1
wxOGhXLoCz88rbdFxPFlqfb9nWrW3aZnYJSPQynTJEybtIVhDsvNT4K9AQrFGg+Y
hk2KDCQO2w5Ugf2S7i8hQz4BRh0oEd6ejXHDQdchonINNSrnGjGfVlOfKglJbbO9
eGjkeR28jImmwDPXKLuW41FWBwWwASmBmUQoC3vXnm30hFDKpnXWZS1OfPfugcBm
cPTkvo889PTZf+YDTM+1soQB7lMDQl+XoabXlH2J7jcX7mKttBQoINCNyH8MjbQv
sHJtp04u3NlSaBnOw82aPdbg5YPX+h+bIeKdxmJSLOpYLTOkGplC3nGg0ZL+DMjP
w7ks2VNy099iUNald/+wtCBkJ9TJ772lWDZ1xmE9sMdQsj/mLCsuwKdcbSpB7LCv
wBTGL6GiW94pjdz1rYUo8ycn5D/JCHLZOto102Dx9EP7isyEBjmzuU2qX+NPBDQ2
D4muk7QZs6OSo+1R7PmMt5R6t1M22ZLy6iyKZTlOg+k2/p7q12yLT64lklEIiW/2
PPK/R83lmkQ9LddayeST4Ba/e/8A6Y1Ds8PC9a0cERAC9mjU9ns1DecEp9rYgOKb
G7oI8ojowSd57RUi6aQoWKSx9T/vOV3UY9xqoPnJb7gEwkRMBMuyj4nFtVKfLJqb
JKEl6yBDkUEQBOq6pM6uzYB9mxLnmGIiuJBAHEuFTPNhXezFiLVic+d899hZqy5Z
X6LsUJiKVmQfFuDSNJEy4/1/MMjZegWPYvN3837waNXf5IutUv2wjI2acQggQkNi
IFE9Irr/lt9Ix/JXPbdkf9ClDAFeoDJxijZZ6XWkU8WGDvJaWLUzfPvdFn0CdWp5
b9uDpDds3qd5Jqt8nTV5+d63B9h2mObV9aHPgXOVaoCN0lw8CfFjydoq38pSyGtq
3qBMmRmbQlgRDMZ4zGnFIkeVqib2Grv4hnuwHuuQ8emKISoZag95VwbUYCyK9czi
j89f8dxlX5Nuq+0vl67LH8CyWBUAuLUXthlhl/rVNjZUj4Hw8bPtE+JiZgWCgrLX
/YtEC/uH34G08KPCugFIELc1UJMfsSAWTSSsvFNq6xzZ2/zeohyjUv3YlI99Q/YZ
dX9vvLIy9D2EzXNTauX/JqCmNDJwyyv3q1CU3WHhzhNpQr5ElxouOA3LAfjUzdRy
KJHlXPT81SN2XQm08vVW45mdRTmcjR+Rkq5rvTyoScAo5f8RGu/Xg1gAhWNddMth
HaO8hjQM95znTox7DnvWKA84nVOS6yhgadWgwFnfSvFMuKmKR6B/HlCj0BI8akaD
yq8cBHi7M3T7QETsEfwSTePYYyKzQMT3lZ30eu/5pu+luXt2jJ1agialBo8ROSMO
5RKW7Ck97Pul4bLMsI7CY9m8DQd5UmSgYGUqRN71LQVQcPLPRUqWWAb2K9APgjVe
yU/XvyaQPWCJOJw08obSwZjtXyQXZLu9mrzfKKPITHE1k3+T/DcCQqWib3bz7EQ6
jxanFdd2DqgcTP2z6hmg9vJugrIEtNfnTOHTVyOLIFBYaYZQYq2wu2uzO9vN2NZH
wbBBQWFKoJwvLgPjeZcbztW3omn8svPY5h29Fshx/+i4riiV+2Ym42A4e0zIXe+y
+Y8WNfqe9S46DskjoGcJxVd9oAPvz7InVKYGRT9JCbtCPcECsh6fuMc6RD2od7Z/
0Y3BGgEZSaW2AYeKeHluT7a0wNo/OwNVdQkQKjJqbQjfJtbIVrALFFb8mr/X3RPk
VgCkOlsS6KqxL1w4lG5r2uj75ZHR5XAxo4LHNjogwEZi1TOtZYri2rANz6rEXDJk
/29pMaTyRC8uNiPQbH3L8pS31JBnKviCyVImoFIVWIrH2fxE2qG6m2xRcAD4fIat
DuY5B61kxRuagZ6KTg4qnL7vc8ccMesmeTQjCi3dfx5wbRAjS+A4p4UT0ZuoaZM/
X8jBa9G1cjfbUvMW2/3PtBX5pzkchUShxawlfa14YgddZQNFFLR+wXiJpiEmJ2cP
2fGs1Gmh2KicA3QWgiKvq975YKjOiRrLj44gKGr/k+14PcYiSmMat4X11OBJrZ7O
Ca2NGkN2IGWsbwJy++HYQbHK3GDHld+ljgcZy69bqazDaPiIRe61a1uc8IhWP5C5
vqVNs2Xtj6W8GzCohiGg+9VHIOfEhr16j5kjJuYSy4HYWjJxkUBYEzfJPcGdwNPI
cXOuNJRramrkwLOIUAdGleHCtSYt9dSqL4m1p4OtPUPihX16lq6Fn+qmrKOeRczk
ut2i0T8fQW5QZmhrEAmXwnKGi6jFE2APU6Dn286RKoI4HKo0NkbkoS/0kEqsxBv/
yYoaYtYK9BW7weyfAK+hn9ZZNjO/Njmny/yvoEl6uyyvcXUgvFs99bZj9ejfRd5V
cJwnhf0kNYACBrC86leVaTtpm8T7czV96/Pea5wiHKTTF4Yl1AXVXMETEkCs2FOM
9B2x2FpYmqQ/0pTRsKfrbzZb5n7j5zxk8ZWcfyRBTaxbBPY8/anYZ6IzIq93jsJH
gNu4TGGRAmewu5fxcr4ANUIIYyj3ZLfWFK7KggMI/jfsEAh68n6PSbAtzTAPjiUC
I3f28YW68woDx3tEv3a6wEwQsI75jGjC4mZ/nj2v3lpvWzPVTnIZFMvzCoifc1Te
99rqgHdUq4R1SlQCjf9lP+8ujZAAseZwsclFQVBYDxJ719ZyPnB+/Sh0SKbXMfB+
V0Q9aYcZwVgahem+mmyq9dkPoqH8+89qcpYNrk6c7v2Rcm+JDWSIP8Pm5AvZlNJ/
TFXVk+O0jeB35cPQI17aJjcOiIuI/pSNb0vXXc1Ks40RqmW/YsYnb6XSt97tOY+B
LShRmJhxwBFpQWtos05MHZZH7i8JW6tssfdAGo730WfAibCPF3HmdpijXzSbfYQ9
lS+28D+jB8tvpdMNJ14BkOo2VzEHtQ6qKNonxn9gpsMFrqSr/oSP35wt98HmutRe
t2Huvfh3WeA8On3KQq2ltP0xvjt+2RUPQ4A3kMdqd5i6ZnEQt6p+KE2LxWWRgXLG
Yf4iOerZZMu+/MVTCQ3ev0Pk6khUb2aV0sDlO+n+j6legPGFF7Se2WtCQSISIHCw
Auh/bb4R8LgVU96lYTdRXklK8Uwt24WqvxqRSlF/pDxJ3bbaX6Fs1+SHXEVlncZ7
/byQFxSbaDmXYIMFuB5sQ58WVCOCZhSFf0cK8e5n3gj3ApQ8mRGaTJloexq3MMJV
8UpsBzQExQ6ktYGOA4WOjpWHynhxYGrZKlTkKKdPJKP8op82U1MwCuQSrsl3DdlN
GGz6tY2DiARGH1zMG3Qj6AeZymVs+ZIaE3Ci/+mDGvIU0HgtC+aWtTN6VQuMlm/g
cqNVg41vMnlhpfKsvUPxtCbePvpnflyOmKHPITqHzUSyTDDKVjVY+V9plgmedaBD
02cy6YiPnJWcKs7LF5QGbbcvOwXA0joXohNG5N9b8IxaZFCkChjlEO7Ua14SvyXU
XIBEB2a8Ic7/v+hCdKmmqiWsDqM9fM1CJXSFjDONnq6XtVRshyFio3ozFBtW/Ywb
C0OIcSqsPqM9BN3/2sTu5BWEB5B9Hy5tbz+AT990+XRhrOEQTSztETXEHfbVHWnf
Uc5Q2vKyENZOIOID/bUlaxO1Dt/ltUO0JlFt2ZlP0cjnWZsS3KleycfAAWcw10BE
tJ7U55W8s0MEXcEy8V98wRWcQkiETXFe7cOI8ZHMgDo8DFo2GpPludt4VzlyoVlo
fBnpxpYkbC10eGdOdV+iyRyYMFZJRceXD4PECTrm1yGQ0/bYIsiOSolxKi5UIkif
DJtT6Bdm3V/Th3/F46N5QU8CFPd/S9LW/CtAKKMcRBlEANTHbpaZAWM3ZlPhrEEq
hMfJK/CQcR6DfnKuv++GxU4wRRvKdDer2uUUnEPaiB2Ey2yEcv7e5iOfsArk6T2l
jJQ2s3+rjn9/5BErjqDi3louIMeghvFkNogQlPKYL8+l6JlLq7j1+beDmsLLXOre
joSSER2o9TB8DeZflQ4bTX/QXIV68OvDQtWAAegM8RIPVW7+5fNYXBUkRhlqGzG6
y8nou/dZx8h/XhWbTcvkVeC/jh+udpv5TJUlicP4HfRT8n2nsuoNnx1t77NhDr+B
DkNHAOh3kTcfA9n+YIKl1GHLRYJv4rF9dwZYJhiVuEaGM8xGQPjGpEGyLqzjUCgi
a/BcmjWk1o8JCs9G6JFEdoXMWCmXx6c4wlVJx3qGUYYRtJFavWBQBM09f7o4j3KQ
P2iviaHjJozfGVS4PhyvI397RWDy9wuNLUX+IVDAWlRA7W3XFOaciSdvm6pAyRUs
bL8hZnfo4Qq5eLQh/dU8V55hpD3jDGWh2XzKa9PjezZ9Pct/+TgF4ehb2WnqIji0
HGSCu2ppvIW5wOW7/sA4ywGeQnOFbK4TuvJmslGBEDR+FFC1JA7bxl8zTliEmXq7
zYa1FCmUmxCeMzWA/SxQKoJ7dKm89eMyO3sm5RpEVVO1pFW+iZ2pDgCZCxXaZrCl
MyyMi1343CIQ8wX7g8rRaT+OY9bxNCFOH+q91KH6oqQJxu8FFmQevrtI9fbXVBMQ
wP/qkFjJ5Lk5BBqnMLJjec5Vo52yvFQZLh3d56Zd+zHILlPRs/rufeVU7/ju3v+c
DIiEeIgKYYIs4Wi0eyDTB2zMJW+C5g0oBCMbxvdh8nH8yva3xD9qTC5qcuFNVGSs
9zIbbeO07BRJWThl8RbsUBFEpWLJdhyte1VkS3hqOPo1wNORgrccWgxd5TAxt4fg
+oAwPPzuiBPP/AEMCQMi//Tcz21UWmSYJiUAf1dhC4G9HzrDdDrBRAyuV/WwRSdI
75vNeczjc87/t9ZTt/0nHMmkWZ6AZrCvaJKrAdENvFqDdQnsrpZm9arFO0HOkvjr
P3mbPzM+GTBENhiAoEZleu1jNQEi3uYe6pHva4OY5fV8arD6t4UzvujTX+krpT8j
26BfV3hYVZC6KZJ9WnxUuUq+wPI9+x0eVmT1vA6tPmlds7EadcDy0a+4pxcPMjs+
5G4930WKDv22ThVXR1IkO26awst7wGsc2eGKnGdU6Nccs8pN849iFPjeXOBjf1Xf
ZbYabi03zPe9V3Xe76ND9yT+qFq4AG/ahkY8u7ZPlhR8eq6se/vEqtt5SwqZL8Et
/waECV9JfG0RMbYRQjUHeopjzq4l1IVYa2F1uBIvKZ2b1WJvPYMm410Ibu1XZtJx
va1YqHoYpuy2ZVhuZtouIe0cpJ6d2wdwCBHTfJFq9D5703zoDMmnAfHtu/EFckwW
3qeq1rTwYG9wl0C1P6w8LML5HT8hYG+NxxESCt5ORbfWWWMbl4yaoCptOikZLhpm
tapns9NEC01BWR4mGy0S5Pys6lRBo4AGbYMAt26rmDATstvXLycYSbk8JUc11R4M
WMnrvNmlbWabHkZM+cu97z97LSdPHvwZKMc4Nh760dyHApkNGrBCk9pSEACQZH/e
Hf7j7Ku7qMzT0j9jKTDZf4afj8+qb5blLlfgHTguWFJgmVhPVLOOn6kjia/bkFRp
vGXZxiSZdIxCq7TgREzcoVab9VrbNOtzCUjXgLthl2CprswTkevKMB8MFMNL03aF
CgD16Lq3rfhftO2G78pmKoActjxcoA7GW5txm/VeBrHi/1KYXkxAX0yoMNolyDAK
2mjOV6LLCnCzMxzOPnFbd2xNbYAC+hAwysdvICi5DZXhfWJM+iqO/qwIGGdPkuTr
bWcZukoYTBgQurpYUF7pOYbgaYISO/o0rFgj3HpKEvzkuvYGi/crFBlrUzGnjOSM
LAm0ePB60cSbvzl7yxkVruqQdYhVYwdS4+3s6mvzI8EbWQzKzs6uVqUObX3SIUzt
ILUz0UWMrTjVyav9bYx0fgYkdHSMIJrFmc2b4e6WZezGoHeMF+QUox0Wm5ggQklq
3QqGhJSWoHXnEfMUir6fwIUgZU7HbVNAEaslDqrLx6orLhdBo2cuox/J8YtnIS5c
4Ipdvp8Aq/mNLidEKcw2C6HRrekTcGTZqvep67nbt9lRJzt4xE8aRISEZ0uUO3tB
Tdu32OQHhZSr/gITCv0MteSUtdaa2b3r247ynaMFQdmy3L62bT7IdjMl/P1gcgTO
/N77IVyHxiQP7CcuwL51vGKadn05YXja2jub19MS9H/qkrD+eSezvZXMR5jhHolQ
F+hECv8DqvPH16+B5+EE2S9jRjPLGmKE74diRnwWip/Rq8Q7OpbHM/br2DrOCmOM
3W6fJvWqUkG7yKGvM77p+L81d93JsJzHaOZs2nhZVg7kvDBOa6fHk9SL7176gjHn
bZpj/9yA93Er3XtyXo8VjpGPfe0pwFYea8wCaG1Vc7zTgDnMUXrdKgGIvi1qQFjP
yNovx6YQu5hDu1rRP+HwZ5wUxRU3j2+4cxDqaHEqvB30j3BiYvgKddfJn+7kWdpT
N1aP14QRw+claEiD37uPkP8qV0+1+fIdls1mIEo1n/lxK/nPhtgy0gwREXbWrKbw
ZJ5fDOEpZg/B9e5KWRfmbOyJMyX9EctS06oIvlgfioW4oUiKeq1HG+GCQvYkn03Z
cixZgID/mxhv2bbJpPw6yOmhfMRjAeQbpgTBv552+3/NajHAh6nL5wHUAlhU3Bh4
AlT4zNANgYKxPpjPH+5hYE2aNmNd/F82lnsjmpbDuoM6LTWPvPbVyCYJVor9NGII
5hWEnSHpBdOmIqVL1QgF7ga/VJn8h1nkaezswoAo+8tyt0HVSknSxCgB4XNdbj1G
vT4rbAX9ddOz1UL6lIw9RY80atwV28Vm9ZqcchmfdIJ0W7P3KOfo3nFehkAiShEY
NZryoMHrLH/9f8N6CR/kTRaU1Z26ZJ/jtc4blNCohhNv8H9S+NWl7WgHtPNEl7De
R5+/AaqQmnJo/F0odHxCJM6OeEg1ckkclmlspDZSfxEWAXYKNyjZqQzaBXGJDQ3k
iMG4njLNxRtc69ssHFQJVUyRNVk5GbTxjpEoH0g/Km1h6LW7FZoaoXxjsWk6Iuxo
KHrsDT/qxT43UvaT3NPqLCWP2/Kxzsb38UgaWFb3J17U7lcslnb9aMfAYNN3o0tQ
zqnuz6Jxdcb613Hl3qR7tWithezYE8vqLCsgj20DWWPzf5j33MsKypSIxVbLV79U
ZAQFeMB7GcqMqYubCVCz76dK/RLGtgaTzKAcUOOFfKA1rxVO6RDKpIrnwTuWT4I7
AeX33iGT/0p+ogFJ7jWLH79Z8BjQi5mk+0NYGDo5aSlXXqWv2y9r5hF7bw/tcBUB
Yz6DXbT/ABH0r3P9kjMYuFsSc5r4VwwS7LrBYsaGAbia0QFbBXwQpLwyZn5EYk+o
rh9EempjDcFdUeJQNsDRGkqVoCfCSYv5hJeF7MHgUJqqQwzga83ubL/hDiPd5uY6
FMg8tSuZ0XilY+5CV7fi+oN5xqd6P9+g4PGWrxGtUxVU9l6Ua6FIH/x68ozZlobk
7AxgHYqA1SHxceganr9L2PJYZ5fkxRBskEZitrYc07LfiEqre8Xbjmzhiy6wWkuD
DmXwKqY4Mwzvbex8GokrcDrcrnuXeK193UFNz6I+mgm2vJwkc020EBV7g31msxJS
WfJSQJK6f82nse+xhipIkKEhDV5G67iUrwbvNed9oGOPRMPXKtIDl93+WDpvkR+X
AXmLQVegJ6RWLhnRgksgs9OiNNrHc0rUKyRcd47aadDNnS0U7KUb37xwjyPljxlu
DCWtMja668Dp1pFj+tMWGkwQYyoOZqESCycUPc2fEwrCQRMjRNeXqENgtgX4FWBJ
FuCmt5ZYfVqbSk5jjt2jt9aMkx+Ys3pGCsU0b+DKN2TA7xlwMkJVPreUTJonAueK
jT7Bnnv8y2BsM7fJBoElIcVL72xcM5DGXqhGUu1I4n3TBZKS8zypFUP8sdgStqql
6kgLuPHakKjiuRoFHhAS+Qq6lPNpV2fyTo+V8j/O4+ulXl5Srdy73nWDEFr3YM5B
Er+4g2l28PuDatFdU+5XZIE7O3WvJf4keST/rXa5kGvgLoquUJDlNHjg06YRp8wU
Zc3ydM+Sx1BF3jsi1sIj32wP58s2S4x2lVSyU6KvWDmqMlVyniwvj/xdUK81xERS
NDOZriHkOKW3aAJP+Ttnxi0tI8bhPQmGhsRfvBZrWI0IqhIV25TbBQunlWLDBH8U
Fs7XPVXVO2rJPlyOncZJGZHB7gnqWTOhJOGssw75zvyZjSDSs62/bQe6sR9Ez3Ww
ljaQBtz/ZQvhJL2ze9aqUeYbJIl5Y8FLOps7OTO8tZ/Vxlg9Q/bIRBrFOLuK3sqe
331G0SEGlKaz+r5laJPX2R4peZZzM1quRePuxV5eSprUePS3mF6hvOivVVrazmjd
W/F32TsYkeWTYMDaBWH2L/pV4zSJyiqSq3PQcL+tdNz9t3UGj+wCt3XiZgfQkv9f
v0J76nEcXF3s4WR1Xy4EbygmoluuDk0psxUPfd34gGy/y6YA6T48r51aOiqUDvc6
M1FxDYowLpb0XHcgnhAplYGNIylpsIWTM8idUgsGS6sV7p88oqYPFkVKUe45UXrS
ZL/050UHtiZSat6ZZ56R7tgZ4eO0yOThb3CaIiuZ/Y0RpXJiXyTXuJi2mp8ATaq/
iyrpaninsZW0Icnge2L5QONatJtjCLl3iz2NJvIpmDvXUFalNsbFr1E1uB6tv8GQ
X9kuSoFJB2DTkwfWLuTyTRIrtdAu/Os8W3/xS7jnLWRFqFpORNiI/tqsz82s/a7g
23vI12uTYuqgTEbpaDV3XefTwIg0qnkF21HBPL6qILf+4S6TaRrSMo5ybjhXX+YJ
rz6OazzR6mcKCG8Xt9r4yGSL6iRN494kFNMXMCTgy+koIFlPM0AOlegAxSs9Qgki
IaIGGunbHl+c+zIriEkrsJj/femRl2EQ8i75US5bZprZYxpCDCYtCY8i7Oq72YTK
UGPDybVJUd0dTBT9Y1l6wbpwMd3v583R3t7WcoSKSFnEufEeYLmhB9gI50qIt3W6
krL425qjQH0RlZU8a0jnEreeQ9EZehIGReqmYyilu3VeUD4Z5n+Lemz+zL1KmylS
49i3DElwWk0z5wKyI6tHX0EfVtbJVzKqtXG5Ik23ik79Ro6SPcANGjqq8fare6M7
/wHkhg1LMMLnOJRG2bvxey6GHUkxRgDNaXQ7pcCDYWqmTcuLB6ttuwEKJKC7hXO+
QXTWbYFOqec88FvAJoiZU4CEqaEmvtmfyGEiFEbDWoHNukJVqPkAIkzY1qnv8Q15
aPIxLc6Co8yiQ+g6D58DpkyXS/YkL9AZHhuofpswndn6dtHx6RHs6JNSuFLNGGdw
zX/euD/JJWMNMJkZhuw3ETjtL/lTbXn8tg3jLj96ZfUqel9elT8XCjjxYoQWet5C
Du/Gi338bq45HktSKZ/ThXFrxEWHdMPBdmUPn6xAaONDFdKNCgg8Cb0xlts8AdyC
dRQ9+aaNpA5G2HgobgvFb/tRDG3bV23xyUhNiCaejGanhsJkGjTSJ7X7RsWHgU+3
7nzua1gOvt2BOLZkoJGDxsNWIwBp+8vbHZ8WoP+ZAOZSyoiOGwTlM6Ryko8Nd6Rn
YRayeJ00OncoYy10uh/W1qQSaoQx7yKXQjCT2DWwnucZ66PTHoyCzmFXTdxr+Ora
NE6sJvKpkAH/UlZaiqcx4JnM0sNHsOW1ky9BENgcsfLFUVTvBfd9gVxAgfOl86cS
q8Rs4kzyU+YWVerJCjihWMgUQg9wBkZ8CVWGKbSB+PYeEUK5GHBEKXnSFWOCtjmr
nE/5U2hByt5DeclmYVN/K/QMy6Rosw6PXcmmKQavuJK1RWkhW8GyNRZS6nv3Yjiq
Q0dk7ht6HEOpwJPNyL8ANEKjzmbjB+esvrvXkPWiixETdFvcfhhFhmNBjeE4+zBL
URjtzoak2g7Zr9ru5NPu/KzYBORi1Dveo7ZhhRGh48wAi6rrTPl4LnWCZ858LpCl
Yl4vKqPLVhR7jkfpGJySVngynKKXTIa0mNCwY6jSkUMtpB+43R6lhw98A6EH/d2G
vJTt997qCyz6m/kojJ3R+KwVtNjIQLvzLYRHbP1j+NLpSkwNOM2w5cRKRWweV5Ee
Qe+RNM+mDlnig5yJJQlcyo1sUdD/EiGxbYmDWkXosiJMN/3arWuFvmaayZCYnNC1
NxQHhI52Q0RTKSf80TXs9tiD4CvW6udHsaNEG07X3eOpoD6W30pWB/zjWKgq4DpY
54NMJPKhFIltnG9GoNwWczv+kTphs49Px/n3T7dxHjRehzvKodrNW+c70k3xnAFA
/LfN2Bmmm4VnnQMEfzykEHiZZCCuIZFuHSBDN6dFRIUveC8v1gNdStRfiMotDDeu
p8sGE9peVTVs8mA3ss1RNg1qyrK5WQ2O27BI9o8/2q/omgeiNUmCoBuzX3SPSZ58
Vke5FYDXQgyv+q38xVpTNQ9ECoVGP4PUd477Mfe+o7eIqgzqMbD+tziYHoUbf2FB
2lIa8mpCbH1rBT08OiAbLbcirJd7UzibH1Ac+HWb1K04KhRbsi39L9XJbQcHyU6c
bpKZYBTic62G0W7aMKqGOeHdM7u0WspQTOqifM9IuB8rvS/gtJR5i9mBdGgA8/pk
rIBUK4n5oM107prfshVHtbpQS4LyAEIpkH4PwH8DkP3VMAiMhRsBei0IBpW9PR36
ih0ZU4Qc9qrU3QsZUiH/tIAW6Hlap0dfVFywHlqaoIWmX3Qt6NmjK2LDj31KXGfH
zSnejkVN4JcZwpGmB+EnjAugEnVTEZpC4wsLjbqSDGfglGMvLEnw4nlbyBz4Gjqa
o9VVeVGYm7iust4atDhc8TtlXWZzR5tD5MkjKCUm7E3m0HsB3sO4fdcYp7S/B45O
oxsyTaGj+UcQ2MwKMmuMFyAC22v7h+PwHvcCgu1V1aSw2wjQd1FuPi+RiZVcUpFY
2ZpIaHAcuwWKGR9uuheWDIDXbMOGxjLzq6iO2oYCe34ram9U28kYHyvejkTnKcFa
laugDYKQbF4KH08uhyuobGttGS28rJ4bR67tooxNMOkrgjPGWP4Jolh1V2X5eFC3
TtFc5y+zgbf65PjfEJQI4rZRO4P1UX7wmqKgZNJbEvCUdBIsJPhsIaTGFV15IUTR
zOL8LxK3vZzyQ7OCq36YgGAWUZq185xOo6Et1POxfAB4AccevCzqS5ZZg5k1NeN2
tYPc+lVTWWh98KJ1s7R2zaw4PO0FgMZa3bifkNoDTncAxjLxl6dUuDCfe+GffWUm
0HS8sUJt5CO4v5Anp+iI1YIe3fXPWAuLizSQju8DbaV5wXvmkr8Ylt2Ou3Iw97Lv
4FLCbTZGbjruEuag6UEc5zomXjZHq2Ig0fEpEJOKBcVlVIqQ+OhIPMfLuGxAMSmK
C9Ob82CD2YTuGvcPynj8h3B9dorFKKCZ/gIXrDoS5NHcYmtncI3MQoypABb7IJAy
Rpht4fVLXXKODo9iREJq/lGFTUOy28Rv1QtLwSf4plArcpyObqSipOkGOBRU+ibe
piuyfaSZ0JaRlv34WsuFILlstlgFVZOdBp2ufDgtyzphP/qdVOypsUXTquLMVTXb
6x41CH/krulNNLEXLl08eSkbLz9VvgBnmFD0FYoamupEts2WYJ+jTCd00uwEVkTp
Kq8xBrUFDVfD5zkpsbg59ty69vRJ0FpE5j85ruMePUtEOrE+Youq/v/4On8nB4Mk
+ISb7kQdXulSYWrXwNTLSoxXJwUet/qm0qbK++hsCj6F2nOAKvYm5pe1SNYl7bH9
gRzEw3j/7SY9AtWvcjNQxa3aqsm3fWEwVjWBGlO1V7M7CQOpgZ0+KgzIloikEPb1
8pi7uk2UcFtYDNAkoI4ZA8NMio2K4E9P/c/m24B1IjBScQAgn5sKK06mHaZDx2Z3
iViy3C+iQLTgeH/byTeEqFEOMwOHrvlidJmOvOZwPbcqdH98rqNDPsjrfZFiEGKo
SXZhCmueKfMMfz9Cus4MuDxpaDIiNfYe3ko8dCRbmWZ3Gt8Ux+Im/oWKQS9HakYf
hEKSVTdfZWF2p51ypL1E8VynRH+/biJJIWLMCkqrX3Tl5o1ObSa09SXRl7MnPCXD
5MCV9+uZsOl+kXB/WkfmEf4JqZ/20KW4/VPWhQG+pDK+LUcXfol3yCO/FhoHdmg9
1GPygorhd8DMCAa0utmbaoHy/VhOd8wKt4prQlP2XNJEQyid61cUcoXn0kf8QsB/
WL/S1je1MBVxTVQ82AsSMh6EMsPOyAtSpfHp/7DegRfFKJnk5oqCTYBasHozg/Lx
o7+ie+/SlnQUjROBPbokP7JXYiLeGJr0SQOvjWOrR1HWFWMg8uN8J/IPUJsjUEZZ
TzqiQM3o9KL4Kz9y5vBXyq5eusevgg5Tm3kFlfXP+x6k0rNwrCqqSMilOKqgMrda
Lp9yTIGvRSg3P9DABfQ80UYnRP4C3rDmAcBBY7tU/aWUluXpqt9wi0ie2vUCNOsO
cC5haaEdx+l0ucOCqB3zEd0Lv9K5LKxMUw26YZptMTZQ8XKkv/mJZNHVqt+IddIF
vof8kdS54YMqudL6Vch1c5rlz3hLE58BBI2ICGwJNS1+wlMjO1wHSfSKW1ILec9C
bfYyYuz+Q9grd67k8loWez23p+IUq/g6Zh7V6BDpnwiAhRL6L/sj8DwXU5phHDJr
lH9xT9ObIslLWnU7Cjby2YsQVXHW1MKjR7PaVEyOy90uTMlanx7yoJbllBTOdksn
ReI3w7XEBNPe6VBiRVv7CYj+fw5qfKxOr26Z+MUPXq4IezPfCUVNI5qGZcqOMZTO
VXApagc/i6m6umwhFc3mkoBM+1v1Oy5lWUq72qLFl/o0f5wlsj2XMCJy45sSxgDB
Gy76OFx/Bkt6Xnrynf9GUu/RzoVr9iuoKI+ocSGT90YfLl2jC40A90PYGomiz8WJ
JUPJu0Yk/ZUJ+wTVHUiL8gmDUbcUC2HzMlZA84JGDax7j+ZwhSyRB8HHrT946uWC
Xp0iRiPDzJDC8IYPPTLnwNLF/LnySfbHmbCAhFrGKfk6szFyCTN4lpy70KBmOrGu
FqS3LxzQjNWtWQFfLX8hnFHUHnmob9quIffjh9cr2mseCuiN4xa77U1kTaa4FHMG
BO5cGnvBlywAY53KnITP38FR59IYo3yBIqpM4lXSMjMN7vcpc2Izp0u7f506362o
qaKGoMCcL9sJ79bnUYb9+guDib4u92m3ghi1uRJN5fOcBdNsAx/2P3xSi0ZBUuG7
ylJHSWWaPl/6tSstUWRFi2vKg8d3qTG5M9a1VZXNJul1zE2NAlYQ2ZsHfPumtwCX
7n1cyURVW/5Mr6P1SZQeiF8g8/vIJqnRCxNbTMOZ1QAJtOj9Wsok6Y9yquQaffui
XRFf85h/cTNsy+CsadrvJ+tAWR74s8uNB4j/i4im0k6N9XRWlng3OCBITVLnIAgU
MR21bpQqAd2fbwW0NZ2y9zSNmBzCzrhhtMjk+A+84bMNojz3u/h/9Wy8SBIZBF0f
LfI1FVNAPFS4yVXxB353DO709cqfXrMoytyJ9VwGUHIIr/G9gHsRGBzHj272/Fbo
qbvtcZUniap9R5/QaiQhbqvlcYMKiYDULFg75L1lG2i3n6qc9dtyBIiK9geua3//
+MKu9Z3Gou+Hjao6s548MiQOTPj6wLfl+WdHcQoFLCtmAxQ+jiDKlezZMQL+A/Hu
WGZ4nwpGmhf5IuIYYz+ozMC/dJ2Y9+e+lNkdK9eLE70Osb4QOLHGSeSZct5KkYS+
C4uUp4Jbkbl6qYJTVe7gx0ih85Ba8HMqv9y7/k9mCmVO5cKjWqDLsBe+/55c6HlS
OsEK6H8xWfwl751ZjWVr/MuoU9UecRaUgYzYC09uH2OQs3NRL7G/Bg7qFCA+Jzu8
RW8bRhAObE6OeJePUvYaO9+rzaQig25d4jEPK6vIidOv0TBVLoUOLJlHpxJh0CRj
FLDqhClVuQi0oqF3Fp5WzvLyQyVJGyGat1MxHJApbBhNd2yzlrd1sCgP7RJmB7oO
CI342fCVUGZ4ZW4QV2CWVyi7V/OdyOJ64SwoS7ExZZ6jXPNOgYkOx5ymgeBDlziy
3DAWGZGr13N0GAI5+h3DrTD7B9Ew5e+Kb7iuL0DpOL1ldHPIwVZXVPRuCfVS0tbF
HxFAHKZ6booOb7gIV6m/CS7R1fLuOfdthlvq+WmMZzEXUPNI06I+KdIW5UzMPgk0
8exFbm/lNAUgld84K/wTgXtU5oIcCreTaumoTBIAvWoRjN7b5bI9GvoF1SpRRArP
voYXKdwYNbEd8YZfpwYX57YUDWQzrq7++EPXpA04RafKfwaQKm1FpSYPq4dx54S2
5YcsjZ+FGabz0U8naOcojVi5xbKgJfhjzXLAW7YzeVQbq1qSBQUbl/Duc9MVdV4r
csbbgwfuzjK5vaFEMS1UrO+3ACvQGKiTxJkPA4NZODSP5yNoZIkfv9/YVbSLwGzu
h9Kw4KT1JkQI3vFtxcq4j0LG9b0z+HV+qMWjRLDy0FGomgFenHYP2D8C0rEurI7D
tf1vzedBbMLfzzlg7+LuxRHB2W460gM6kS/kbmScF+7RvN1m0hpeVy8sakM79qX5
j1viM+nHtlwSYlE16SJKvhMeqY3h62yYSwNaT3+lFjcUR8prD970PxpaoXYWvCF/
t5xRL5gsYAh33MUsKmO0KCu+XZat1eT91iHtjiAifgAkeVDF6yI8NHyWSM9ViMWM
GCmQeE9NGA4pYEtjSTjM0fqnCu/y/HUu5hEUriXPVg2GyDdOm0G+/BYfTY5DY4zh
ElqkkNsCpTDRUW5CzAZAwk9d1fs+6Qlogg2f61gUWqaq0ffDZf+3lyn0+UiE/OsJ
6odT9bnWyb89vaMheXBYZ0GzCItSCu84PwFtkc9tqXR+I2O/4sFxeveQh4FGDxsf
UkQeqFOCNzUPrhotXDXGu2UjHIYYICwdFvzV7VUYz5VhsPHRWAqLn6vMtn0kIc1b
RfDh/YIjunC+9mQpXO+Uf+dX915HQYN/9uEqA0s2e+P183R7vKSAbflDAyo7CoYP
RcWn/5fzsUPHMEZtZDehCrqOWt2V9yreJ/dYX4y3naEDdqsd+FSD20Rzqo60ekFA
dhNZ0llPdv7jWpuFMP1wnfOkZ14KThRqyK0LHE9wE2cp7dO0tFMYfJWV7iwId1ki
Bz+FRvG3wGUxtgjoxpdHn7MrGJVluhoCg5z4wmBt+FtKWNIYeh449tedsi7pRptO
MW31VC0ciLRf6mRWUKWI0vNIpeaGtHXtMGfSw3u615EsTNfJMNHToP0L8DyodP0W
M+hiFxjbVMG5/me/ZpyYZ/CX0S1F6kl75VSvAFQ9zGtbvXpk4F8RWVE324iRSZcW
rOo8aGKANIZnXtGaOkx6X1+oqN5Z9kMo5BS7Ub5xa6HXKA1U36QzqRAB3hPX+FWD
/vZSjytESfEDHaaQ2kPtKCy9qKeeBy2VURhvZNbD6xQJoYd0+jDSOfFVvI4xjOW1
ywRptRysg15PUhgAaZYJmJyMO/kVcEarfwqOGIItuTQ4aNYFayy2dGx1gXigOc9B
SPpxn91aDXYq1xknE+xykDMYB2eZJU10yhyu5WANLf6Y4XRLPV+Zdi1wvXOH8VgZ
9O/FapVXwg/55WXCaJX8gNi00DsiyoNwPBkcy62j5x0u7CeJiiZjxiDGNnsY0Nco
3eTNWzQ93eJ9eA2TIX2aOe9x+MypjQw1sCMkx2vJTlp1l0pEu4iD1y0aNQ0afJ9Q
eGmSKCURzn/d4fIdhxhu7EqvrbJMJHEXruSfhdLAer7nuJ2iEdcH7lT7qngmRRix
jKsdJfSPlXqFHSdIdqJADq50LMX1OvsQWK0jqPb9/NP4ZEWhsktmwPs6wPmMSkVR
og/sI1maMEHQJXvWKI8If1GmZJv6XTdXzNkaDkRem6/SmLaLCDK4uUN/trHvEg/6
KMT7APc2p4rfKMkWdWIHjsgYRPbdggoUrzcrZdSXdHzvGds70WsU8WmvT+mz0YnT
TWwADta0edBOlYB6UnRXX0jdKobtmSc+aAh5zFyZ4SWtQ6gnPoGDAxeb0SSuAFBh
SjNPTHYsnOPfpm3Kyo2AaRLst/mYDGGCz/vlvibwJyuf3g5rIJNZ2E1L/ALBwAcC
0PLUsLtuG+DkctnC5MQAEBYVejmys2DNYMOGG6BFiWMFmaQOAVlz2XYRA301ol6S
iGWdEH2O+WKJ77CLwsSfBu9PbDcmWe7SuEv9uNVrjJkQAd53O3EZjjXeAA8LZhE+
pbVLKLiVkAveP0LNDy/5xHc9RKpmMP3YVoNsOyXkHeeZ7XyHG9vnVEg6mShln7g7
H0xrjK90u733Cyg3HulPHGNZQ/cU7ZTuQAYflB/+ZBZpj4bxRC3Yfejd+FFJH10e
qaLCzGQz2FDBmE7K7Y2JT2xVY0NqKTP0S2piF95Wg2Dxe1IB+BbCsKJAZd6jEoAR
tR92Nc68AN8ukgo3X05iKjE1sfNhcBqKhryi+CUqpHC0iBhkOA8V6FFwZDsCSRrd
x9rnL+A9CA2n6/L7v16j9WorHgR04sqlIJmb8GmE/OtQby9izRm1blouplV89+mZ
NBCVfaoTqWpp7uJVxnl/4uzwo3q3tE3EV7E60v8qeY/+mf2y3r/f1deglKwgV0k7
i/zKR8h8UhOziMMHsTgiuRIyN8GmQuPsz8e26Q+k+7p+MVD4Kq5OsTMcWsBAUGoY
uaKZ2PPgb0MrHPTFMuNq7wswKapvkDqor4J1NE7DunfEq1u0saPFN9KujQYop6n/
sf7ePydREZASF3ozZdE1dZKuzfkVoFjQGP4DN9IV2V3o49WiUpopYE44lcSEDMjP
5HjSCv+cNN/nCDNeMlbtdbzkg0Gorih2pnGD5dUIuautRG3zv9+Z4691CMz0Oh91
4XMp4fHMKtk1cEf7CuExy2fKuq11Y9Wg+32FJAFGCjgq3M2btyABy4WNCgE4do45
LE39IW/Aw5y/94UmewbdL2h5tFTQcgXCnkpkbAimVz2inlklfU7QR7Eel7z7G/PH
kDdXVHUShC2nl1700e9DifhL4vUsEgw6/kYEf6O5sbnZ27o/3iny9ZoujFsj7Zsf
w/A8ky0nuwYQRJqvOfEkxRIrze7H0xiSG1kMyW3FFF5MlHfblyGK5zAgmVFNp5OI
81iWgK6iSB2V4xyHmUvIF2PegMLWvaFA6GUKlOxX43ziP3LZJ98BNnkxoZ7rqn4j
qkfYhH3dMguNF72Srk3eeSiabKFuNBw3ICvoELwWWsD4kG6m6wh49tALZJaTJZpa
gCKvZkFbXW6PR6Aq6HMnetlu+UUnuvfQ86A/27P9X/YhC7bl3t4FYNrteT4/53tO
tUo6WAvxTp45huPPfjrdB5Lc47nPJ1mLmzi3ypQVG1cK7D8QoavwdlZ/TYJ/PcoA
rCJetK88ZurAGPFHCC1OFT8QZt9cTKgyLKZrO6S6356Z5A8DV+40JwxL1J4lEXIb
qEHt+YnbfsYoU967bQf2JiIaGUUR4P9sh5hBxVbn0ijiSOz9cc+svVsv5kT14EOj
z8QKNAUDPuaD0AmIUGJoYO8tvXm57NW+M6aad9aIoQ0amMnusO9F6PyIsU1CsGbi
deOke38g6ucfkhnP9EBUD81Eb6GaoOm2ei/DK6sfQFUY9RCm4xFBN3h4p+T+mrML
ENn/kvGZplK/UZqks45ZyeXxt41TBfuH7whf5PccBJXYRAZn5WyPFRjIxRyxMnJr
lXcptYMBRFv8L7K4YpM3grvtwppmjIFD+zSVaU3lO89/zTum8uQbtmTgeMNPoPYn
xkBQL8LFsBR368M7ohRl+bp/gQh8fIIJwIIew8OTqvHqQfWodOSp2BccvFQC9WEN
i+XZEMlHcBGak/gOZZpZeqTasdRa2jnCUNLxWz2w36OZfRSdflsMYPMvWpGMrTNF
B57/BLjvjvtMdG2GuyRMSEoYU5SaqLqXArU82SBz0ry9z3374CC7hPpYTYM5LlnG
Sw8IxekQrOmu9uFCfZZ3p+sBB1jQ3utnWSqc5XUZp5HZBlg2+1b58eOUqXo+czuO
VeekXKgI/OM6Rr3vTvApvdjOgNfEzQJjXThKIjMrUaK0ctoh0QcgNw1qG4JF03L2
NJrEH7D/u/CqUZL5EZa7NMsgvLHkzKqZvXLWSij10czWcHANl9GKGcw8YQ8w6mTK
8aZARYzVwtdM9AmgqFJa/sO9G9fKLbWJCefkDB5OC06UAleEROQ6wl3opRZlp7Qn
pFK6ydaHuNxwJfGW8xKjYu+kgw6fZ6LBUXqy5NvbGEiRQfYWQPPTOIYwoQCr9I6A
RchcGqsXtSGMNdqdYR9w822r82zmy6wA6WxLKfq+ZNx9otuSoDcDwxFESe+peMNP
tv+Jgxuq51AAdqM2gP3lsU4UkGyGUyUTI46ikEaLtHmgsJgKO6VXP3vfekjndmCj
s6kGl+OaWZf6Lw2T5d8k8xowGzPgoJwK9dkKBwKLxVPyjFCUClMtcZLGeEjz5Hmk
gHTO6Gb0WgAjlXAECZpuII7RfYEcfDlABNgD7nbN/an61zjqi179yzDUf2aTsFdM
rxoQdHHQ0EH6+4iPCR6UJa/2FMHTTmPYUbLokFb4VL0UPrgukYVvgQsyUW5s//+N
+wgWFtxmbOamgpBN9b8+gswnFi1OPYaffh16xb6KZwOYFnBVJwRaIs9h16TxTDoQ
8qCRTcC70ys/xv0P/MUuoEaC5yEp63NXZ2Qh2TV2nzWw9tJuNtdx5vyHvh7DPW4g
pdyaUqgFkjss3PAVux7qKV2tUPlB4vsrArR8FevMyF9iFBQz0CeKsYkfHk+O6SBE
VcNcILYbXJzDXXZ0zrQJbYsyl67L5xqFz8VqFto6f0kgJzvhJgnMYRUalApFeRIx
IhOkNHeFKbmGkEOddmkv+58RaWnRy0kNyJ91nx0lkDV22LImgF9GwlAzOHDonPD2
TKVqKgzKNO50piupfTEIHLu6w+uuOpDpwEJYZjb/aMMktmBYIfhjxJWZX6FiMRiN
Nz+mjRoeIW1QbXxErEJB7YvSMGlTn6j1iUuNXZIU3O2O5Zwc1zmclUxcqywX5kaP
0biia1LtFJVxbuku9UincpYRm9yakseYogB30E89OHXSor1JI5LPK8uX0gSbhu6b
27fSjHsWPRyg7dHHm1u93B48igN28sMpjdbcqGdqQJPZQtwBdGd49YSbjJad0WlM
RCvSXH8ahPdRQ3t3gIJdWdzp9Hdi96LUNbe4jUo1CQDTn/G/6o54DooM9hFSg/wv
9MWJsUU/UU0CsFFDtpuKhh61LIwa1xYnVUot9QzVtS3VjSLABU8BW5LD2mxAg68q
ZIks878gopTRAwpZFrFv9/dbbAmA4je1A7dTBopohp5tPZrX9bShp5oVow34Lz38
qk7PjyXHYoB2ru7uv9qKmfCwFijd7ND3iok5f+Cg87I37oEEcd0quyUedbns4ILy
qIQ7VnqNj5+PcJTQBbf0/p/Q4FWxD1qLnuPEFfvQxIUyo6JD/sKHVXDizEkuNjgs
xxhASVaNWwKMF02K7n8DhFSjei123uH2yRd3O8kjKHxP9ULeIfifly+MGGNU5MEu
a2qPwdUVTxkRZJrKKOqaJXKzoGnMGfOZ2A16khoXoyFu71dvHAOImkAgHhz34JQt
dj6jmIkNE3uTbraPE1t+Ex8pgHxFR7kq2eUpbtQ6i/4GOgaMAAbwryszvnfaX584
m+fob/lLeyLIqX6i8I97sfoN0ubrNaDMXlEmonyvpT5cxHWWZfNdD6KVnQONoN1v
GAYQhnuneAo6Y0QtoNOvYFnmttQbMeEMZAf0ywRSMeEpA9NajOBdodhofQerdAFD
RdbIN6sHzmGrcOgoXAXGCOF9PFxlM2KtUqQAef3WZH/4QQcpmVVjoLdn2oH7ur9H
jxcoUpcz7kxvanmK9+lH9cRIdMbq0i3xmMzj37IDs0dvN/emCUvwa1N0UcsjN1e6
VVB0e9ez1BYGaxz8basM+5mLcR0yt3p54fhnoFPi0l8SAOPAwAcosZ5vgKxyage3
icuqhRJbGAOgiUcroRgZoZjb1tAOzV0gyjU9guzHnvoeAz9ftzshR8fEkt87jApF
3/rshtNfjJZ9gHxOHrDwPEcCut4wWm5/9l17PXR5jUwcDgTKg03X0YSB62bb8Vwv
4/NZOzvllYcoiaSRP4Ielxqm/zoW+ZWVfPrUJs9v2AOQbjlPpsG1zny48KG9DOuC
aiUZNI8JRmbdwMZCFGPrImLzPqBsOtIlxrvt5bzDq7RC2+NhWYsHzadULL9pOC3Y
9Ihs0ho2MSp4y4YpSjRWTld2PQFgKJXTMmQYf7GyKV6ligzMhmroYeXHng/rLjfy
MYE1SSQVa40ETQkmtZ85TWVlkMONuENcJGLkAYFWDgq9UTWBZDPXsX9Yk/+HcqX0
m+o35iqa4jfpe3iTb62Jq9EjVCvkY0L/d0dB5iAjmbJzFzWkErIIEywQ1cUa5Ajt
9ZAO/91njpz1KnILgUC7Z9Jn+jrrLLgAZO5VqGQN0I+YntJZI2SbQ2POZ9gLMJp5
N6odkRKAyAQY6iXAZSyrew68JDbaKTfPWpalvqz8yrRpaZ/QdzrGGPk3JJzC9tBn
M5gyKeR3Mm+LEfyxsa/l1BwDuYGGKb/YXk28M132IuATEYP3pdQwFOHy/QyaLvx7
hf1JCdjDp+Y4IFn2KddMmR7+XE9WwKSdOfuLNxsaKBJEe0c/nyYzxX7FSIcgB754
xz8rMsMS92D9PiFefe4BWCXROIetSc2ZpfI5LiFCEiVOhSBns6PCo8frOUgEKmu8
RpkLG08M3mxFY6dCvHT9zPppg/Ia+5zARxzG9TKtocYdI86L91W+XzvHjj9IIvwZ
KNdGYca+O1XRC4wZd4kC/sd0vnoEiqzEP67yQdKMwZeK3zv5RAMbyKkQVEJ+nrX8
GRT+3uWU4+ym5GdCmWheVa7erJ21ZbbOW3YaYQr7DSHuqrnlaR0lv8oSzbq3CQ5+
Ec7gpWoafbjou+Ktf2UBeqmv9a03OjJKbbiJvaVQOzWzgRv4wCpNZKiwByzt1oLA
FnblX8tvVTnZzVPpWVU8Szky9OnMQ47ZLgpMhzkwwfuloROsN1lZxQzzEUR2t8fv
IQ7/lR7p+R3kPyt9ToIH/Jo0yYegrHfiAGemK1k2V9/RbWr89HLp4xKT7O8Xnnf0
ITgxzd0uNKaMeUk/bU5eAnChBxoBCXlCG2EvZ8x77bCki7fO5iqH1rWvTVnqcTSp
2MbbgjVKGlAlr6ubQ+koUQkA2YG7bTusNz5FMivMh6wQbls9p8+QEUXUShR0rUo8
tT0B6BXE37NRk1c0DB/98OYT0ay60QNVxzEF4pR7q3J7/ZLtMf+0HR3xe7OO1Qk0
/qMK55QYbR210ioT20NW0TGJm5SPf/Z22vRyLqEwPO+zOiChiFEw1+arYiUDQK18
SUcAm5HHVJJe+1yKIoNoUk4T8Lpum2laLdbS3fK/f+KX257SjW3JHgEKU8B7jTR4
gXlEly74MKeX40ahgljbuGqpC34ElkDGBcRYkfdsVNWrKDbhumEhAVIJrDH96zU9
rHF3PZzQQ21bsDaeyCyEpUSvWzfb1QpHt7LTxTnnp8bn4lO7CB1oB37RISDSpxEb
hRdv+N6GguIl6/hHe0G/us8ryuMHj/W3gRAYd/GJ/TlJrYnZMo9/5zLurHIf/x0d
Jl3tTvXl0LyrFehCQEYf6t29sWBzQmxZeRTOWA+puTvCKcH6WsdfHksjiXlzssGn
WqbOQ207KVoJLjPI+VuxRbCEXbcfuo5IBRam2iXFoQMSGStwReDHVGgd3kIANRra
NCGS4tNynfWS8bgoKyd8aZ+tYg8CbVmMMlHES3EkuJ10WC5BEK/6Uhsx5WvBHAVA
PhDqVawpV5pSk4sqYq8nvb80HPDEDVZUaUgXiGyvNpi4hEvCy0SD8IJMtgeDUsfT
b50DYz88aOMF0x8dZJOVX0m5LXkqpK1TyQ3V2XWvo3mwhWxTuMurrXsa/zV+3M6O
dvAdm1Oi1ajSWwjxMWSL0Hs0HjOw9YqJJtI29e6IUOeFCeRLYEugiLSz/4JfDiL/
zUI65QUqmd8UYUul/E5zW/448b2gWkyAx9mnms4UX564MiCFlpNqJ4Q8aJ/14ZQd
uSJrWFVvCC8TM8mtLP7ZD+0gDbvzqorqnUFkOHrav79BFJ8LbiDsYzoH+cO3ctP2
riMCxOyTPsmKp7x0arPkEwHV6cLK/BSxwRGm69I/63KO2ia8cwPNzZRs479OafPi
sCj9oXw40NM+toB+WJ08zH7mjel2xhU95nhHxVXSQX00mQvF4cAWN+AK2UwXCspV
k4WivMEa8/fJE06Ru2cO6efyZSrtrR8GUhTXXeqH8p5YgtbL4VGoMj++4Kp6DT4d
i15dvxKd3xHBn5oPXIOJe1ueqMkgR+eaL0f/DiGfW2Mf86AGOaXB3eMGZXcnD8hZ
uBNNbnpD0oQIpNpOWzfjTlgfWUxPAXwszdrhhn+PbgCuQdZWhDYb8AufzmpXqlY5
vxl5cGCBgy0rqzAaU5yzgXAly4zWeJlmKshMaVZekPuVi97DsrDkrELAU0JJZW7b
DwBtRqLEWaNS39u/q6jNCgx8nfpcAL+O9tBsrKc/gsl+2YuUjjDIqX3DuLjX65Lf
nQ9f1TKELGUrJrsenUqTeVcU7vIgBmb2Q5nPh4SeXq+6IJo+EcX8KKwdWalJjOak
V/VqYXDiRoRsYS1WmYWfSPs6ElZrXq5BTSFHxZmtJFEyzweJd4Bm5xVG12RdYpwE
pPfahJTL6xpZR+lbvscNkG+kE+8drYsg3fY82iJj7XoNWAhGtwVkaEi1zSM37fAU
Gn8hsYrla1mDjF8XSia2Uq7Bl8DhduG7WTT80+ycAuVjyoALtQGkU1MTrVrNbLpq
AValIxCn7xXi3GMpBzgM+i7sRAWc0m4/+4YR4/irDoEMNNKYQ7yBGXor2fDZgZi2
bOe9NpN15MaTuydraOsi++fyrmghY+2DQL0IY0IRKZff9akyEfD91DiGUGvxFt1j
gI03FEm8gWtap8+Pz7TPu/FUB7elnn4hW3aIrf+uV8/D5QY0DEzMhZORX0YJakN4
DzpUzLBsMlimN0FLkNFkTcPjCLAAFcJwvLIOa3tegkgmtTFxTladOz82ojfNvR8T
tXwd7mNvtOW1yRqpJYeQQ1obY8XSz8svwIU9xegQQ1IdivddtDMyMgSkXBdhcWCP
YMiAJSSuVRQXZSWKY5eG1U0A7tXMzs7S51NiNelLKq1ve4J8W8vW6nqd3Gs1SK+l
NIoQ+Zsk8hnfgMOjnh8eFR6duJgaKKkUse+V/Ew6jlH7TVji3pKcHPSpe156nak7
y6xeZqBxd7iOleq9/uzg75em7paFRpzj5ic1ANj8vkfwRPt7DGG2d47fmOTrfOnv
XZ+CofYtbZEHHjGlbHLN02OTNLtGkSp4PEo8Po3QzBgO9jvzHa+UedaeQRcDVnQZ
TBo0xt6oRswra6XxspHzyp5bvgvaOYRWlVy6nYcsCALA4HBNfQKeZO9RxN5FaB36
N60f9/1z9rDas3r9OoK4m0JWJjtuQGJzvawBDTegDxvWV5ma5HUX1FIAAriv7sFq
/svbOqa3/O8k2mWaHuve0Q9gzJfgwX/NxU3GY0xaWEHPdU1zxhzgRHetQaxB4fYR
lwPFGb230n7g+Hs8ZydaV6xzLsWAzEL2sZYCaHM94pn+YwNudxgzsfRBcVXxLC8X
BXRfabwSyRKD+t7Qtiq0Kurxm9Xz489dQVxhPpaExULLgSKp02AMZRo9GYpdslQK
QeDGDZocuBTQRlxstCAmEjh7IhqdQYgAZyecGVT+9RM+a810vabe/QZEZigGbjiL
oW/DDJB6Z8m2y2dJbQBa0xesmQg7hejB6bc5zsuRqRU7QyZlY0YonVjj9Wp1z37/
dX0C9ya9dSN7erQXKPWP1ifMdm+gx3rRoYyn5toTuhrNuLd5Qd5kkSKgZsobwKsJ
s77b8tC9x8P5DI1+B7ReiSQ341keGzmWCtlyvqh2WfBSUJqruTWca3TuUpV9h3TL
ubunLbpksAxfkhKTLKMYlUMwSynU4wzamVDr8D10hJjVPa1OQzX1KP/VO6WyVhHO
hAVzGEzDgkVGqMyxaHKoIBuDRE4pUi3VnIx3Y6UqlCqzcgz3okxjg1f2NIIpobbz
nIbPplJDllKiDn1s64b/6g8JF30BNa3TOjEO7OXVhdcppsdpL0unMVhNEZrPIPT/
hwaWgxLDSkacCqwPe5wNhwPXXSWDBoOUWQee+3Wewns6uZqSIqdXh5sIcb9fZJoB
zJcCeScLj4h+NnzLFjgTNodtOMoqRSNRSXeCX4HctKaMRBpZ1SXO/rDvyHqovkAj
0iJs0FLgl/lu0jNcFGILSsvViokx9Gf6hbadViwctM4i9Sn6qm66AkgGSSpTMhqq
WHaYUA+8HUBoHgeS9Eeb4Z6KhDgBB7xukEY+OEiQRLNCiuY37owzoDXQHAWr9POB
wmW7rvxcR5F2bIap20jJnxp92ELRN+mMy7ZSAwD7TdrxM35ZJmR2MKyvW22OcWP1
qASDunh87kWlwF9bnEsSGUORJOX2i05LeO9V4f4Rq9mA2zuSvs9y64IMSojNnrJW
mLETXXVb28qQJkjZXr19eHBMk+w21830v8joEjY71PR2EQNRl5i9KMcR2bigb/JV
0hYINGtbCGIhZfDYvgdk3hYnSeJL3WfnJpf9jdz6pWL6O4wAzhOAani1n8/9AGwb
l5XdSXnMQWN4/91Y3FZGe4sH9d+LJBF6zVpCEDaVrn0knpqcUlvNG+MO3lAnIR2z
x898WYIYtuoH3yPvbPK848DTcrs0NDOC5wzWZx+QW5fTIcCbitsyNBIyOYiylQka
TZFsPtdV+RaC5/88Qg9xzJwzS29kUNhOPI8aMeE15ODwZzmH0tgf5YEo7smuiUZe
+iZgiyjeJMDVm3FTHRfsIm+hP/r801uwbZ2oItXZscUbbdHISm9p/tFU50ZM5ymu
UPIyHTaU8+y1COdr+cA0nn9GgwW9fic3L1vEWASgkks8pr6tEWG8VP4V/j1m9Lzy
bPo2BW4FcCNfZSuIaFhzsbzVVIMLz9dKGFq82TkwVg7nFa0JttdamOtHsPNBhEey
voLfGaFAuvoe9BcwYml/7RO0dXSb2/+A2NQTJoQmSDwwtNopOyzc+V37by2trxJ3
jyAy9HvqeCKgKFpuyd7nPMkf/8gf/sqcXgZeSaqpikiP8tegZGcjd6nEW/QKF92z
YQ0xI35WxF5hExEd0spcXxY/GMcHVA2/pRFKRZrr3o7mIwYAPK6Hr0PkuD4eaopD
d6EfI/+0Rvsk6vdAsZf/056OZHv8xuPXFEI0oubHd8J2MWTbOJ7yg+EabgoyUiJ2
Rc97ecobkJ//XxAByE+TcPbt2cCG6dazcPbByfA3SNHZWMSMVy2DqpsW3WtK7WHT
GFpYYBq4n5+aDIR9Fvc7DM7v2O6XcjGA4kD5NAm5WS/TS639Nmz/9cbV2rpcl0BO
gTt3nNXRC3kAi4lCJ127ZXEm/8s4CzFnEB9QYIXF3SxP8+ONBEsUbeDi4q8foRTU
3MAhTfgP4LDzRUexRyi1ZvfbhzdcqVb7cp4siHPSfcPSz174Q8OOLMqxHv7qV5vo
Bx15Zkoqn7Dmz6smFYG6rTDI7SQgsZwZuJN+UlXadx0e1OYjBbZMOOZdvkCi//36
oLS78d9BXa0onvCgZ0FYTmtLjDVKY9+59JJFghoW/+N176PlqWiwFNv2c872mdKg
xx9W5raNZEqZGpgi53rKKQaMRZlks9vVXv87Xb32otj1GGeTSHAhd1NGXki0uCBN
TvJAMIoin1VBBlPhoYIxWz64G4+GQXMMuramgJ9SUuRtQ1H6AKxMD/HU/AdqA2mp
FTEUFgDIOiTbxb2L1a5gcWsFFhtBgqDUj4xwEiYQrwUZDYB+kZ+bHAw45Kd8qtcn
bnhoUiLOMT8hGrT5WP0BW/GJrkWjjqA6lqGcPycrwuqlU6UiV4rRR7ISSjPj9oV+
RKR+pRPsoxLn96ydfTcnCCNZHYHVl4TU37UMdddX05Ktg2ZDj81UsmqN1fwoepHk
S1dgBQOIKUkKfv1zHpzCaMMBbJD0P0UVUVnCF/GhbIYUl8+E4qE8GjYghChoNn2m
xw9N8KIsKmCPymi4sUXIBBCvGDevU49ZAwEKdHWxNTo7bTk3JxqvWFrRvUmrdUeV
P+lREv1g0IktzvFl99q81Mkx9cfQUnxBM3AXvDQ1POC/GvrbcMU0GHLNNIdPlGcx
OQtQAFwy4Q9wQEqHxXDXPh564YdPWW+dLncauaK0K62bu8B1GLYnFWJMsKaaTvTJ
MUhOrjj52mEYnuZMF4F+RAXT3mnC3AZ780dCLY6t8VKYbb2jCPQCIyfufrtip26V
GP7KfMolc1jD/kpr14YBQLRiYiN3BNXpJDEEwnkRp5LOjVkWApzXQLFW6mfyXER2
Rzjfh5d2Fodx2I6dstR07A0Ow4xEDHdLl6cjYIy2lqU8O1HdZmdGC+bu5nYzInT1
wyqTWBpHs1iLPR1h87la0GznQTeocqY2r2FhHQS4X81U/YiCfH6JE06vNTJbd2z9
85l57ryuyQ+tsto9K65uH9pGhuZKWnbPm+rZcGXCd0w7i7jbd852UZhOypGwdODD
GwlOL/yVxmGxEGmQ1EtgAXCM99otTlHShwPk7g6CLZhT0Dx0WUQdwVhcMq7oUdzy
d1R7JNKTyRVYfDMpoMpgc0XI2iULIVpGINRPE66Rst66mUOI/GiPZnqs8OprqnCv
C7182k5nuKYBGtGY1ThycSOMl6/fXqBukYLo1HZEYCtNEVG/ioLWXcvmjnmNJqwL
/P0K1/6xN4LqA4Rx1A4JAX26cW+D1Y6D9O56Vgl4Ecu1nwtHk2ms60J7pTYLKc/o
Z6Kah27N6zylHLgrqN6Kf/glNOUx8+r3AWdqI0JCUR7pAiEpAFBC6oRSyhM2qsoH
PbUMMxWtucbckHvQu6vjLNphlDi2ys1RkBLLz3I6mXfMpK42cbcotYyICbxlnpMb
NkONm80RIu5l7XD1bs3FTbgGr43dEia/NQ44y+ITmM/V8vwBciTRuUY8u9NlQI1k
g1Hpzb/o8WOQGpb0A6HCu/73oCTMTpI20LsXRENvYbKUdEyWyxk2T2CV/4cAeeTe
pUxAYc2RTcOMdSICS8Dducax5BJJHQFsdRvBNV9gS8B5/EeRVdXcC8Ice/YgEygQ
6yVxPatjLorLM123jiuJMYpRzEfrQHimooCyHfQ6bBOuU36+xAtbmbffV+0+eWwk
9tozFaERTfHWEiZ/GUeZLuUB78rg3UOmUKq1lGhafp9lRMiPNzm8NpY7xfuq+Eqg
7fEjo6WUBQKblrRbJGzh4/tXNcYYWIC7fZL3+OcMhKRmrXc/rNAy44D9awIKHbWF
IosUSKl7PdE9Xs7j4pcjvJIbX3Vw/OmK9wizaPq0RmgP/6cVPidV59RILIAL4cAa
M0LB+cLnpbtohUVoJfKy+l7R8E3617tWASS6X3Vkojx17jdQW9pH6LY23ILutxuV
tAq0gNPMYB1ytqklHRd21zWTgXW+bhHS1Vy5WMJ5sss2dvZpu79BpGCffkgIV7sR
igH2I8l+HsVq2L00+19Q6GcAkKmvNyys+mkGmwVUTROiRvxF2zP/q8WUkKu98NZ2
hnIj1P09vMLFPwmI5rVIJNBIQ1Aisa9IiMMUTXmqcYAQL2J1+m1BqDbaKbaU9lIv
UR8BpyDDIWORmqCDrqkQbaFllMLGlwtscvw22fhDQLt0fvTAHLlCZT/tQMJOueqp
6NKnUbip+vY2q60J1xldJfpzm9e8WKjdLdHP6MPqyGcLdOhZ5+mRZwhraIMGuGgD
xcMHzZ0gMtCMUkNIRyFevckaxl9cDsm9dZCSkNYGVhWkb547FZ+q2H/iCfjt3R5W
yuiZsfO7DuE/ne7kDFbe4tIll808BlZj2XYoUoFJ/wOLiqFgLA2mw52xaPp5ZIRg
XPiWHfqU4VOmKudM+Fgqkt1KOlamiw4DKZRcEu22HjF+9sXCq5ToTsLUKOV7CdC+
o/aCllOA3HsI0pVFxTeQzYGUtRaznxXpJKQO0G7zGfD03Czg7W3teq1JTA0ixn3Y
MUwpNkjzSAXOOyCis9ao91R/thtkIr+LT6ckYg4XRvwWL7ql4BYfpLfhEUnTpVwf
GzzphzjdiroNTkkLhVB9JIb3pa6y4WJWi1+oDTlL25dWVPw9UyPfEV8AESTkwOl5
pDiwFkMfqjBM4TvEQs6iN+Mx/CKQpvIZINxdBgH4LfiX2euzz1ioZW2uaJlGCKpV
dMtXvQRURFw0F5fRnXss+UrJwfe0WWD0G311kR0g9kQTxFSVgTpgcZBDg8qPrfQX
Ej60vaLQSYy6oJSp9Bp4KZmBT7wwQyQmr521vXSdQ7Bb1t0B260jgbg5laeSxqTR
yTZRTNjLxqjsolzT3gcTbooc6ZmV9xLCvaLyFd3aG7y0Qo2ZUnzrfZKbugZ8SPOg
Vkhi4FzfqLHqY4b1ojYVtTJWqNNmJZLDgu3kZq45geG6E8zG3ITvvUkil9pVAgu4
gxdEuMRTkW6gXqSp6Ycvj3iUOZekDwHdLB/7qZMWwuA0J1f66xTzwFBbIYlEOfKF
VB2AUvBaZehA4rj1lhRdjrP96QyenqJlywHZ7cXWO1oUrwjvqjiiB5ugz/qg/Dt2
YvOGk/wxtKzj4CmsI8sgutzrB7sgk2lLA8v4jqlcoX1NeCgphoj2pOVmQHu4MhSB
oJ/CqLwTUSmZwjMXtenyH9A1acSWTpWq2lHEx80STi8WqeaST8pOiAUb5nIBA4Mh
j5YkSKXiecqlLYQan+UZKYPcPG5HKSCp3Th8ok/ZUnPaagiE5ETIZQeK42CdeYv3
iDHBDkHMF+nUqNW3RA3ZC1vYZULQJKk+7B0JnDVcepQZW8NMORKurcnvCZYXuW3k
FMgRyROr/k0IF2gsQa6241aCINEJIK3awUwEdQTpMOaaAuwxZkfwHqVXt5DIlMCU
Acb6RhujYVuOx8Rwcl29Bs5fdjzw3CV+nUkrcJyxj84uStIyy3hjtiElLIJDuAye
gJwIxdzFsGG4+F2C1Nr0Ciz+ESl5Np2ZhA8F/Mn3rKa6E9RHVkgmlkuyLWHRNUI9
nexxhQQYjx4bKKkZKswIT4eiWMh3VJbwpAFdPZXkwsW3KBR2NGuueJHp1Xoadgtn
0GyFU30l26nIq4ROQUfokWk4mAMQhofQxWr3cyhC+pTbbIb44Hwc7nyC5TeaaEh3
wocx3anvC6xGVNQhMruB2OjcKNkN7L55MshoYuE7e8XXm8Oghd7DZOiiYl2rUbgH
sM13DnnaUdbZQE4HAMSezKOA49Lec3fn2AorbpkaR1Zdi6unzXNbafXkrIim3Kft
rM2H9Qn/Aw0RQw2YZNkULt/3ZL+HyW13dHYZrHoQzwtQEgubO5ntM3zr/XWoSbF8
p3oFGO/+r9CGwAFhYa19PpRD6DWUu3VgwYdrt3grMrlpxsF+YXED/ZN+KEJd1w36
huzD287WI8HCai0CItQ8gj5Q1NGhH4wUze9VSoPZubXG8xkbq3oY9wBoB1JmERiT
k9dSmiwLbGhqVzbu5YG1UAClNyOUoCDxafZVBZYBM0ElVEe6YK2nW/jkfuoVp0Us
/83KbpuV/Fbjg9j01hz+Wp4cTB2Crrx3WueO8v1sBFhBpcEH06xQ/xQX3gndRyI/
q2zKx2CDGtuCMBE1EWhu/4b53nx0n5nTqV7elsMWfj+jcFQ5wA7F4dxfmyOwirXL
/xbVMwp6w+FzU5e7j/jiyFxmkpJ94E9fVENxFNsc4tYdJvBQHTFAd3G7HOwnNt0P
Ubkq1H0ELParbVB6hrIl1mRaIVYsuMpF/5RSdvNPpJwoQRZss7bFtGActHLxp2JE
E160OfbTH9EpnMW+Es3ad8atD64mv9l45v85Wkj3bfhHbyl0wxTsZLAnFiB7KCB1
yLFi3dkVWSoKJhdzRfdV5FSDV/iSA3OniKcoQ+GG/8hxyYxAxb+tinmPABVdbNxo
EmiuqD+B0PKXfaRvAdyFCZtVbb/cru7AsOBWZjoYGM9WOJhs5wFAsB5ncaH9jR5m
8KNpWkiFnzkCE+CYpd1GI1R5P5yv3PPv8q8dXZSr++C3dStVJY9XszLIpozPjNDx
owjumsgR2mN2/Saad2h+wB3O7MovFd8gQT/JpRoFzAPSUr81nEa4yLqrGOrDvK+t
GxB4JpQyu8X7qhqp7UuuyZgutqtCK6sySXEpypXnbIDXpsWvPzYbxXC2EkVnCqkr
isOuIplnoBZuq/ZAyQ7x5oauiM19Vc6ECslvjq5ecFUJ5kxB2Kr3wMMTin1R93R6
M6uGuOGubRc88C2AoyN1+R9b4QyvduFyuSER0tbiKZJgcQPo7Pj8DTT690eipPYy
hhDQYCbv3p3rJgs7r/YqVRS+EZa+QUgwINyQ7fJVAKpzcIo6L40mx09ES1cTDKFv
yjTOw9Y9PnfjBVPJMRfZd7ufp0BdfEgfMafm3E8XQu+/TVdYmxIYhGLX+hJo/4Ll
uLFhp0GdvrGKhjuWHpESBIVC/Z8VD7PE9SQigma3i4aidomjCAxdG9DxqXRQBYQ4
yZxbxVDZcoCO+ODk7RNokWfvRhThDrjQDT99G+jwcpX+P9ind93d5WO77BHpC35M
Ac39daASCJDBpmhJLiFCCGx0/WyoHgxq9KhgksPCbkKHvPOc2utqt25gnkLsMnXS
887EAfyvUu76y+NrnNLWWywjMrrvw5ggKYqD6Lb5RY4Jil7otKYrtPWDO0/mmG0M
Ms/JxGRvwwCAME3DEeAr3DdBpsVQGTLjvmhtsG5JsD/hhZsTH5nHj0+8KZ7nwYII
ucMdMEEXM2KIDmk+dJsvG5BZ/lnfyUwdRx7BR35/iRv5hEP3fhpBjQoxg0xYLj6f
o7HNVHX1XYj3GFYYto/uglCOxNXnkAp8tEwF3Q9izY6QhJ+BASIBBl1WwUGZtpS2
nhtVIRw75tJLwNn7HWsKQP955iUCG/zTCE+l7buZisQHR40VkRnXJdKj4utH19Ws
MCDz5vS4S7FWLfaN9Zq/MQfytC5c2/0C7tgfLDoZkzJwgUV2qsk5e6w4DfW68g6f
Aq9rl71O8fbMQwYKBXJhIxjESaoTGXQaCzA+8uaaeC95z7vyWG/Fk9EPJsAFd6Q8
RqohVxlNl+5miAlQsaxt9gTbnqFjRKIl9sMy1mxaJsPZf+vCByhCZ+EGwUDqiiEB
XEJQkpsJDQSRnaIGaC7UFkrvqcck0854QqCmE0GiirBzLBtwiY4AfJnzzIpYaZOn
GWbnzlHaeeI4sVPq+/vvpYWc88sCg48Mc7u/cHiVp8SsI1XXJlBJK9vRaWftyqv1
FoCvOruvO86B7M09iJW3A8xFeH2x4i/FyOKkbFiHw42GEgQlI+OBm+LUvNRPXEJY
uRK7g62h/zQAcA6RqlwXhDnXtebfaZ0bjcuRa0MDU4wG553J35fAQS0XhJ933pba
JhxByG+CGPNQqgpbizDfroytEVmgoW+E3O5obMJna8VAthhlh2kqVN7ZnzFoRn+k
cSwH/DBW9jPrcnGop65h0w8ShP4zAZmOfvS+5JV1kUE0OWUjjv9JL8QRl1e9OkEZ
rzF8qy8OxYMqamgD5dElYqvgx4b5jzOs0RxcmS4epoV9VXcolq135RnfoB5djWak
oLPB/vBt7j4n26ZdDcjgut1J3Rsy6jqwzrGEgsd6u6p86AdAkoNHQuM9lMnA+JC5
/Ah4r5kxTTIaZtex5P2ZSVjWRkT45gdWrb3IjnqHLJvzNKQF9hBxWIft6rhD5waT
Oln6nP/pyBw0X6RHURv0qgdkoFLr/GssROZMi0dhGb6HLU5IQCE7rI+1iXtGVgsk
WFHhOxF3zK1nYqStd1wm3+ocUrSwvkR4ogFofIYGdKG8BUzYfQCxm4K5oay9IYW7
jraBhaSOgjbQHdq8Ia9B3vliaFMDZRu0KpIL+NtlpHKBJac/To4Wuf9ojeSKHbpO
2kbTwyz2diODW2Eso+jEqo5vl8OLMcyTDL6g+9ribl2nU6CFBhp20joWWcG1x3qJ
5aA/uqz+5i7bBZzP2dYUI5RmIpQ6IFjFy8SY7aMKLkJMvDuoiHbXgzurLTwdhoof
Y4a2BBRMM70/70GYUbZtsp8vZIZu/uj5SUvdPVaVizgVB4ZaZBLtJZdReqUf5ctM
wB86WRRzT8SVEIpfXRJ42p0UaOojfu+9yga4E0MO41o9S5sus70xZ315ixhWraa5
FuP58oCDWd1Ok43Az7VPJJHxvkoTkhi0jZjTVsB3EopVavtsFJbsOxIJIOLJqekj
i0nFhXR94nrUz0lKWgWWhMDIlF+DEtwJwsMIbUNo7VFkXJ05VzuQF+Gt0m7CB1ke
2b51TCreJ5raof/odsywR5G+JeCB1C8WBwuCJdAiTuowaaTI20U1unRb+2+IPxj9
+0cmF0qD0KkpwVfgZQxhWAfdQIwn2d9K3UfLdYZKjcRAuuxRw6RDV3OlaIWObPjc
Gib+pSlt2HLMg1knHiV5xic4/ghLixr44iT6dz+WwEs1CSoPpQHAEJsvfCzAVKb4
neQ4lhFxkm+EwmW1BMo3xGO3G1u/sFNYRnhmPKcdsIMWSxj7Ff81AfgBXAMq+RZm
UZp4pW3eMvIsbKI2cgCNsSnWVjS+cl30kpkemQsDcHWMMpnb+0dH4+W45ymNybnO
VrGKO10DhZ9guzyDwlXDmfm5cHMWIjEKly5025/QkSXK8mWM8cgLF75yVdcFZaJ/
m6oMNepZwZAg9UukhALGI/uwrg/hKmeFHAWoJsorXq2NjZWeldTgddduKN9FkAGS
nGGTPXh4iUfFbb7IWDWV8bROnzDjF6i3ZRemXnjQ7a1iGJ1zlfTDcd8QTST1Xwhe
avwb/UqVkYZSYQgZXtZAwYMkebjhGArT50gtFQ8coVhWKK2NULQlLiXVAA7b55th
R0NNDzUoDFSuCdgRAqadYZ87bdHW0muX6nhiTn9SnVXHNnBaOo4yFsOTB7V2u9XN
a7tPqvXhwr5I++baa+LWE1JXPXLsmXM1dEmq9+WNPbfho7XFddun4LLg2ME6FkHd
LJImcT93jhEb+mUFHv4SjBwlNPkWxy3s9mGUcoct5BKS2tuRJE4B4ApCXQyX4D7P
TXyVeCtR1J3ocZEDqyd4trLMu2rQ36XYvgalJxPKwyKU1wjnE80pug5fDt1Bhhyi
fQVWOmKUSRz7dcYf87uUuPvSprIC8/0qyMSUW4doKAKsoeE/lEpxlvxH6NxpETQr
sjXdfCy/lwyc2Qu4FZqJ41jNEDqkSNmvpXZZKkl6m+zPu10b3UPMNQxqsKYcAcs2
vCU9vfX9OBiHpXbutwFdDLe2D6SRGi6QfPdsYtpHmd0JKDdhYFBJmd8Vu8xGxPiN
zMNW7E7jSl5WZ2NSl1hQxtDneNP4/Ig+OjvuTv/ty0LibYaYqxOBiP4djXjp93WE
DD34rydcdpqIedrp6lK1uys+zhF1Z10BLz+mzfeTQWcEthkxjuN2MWinz2AaQ9fo
AB9qCPqjiNb9Mlp2Pxs71mNm1t2/PgxSAA4qHMWEKH5+7qHQzlWWxkdY0a1eLiqT
7AaIxp7/ejzVPyxX2hpZ8o7rLGt1PMkhfe5qv26emgr401k810yppnLSBQYMefm5
gFmoaVOpXUJRDD8vZoesUFfQu8cHw0tLelL4/0SMytujeqaZSr0tCT72qv3gUjtd
D/RPaRlp8D0IjUYkJiX/dnmkIrvwGGjhCKjaf/VkKNJKbQX/aSKv3Tml4tGlMXSt
UAsopxq9glQNc3KP1it9y1yUX0lvJAFP5wwFb8KVKfqZ/itBkgFZTGCd7bPaSV78
G9QysRVTTrSm8ow+PaX5RQ6ZIi4lVCiPl9vj9DKwhx7HvuWR7rQLGVtCzljH5dgJ
UdMQd/l0Nxs6KtOR3XHjUqfluGI5gXlvzLF9/MZ7kZV8QiQ6e9Xh9RH6eeFiR/2I
6LSmITG/u7LvJOVBBd2ikMkHdiCokX2sSHlqsT2h61oAQDyveRdbXZ/YesE0HOxs
8KagbQ9F3CRVHWqVKGEtAl2Y0BHj9LRGoAxKf4iwKd2MR+I8gmU7m8bCR18TcZVY
MDnMokupiwGNhfAcGrBU8b8z4Y4XbtFuDmKOQ4BBEjgo7cemn6uLaUuVv+QLRpuW
QU9ke4zjd4tYonYNaApKsklhif4qyMhYx44VuN+XrdFKMctVVi30/qsQFO9ySS+R
SahMAyi+AOOBBasTSHjdoMvhNfxg8gdDp7qGTBlpIJr21T4Swt53VEoYs6Cqkeqa
VXnUalkPwgY/6E1kldX2rEBxkZz6dKjp21n2UevBBTRRCm35fRklJ/EUNkLmQGia
0lyRXfRIoN4BjeBEfD5cfwOmUK6qRtYHXGM8O41lxO/AAS/66eEUA1blEaWKtalv
TRjGoN+XcQTpFHU2ZCjBMCamGbLuQEpQSja+bS2mTiNBNNPV6+CyQsnDdawSCKNo
PBaUcMXagVU2YEqN3lEBx4xVmjma+caNm8VoAbhjq7/EGYJTdNTANaesF4ol3EDH
2VpkJ2FKYEUH6rzXh2rClmuPbH+5/kYrYReNsF8aU4TtwUG9ai64wcaIDANtBFiV
Ry4fnr1vMpOKMZFbhq2Dyw/+SkdGj7D+HR4Xx3cvt2gI0bqbTrTUkO2H9aNOHkZw
XJG0+HUnlXWiEGa2NS83S2Gf0Fc8i2dQ0zJJaTBZGO4L9DIw61xJxmXPb+E6hNZJ
muPWmPvUzx5f9DPVZlZz2zBsoV+FUWowuX4Uz867F9Y1dTxL3W5ARDdn7XxVTwR9
ARnDKenMfOxg+dJYKMIV6EaZRQrcuDYhHACEfLwDl8FderVTnQ4LzUyJcr5hHQ3l
128esrZl1gQ8UgFWEX9v9LhIwuchmEqdv0AGMj3jYnUQBXGwhtRy8yv6gusYbUSb
w/GFJZm9BwgyzVDtDmqwfoSWSV526XET67Xc5TvEZO5xcEiNYHPJoXzcNSvHAaPP
X78HAYSNJ50ZtdTubIMTDtaEURWO7gEcLYjb8eVXRXCjF4eOTQrxC2/JMq+DyET2
rYRHJaZ0hEqqe1eZRmr1shkz81QoPX1nwH6IXAKT8X6fCKEymKa4TnthQSv+DhPg
oNNlOViPXaulne80KsWtIPba3aB5tewLkkSRlVLVZYrsa2RpOMh9ONWevBrHMQNl
d6f5KpoYCCENtKumxru0zwSyuiH2KV14cocD3oDTbJ4LhFzGdWgLV7pBss99HPLm
2pjFNKcFmsg6VZTmmh2Hj6+qO5jR823zxH2bmUfZXc8c4BP5UZ/xg1mHL5okyYT3
3hn55i32FyQvvr5VOLR6T07gS0JH6A/9PLY8e/9uC7fRGB6rVohf/LOrpLIC0vdt
W3xRnnVHe1MZc/VpNCNvfQ1t6IiBeh60I8qUxydhtvM5nbUp+Url2wyiHaF6Jgl2
mCz8mcyDJKV6gEbHhMeSEy0GAekzSiR1kPGsmMjO2qaS6/4tkLImHcBTz9i4QZhz
qDaU6ZtuhR2m0rhYVqX09bQCvZP8C2/hUCdkkxMpQiY+UKEMmO5Esw2QvwAoGCir
1U41kF0B04VXUxAjib+Fp+5tmf+y6Q04zLJfcEQixnDUO2rllUAZAaPze8ahf+/r
40lW7PrFp8qurg/ZoxJfiLsqeGoIIpXUXMy8CxhgTAEqfjwMTp7yaT0Cz5coQQ5J
SXtEnfn45KsTqn2jwxa+KRVW+EcLiIEbMs6imx5E9+dDvP/e0IZrPQ0BETJYGoK2
gHMe3x4T0Hals4xPByaxHR2FiR0rdr+slG0VlX4Xdo4xer07ymzQx+32w6RBX/4P
IPyru7AS9Lct2cUUUkKDhBUic7xNOHb/YfZ1fVnm7wu59a/5maY52VxUjOHb4r4E
CLhVSQ27Znr6HOCaXStoZaJLLdrMqjnYV1nDdF0YsnauU+ow9TwDqTA8XKgZBKLK
dxgGHHsvqHgg+h/2yLwNgMCTRJRYsiGiOKnfgk5RCKYk9UusmSuWOg5kHSOsyThQ
CurJL7ybT4N8ujnFfh+cpYXTo0vZFfjaGCzNJJpQhD3EyHhJBD0GTAWTTQ5sm4Ks
zDOyV98Jius+GRwlPkn/JsH8Mk/+Umgdh2APZOgm9YG36W+/EkenOFM6SMElA2GW
9lhEGs9txlbYHlPTOFd+RrCUnaT3pnqD1EX2R9J/dCx3hiKIv+fWxzc3jC2MwSgM
FkEdVNhCg7Q37OUO0CZUwowkvDQdZy2CYlS3vCfIsxWipbNer3MabqeIqkouK8K9
AOCrmtMgmkodAXb0xlqREPAOFIwIiY0qyTccguNNFrB0Ke2T6F+kWUElCVt+1Cls
if+tYeZls+AuyjE4f7a8VxVmq8+EpuOhgdXdMDKy+RDJTS71dTwUXEyr1U82iCdI
1sE7aaMZ1lBWfuC5tUDIoc4PdLbNJtWL5vDVgKFpaUR/fQFxnFSjt6pZ3G7eGTPL
/QEs+m8nZUqkeTWC8WMBxjb9VGHPApZEkmb977DJqUr+8qI1dpElE2KNDb9bY7fk
AQQaSxtiMhh0V2U2zsUG/IXq6rK/Z9k4G70uhvoVgz2hijWKGw1E2hT5Q547MglR
DjSd3QUvPUg0zwl5iif/9SsQy5ypEqyGTaRnWCHcL84mDl74CYFnCVt+gXoDW/SS
Xv7RdSuCPWJAHViG+SofcAS+PWKtitYjooxQUTF4otnWsUCYq/SYOOc3JvNgVNH0
CW5R+fyUKd6ErM09dpD+4zy0kaZLKi1l0mACzkql/wPID03G/3XVzqg3g+9vNQWv
xlKVloaoY2s/ev3hs3V4TMOwDM4v1yYcGaaqq94HvUl0xqQBujwoc5fw/pXPq3/e
b1wSu2YvyPSLESxfcyENIOjjI0WeM5oHlAzQtLlTE30mbd+hqMDORya2dfvlbqW3
SDpfvwPl7nb0SI5e572dGfnGXu3S1ttvp5DaEYMYRZt7IVxHQ9VSxHod+tBUoCTH
BVw5ULzWfcr8wShjmivt/GXG9dyVPRG0IipmXiUtDbLVz0bTRk3GskQNY8R8VNJ5
b5ScyAMohvSVCERiE7kYF1x4Kq3jZUA8U//cnm92fbtUPSove03T5PVPPSHGE2cq
j+Ms7rh5MF+ZFKMLEVPB/Gy2yxUl85TCGtvJhq/Ud0w2ZS42ZsDlYF2S4jeEm/A2
4M78nAs8/cSPs25VSI3KV2bQezqc405yvaNj74N3zu1LB6JyASv+JgU4HQdPa/iA
7wM4aUNNcLVteh8De/ssEOXcmWWhE85n25cliwTipcI2BBYIlJfFRSREHKOS18eh
43It+Ci8bKRncDnKtH1Ce8CMS3lwaSKD7agbZvBUWR/Ts333vfl5hvRet+MkXdnW
Tr4zaLDgYDoLsX01UwQzOl5hEYxYzFVJKkSacCYDPiEoevWc6x6hsi6aOAwkchKd
xTuBP3wMYxsOg0BD9ZBum7pYZ4yyRw/OW6NRO8jqEha7mknNTtOP0BHPaj7q7pQ/
i0vXf2skF9Oc8ft35gaa+3iBAP6LyRoUfQslVpuDJTbEShVzN80OmKwFjIQXYgJ4
2JWmtKtqYhO2t6+2M/Qp8Dsn0OXVLTNnRrZ728z8XpM9lufOsoISyy++J1PQq6XH
tsetvCSQrDLrAthJn+7UPn4xhvdgQgsIjdx9FU4cf8e8ilb7LtchxWZTRqNkscBF
GbXfQm/BMZin3KEaURUY0qt3j/2v7U1bO690bF6KI+EOXSMYRhesaVQUTGQfMRQj
LZhYB1R0zF5INAfiAU2qzRdVLzL0h7ATKQz0mEdKDFucL2usvo9Aq65xKTmpZuGR
fvYaCn1773SesEtgpODOqkZ1SWbDZB8+7ABC+abZnjuQJ4zXG9i5h8fXVSbhScTo
iMfMM4M2LgDh22Ql2TJ6DKUYK8PNDTbpF1hzS0HuzkIRvGvNHURgcjymsu0TTR4A
/Xysnu6p7KERE4NvI9LrIHQ68hoCGNLkj09oI1cOWFnAfFcUH+pzgrDzIVO4OaSi
EhfOECBww6x9l8aGjf/FJCa4FeCns5FsYM5eT4jlT43BNPZuqC9BUyjnj/cgYX9O
bCi05n1BtcOL0kR4DnnTSf7ZQqdTkpff7BccBTggo378ptQvpRhTQgMHGEvhh9h3
VhGHFjdUdVOaPPJIwuqnKvf7oNHe3qje9AqKMsyvm/ThotKnaWJNg0Q4IvGTmfs7
FsXXod7dzh/+2GkglXipdZB7TWaIOwvkTdWQkNNTe8zes6Hm35uJkbcpPLgGFpyN
GeBPvY8zZr+VXLIQ6qS/iLOlpG1j/bcsFEExgXQvmPIXUXM3jYP8qce3WMiakwL/
uIjTeIqVFkxT92c5SSPvIDkd1/gwl+jHT11hLg3T2gIdxvPubRG59ptHZzIyDvTw
tUoY4W4uPzmXR9YDo28OzowDxMCqvbpv2hvoX5fnL0Tf23U6S2gV2te1kTukrCst
kjf9GOQKnzJKiTbMclX4QZBM5ftZG6/NdkZoQ9vAulslNjY5XkbEdMNyQNOZ11sv
GGXX/LZLCKevqxw8zN8Jxuy77KDzhWTMnM+QKn5nwRR2NgjTzsQ70VevrsjXhA1y
8hAgE+rX8+aVW967FD9TECpVl+2GHwJEw2NJ/1rUlIl61t6Ae7vnFgpo72qKghpM
33a+TCUBvlbLl4mbdOUNctVSHpwp54jK1Rurc/LOBjuYyQ/c/vBlG39usX8OMds4
LzEph0rU+OnlWlkDaoHBjXztE7/nUogueRuGb8BWnsOUE8lnbPo4eKPrFCw/OcRE
p4IIsmIc0jOAoN3z163x9uTO7piFSHnneUwIhO2MVEk8vHYxw+WYsXhj+/BC9H0x
3CaA4z115enHOhrSQyJt7ZjBJei4GELiNUqhfH2qQWkinohYzNfLzrtOYeQeQBHz
90yDfVLu3HGOspXPJ+xdSanqXFRKJEZnnIauJhjpcKHwoVyPfKkW/xgmTbbB49R3
MSnGzwQu0xKkAPzbAkD99qhGoWR4KNb9ysrXoJYx0h2dftHDXxFvIvIuO/ZbTlPX
xyRycefkZwwxv5qLeavLDqDR1KTjUEO3fdKK2eLsc8S2HXLDpskRKqCsMCThM0Pa
v9CewmMgQQvHVbgQmzxrXJFH4umR4EpsD0V0iK3GZCmirCqY0dGRjdcAT2pBCWQz
qRsdYPSj4kClp1mFUwptyLLYMEWuHamLYlEE4asst1eoeeFfph1xZ26CWmXYky8U
eO1sNcTH8ajIsm208Ki/pR73emy0ESwR8nm8aD3l+i3K/JuvFIh+dJbR3Yu/kjCU
NoNvT0Em062A9WevNZnAtxwfn6ARIi2LNBGii6IwROwFC/3L97B+XfojLhVt2GY/
Ku4SkQ51ZKRAU0zy7lkQQoHhi0OiwjcZwdgLYMjieYsHtzHzY5iQdbAwIkQelmvr
0Q+sTbnV+CyTRdLflItcVUpPnmhKmf1IJeCckxm4XaxPx6r8Ae2HHpQuRpUAdwbD
oNCOs9Jpp0pipudwGGNic+pG1GPygyTg046O1tqRZwYlRrEMUMC+tL2q95yWD0AQ
KtQpYaGqgmF1/Ur+V328rWdRVQOlYnsrTf8ZqNs1dEyShRAMb7nBOtbhklIlfLFp
VeKF66/rnfov5W2OB1kIkdIe35OXPVhBzQb59hv+EFzwuDxK86Ed7x5FM2I48oxE
MTak5NBy6OuVoNLWZG3tLMvLxI9OV86JvwvhumpuT8u8gqjDa90iDrNYS39HV03G
ofjahwvyCM/iloAifm1OXNdn+QUCsC3O17pfyxb4bDzCzmCOamWUEb9XxOEoFS1E
OPDxY/o9nZZAuouLXrl+7hBK7dtGOJKMbFNBnB0H9tDzitLE/ErMhW4F9mZvsCQz
NzGTd37DroJjhoQXAzktkLaV/mhT0dD01n1WP1szMK+bng6J2yuxJqpQuF0x8GrF
2Zh+/NDH7+2VRnSVQO0WHBTkUwVwroIXEi9AxmkNtEss3gzSbA8bW0QYfmk4KBcI
yNPmatR2rbzTXN5KcatiLPrcEvNuphxzOPY3eXsgHzkm8c+BrpYtptnoYqLujjkR
RNj8PUwqd33n1Lnhn9tKMIZLPu4tSe9FeaXMk/eH6hRgpYXco5EXZoFl9moV+Nfz
9DS5sCOfmEFUnVIGzfBreglun1ER8LtYG2oFZNP6KDr5ZfQpWSDI/A7P/wJJzGt5
gGs82AsL2OQ+889dErNggUc+MS05a3bqmkNd49GnSUC+TMvCg2NUItbGu+P09D8P
gVuooMMp9dXBrJxiKVKcEeYal/cFhuc6MOdH24VwxZvL6hvzOhjugGC104kDvyOM
WIgj7d6GdERl1kskhTiuowfgBGpoTOLsTktPKhCtxzZpJCT2hbWthYuIBWKwf2qt
8m4QMhOYZmggqkm0AirBUiLEX3dLLFHAqEFE3g3i9O6XBclD8TqN4hu9Slbpw394
Oe5MwteST1DNYhJPIW8V/1QI4l6EyCzoYkpKt86liG5WocPlSHeXBLbtokl4ctgi
j7Lju3M6R/x5SofZ0ZdAL5xfK4rGq8BJLzdUkmYGYa3ORh2HFxa9ShLSeou64IKl
sWZOtz9EXUF3ODYHl+lZWD6Nj4fMBFoZ81gTLqMUf4nebeZv1stgdLsUz4+jBqzZ
STZ3CqjCCUO+amf9d0+IF3larhFwo9Q7EXTxur7iQRrxx5CoFlVNAnbTdkMdkGjr
52sffYnLN24+sA7f7y/mJ8fzR1+hQX6t3La/sr7XNUQFEl0ohvRKlzlzebwKLzIy
ef+bOkTcr+TXykc5D0ZB4yGI/wtGiBY6RqJ0WZt4bvxzzQoJzeldzaTN43qU+s42
Ul+rDZbIQwlK4QxfXa7vFoQ9juQ58Umrr6m+xTWjcCd62q073AT0teVXML6DNfvP
Xqt9mppXRO9cE7ykOt7boX8m1PZPpHVpiSVlN1u7CIrj73Uvp7w0vetTwFhGiQyf
QH0B1bS5vkvsrX3JOLsbNXNyu0gN3QbjLS/ybBPRza5GNMRvR8TOoSGzkmDUzAfz
/DKjmWbqLa3B4BHj02XVPVKKsatjrFiszBnLA9JpPiVlkGvV+S6ETpb0OEqvKN1o
SfcKcn7CNy4F24kO11m8iymwPg32wHV9OqwKaMZ+MyC+fCcI5RUDegbZE9aITWHC
ouJEONdda5dDj4Fk4RPTtZ3PSak+uZPDPY59L7sSz7Q2U8LRvxlyVo7/1vGhm2/2
AM2z7MEd3AaebUmDujIiTPxKSQmjKha1VF+PIWbd1PKWSESZC+WP7vQCnusXzeBt
yoC46330NUxkvjjBfHTP6uTfkROnn8go+sjuIF0Ohxpo1PIkOmPDlJEGjWBYRlTa
RKwjoBlbrGMEp4DBWlPhWaA+mm2iiuTT+nGERTlzVBUCOQYbBUl0jOBmEGl6a/+P
dyN1v2QOOLa/dNccm7PgX3e0uprPn9wkDydWZTqgFZ8HQung+fhUSnl4RRFj6Qz4
nzA92z1g7yxr+FSnEWMvaU7ZwNJH/G8GhcpEQeho/YkrLlfNEJS6QIATWwsSTrlH
BNryQS1gkNufZgFDdm7GDGKXCHk3cABBW1AuLR+d8FHOEXqqfEyAaMcnbo+w1kt8
zBC5HDZju7ikQii5303VqhF7D4E51JGrjpd7jiEQItQYU2NCEcE8yzdOl8QMJR7z
cr4OU6YU02UPCAH1mAVb9OC+JlKqWm2TuBRbXGcogCrdg1RP9MVnaotwfUWaZ4eQ
Vay+EJsrG33iFd21P90c/CDvHO/gcYRXrbFKbo0G7hm8xcbOyQsf+pl2KTqM2cX7
+gdj7RgwvGfMHkaBBj6tVBJ6h6MpkIyaXOJ6DM/SQTD5XBzni0IQBeu+HMlM708d
DwbUCUb8rbVJZatPHlu8jPDpQG/UBpOABznErsFnKtPfNrsgBSKlIcw7iv6OdsQP
zUDN4vsiYPWN2GS5wse9BMjYLfL5E5H5fMaNXHLGfiR4j4LJzHegbsR0zZL4MCNF
czkHMexjHFy0xpBy/ZnyNnh67c5A4QlrfnJU+UVH06P2yZgf9JtPXRf75sk8MpKZ
7p4p/EtyrX/2RYAKGMBSwGfkSYwW15D/biK8j/9KemmmayXhG0eQIYVCWUn+q4Dk
IkC0PsJPnyzGSGUiuNq53linEfxiHifDwxnMxuXFFNHwSJ7eEKfHU2do0gsgy6xr
HkOfmw4F0rV05zMFhTjMGvyBBiRziSZANgWCDIvKEMi9YacLXhQyfvmDN6ZQi+tN
Lsew/nYshQUQ+yvseKFa5cXLZfGosRG/+gspVhqP+cFruTUgmtXU4/LXEbseE7L8
SdWZ7MtTluSItdYyGu0g9NB8T5qrrC+wccE/49MmaXUwBGXx9J6MCOvvNXBxzPLe
YFdmz+P8LAMPgEx1WUqBBP4kjkBGvehTqMe74t/bv88To7wWmrmr/mP1CHEyu4DO
CW5nqYtB0aM/YOG15JBElQ+QWxDqOwbDQNxY6149VRLvudzpgHF44hA/iXs493qd
qASvXgRKgDU+whqAZNz7KCHlDdabmGsGPTQgOkByQqJL4yB3cOUHpOPoJBjR0Xog
/g8uOR23aLmOlSzHS6hUTMbNm9GdSt2YbxG+WQbzXM1RxgltnmwdEC9tIWg6Ho9M
el/wjWSPkOGXZgFE7heICAVPu3G8MPnDWBefmncgOdsJ/Q4N3n2t+GpZGPv6QTq7
nzJyezHBtH0FVSeUvfDD58vp4q2wR0aVBpirod/gUy2kUEXwMqQKljBreUfmI2vI
NNlLrQrwL5EyCNa6j5poFHmguRiw7CoOaz80SrvsXxWlT1x7LnQ4/vlCT4qIuFrB
hHgH9njTtyNlcnMna4KdHrN6jsFzdJbGjiuI5xY2e7I1eN3C7qaTsldTz5+duMvs
4jINJK8wbzuh3kjHU0IaNX9vVzp8s/tczcGLGgFwrqFuvxBXKULU5sJvR+GLg0cw
dTZZY6J6c8MhJYWJJZf6+5VWJUNZ/AcCa19hq+LLxT+jMYdLonko23ylZVngPWUv
xUx/G7Si2KMOwnC7PkgxyieGQ0LfO4AIS+72zKlZzwBUmOylMu7Y5Whckmt1w7tg
M0tDw9mI0q9/F/U/ZK+1fIJeI5nLNrvr++sbWUqj3e93k7NjGO1ob2hLszc0meT/
Hme6HYMLLYBiXXoke6vAuAYlFUQ2vRdxKCCC+nZf1rhGZM8NaD6vrneZtArYIwSa
Rbawos5IeNx+m/WC9WB3vs65LplkdrojgNMReQWZrzD8CaGPvuOuIKhRO/Ks09i1
ZMEqqHHxEHbhrN6PirLWnhSA4lFw5oLTMU8t/dVD/ALvl8XsyU4dQ1wZ5D7DQhyu
qKetU3LKYTuoK7UH40KmIMaIe/2cEDahzPJFz6n3LNREVpDVOqXBziS0X9qpLQbP
FLMebrHdeZlR31WwXYOtRdAz7agnvhg7TXo+eiixP/EFzxF5waQpj19FFo31nq7K
q2gl64aTLa6qDNzeDcwqhaGgT+awDamXFFQzD9kzH45+toxLJJKUny7719aOmPBR
XSsrclkdxNk+U7/4IR8n8p81qZetQE7FtFTnJG6epdmxC1C6Q1DXYTSyzkQ9UoQ7
GhinZlr85+heaoMu1JAcnpqY3AlRMrdQjZqsPYvPY6ly5QEGQeHO9rImFSfrjy7A
ni0QSfVheCora1RvPmPwJW3c4zbuG9Tudgk93LQ/coz9FJioWms5+D1UnnNFKO1I
5R10h95CjjLXqJSTj0RrEOBOFppZ4uvqBH137uRGHBixm0uq2XiUIY+sGxbywOf7
QKsFq72cNLqj2snUENMNklfXbynCKE/Zh7YISuwvK1IBIg3QOxrWB61A/HMjDPMc
0Mb1avAHzupnllLSIWVIepR3mAWYFB11QsZ4rWGu7mN2mvntLWLWCEX9kYO6a/MI
srjQLMPjMfJ4n9HEHHNusMmWPsNEFy7udzexj2moChAi8rRwzXnPIYkmdN/gAD8n
ysJrM4L8A4L5mfdnHAEKedxaD5WdSTwOU/7F9N43ZlTYwsoViIW4xGnAqv1a3psM
bP9NtW8wRGEiBdvq8pazNm0vQkuwCocf8CzBZcAmkOiGAe/BLPRvn3VF2CTL1EtW
6QS5xt5SFsGZHsOycskVHcfQ1y+cvgmCYAcOlNkAe0WC+KfMR8GFVaAXOQOe4IjS
N+KXfZhABguwOu2ShBXsBxGPoINDh28CZocP0zWAD2MCfarMP2l8IkmLFEplzSh2
dBktg0mQ8Ce7vKAfotwIZ2YBCDbHe0tVkLGglFxf5jcGbPr/llattequ4n7EMNcM
XdCcgAH8d3cHULOJg+0eJLDPV6SqgwKajxxE2Gh8o2PIyxhRVOXUROcSz0u2AZm1
Kt2sa7HhHt7d+JkSgSBXEcTH5kYRJyXeZJU2PLR8s36oWmSWptENEUXjCeSBLPJT
8i2+x2693fxKxEOY4+aXzQd55hftE1ZlzPzTc5Adu00nje+dJgqprvkYC7NCZxhs
HrfDYyBRtBVWoiTG66aRAxyAqDbYxA0GGDO+XHVJHclK4mSnhrhTeWx7QN5Aw6SP
FU6e1m7B0w5C6DU+9VjYAV06sKle3/5gSnywcjVqE3kxvEzJ04LU88IpfaJ+2Nxe
DIXVdWZcchazELXKcabspUqQjSZofCq4xXV0ZK87NaK8cG0BnNFMbD2yQPzptQLK
8tNTygtfkGLyY4shHeZ+EAsvG4Fd9ial98g84OD65NwdqDQWPcwZZ8z7H0yok3TJ
jRTiDDJcOm9Tubj82d9B9ilf52wr8gMi0Cxmv3Lg7RcVFgzsiWjbg0JYYJoFJNlZ
+h04DvEKJBZxr74OCAmPBzGyrRzZIKjgPJSrI+yqA5Fsm74QYveXGaStSX63zwmE
2xAT4JNvl1lu5OZJO/6i9g4cr8AX2s+0L7FCdZmCOb0B9i5u0hQC9h+dMLWuQQtm
KX8vi0pMXq+NhtysvR0fKNQnk3sfiw0nGr3oYekVZ6AsK69rtvr692D74L/esAfQ
icpkLu8JMMueitOvKiNgbBR/Bhu/dfvpVHnlZs3OfRJ/Z4wMsungXNeP74Q6z6sl
MmhP/ITrgOiBQM+MKQY2+9RrcFHZoR/FysaBDe6iHgoRv8P8sZD7qqZmeFWl5zGJ
9QuswOazOgwxW2AKe0mlD4eP6n6NbZ41LSo6DECytiAVGD7gG1xdYE8LBUxGaPZ9
P+GPO6XOXDc6Usu83PkGfMqOY/rInsAyVF/vNMtQ132rFSwiHfKN8oq1XF4Ct7db
020/8okobTZ9nmTgL6vhcYLbN37yM10H82Vi1sN/cisknZbzQzydJs/ipig+elQA
1iBkL3XcdLvdlWuRmN06keGMxJsL9rmR5seLAbpzbIpB3f3VLTQLX8wCH++ILFpT
voDMYQRD4zoE7+re9PY5N+tORLbCBUrqG7WuVkDIjiB+JJ0AlbVPfySL6h1SIjYs
1jyY1Lwd7xzbTnkgJxJre9NuHEKH9WhhWIdRUG3+hEVEKfItcDjB5TOn9SW5V1L3
eD9MW/jaqhCfAw/HEp0ce/pyyWOpaPRujTl8O99KKmyUd/W1zGNm5MWQScG2XX4Y
L9X4FDZ+eYUFx1TdI5GRU31ISv4oXOgW/nV6JjfzvIxG4xCyOU/oNeGiivXXRWug
4kp0LDin5A+ghD8OLlTFoanq61QZ5+aNP1l5eA/IoyCGPO/f1XJrxEIx2q/0RFIN
2/EVm2JraQb78tVjuYoph5NkLkfUX6O66jCqCAm08EDe50P5Om/EZxIGgtgfulSK
UJHQQfX3uNm8JCvoLU6nyMlH5if8GePEZdt+fXd6dNcpa/RRC0kDOkkvMyD0L8fe
wU5qHKwSAiRcrd2DfajnPLdr+czYnIW5wqPraLRcTel+RhpsEgbSRfYKPp9eLgkf
a8RUIZV2E4tTp9WAmC7TTcbfpTyq6ExiXP3mg2u2aV//fmcuscrDUKOgc/o9b27r
kbu1D3A4OK9+P2D/oceMVUmhHjoLP5F3zG/qGxhkNQobPBOVF2UW1u5k8adOk3uO
2xcoR4OhrVCgE1DYsu0uoyl29g4PfAR9cU459YDKo2HUXcj1wy8u371L947uM+0F
BvzhqUW8tenXLIV7cNon90Vw8TpY6O2hHI2LLzp4WZFTsafYhHQuIyVoo9mEMVkp
4yorqZZ/K6gSIwkjB9psGyYlU1XhdMaE2y3AEO+y0p6/IIsVw3byL6hunXQcr8ZR
S15Ia5NAP/Pl6NrgtwLcZVi1Wv+gdsBY20Hu6ul7TpjgBtQra7LW5k0aUhXPCYZ3
vwoqtsSP0DPrsFR4mUnCvsCSq6Jm2DwCt7xovVa7pPkkmvNn/N919IrHZnv9stOv
AjT9xkJkBhidGycSgYu6is8tgmFCHnuvuOOrRkOS8sNJ+xsuS2U9n58UjvbrswUZ
MdfRlHw3d6iEj9UpsWE2JcSPuB9prMAw+TZv7Qu7AvRK8gDemVkwCLM3GVowN2Xw
dPagFVA/cc8vzrKVRwWy5r4FP6Ug0EAHFUgpaRyT6Nwjb+OwhGQKRSOzMCSYYRlw
O88nyikavwqah7e3gC3hU0T6RkhULIVNON2zn3uB7mt5z0ZXePunEjTcFhTTPYP9
5kBtSOUcdU8lUoDKeHgR2xQtVM91NO6owMHn/iLdu6F45nNPzfnXIb+Ek/89Z9sm
jUM5vUf7fj8FaLToL7+E1bqLDzhRgDQx4W6sXG+EmyYUx2hdOGB+6Un+vSvv5/TK
g0m1C/gr6Dp3+cbCCQTVB8HSYFjA43BVWZ7bBDziCoKXJKYre22MWAKse8m8eFpf
tEwY9hrY9yeopEpRiydu71l5O6HeoL46iPnIiFGgeWKDhZfHFpuXVrxrayM/fU0N
X5D60rx8as786RPgRMvNxbmgxw+z6F13hnL++FX8WGKIR4Qli0XfriSa8doBh4SA
hJNRN/tgatI3awYylwVIsrwa1CteL3NEf+uf0C4Hj539aHnU+aitoIzgNtyS7gMi
4pqTQNRNsnND3vPLzxOMbdbjFLK/3AcZ8v/N8km/CHFWCwyaFh8PrWlIhezb+un+
diGhFXZRLs8fws6uza9XvEwWRFoDj7/uawXq4Y4FZHQKybQG8QDjFRBzJx/OBIhR
giiOn7O+lthSVPn6pMMBGPxUI1oyBoqnf5hoIRznr5q1sbgzn2acp3tJoIu/6lcl
Hwxh4iTP4J/blOdPj1mKJd398hZEt8YWaxWQEyTMtFscHBRGFl3aBlXayzr0icks
D2J/vJKjq7FriQZKktmub0MWJb2fiBiYpe+j+6/VisA2Sfl6darnFioQvunifcjr
vXwmvQVFzCvC7oEALIA3fayoIdiPKmZ+oT0GIO+yxP03MdybNmKdALHalcz8xw4N
uiNFkY9jzT4FZvpX1vBVXkoqzN7G0GLLziCbZbitO/HXYpcnil0x0YgdcsXuJB7B
OdNXZ1pBjBsCwLOE+FM+iIVOc1TA44Sch8D58G9l8L4H8JMVZxPtFd7ImJFycsx2
ONcnSb8Q7MKpg8borURQX//Czcn7PD+OqKukm88gJ82h8lmDSnBfDmnrZizlzBDx
wi6UGVGsFtHMiLUo7Xl33PxnfAUERxCrTVQ6mmKZg9dnm9Bwxn4vT709avgTwhWW
epM93wKmkOxSaX4jxN36F3qirXqJugvOd4GxDuhWePrPxCfpIR5EzoHfXjhGT7yh
vYQE83np/FbjNpp2Krkxvt1hhNaPbBi439pp3ZHO/Y49lMcEOb+B/ojSShs8zd+S
Pr9p0Hhc0zqMhMAMnkJ1vFNc4oEUFwczcIQJdI2f3gATgILKGWSsNuLUablSA+ZX
9m//UW+I7+IaDa3HRqH64v69+1nrmBlXjfhM62s+eQzjs7V4eZcz4IBVcMPFurBL
CgZRlw37Nec9OUKZNjiP4zbBLcuFzNbWrANFq/nY9iLaVDTr1uLmlOwQfDlZjbSm
Y1LqAHGnPVhaXII+UjDxMKsTjTwRLNbXfom9KJkrGa29NI24pQBsjwyYWWznU5nF
OMjKhSz7Ibotvkjy6ZhrZMfRWAXpVJFebamyRMualktNDoZg1f4AdP3ZrAeHPCWZ
ft0yzy4UvNhSYqGUBIF0t7yHNg7hVEEJUbvkIPPDTBGLoKL+AcwygTDPZkL4uZTi
Zt7FGTVIptXj/fAJSUNzMhnkes9lUlfHQc8OIuezv1JDVQwsApfUEShFAgZEY2z4
NkgwKWsNOCPQoUB/fzoO4XN8CvntdrFSGZer6uqJL8SCqz3qZJFwz5I8eThTbjAO
0PU/9TeiiehurOX0k08gwZFGAcaV9l/8ZMTrtRz0oXwNFurFE1vpiadVLGziKWCr
jZ9qmO7262cT7I2xM7dYOCSA7X0UWhbuxde0/teZJOHmAaqyqXoeNIsCuRd7L3du
XuPSlt3WYrancQQODLwrdFQ90tGYRMRRh8MxTqjDO10xNJoQcfg++XQFh8qhwDIN
+NK+rA9HLeYHCoARTIP2F1XYWr29nYEbg5KX3GFAbeeeTOwg4iVzwHlwlLB29q2i
Q4xak27L3BUYORof4EuFWbFn1uQkpLXII7bDMOT32+6Q1CyFz0D143QqfoDn54wb
j+enEkYHEQ666gn4XkyFzs0xi2opAHixz8RsdwWeIn+5siDEOOUyBTPb08TUsReU
FSf0PisEbqnK8wdfDMu3eSqs/1bWWYq5E3ZiWa4gJ3enMC5xMqSGk8v3rCNrjPSQ
ed0oBLjjzpoD/DGVx2Hj/EyTkNkP1T5IJ5ovswAShy5J8/ZizZa/9bU1KXANcIZl
48c9nQtpjprNY/uZ1nGgVPdbWLtobfNHwRZ1Vo6LELyWu1JDAV1pLd8GWsJYlHca
+4lTlRAwWIAXLtBiN90TUTUCBI9ON2XhtpiiE9m81tFjVGWrcqLgFIBQwZY0Lq1O
+cbVtQmu9e5aQdHNVJjxjymtjEUIzeB4gcV0zaIaqfLpWyrq6JuQwFJA1hBPwAUz
fggQawZHIEvs2eTi9Xj4qx0zaKqjqpVg3UmpSTb4cr49M8hE42N3OKeDpA7m70d1
FVrHEe8m3vfwFk6ZNdc7v2h9IOrxfpfzHM7lxfgzleZwtHVsueLgq4buzV7HArVU
XnvNxDNWk5j+hWBreCTDmXurCds1cilu6Ghi0idK0Vh0fefShxDzNB5TqTViCBoU
8yS93Y/4XY9iOkAN7PuR2d/HF4lzszYDLQFGTvKA7pX2I8N4XRNx60Ez5Aet5wLh
5fDhzw9IF8koLvtRnfb2SMoIJEsHU3oBUdESD3jEIV1qMeTwIXOV8jiCjDWlsI6B
jaQW1ItIoRuP8ghKOKebOOpKaXvua+AgLBsm2xEOKtucY15kca1XRVZVsBfTWBKT
ebml/tquU2JR5LuQtemCKki18F4NdtHpj/38o1/3+e9Yc+IiIurObtmGsEFdL0+a
AaZe09LrkimgNp4/8uviXyJNAsjbcgmDigms1EjsU1CCvzAYaoOcCFw3Spy0R7R1
+TVcJ4cTrmrXVMfvwEtsVz13EsdhZFkAF/GL51jtzBZN2oXaf054IqDDK+G12dIz
LWd+67127PGFzOUCuVpH8ZUQlOp3pVHhVyEE3zHsS6I+E8BMhPkiOGt0UV4ndL9B
snz37pY+Kg6K25Tvh6K7NCcjobY1vwVSC5UsZkZY8Hw0s9WDvtPl1+B+biPuq4BE
RKjn7e6evStEEODzX9NtXyDmWJ/WfX89ykqeUnR4521GDx4OU10JbPten1+JBL2P
1Zo5xjS/noF3wQKf9ALzlux5Tvpuk+Z1wk6HCKMz6MT5oBUDNxV0AtO1P5n4PkgI
DnkDeUkEY6ir9IWgC7My05OODQE7Ebf4MH/vANtM0j+e4rpRWOim+X4XXe81/l9C
zjLUgXVnRDCNoNGPjYBGb38VUwFLIuBR9CLTaG23FUfubGwkshp7evbwvh6k5Kac
7IEfuw8ooQ9Z/dxd+ZKjY/WsgVUjuXzVRXAY/DRVIJ8RvVXcXhgibO6MSHGwJqtR
b00N8fUKDCg9snXZ9YyU+kK9/yM7EUUWWO1LtZdUDdzyFzTrXEhV6IPB4bq0fV+y
hzVF4vMjrj9HQZNDwivcX8S7MtR053MEpTFj21ATYnofFBDZzDxdwjm8EP7mvzBk
g9Ya9Pl743IZS0eNQr20sXoxtHsXtpZN23AmVcWKDwGd2ulc75BXo8GDnDFhGTz8
Gni4f86Tb/kZG+kLZiKlFK5huMERzDP1+IqZxYU5UeApGPwdUtDFCKWkFkPkMLQl
cIFPs3HV/RRWoI2EHU0iDWMG/NR3OiE4zxSR/nBvUBDNPfy1S3QCeUYMdaQYjABT
Rcg7i5D1AWni112ZyMbmIewOR7JlgeijxIE1KI947Dys/CIXs9kEmJA1ycvsCzdK
OE+lp6RmFAcpbERgHS3WJTm/qtXYGkuuFZmGbsjUNjA+WQoqbdFsr8mHxz32AT3I
zkZWB00J4rRaoRr/YIzxvkObY8Y0TOZVGCHDNhTDLIQomY1vt6bntm1t0k6cne0v
ygCcXYLaaIwMJ3WjIGGUvK6XzLuk1ZxYZ+XJz/fUcw76B2dZ83c8KRMF/33MJA3E
RTphgDgLdjd5GZ1w2zhItX5hMLxKeD8QQn78sg7SiGewbSegkcRd4ZFFqEt3dO45
TvEIMNL2c+Ko8vQzHVbTRFiLKdFUyG1gfJYvo+2K6tp2oNLGS2yWEO0JKQdzEfR+
ncRjijn5Z8soS2mZEJcoGWq1yHfIAevC+WUkryD4/gG8EgBhFjAcg/bDtXfj1MxL
/3x/b+n6FP3dweNz3gOHHGx57W98L/O+qu8RI/A5Iontpy7vvkbfIXrfZcH6GT97
/7AA0H2jCGv83IfQOb7Z3Z5Q06B9CzMYav6xJGpkc6lSnf4tm0oHUUZQ5geQvdXa
9Dl+lMcJCSrtbasNgRCfulUxnyYQlKJxXvM+MkK50K/Enu1oFf4K+74iwaN7Y8z8
TU/8Uh1Nl47OSx6dvoGtzD7NjzaDPPmbcv3RbgKVAevwPzRca6shGiSmlisTh52g
W6vd7A1OvrFv9x8V1AfUWURtjp+Szr7eHeeYMeZ6QA4TtCSY2KwH2k5vpOMCZ7e/
0tyZY1MUwwnReiES/UzUx1dcfM3gyfLH2xFVI1fPTGLXUm8zqGbyWJXn9liZXwsV
NFKPTvsDJxVjRorVgGaCIGa9uYOwh8kIkJnJy3FK8G32BdwqnlnsdMAgmAwmVuDg
u7RHcFpb0rJiZMo+qiDMEvXk7ieBexJNU1cuAdfyIDStcxjxN7g3hNDULqoOiqq+
AZ9hb24ZHHEa8vpC4QY4XWS6y5xov+Zr36RI/NybQN3kTu5m1uyfAgJOOnLpdjvb
IDCBlHBUNjqXzaIAmrEyulUyaQjVOUNoq0NQij1rQ6cr/2z6NOcEDmDrvhAc1kQq
yNVrr2ZDmUdC0NtdiHeYRf1mQiOQbnJoC1gAvwOBOcAyklBfsjvOMHe+Nc7uhJ2Z
Hsx05B5VGxcDjF3m6hKY0G09yinGdCPZJT7d+4XA8/+bgVHUyTqpwzqFR92cgTLj
X7hY26cxs/OX/rQK4DknyeJG8Hw86njISk+2FKsf0jN/gktlSKbivFhjoI/6FtXn
SgQDGUoqPnEcha4sRCP35esbzffWCigK/xYGOP6P3Noxzi9/xWLvVq305LPX+MIO
56MjBfbt1ofLA9HZbzyG/8u76b8uHhlaHMa0wsgH5RhYrm2gJGzqezXytbqeUqxQ
bmix7iuYutnxV9j8tx9njwahvFvhnuBUPGbl27Qr7pdDNV1Hm4sreTubDxZO4YaG
lhe/hFqjiVDGlV8vj8LJhpCULySXWDK+jVCwcGKxvkjVzVQTVy/DqRXxqVLsKIwJ
ZVyIaXYWxY20Ucq27Xez7QwikKtNWHGazRh7KTHiqIBdCO20mSeNev6nFL+giQSL
WlNCmJoGwpUZw6Bdkrrh775lh3Ga3KGELbQfzpY00aH//xuRv7tUppDJSvbozmX2
xuiPrsn1KmB3RLvV/Vh7aPMZk3CF8q3rGsLg42gjHRJRKbVQFItUSpOF923EZvL3
7lwJe6ELoFjrxL6Dx2AntrSWkCWO6CSGTUtCLwWRpBdx9uEbkHWGh4okh9Jcvdqk
2jtqLmXb//tAwFZgQrq12omz5YfAYyWOsmRld5lBXVsJ5a+ayqUGcK5SPi7dYbMA
zTIobU+duXsxZWd0ZSPU3UBIusCEPxRZuA+Y34bcKtJGo5A7g1oyE8hBoi5RVzg4
ueU20YBvX5apk1L2NEVh+Qaufb1IJoJcjsmLeR3pqeFW7DqJXFsnjnoaaw4C2zDC
cDdIs4yVwI1G0lfY1VHFc57KiY8w3Dhy08XJ0AIYOrHnu6oduWNr3qXB7XBg7TRW
RH149BasPGXdzEu7uLqD2F0YdmFtFI2NVkPxx5aQPUujQmuG5OUVcDxwgoTh6Osy
242Ux0g5G/QjPNjPfymsPN+GOSbsApLdHgb29WHDp5YPuBsaUjPAcXircR4RAWHi
vh31zfA2NOwY5pmxTJFB6c61x5w0L8HUY/d7iVZOxuEpon4KEyXr8b6QI9tLFd0Y
/K9OcEj0afnvgswAoA02SyFRTf9n5ZzdyB/bsvt/YScTHJE06WYQSDeZ+DcW4qf0
1ltKalY8FNOvKK6AuoWvBzI5XGSofcU4I7Nsxk95D659VdSiTYme3rtZrM4bYCIw
+xXnPZQhD/p4S8mq7Yb4Ho1rdsQ/c/BEsWeRgWdRHgYk6L9DInUnRKWlMX7kaOMB
SBTwmVFUzxUKMNhJgnButg2nGkMfA3iFQG3MA1et8d8MRE5ayduviws+8cT5sKfX
lziO9O9ws5tAQ/Sz7sk7+ift0IecJNEzmREsC+W3lH5a65cUjLMS9wqqoVKlna/N
g9SxlLwzKvmMx3Mk0yrDRdDkPnE9n8oAML2iYfkMhJsdmaQytrqMIHb6UFAI0s+F
AUotCk7MNUlz7Q+aGFycN/0z95nQhHJxoZyQds9i3tIcu4dRsmNPkvnIC/BXjSan
4iMDB5d8Rt4f4uuw8XLjB4BDunlTSOlj+yMpdyx2wFeMPxutuZKLB0Ppn2KJsYue
LT2GNONpcdtcSEq3ZedmJOEEdaA4faVlcZVtw137iP3QKj5Ubecz2HcMx8migjzY
WO0MdVWfncy89FX/HlFhvDoUlYUWtTOvbD820uPBe4TOSvubYuc1oi+d1/2ydRhq
SGnWogHK12xqzpQmQOnXjsS2Exh0ytC+8/I3zMyWLuoLLi6y6dgkZBxzdRV4+8rY
yAn+x1Abs9/efrwbAcrMIFJSzoBNEKjTHrcmJ9Y7AZpGVEWySVFe0Tf/8J/7OTxu
hO2jZnSE/m8dpzwtKGqjBUBoJWbTVteV1Rfo/Pv+lTGCP6Dz5M0h5Z8+GpCVZPsX
fy4BcWYXQ2EMJTOo12vHXfhuAWWzg84PBHrNfp54K7Wkh84tRD2G/nPhzJG2Doqm
Y3Zq3q8G8e7t5b/zuzgqPPp3/me5vAgVJN8jXzmIiqr9gCAnjgTNEUa4AfCt+i2f
r2XvbpO4n5dkZ3EwvcYEC6sMX3mTFPTKI+B8nlr/x1Xve3KCffBtanfMOR/Nlwej
K2IYWVvwpoSZvSKx+ozW+rTVUO9Q63217Z5C5OfhmEouOOgj/lEL7yIA3ohAnE0l
zGZD87Ib+w1y4iyeMTH7M2+goqxTvJO43iG2SarWdphRmHpyOv12DdF+S66atmKO
NsiuEElEM1CCw4plxgZ7Drk+lPiSouL/KJZpEOMiosQnh/7nQFpqd8amulZ5EXGJ
J5KcYKjVl0xKZqOiVa4vEp9YfFWai8rodCpX+27FYAHZ9gtzvEVp6gXD1bo/ZqN7
MaRZQGnFJpKd5TcXqlmZZ9jjHSRt3ywxUSOFn/vwbvdIEL7Y+gx5dWeQKi74p/m0
Xue7MemitR+aBt0sqziKJBsA0GTjndDw2cEjvRJv3eLGhIGtvv49fx/C7y/tmA7+
bm6qkra3NVokN6VSVBEcls4qt7gsGs/1IcOmXr9pRIY4OcYrU6D+6s8ICqzXsbBU
7zEpfGBI0x3hUaHYqLSAgj1thCaHSsxmtzNQ1LEqjpkn/EcElx6e8/9p8SzFTUi+
htz8ZpZDep2mddM1TYnMPWA/RUwY03mhEvbZTkbeFCPvgujRcs+Nc6hB7psPEw5i
oKq5vXX8CCYNKaaT5UyvQXv9KB9wDWOqrRrN/tvwsDz4WBstK2u79mipykzosWLa
PJqIswh93qd/LkhbtZrtPRILrVOy04PeJC7E30sY1OPvimEYyypVgSnMfjuL9vXV
da+1Bs96tlbsIwIlJ7TJR1uQrjaY9IULGIgDUqqRbffAd0nB7r4hWSfZe/Q9pcaj
DmlE16U2LogOt7A+3ZDLeHqOwjfMAy2/43LIzauEgPXtTWELkuzV0vNf4se4zwHg
7z5o+8h6agDkfY1tbW5llnr9dNlgZLQ8WWMexGU6Ojs5tcL2TX+vQaSphAcGeVCI
2euD3Y1Au/yj7Y4o/Hd0dhqMJ6XK/aedUPVNv3g28Mz5jCDB21VXcCOmPiXNaiL/
A82Lgk6hl2snTE05qw1IFmoYKDyWNetEoEzGdbrfoF4J3aJoGQ7IEstEi2NXbhda
Hd+5XYK5muAQk9vNeB7sjAgGPowLM/W12DHrs1QgatbxtNMgYISsn++6M6CdYz1e
MIUrNOiBTa/F9sCz/z4owG2Sg7+ISVVE8tFFl5aF6NTvNL/KnPqZLeC9Pb+K+Egy
3vwHAGnCpHFHONrBhniHG4PV3BylyiNt2vf9KbLjAxyB7Q7SzgI0DOQJ01WQD1D1
zuHci0/H1+pClbfMxWqJBMkeGRTJo30si6R5waPsbwSlCL+zv/FZl6dSVuaTHi6q
bDuo7pp3vQFh3s91UzbrZjKs4oD6xld4/9tzOlb8A8Bly5OnqTNt/hphhP6yAQ9M
8DV11NLY7zDkWLwSN/vvvrXqIbO8ydy5iopSe2GpOQy2bSLvACl/aNXTS6CV86kD
+dHlqpjLVJ+6vxuxxCXSePH6MeQrUIbQ/4YKV2X6E9+GRuc7rdXqhlAc/9oHiBbb
3ZwcrFaoIhEi0hJzS9eq0O0KARv+JDuydMXabeW2tt8lLDYgPqwJp+iWwW8fNjMY
K0JIav/rNMXeYFNOaWorxDlAqul4ejf4ZvRmEFvdl2P15plQt4J3PXrkNXPDilLc
c3X0LbEBfRSInVzPCeDD0QGsPHEjvI6Z1vSUKVSqcuRv0xikcbpsSwD73C4rpx3y
tmN8531/A6q1WY9HqbP76ez+Er931sKPpCaxA17gVOI5Sfgi0y1DGUkoekQ7OSLk
k5RzwiL1mUBwzlAkuWSTnXqsv1HiVaGxz94adL052J0bjNPulZqb8O9J7YTW+l6W
ba/sOnnUxWklb1G0H/xcQreCs8Vccq0SJYsMoCh5b3PURevLcmC0g1i3yxFn0g0z
LYP+MPwYqHsx/I77P/aMS/7q/o+GL1KiwvGfyOy9TlNvNDEU6TnvfHIMFAku+iY8
vndpUukIES7MhIhZ8ZIBgCBGvbBzRPJ1nkPq3X4sQWW9GqWqe9wWXQicUlIBWYAP
7JulpnAMg6Dtj6WkZB6avUd6NO3aypkGFFPeboyXX8pDRC3ueA/DKfPHUaHAvnXx
rz0EiNh111hWNQ6p3y/H2WkFFUOG6fsPXHmeplbZ53beo1A5ATb7jtyxQ4ZxzC1a
pFOqCKD+tMEMz9G0eL0/Mhl+kG4LNc9+912F4yW8oMIGOGhtdxESeP07O/242x0t
Reca9Qn7UqsWiL6ULLLOqzaMtoL5V/9fqp+PaGicxcyMKiQqz0qUFmzbcjNFi9nX
Su5dtAYnzD6+FjF0l20//b0quQhJIeFES7mQmlKUJBC9dq3IHMgWeSWGUCSkhiEm
GHv1REXZJzxPY6LeLaRQJtKIVT0yB7TIxhE3ZTifIVTLU2tBrCDCirzDaVQdNGGb
TAXfLW0oru5Ni/Z0W5pKMKPGFEtBgC+zcenauHTMfJ8DTiNTU4Vu4YVFADHXQclr
7+Ks1uy/KnfalY65QcL/ErHWmOa4jh1YFVUwt5fScZ1bxDnSF2Qh1x6vgkFjct4G
LLg47cPA9CWka4lsBHy5+m4tvaKfvk/7fWSmXFUj96YHXt4J1jhx7U2NMNnzfRBC
cW6VfA8f51CNvOFt6K+mq2XMyIXKFTKK9QvCZ3KpjRBdEYEmqRGuamL/lk298YIk
xnmk4685h6jvyCs9spOoBkQZoNTBNISrP30+jnq20JZYCEiqkT0HVBqFXWyUj7Ax
6cVGBSlE6WuVqFUxjvtS9gdfhuWIq05EtUEYRRdsfvCj2dzmpdbOHfkicCKC3J2j
aRnuHRJPEXgg/h400+tXUhmvoSRmVcDHZ34X60A/5/VLPmoA7uXFEUbIY6imqdmB
YQOpS6IbTi2TI0Wqkg9IJdMDvz+XlJ9myLSeNjtBsEX7V0RoWfTkzEmQ3dNyHhEk
o0C4g2PLdSIPWNtNSpKXmPuhG6zQ771HAH9JQKGWN/MErACUK9NJUzI2k/4pLBzF
4l0OPtzNoLADISKvFbyeclNquoeuoJ/BgQ8ZuaCF+8cggvlTrcB7IrPQqJdAuPfN
QwO54+XEtmiUSpET80k/jRAUTX2AD4HJePHPSOcCc5skV/H42JT2Upr64Aar0CHM
CTPvZu+1V25yYqCumQMcu4iiV2aejn4T1ppMgG9I9s66s1IxRSpoNIBiJPvaP9Jq
iQ9o8oSeG5IizMxkoMfIPwJwdeYkyK1AX3a3jiItPh1p04Ca6RgyrO1tSmFNKVvC
G72vGqCRJZqI+w91NuL/8Mw5MrzhAYUH7iFgUYtjopNRxX+KDHtzy55v/8W9SMa4
lcVJ3knaZHNJ4ASHOrbNcG+Iz/eqQBlXFJWvBpQemS9lfVoMc6AND3PBCc8Gs8go
x4K6o9ULEie2Bdd+oEurCdPaufrAcMLJ76n5o16y3ST7Ah1Wukjl3mvoHx7Y1Tx9
CR6L+titlU8F26sfr6ZTdUstAC3rxRXCte6XfgF4qLNQgCly1lDOVuU3WjGKZ15B
Bviah8S80ejEnYitzNeS2Evn99080pSlwvAUwUW9DARTvap4HzbKgrS/hdq/NBqU
q2r1WyYTAmxiCfiH1CqFGPhjLEb9UxTX2R4AC8QUZow58wJ9RkWbcOon3vBp+jUX
eO8mrez6XI+idswh2fGBCLOuc8eZEZ9WXE6ipF3kDMjUTMbFEZT1OS+yGZFLPi53
uuYoi37TFKoiMjEy5ZMe1Bh+omWIjD0c4cQ9t9z5/Xhw6sjonngE6cJ8Km/+gBU4
5AckqkvWRkTc9iy+NPfePdppKkzgOzndCriCIzWIZCVO7pH2VRZ7RNdkqekJRH+k
2BIhBIu8iNaXuM51zwSOXrqKcGFYmTFFkBg+YQ0yJ5z1h4dMKBF3zfR8j+6gkwp8
ZH4PUgiClgMVzzcSs2G3LJY4gg5Z3RncGZE7+JBXx+DgS+LNkG5lo4fg/j9Nuj7r
KwKMtpifZ8229UKVcJge2s8bLP/eKUMiN5Z128d1QOUzmeE5mu56pGawkNCwGVP8
uNQNSGjhb0YvLMee4CXR42T5jvuqa3iYNw9Wn4t4OuAdca2NPSmbR/7SUrh5MWRf
3Iy1Dty8z+++jLOGnkicpWWDe/7xn+tjQBdXm0OGhTUTQdRaDvLlASdsIH6SdPZX
YEN44/XhFgogty3lEbgKnr81KJ35fZGxu0m5hp876uyzPNzxUNGt1widEPH7XOqh
P8p1IVc3AcpCtNR4uxA5AJOrW5t5jiGBR1roHsQ9Fii2C0y2OuIFZNIt6tZWIIJx
3M4F776hiSJe0fNyXkrqAf27GCDdWhOwrbs9Kio4fkNkwZgZQa9TQ6dmrNDvER/W
GQHGPj9H6Eh1OU5exba/vFqPAoI1nVziZczyGOX0O8WW35m2hUMe3rAOjaylAsqS
UHMPLWCxApuKvKIO/W4QlJPe9OiIfBLDDEzyKcmU/nPgvkd6fHEH7DMalsibArrW
xPWGoD3AuNPVdpygA0U9ZY8+njx1TK3cCZyYQDRipPAWQOtwI8MvxcGHVZBbmp/x
NzmJteDyWs0W+mRGK3r1tYVWXDE/eLdetdDoddKIx0VdiE4bdOJBI90GO4V7IjuZ
oAMv7WC0uM9vMT+IOIJeGaPTSs8yHYWWMKCUF9q86omXYnaTiEnMfYv/SFJ16qQY
ux7gsULApRIMbzWAd3PoDWptqh6h6d5U1NcMn25zBgl9uHrFfCDwaKEEwFYZ59Fb
8WHjMBSO38IrRJRj2ZjyvAHMQmH78RaGsdsPCo/wneKdJ7toty/QCdcwbELiS7zj
xhSTUK1N9sdA9XhhaP+BWmwL6fa9eCJJG008zlM/bjP3Hi7y2t3s4fLNc/L9RZds
I3Gr+W4Y9M+TtPfy7Ey1l7oHFmFwpY+X7vtUuLsGii2bcuDkfwFwCaZvtD051s+y
CXsb5t4Jes1FxfyGGtAimCig1Okul3PD2ChH12t7ATIGgVQyzYL4LSYlpWG/aZOj
6wJRnVslnztNBUbYDdJWGy6REvSA1iJ1eEapRRkFY/nMPwVmsMj3U+WBXj7o8UT8
WJBQN6HDuJhJ96ens4bJOMqqMqP6BVaW5d/dVDGhYPz/bTnuLp+dB3ecJwTxE+dz
b3/YF6E0Fdd0uz6mNyE2AGISHtEur3EFdeFR0FX1FXruPtQIVn06dmO59KFeWSfD
8eI2RaY73XBdy32/yQoorv+Eck48XjDh/MR887BeTt0GmSAOSFOMRs+fXgl7Jw4a
aQ2B7MX/GCQUWIlPJ513yji9cwWr8wt/zHBW3bO2rinM416ojh2Aq3rPGYJF/jXi
5AX0BJ3c/nDNl81FuGxQqfRwzShsrn2TNUrU5jR9T74PfgTfTaRtGNEv3KZ9cE0v
Kng9x5uhUqUz/m7tOmuJu0MocgPzf9fi6ZVMziehqw82khq1lh4NkR9PHGrX+0/8
e0nVomtBlL+fKOcSMhLtdPwZ6o9uc1fnTZxHCITgwmDdRcax/HQP1c+Tj8LutNnN
Su5RG2epRnN9SrMV+aWoNiIMCBnKtK94jP4cJjxKwga9fca7gXUjmUPq2shoqMWo
HURiTeZ6Ucm0321bu5xrhvHmgvp/tFcDItghTQJWLF7fOR7Y9fVsMSTmhwhwoLoA
3YNP1LccGvmp8j7El+F49qQfb2fy5xnNfQ5IX0h5Mr+4rKTw/o6K7eh6BZYV0HfV
QoomYNt4w/ArF2nbCNSHX+Vw1eoH+fbM6Vsdqxo0GNZOWivLrMrKvnzt2ZWlLLmp
rYdThJoIkKcgzOBC7eleGA6gR/hRUwtFfZzbLzcECmaLsN4XifPX12bHTBhJyKem
EMiqiGO7YzU420MLcuyOjCziwWUREQo/UXGURYskFqYtmy3JmSIXcoolY/cZ7tsX
BEFZtsZjpxOt3oBoxnPO0maRHBfbTIzcO/2Nispfi0C0oSq+vRW3aiks/ULXcxLM
1maL72pOdQskFIRm4rhf6eOpsjHyVPG0MUNPW5DvPQ12r7nO5oFD7JpdSIiOjxSi
zInkPHghFcQ9F0esFUXn7vqVGToXNJeIivybQ2koRzXZUdzJLksxFP5rzEzdukjh
TZYcT5cEOeru1ba/CJZexsaNVg1eiPfB2YcBLxZpDB/ln9zQTVckSDx7AIG/68X5
9F9KPetY+UVlaSG57PcXvJC8S22d8juCmx7Qst4GGswc3dsNegToHvzftQOC9+VW
mEA8i0OvWzuK1o8r8xf2mUrXh9NXYb2IoOjZeN4To+DGRVBfagvLsBCOPNP7SaYn
Kv0VWNV5L3tbxffeqYZN8DIXhrJJ8IvS0xWk5z04EXF+iNkfQjflEk8ggqi1xSXx
SyHu3RClePdfCidbMyu3dDZp6x1T9IZErePAx0Iwmlem71ghc0ywpcUQPjAielVO
Q07Go30+dygUrmTYsYTkLF9E+gC2zlzQS19R1X7sZ15L0MwROh3pEw9d/I99cDm9
OoRvZAWpW7o0VoqEoLk1pOoiAyS4mSAw8fRzBErsOAo5H5lcI0pyMAwzBfxln6BG
Bqm0Sq/nJSUNQqEEe8MEe3DsSXIdcwc7izNLeURzR7EBtjIudvIDr+gq5gs5e50N
asT8Hu+Q3Ztunm+rAExwum8WXWRwU6ON3yB/1GmbXm27jJaHpibhJBDZNYWHBb+z
JBb/CUC86upjjH2ojpoqXV9BHlcOAzbSI1WsJJi2f/rVLGnV0USeEA5Te/g7MF2J
OK6lYcrqug+Bx+OSJRf28jb1WXlLwJhRKcDgP1sqfJ16JkxbaROwAdUAWQdW6Y/x
qtporcbl1nNFdzwz//dQljzQFCyVCKMs0M++opWMqpPN8aazS5nRdwYQGEIZoSaM
QXVVsu5nuledFVAH3fk7BE3gk+zUve7F2w/QU45AA6r5ajfIbjIQ5HLnt/lv/Cqq
/sAAb2oD3mWdgZdSr2bL2YJ/I+8xjy+HaoQ3BKZ9gKuhRvbky/mSjy9vYF50VE44
uk4ONI7evh6P1fpGJjesbJaVXpzWgBsucUJNXcD1H58hPZ+jKPAAkvhNGqisOpMG
rFfNuFL8PE0HvTqyDXbzsrMxoQpHdVDtNbMctqshnCplLqQs1qokcyJPx5N2Ygdh
Pt/nq1+AIQG+Z8QgGLadfreTCwZ21B388Y3FDDa3FfzAMOH0F1VgBXtPnl2pDvpJ
9aGyKG7nzWwnEDfRzSTXWViKbmchG5UvLOmYVFYXyF3oEPGWll2X0/nGfnmrfdRa
jGvJF+mF/XpZW4O1HlFVmThb3bBHhlvZcOPU93hcallnKgjf0QEZT/pPsO0g5XBH
HdsMYj/7UXskLXrUlRIvYqKXNX+mQw95yf45INTBh9a8098N9k+DMfkFAL5S62YE
N4Dal632PJvYWLdfwBaWVQqS4HBD0AheLf9Wzwg2KF0tIC1G/Fv5j37ZkvT4aCqC
8NFsKQx2Z2oDZWuMIaMiqmrB5WGiPxf9Z4rDMsRd4rojeOXEOLxMv2xZg+7TzwtR
at2gcT58RNDtgE0yG2jX0ra0VsBbT9b+yDoCTgObjbqNDk6gFOKZrLomgX3x0mkK
yDNafLxLhYqQmSPaBxnY/Ou7zkpVbEty3Ak892bjFyxGfq4zBgJGYRr/JjsK8MkP
bvXSUGv9iTZ43EjRuub622NHEZ9vxBviaRYgCMIC2Gms+s734scuEHKYRgLFbrjb
o7lLesZldx2OxEgh/vZn9rum5hImXOXWSK7EHDL9VzKA4b0I3NbvydU48B+G3gMP
Hkg1BTPV2kqreEMgYcBa1sNMgvF+uov1k3z7xda3KAVLvRxxI3va6L+61bNLCTjv
ILtOuoT4Y07WVIgsAr1vh0SAKizH4bbJK1+EZTwGUUuXdCGcLN5bDCE0Dr6oe6MF
mQ2YHYnOcvkLOJvXkEhSz7EQPjt/B1ZWukcQZYGA+93ukzT4hJgekyMYDC/7SqXQ
W/baIHt+0Bs4vYo20KkSmCHIPV1F3PkF9bWDsDPEiYZ4FDbtwOYSGEkVbT/169n7
SpOW8i3G2pO16KB+GMOmuNGIIiAupkF8ZB3TM9u7B22wnGSXvFCQQrj63RmzOvDV
yd41QiGBnSUnVaLBdS15H3XT9cyvRu0elpgWO5qjsjI1fAUpmeWjUqLEcKoWPl/7
ZkOawIUfrbZnnd4tuRVCxGPLacR6v5jXa7S4pRefdwx6kEStk88bNRwlOjXtNAuj
vvIuhprYaCO4rEKnHLynoLcjh/Ml4RnHNNRDbYMLyPboYIiv4Ur5LfQpQQStcIKK
8WA968nqbHnKYV5issoxEU0q+VZrvwOBTAc1/P1BD/pZTliYgEKdNRb2elIgjPWm
W8J0trj9MBSjB8j0dnY2mgEf9xj/kbnVAg7T6k0rFkM8oHWwHFCHfyupiLC6Jj6Z
XdOnbHOsZboxBEzYozQPB3v650ZpX+SuDFlFlnoOWUVBUHsdWouR7QfCltBs+rXc
vtWhMV4PFAzahdY5onoO7O8zP94wnvXaLij37z0vxWbqoa5J4N0Ex1mmRoJWkfCG
IPiPQNtDXocP0OR96asDlGTiPNMs38rP+2NuLHi93hygG5NzxeeGPUaUatnceASZ
EJ+rD94oMCJwyls8TzVVOhPXX6Tr1qEBrWk7fbZWew913kY4X8MhkbK7OvS3BOrC
A781aDEViQacn2vLi7F7aVItrMEu5E2U75zvFcnDNIruTX90uXUhg46+iVDq6hVK
84qIpE54ly9nkrZvyEgo5u8SJE33hYFR8LYfbeEei4vU5m4uoaTSsi2MAjT645EI
6HPLclq9duynOEcVnWR+8/L4pwIaP+nYB44ByGRvnWJNmzxPQyuY9p7WaJRpaJ56
XvYWc1JH4efAfkVMBcwbZrvRTcpYf3gU0diANZx9zaDR5f6Ex5bQGVGCeNrerSvH
i/hRALHLpGJ+G/gswo+mzh6YHx6Cb567O168lIyAzVYz2jeNIx9XSaP7Cpq1022O
3AmTeUPuCuMILdnOa8SJp9AQ6YmDMjxY+RATdVOnQL6sw/0tw7VgSdv7WT6yScJn
ESOjW77rHZIYrBelEHOMajbvgb9bSHpyXuAozF+cezhT2bH9zgTiPMF04sNfDNOf
EE0dXvGlhAP6kFz7eMuWiUg/oyB8wmGmUxqImLczYkbShteLt4dlkWRBmqk7Rs0J
Aop+QaDcYJYehFHmm54iFfB/wAcQLtavfXh5d54J6DxDIJcERVoWryC/Fz93dEPv
Z6MZfv0XDtQhxyrZQn5iyTdVhoRqOFt5IyZpDNJ0qxbxukBGT45iefCXZhXPruc1
VRuWinBHATpQQOkTNgoiroNM0xPerSJYx+l54ZpOIwVE9OodtEMKfK1xceJiPZHb
dBNOA6YzxHA1MSZOu0gEOOLDz2H06fsAAE28fy+nfJOJ5U8IMYoQcePKJoUvMngW
JgLLAn/Cwk9EPRgMG3PYLnccbG4bPwQSCxf8+Akt9TUz9cDc3zjZdsY0LDIVx9J1
AgiJIVgx2bvFW1UDmQCwVxgyiBlpNeh4jb/2aUd1E/fWWXOB4cHr/IyYhBtax845
r8Q3Nx1Q1m4av1s//LoZYwqqMV9dgvciD03hmdh3UpRpbDC77muPS1gntJjtZ4OE
3shmqK/Ys+Aa53OjG/LHkDTyv3zYj2GSxVWrI4USFPpavcpjEfCzsgV7sutNc8ak
w708ib/NjF7Arpyl7I0+gC2FW6pFVZQN/ixSlruR1L3Jpn+d3vgQRz4fuzsGnB0g
mb3EhnL1kEUlv4gAo22PQFux7p5/htAR2D851T4k6hWCGbCBAjebAC3RkSdAQX1e
Z7LvwsrC0jq4H1KnEH8uA46tuYzQR7saeCq34veq/4d/M204KX2UbbCOLnfrgiws
/bln/QFhcOGNO2ayFHS27x2YdKwkIxz9RkQsyT8lq/XpNVI+5PhF83CEci7MsJ3d
pMSUYuHtDZCE1zw8/52BF9CAWavncIk5elQXHL+OMotV8nLN0FSaH9a1AD3tyeHd
hlCr+cV5F+wYexx3tGIGgq29yAkNDFdmFYAgz4HDME/Syo/0xbJ6KeDSDx27VolB
vnhvN3lFsI63zOwCVc/zSKz9N+8bQc3b7FdtgZ+GWpxAexk8KYWHY8OZ+dL+05yM
bTU/z/GMoQdt7Vv53gBKsoe/Isq2vs5gxg0hjmKTrydX8Gen+WNSzfMDYtL4EyYI
L1yrdglVkk/NHguSgFLg+Z8fDNl1V09FIdaFTku1NV+vvuL/n3cBOMORfRLZIdyF
Ju9Xe8wi0KPOamI7kx0V6WT1nzZOGJvE+sfzcSWbanrFyscQqO1Zu8uqih7P3Vin
fvnTsG6NlC45zZ8V+ANmOYVzxO7dxaIJi2ZtQiwfcwZyh1ak0wt/6bkDq4i68BLU
QWUNBFQZ1XkbDolHZS19JSkzERIgKZqihx6fBQ6RSHvJ+se+4V2pAzjrch18KETp
3KK9DPI5dbelseghVNJ7LOdLDQW3z4Ga4B5srpQpWrFzuzqhZU2au2MwvI4AZPxZ
zRUUTB2BnRpySyIcoUGKgJaEQ/YjrB+rlLjPAh/+9/DEqP15weW1HKcekFRO5qVE
e+7agiLWNsPTASiVzgLsNvutrpebyjSKK/tgNuTeKb2+2G93+y2kub0dWLvxBxOs
jfqVr5Bi4vJD2yig7ql5rM8U7A3gMyFwL0qTmLuaAKl8LY3uEHctCdxAgccVKFYO
FoYSnW9cpPq9O2KaVJwAClocIv3MTzEBgB8e+QworkRzlOEK1dTq9uz7Y9q4GfjJ
KnrdUqavwZZy3VzsMDnhQTl3afSO4flJWaAP0xFzTturvfbCi8mP88ihiynilZr4
0ewMh9499XHk0VhHWybC6nryMi8bKNzcR1cWQHjZ40kcgcAKcyag87dHT+JqACZe
Gk360zNc94YXMBTXYIAeEiixwew5GzNfVPpSurBSRzknBDSCYsn3xADia6D7A3V/
G13boTo8OTaASmUD7iVpZJCqcgiKMv07QcPOJqzLgrPOXWtfzBJ0wleNgFd2BZL1
P3/JyvGQjTc2vSRIQ2zowqcK+C1kliUT6XZpk6es2zg1wshrIuQzvpvbllGiqAMk
AiDbWBsUnic6BvrM2jbsdEDcCdeF+dN5qOdBc9Z56BK4YIpTB9VFkmWoM8pjCgZ/
HYG0Vlc3AXs6ER2Yo+hr7ABvqqgUsU64mvE0OAjJPG8fZG3HVhY84dA3Ze62BzFy
2wXhvjSXUs1B0oHf9vWMmJO6z2vIfYjBgWKbakImkz4hsJvYY1XgCklyB0XVSm/J
OyGvwxtComiBEsg691s9lZ1HzhyJTuiUj3Zo97F02JyB9oypzifUBYU3O5wBKZeH
B23/1ZBy1jkd9AklvJrXxAh/n732kKrBpW6ALbnVdCRFtYoHWy6+tavDHXf83Xtx
Px4DnjQ053lmQ6jsWCr0uYxHQWVjf4EsYAvvAhB7wjdkX/S587t34YhiiL8UxPkw
fULOVfv2LiDzOSthDxgmahjg6o2hesFeVga+wZRzu0X9V2/ZqskGsOnFk5QzOPhZ
mLVxzJ/2Tgzb2hsQgSaZSizeHMkd2622iwZPM7xzERIQlK/OYWEv9uQI2WBVAh/X
wZkycpx+lsdOtx9tU1zvmjjVYVds+S4PSCM8ILLXKtwQU08b2tZKacWMNIRJGrwy
w7X230zZmwjdNgJXiQSz6ib4Z+8cPhTtJ7NuseYemVmsMI2qL4HF8go1YRaRgq4s
ri1MhDXOOWYQerjvR6PhEOEi9CnOguSLgS4A8Bv7RyuuZPzYmuJg3vsUCBZLl1gK
uXVgTmXvCEu8XSOUAu5gjjdXPGWVWHqqZH8OAz5o88AcpKls2yzAMmiEgGCxvpnM
FnXXzA/0bdV/M0OUdag8vOaTKPMW5BR8MP53JspjufI8Rvu2kmrFFcfuyh/MRucF
Fv67asvBFpcq5yfSGmEAmh6/EAVxj5S7EVGhLJ8F2p7x2LZjRht1SMbS3x1uO9Wn
stnIOuZnq9riIiT7a41SpllvzSMCcki3iEKHHuQ2n0col75tW7hx9CQFMlJTRKp0
PJZgm9qplLbViSDLOBVVen5VDVtFCEh5hzyB21l4cDtVocWTjMCwLd7EgiwOtBbM
USuSY6tXOpifZP2F7JPMvSV5RfmFjk6n/+cMTuKgtD/clhBj5i2w3lpX16Gh3VrF
WMHk1yKmjeLCuPcmwLzDMKui8to/jFQeUh2yIxcrtvPlZXzUfrnVPD0/2akPU+HE
C+519Qls3F0azBWyxN6lsbMHCrpAFm/CFsEBPQ8iXXkH3cTvTZZUzIKVC6+KmZ+e
gIdbVcl/52j52aqoq0yqqXU2tNEc+vbSCLPL+4ZfA4BHKX4ugB+eKLdA+3RcUXOs
rgpld/06g8vTwsgWtI9uwLg0UH8x8EOL/iNaAYtR7G5rtsw2AbkOHd7e6mOZx+4m
w+sR/S3iaRP95vO6ZzhwhyKmH65bkExayWnSe8BZyNemmwXDDXCEJxUMPgjb+GTP
rT20tu+3UHTq/i25Xx7BGr8+jES47grhz4Rs19DBDNt2wzfoCyj/AYMyvN0a7qAQ
djny3Y0LFSll04KD4v4euduDmIajXVgu7eNqbWBZY9YhbiYzIG3UdRW/BT+wck2H
Z81YgUJWh8O8teGqUFbdg5Pp2HEAfJ8g0R+YOaLntelRyEOYa471DSnYTRdNQ2Yv
5kIJX8WkyBLGo/wq4ju3mVm1fv17bxFqOzzVLtsnonKtLBcW5bKrug/yAes9q6A3
hmmWW94CMkCWDj/QDJ/oSYOqMBH1kTmW5BMkahc44Eho4L9ulYrYvUoSsgC4r7iJ
3y1FScjhCIi4lTCC1JfB6nydCz1mAdx2NeptRc5MPrdWYUq22iqwIbMPoO4vDPWO
rozCsYnFUr3Q//E/MyvnNhxpB7UXQoydd3kQyKiEaMc6I6vR3g32WtJU8cQQAoVH
KD2YyScMW+cSdRAFsTbhGXtOPbE61FMDNaFBmdKrLmQRXT4zJfwV1SPGytXEH1Pq
4oFF74vfI1nVptyXnu99zkiBVayil7k88cj9w+2acsqi3RgyZzwMq8smwW7+Als/
7kHDT91ikGxDEzSrszDsADqgZdD6dwwLt5zcMG0LFxrt/gY8VhnmxYEjz3BlHRWI
hgbdL7/Nmoce5fx8du2ocUgfzdR3qMBcUNYDAWRtscIXKtcRFUs9X7jfTMCO6b50
tHs5rEGD9KyU5avEwNHy9DpdiBBt5DjfnVI30h4UigUVv4pbeMB0Ulwe26KVC8fs
Jfgfboyc+RqeF+oEYaVm4aHc2xY+B+bxDC4ZLfzmAHBIDNX/M+m6EDEM/6MHQzbc
6KVZfdxKxigruGFc+WaN1TFtpfzmyG0+rcslSBGWm17he/HNYQ3IzXWtVXoexrk8
QXfYGr5nt6F3xLzc+S8rEBs5TZZ957F3fqrdYssLe/6uToPXX/brVbnzysYZKtpP
6YH+MZuH9NWDbnl7JHCRM0qfHi+LLAsenbglHjbLOltAIU/xTQwlZMYXi+7VfEmW
gRWq2KNILQdTE/02v+6+sg1rbi4rptt0o3EAuc9t2VYAVjgaFZaScUiDqsY6+q2X
l6qD5fcPap6qw8UXDDEWCZ2NbHURHLAjSoeXDQPI7GYsR7Qxl9QLhiUwmWO7Xkm6
QS4IUN1+5bOF2px+d1C42e4o9oXkL2tHC2bCZOCojrjZW7cApgV7FEJSwvmzlbF6
YfVJKMSMdrOhf9ZZKUsVHY+PWaaZCUv6yneyFrFiNcuff/rdhUvXE5t8MFoRPi66
CbriL9gLICm+74QUeKGKbLQuvHzy0c9XBG9X6/QG7RWropQKFdd4wHY/CD7j1z3C
7AUBHmmCp/2Us2B39n1/2v8l6GXmas7AJiIPgejWlg2T6jYttw0jYgE42PcCHc6M
cXW7TzFpGdXXP2UU8l1ipB/iLYByQwbvEtwA+Mai65CwHaJvogTqKuMiCxc/7CEV
RLx+45okvobE1Q3fuavtp+lwdW6HLGKyZKBuLRbiWcoqvLkO1uTbafjqrBmSgqbM
Ulq83zu7XZBtAyN6sc6nWLIOMoiTy/5jeZt1/6nhexEkRhs/mnMxjfAuOSx87lJ8
uXYl7T0sv0MuLj9ug6njRfWOLsgFFBQfPZ32rU06A3Uv/EwnKpdj1o/Hsc1yBNdZ
ys3SS12HeqkDd91a5Wrfh+ODTPf0IRSm/qxxiuOJF3E6FzikfYSgrDAK3i6BIiZ5
5ENVWxnEq+Xh46lO3ibGPkkpNSLlRAf4nymjlACMEa+E364C4D3okoEplghYaoqi
8SCqDF0T6JWCzJMB2qUug1YICYIbnsiAwZ9kMyMSD2SGP2OFyGVOOq+0gg4vEFL3
yXTLYGXnxtXJjUF2oQiuhzChUh29mDmJoYAMMwcAD90kPk/uJKTraG0Pwt2LciPd
gecnM5wa3+SqoFMDB6O4YJfX92moQynnG6tXX03vULsOkhQjhxMa6Q8EhjAraaBk
LTFj84/NgqRBDZfVD6JdmbTU3ZZA7uYT7oy3hv32obYsd0kPoXnptWlJQEnFeR8J
3r6ByYCWYFRxneV4X+IjdQ8lU3pW0MbXW4Px6JAOGf/uexT4Ce7uHZ1UTFmSYmmK
dnl80zFWKfXWiX/fz++QMzWyop5+CilRClS8p576+jkPfisgT+olx5+P5wG2L6nT
SR0GtHRFZi1lgG2adTTeoo+9OaqO21BZwSI/rL7m+I/AHUyMnxMYigunrAo8AquG
+hr6AAZQDE8+JHKwroZ5ewd+lNMOC+Xik1gzYWysJ3kx250Fq8+INC3uj+pVz9h7
FvUR8a0paS7zEdQOTXWFvlcPquwfLIzWZdBsP9UKf5tO4E6ZJz3jcp/ZzGzYZEcq
5Jql2KqGWxNaYDLAbUUT4DgYkYVaKY3JMmgn7k31krNQO399cJA3RCYwpMUl2ISg
s2BrNNuexfHORJFRMucZQQKeSy85RLJfT2bLvIKGTNLSNUExNh3I4TQTHKPvsM9B
NYTJeI3z75PTp2nxEDmzuIkPFwfcph+xZ94fL7b535A6F/oton9dgqJZ0f72tAvR
k7mLm51KOr3irESVia/lAsqQD3YsLn/3FFIzILyjAeceaOkJxZ+DFCaVU2JUbPkM
87Mb7wIMu2K6tyPWdMihYpWyxSWMNGLgFL3xp1l5C5EmP1fUIVeZu5fsCYBjP3T3
/Ryp7Q488iX1CtSYJd8219H10pRLvbV8RU4B1e/kXt88o5Inq7oMiIvQRLR4wOYW
9N1W49uJ4ZhsqQsHyagsN+rfauXJiQsnQ5/52baRcLLiY3u8P/dQ0396558SzyM6
Bo2GsH9TCkC/PAY6Z8pbSJcJ8XPPov02XYZmmAmMCmzC3mH+CVJ8ZCj1hkYCemuC
6Tw+xzd65wUXMaY4uxznPdH6Hz3gJxVLUhZkjIRPvmDH92GZo+cx1FJpE0mmfq/m
0wVx36F15JVK0IgJJxNcSHca/kiSroyZwGCWK5cQwRj+XcomQE39SOvoPnlqUWsV
PSzcB1dsLkzJrE9T4DZpA3mSIbQUOeWZZyEHOVPm3t3dXh0u67SFtnJ7jeFnA4+6
zhLkLtXQnpU+BRR8QWysLyccxK4alOkusOYgi+9SE+LZ7/a+xoLs+exDdvRYpyQx
VGMJpvr3KvpbnHbqzULvB5/Snl4KRW+hNizCofGc12+VOAU4Dc9rS/cxxancHNUz
u4KwtskOGkvIAig+tvvGigqoSBrJ7D6BHcJ4P0pW1FQBUNXFseA4wQT8QZG+R/Sg
3Dg3M5AUKe0zNKc6x4mzb7uVErQvyzzlgBJW8vJfkfAvyuuWS7hXF7UXmmKjawLf
B8+rCGWO0gKM+eKJuEn6VFBCPG9tXxUhFpOepNRU9moa2BT4URUhoyism1iRgck/
MQlqkmLtz4K4XU7bfrZj0fHyqNqxhi6AWU+A7q8fjKh9KCSZEwhO/j0wskfMkWAx
0zitGi2GmoulBHkRU62ynUpOBEoCsEzICFMSAsN/f8DIMz85FS5ICn/Z85gs7GK6
+vBXjECX1xoF900Hnjp9EaYSSpuaggUMGPhvFOFyYSX599/OkmEWGvrBpFRRT4j9
rF4VUOPKNRLSu7JUjj0Jl17NKXA//DQ785lS+cANMLniafZTiwe/UDNjG9Yom7Gl
juMG7pXlBvGCfhTN9pFprqCu4yZZyiAopOgubcBM1Byn9A2MRxFnp9ZulyENAARs
MSRhaGQKMdF4iCFVU+lrEGJPJi1jEIk8vwIElOh56qEDU25gMAjDByvTO4M+iTzE
pujzXhbW0+knCV4hCSBUL4PTuy9xAfkQ2ROHqevs5y/RQIs9YLQYFFdMpqIMH4IO
Pvhm0O9IWvsRsYABbZDpHk0UboLV3k2V8Df8SOM7TWjzi1/RYmglxAPzWLnX+BVr
yANkwHreIIIFmH0FiE25OqP0LdFzXB8n6R4RugRxK0j3phHrKZSmb59pk8rSUNMC
xqBpLxm0wcDNEpIAN5xDQjNQYVIR7c9k9qJ2QGEsUC5yv9TiCNzjPXq28TV+JJ2e
mVNfzZJEH9VDWEnOf+2aTR9MY8wF4BdvjYtHi6H6ggPm7KlMGzTKWr/9nLdDzKgr
ib8+g6wtaJ57npjIlolg2zsZvgSm9kFtewMjUQO5FUBkahROWfI05z83/BRIW9lK
Dt2N2Fap7m1xfFj9L540zyizc2hEMbkYE2hIISpvZ374J1ygg5PV/uFH8CRg2Ka3
FlWiZO1mLBDSyZaZNEbkLDt1i6P3qXig/APD6l5Ly2OMXKIc32bfRvZide63Toy+
jGaYDW5HDocz/9sKrYW6zmC/AVVui29qekvLgKEXGnQ8ufvxGE7dslDTjiPiZa8X
4BCZEmiJ/kaEAovvcifDlalJRYiLxSdzHo11Zm14OfT9yUfbi/sRbUFFHiLafVu3
PfiksMMRhkukXV4EQxebMw5CxnrnjPULrJAO/bgMELmNFrTk6/UgUxSnWaMGRKaG
c7jAtQPjN81tS0ZAuVG/Zb3yYB1YmyyZCib9GT5Gsa7TzM2hOqAOWZ76VX/NyNXx
LNspiY/91++JrAXiYvLWFCkSAmBA2g73jpSSRA4tSxo9qvMI8+1P6KKfw5QsUai9
55dK4KmcVFUhlCWs3Yb+28iEZNdcUNwT9qiKxtdKS/n29jq6PSWO8ed6pmZI2og+
vye4yd04Z3sko7+YanVAD1CFaZYrF5BcmytvMondQ6ixgKq9zI/SCjs2vc0fetfm
ni3jvdI71VmYsDFk988hVe9ATtTfs2q/TTND1Gp/FMkES9L2iZJk78At+LcFuYcc
dfToiK41GX40kyncVByR8Z2d95wwpRECEzT4jDjcNSKUm3DK0ljSx/U6OsLaGuX7
/fUJ+lHcBR9n7OZ2IKltzAa8j4gGHSKrLf+i1nbLfGJm1/6aEMdi0oBNjpC75Z3T
6/oemYn2XoFYSHFocaN6KlvR/l7tBNPZcEGcwg6yrZVlSOX10gdnqbod3aoo+yT+
bX8Az3ViC+ROhkI+jZ8mvmzKKrZeURCxRy5+yOBiVo5ZZmIkuts0eZYaV2WM8yaN
hQo9XxRFNt6N803iuf/MpEzvJ5XDK7AOTSBFoAQ34zWGpXBSEBfRNxIbzEMNsNni
HtVa3kMgjfOIwiqqwvjMzE9m5zrxmOFeGHdTkimdodndvFjodqAv0yj/nlnrg3M1
w14tISOKSZo/5eoH0MvIshSfgrKRpzvhKDwCxTbQzpj5p9o8xUuneo14ZD7q9Xan
r3qfI3DQtYiymOxIM4ufzrghN16EVqMMcCikCNg9jRX86PQVA46nNDDS4pJWdAJY
ztJTgVOAzCl5CtfpJzV1gVZF5OTXDbJMP3W8dSuw+QCFva+673V9db70wZzA/qSh
9VFSsUOBfTbJ2rJu1GOgSxWP/g21RPlTSGw+sXCB9N0ndMzygNBWehelfpI3QPwW
E9upZnIMi8poGhjR1gWXEHVEBHp0NiGi3GBrT7a2cNlJJuHxcE4LD91r1hpBdyS8
a0V8MlSQMQcQyWURuJ5I8PHSF7MFs4vGsOHORbQSj63ODFzNJk5z8OPh4e8vUmj4
WtTPUP6CxRpJ04gRtXxKeEHwamQTgjGXGcOXFDE1xqlRmSguKGx8FNp6IYZ7DK5h
WVd9azElhVsZ8PvM3UdDET0oO15l09mu5lAB1iyWQbpj90KJQsdVvcWwx8iTxtnI
ETOWs1VUnW1mkbaaU4neHxaNh2AzRudq5AmE/8GNgfoUWeFv4ihbBwiAeOWOjuT5
4M91aMpaI+shegijPrS7w7UkNXEoVTBC0F/xEc/HIW33c5LqzCnayTKJPcyoWUEW
xatEH/VIvAL79ymPoLb00HkGhmU7s8mocYbF6KW51OKYPNKhvyksg39ldFty5JfO
DjwwBY8b/sprGoVSlTbR+3mBc1GPnwzZ5GPiN2TBE4ZediZXWYDRWEF7JOt9/TKS
yREQ6DQw/7Fz1xuNCXdFKilHVpI7uhYmFwbMfBcfOYB0C0iVCp9+s5v0rLDqXN3L
rQfX5ZZjF7AhaXSZwUpfsNDQMoWKIa3AY4ajglGtAsnp2oHy89EcXrrhZha1SSAp
97RoWkmxHID3VJSDYEIoVDwcgCE9XENoGca1SfH0mjKZO+0FqqbSJgpxDAk9RzHD
gzvhrklFvW68Of9aUX2UkkX19hnNNdKA9yKfvjvY9LoiBBCo3LVQLWOEDYa7Wfn4
8jrfUhWw+v5TLMoxG4etM281gYdEi5MdjtU3ggNIpvwqLdTd+XkSfvrH+zd7A2Tr
QRHBFG5ANSzgIGAl2ZGN0VwBxHZOd0UNvbbUrX+1JfkxBJBykIO7JfWz1dWX4kBi
B/mM1ZmMSV5UuNGF2to/pRUQj7b8vWm8dxFeeHMPByirnEEfx3Om6sP4UPpe6W0E
qMD5qsYbOn8p2ObY7Oymd1biv1qgO4JfliIoqV8Y7W7Jsyk6FsvWiJPD6bhKRbRN
FA8GlVV4Kk2m69CRwkn4dlJBbySV2WrngJV9BYJRPA78c3yldSoqu4HnJf3vc04m
ExizXm1hPYajnHhd2C+3jFYwBSLdnfvwIETO4YA+vmCuR9VCyWgG31rMJR5v01c/
hqSHce5QizRUtl3iYoN3UhBsNnjg42UcIQeTp8003IqkGm6xXJiB5xNdK7ESFzlB
V8WuPRhEB+qUb3V7mY5pm6BS/pFXIWHAqL3gWR5ICsY2V0FYaNo7rm35HL5O0coL
+3nRgjgPc9KzW6BofOd/4JjBX1/KTH6ZTDuETjSxYiTZrLdDl1nCdsn1KGBjDw13
YjQ+rcpElZEkNEkQvfLIFkCVm4UafoMbyAeO/6G08/yy6TdAXJY+yuDda4OOka6h
0ErJQakJARgyMEpZ2QR9e2ngqiN8oXGHqaqJyExrp5shnK7rq+5Iir5Ks3HOi3Nt
tx/F31gz/8AwNw0B8XaPAFU1ACOdy+dEdK8m3C2efpNa88HZYVSB8g+U+emV3CeV
TCA1sDjFNzl7PNi0H109kdmK1BU8fgzmPjdraiTimk8OwoAS0PZ0bDt/hPSDLAIC
qotZhntWa0h5kpSugUKSwRTOrYLjROoeUJAzCHMbCNmfwMUUlpg4c4faHr3mlAxZ
k+RfeNKpkmi+G99tIjjMyWJ2hf66e+qdwjqKIZqI+F3zUHDagnF2gOtlJ6i7RqK6
njjp/jaHesAJm4JMZgrcf7nCm5Eu22VA7p8CP5Q+r+ZHlbIGb18DMrJIhCFLY/39
9hfC/BlsBIOzWgbwoHIhl5KyESWxLvmP2FWrUen2tWr6YbTawglQgs7MOWmUf43S
d7c50X2bee4nCJ7JoCVKOD2G5LIk/yj5YLHzffwP8IKDW7mMgPtwHyxCX0mNfdmF
wMcraw3PkNIYcF+5PW3vRpLogJaWP96nfNDhehCdIF1X+FtE+UmSlIX7QROLyMnO
RHfnBwvJ7X6aiseMbvpUAIkr4SWUvqM3oQ7qBik9L43EcLZ3evSUuquSHjHJoLay
eAzoIH3BfGPVgmqvtc4uCCnGeGm8NZJNANsH+X8jErYkqadXE9rLV6yMoNF+dTlE
V7qCYc2LjpHiEc1v8OgUR7HVwxOUSFs6UJ2JH3NbEacx6pdBSta6YdW0BXdK2c9n
W4rCRd1PcR6LvccVGQ5xuqPqSz1ftWLjzgod9wII5Z9WlOhVGdRcTR0oTFFtqhoZ
3U2K7VSM/p0IadpKtoo5ELLaIZokALxOEbdCEzzRxqdtph+rMUqcZlhbAkESuzMI
6MQFNz2nlwCyOBn29tDpdaQfn4S9trjvTZQ7nw6gvXWT+Jk74Qhr0jCbe9uQtxK9
cT8GXJgADJdECDU7oDCjtlO6SaMkyodnVAsUKbP9wb8uf83HY7erZrbVLfPvaUWl
GU04+RIkW7fMFYNcv2zjXLMh7/wMik1Z+E2Be3HCvAKkC5zYScmAorBxhqPGkfeV
NjaImJm2sk/MUiOwRVQAIj0dMzZDzqr45mCJD84meTHSbu34uETGcsdZ/QW+SAIH
gz63DR3788JMuYXi/8H3oeFSA9ySG7xgSQyfbXrgacobfGCEjLi/w+N1r7bztqal
r15DrciCmUE+if3lgSmAsahsG9tA97V/ZBTpXSyuGymQjTeE2eHW3Cc9cD936z2x
OirUuxO9ksywKx2d0MmlfTbEB8a86FATcG4eLbk0DqdWrcjBeprRP2RZ9RCIWzSr
f2MKry5A/nJh4XbGIjz7x/Nljr96o73en22dkvv1xvG2Pv+rvsT4vVXF1TDbUp//
x/vfPXEzEvRjYknv7dmD46D8mI/4xFAqZZ561JATRKTkKXvdHKR2AeSum3lE1Sal
b8QYaDrf0yzeZTlIAJHDCQBXSOdXksauz/LkTo6S3jbU0HGWZ4q4DC290ToK3qvE
aUu2ugsTZJVvmlSn6/A+fjiXzTAs7IUNqKAnzfhsXZVWhkBb1hHXKaWFWMMDqQ0I
2FVcDzEuisNl2lyw8vjuhoJ4RBVasc6vAjQBwRYy+W7iJx+nN/37Vy022suDsVRL
6M/zTSg7wse2ZyUYmYD2bqYs2KyVUitFIsFcAeBUDGga3mkZEoY56NVe+08aLwM4
q9yt2YO/oFY0Gqa3ieuPosOvdXzSCKi3QfuR0GveduE7/MNsvuksjD4hmCQEpEoM
ReAT+7CijvvppdKC9CLvqD652d2YygytQ+PIIELIa/8tzwzHi3SQywy61rY64i4T
6hfa5V+fKeSdOEFwKPb5DwgZmkNIJ4vh+MKA5W8YQIR199cSf7kAh0q82DQgZn3I
m5Y+diHyvap3v5P7DycANtqe2f9eRkg7Cz1Yl3C7GDV9iJmjlMdUkdY9jNMQcKxa
LS3yWgttRBgAoCkM98BkDwhciL0+hFTUFyj+37pxOkk2AJfWeaNmV/3mXLxhdZHA
5vsNPCw7QJs21CfV44/BqZfWPR3Ron/sj1o7enV5wSoX1hYVFUoXowPn13JKum+c
6RVMR0FSTYIVsJrJeF1nbo608kbMoVu3f6Z4rBGr5p72t4TfZOscSFefQF7NQjsg
2ACt+wBFSKR1NwA5I3a+o1wMOelZoPtzxOsKylH/qmCz8FGHtET51tEKpej7VgwO
uorodfKkpg5ngV+Z6pOmls3tyrsnRHFj1baozozd0SDVMm+OHpbmFIM1ctwJu3U/
ItOIx02zy7fHWxqffjFFiYZIa8dEL1twoLd2vC1R1OPKOfDHx7zw10TW6rd56vfH
U+EMmP9PbGMlTMTv08RNMQF82d9Qc609wfM0v0jpT+fqZOzbm4Ane8xij7yYHdod
kXExJjBQ4TiOi16wy5bc8tZwqRpJp/38jg/U7S+mo7GGX+eY8EVcGB1t+3kM628i
ZnaDKV8W53/zpu99VF5jyuaKmJYrTiZ16P2ml108BPEENKXTvSY+bW+uzM0pid5Q
uzz37hrR3ihBf6KVsdeiP/JAqXS78lkrvdZZxKGVxBbh4BZEEqtad3Zwspx2dzkB
wU86yjBZ7LgIBEtWvmyMYr+tYjEm+DS1c2Ze7wcIBWQa/KC+pmXu4uCWb27RTHfl
QeivUYbwetERaVCBaHkzcZK7ix07qkSnELLmL1gF0skg0G4bFOZMS1753iOJXaMG
KPRKV9kZFjw35+ZSwNXXGFMb2Fo7zfNcn4TzVmcEh98+tKHdrfnqMQGkx1W5F83Z
6ankUn95iy87kcg69G689UE7qLeeYlyPITmxltvqv2LPcGbYlvqfJxYo3ymHUi2Y
5ARDJ/pE8nF3dniWVtD8uEw0uL9MTAIpdvjAljVv6iadUrQEVYrqxJA/ov8BacRH
1ud7KBJzA4mfiUBHaQZ99PCdKk0V3PbpQME3sZzOxX9ds8if8wWsDtrXgI0X5JUj
7KKvlQiiyYnjeOY6NW4Kc6QgS64BjojB0EvVDwuzeny4GVNr+Cg04hhWFXL1Tmr+
otQN4DwLhD9uPjh/gasab/RbY0bI6CuWLvuKNExsusETufMA8pvNeKpCgavGj4ok
vYNkBidaGH8zmiJI9A/fnQO7KwOSpVINckXlEzIAYifZ1WcPYeAoLEQQiu2Y/WK8
sjGaUtyHhU3SdMU6sg0HaOADTtja+H5Ue1lCoLczsrA1CcsQ9KNco2F6nK5XAo5W
3qYUOC+fr33JDs6T4NO1UwunydsyTiIvTJCtYEMPBtLvlxjHwIDuvi5ThtSivXgf
fRiWpSghbXm8RmoopX6755XJDZayGYeKcBB0o1PobR4Rq4ircrlLY6k9paVu1KQt
Q/aWJQHsJNYAwQD1jT3Z28vRqKxrD3qJ/ytctGkWlxyyAuZJr2q1SelLc4aVt/tV
Hy8Etlp9eV9x7WDF2rpZH7fk85AdcDiu2CF2O+eIx7xrXC2GsdDD6z9Eky2LsvLU
YHITzoNu6P0vrfHezrZhwzSh8aGb2fXz3nnvxeliecmIuq6mhjTmLdphD5gxlLHC
9cx/cYFJRUWLyaAQjOrguAe/IKbfxHlTN4PAzSS5Saq2Jvq8jQkODB7KMvVOFMtb
ckp0ufvj93c9sqQrEbnjJL3ZehgEIJvqWdzIPYqBdzaEU2SLu8yKctyVLZNS01UW
U83zm7HOos+3IO1SOLIzl7SQ+Kd2edD0di8azanV0uNrftDUt9H0Ln9q9+yMpLb7
ASkoud+v5YUddUfAei59YhFSWA9doqwQvKhQWCjXPymuy6816IKdODbIux53PWIG
aKbX3r8BkFwIGwCuIR3/iIvhw3cUJZc37hf1Zlc/RSbxp8Gb/2nxThgAsfT6HJwP
yjG87HTsc7bb3aBJHUOvPx1lWwQhpnQQbKkp3MMtOmZFkQLWqoyT35X39pNpDzBZ
gjWmsJt7Jd9N0ekDZ7mDQzLHnSHUSREbjQOvJJ6VDfNSHWihlfd3wpsaONYcENmC
MxqsRHCsmjJ2+KztYfrY+2O9g4VlT3SeJx4L8jV4mjLqQatHqTS4FdZyzg2mlkbr
V7Mf+bL2LlUVRtyGUYUovkvWJOme8sr2EVs0BBeEozLDxz9PCGA+T/NMQQVigl9p
NcEciJS6LAnCC+0CyqfNGv9Xr4eDC/iivAYkI/SR6B5GCWo4vGT9tUZAxzb3FkhK
XG3jJN+achZ4DtrNYd0CGdWArgh7p7agFUnYpwzw0c+B8J2QJmGF0p/PV3VC09eQ
MMiSYWVo3giE9oFhYxnAYmrS9XcDqL3bPw5L7nTMETvQsIrGFGIGMplihjAQc8d2
cql1eX8otodVjJaQbMgebF/JYcDKLQVHc3VgR3oQvuKhjJEKi7xK3jN31Ejis16x
MwVZPbKfZdAflLxyeILDlSRQXb1LkfC4ye8JnaXYcubKDuH+wYR72arsrqrXF/ha
WlTny5nFlO+xYAMGxFrY0yyvOzSSfEuLVmKISB9IfOTYuX+FYWfBCoWz2c5phg0S
esJZ1BZOUI2uMYuso5SM+KL/Xet3nsskHjMCc1r5rc3CmpruA9qnVzVu2z+j/axq
JtXlc+5pn44Eeo/HW7ecbxy1kf3rOqt5XCA52ITHWv1Z1BZjX9zmk8pV4wACF07L
doTuSX0QoCn9qQ0PYhMII/eNlkHUaBB4YJPiszfjD8JaockU01l6+H/rly/I3a4U
5Xzi9QR0VO6wqhcPi7xBn2KNyuJKLkCDyv2jF1yxLnjNSViWmRc8hQ5VT/AKrSUF
WT+RZtTYr7SXvyDyl0zSzb0de7R0mB921G10PsfHoVnZYuObanj49C8YtDvZWvFb
z8PW2DhbsJwoOAN+sXWZal1OH+LEDvJ5VrZELyeg72m53ZVOILMAJj8mDUBZt07U
rY6hKEBp05fXvwLf5KLsAk+a3goTOpiHmODF22RBpDEIlBJ7k1RvJpjkgq5U3GQQ
w9FLO+L+KJqd13MtCVm79zL/V3WrkclaNAMKAdj0iZ9KqeVJUY76oVXhbdza54iL
eRIXIfPAOJKJ7wKLb2cnLrMY+1hr/As3/2crgF7aYrRpTNQO5Whpem6LM/Kf7wH6
TSaNTYBRr//Y9waSsKMttmDkR9hFyHI6waC9dUC6Ka80KmWTFhGqfbSAgC1zHdiM
`pragma protect end_protected
