��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_%�=��� ��}��v�����L P{u3��_�4�]�2(Z�kB�2�ׇ�T�fay�b�=n��p������1�w�L{+�+��b�8m�Xm�eذX����☾��5�a:�4RDçu�n��4m1nMD3��d�;��b�lڣl�`f�o�:y4y$�_/��������0�XC��:>:����3�_�SF��@�2��S��f)H1��l�c�Ts�H�2W�j�6�U�#ZM�Y�#�cݴL2X瀽�p�
s^BM[�v�_���3ðc��(	���ge������yx��>խX0:Y��x��;�a?8~t��s��n��E/�����ެ��&�*���Ha�՜�bH�7J��)kp���X4��U(��q'ǃDͤ4����#[N=��"X^��=��z����j�� 8iNj�>צ�Xq�-z���0kY$�@���@�J-Ly���� ��Wp�$V*�=��dR!5F��>R��>烰<FÙ��$c�;��:�!�.�%����CrEY��ra���&r�T��bx���_��SE1Sѱ��js�m�kc߯'kؕϞP���\�� ;+��*�o{@!b?WAӝ��2���3�\�Ziec��22���#{�%b��8�;�y̪���C~:���2������.Ľ��������o�D"����_$����zt���G��Id��/@lg��-ҵ߈�cd�����Q���_�v�����4��"�W�N�]7�0CS�@Lв������!�54��#�O��V0���W�N�x>IA�j�`����x�M�B%mXrp9/FKcVL{OV��PH�۪��~7̍�� r<�xв
��s�E5���핾�e���#�Z��o��̍��Z �]aɦ�[ټ�&��+��Ql*'-x�y������o �x��N�۲r����z���_3 T���ۊ�Lvo 2�A�"��Px��)o��	���%����x���ە�)!�=��X�3�m?a Q:8 �V1}RƁ��wE"�ꌊ臗��֢�x�ڄ��rPuI�j��� ���aEJ͸:�P=���������S�\�̪���9.�4Z�p39Ʉo���
$���G�cN����q�%x�y��)���� ��"0��2zu�Mx�0U��_�i�����������n�&˥3��%x�(��S/�Z;���.T�0ܻ��mn����R�+]8�싄۩��z�	?�Y��U�!WV�+FR�O\�����*�(բ�@R	���J�Υ+�Lt�z���7-^cW �I��G��\<�D�3RS-���yk����"���gt��Y0�D�A��b�/bVf"����D�h��-3��8{� v������l!��ޫ�_-�/��q��~�h�����M��,�"dk'f����.瘓P�
آ�0>��Q�)��do�U{XKb@�
�"Πk���{0�Ýb_&_=>�^����m����8�G���˝LU��M�)��zm\�v�S�I��_f�8�M��T���?8ݘ�n����5�p	؞y��bw�edX��3o
��4�{�_m�z�Re��ىq�cqe�T��tv������ۭ��n�d����0����Y\qe	��pL7~���SE;���zU�Tv~�WD�?�����SKex����<�F�*��-�i�������ڭ��]�E��A+
��n�0̦4�3��~
�=m�'��Ǘe�.Ջ�¶Ơv505�)�&rm�=J���;Tn�����z��s��c�J���h}ҀYX�)R,�T���{�l��3���C%C��X8dI�tH�х�a��3�F� �U�i�K`rR0��&�m}#"��3�o���t�ʤC8��6�.|s��{�<hSTf�o'xN�n?�5}@�w]eU�`��q��b ��7 �$2��qp4jZ[������v����h��~/_�RnH$���q�S�J'Ɲ胅���+⚂�T�𚻅�%\��v��Jk�l�CL����f$%ET��'�Edٍ�W�q��⠭m��TJ��/Sց!@6�bX����TI��h�	d�3�2+���� M�i)�9�ᇽ�>dR������e4���s��h7�5��b{|k�<�]�%��=;ܔ��5ɼ���;��5pD��bj�L« A���L,d�](5g)�VVcZ�ϊ��;���H|���X+?o�}�TAMj3Ȧ{d�XA���K(8�C0?���xbvv,eeٹS�,�52Q�e����|մ��ɂ�2��G�`�$��Mr4��o�+PCn�l�{.��Iv����y
�������Z�Z���nJ�?f܊q0��Z�{hT`����?��K&Pt�����OSj�I�Nm�f�>�C&Uج�S^����7�u7��H��Q�ͥRY.!i����Q��R[�],.�(-}�x�h���`�7��""e�^&B(C��}6����jA���GINrטY�KPǎ��ѳH&+��$����ϒ����@EQRl� qW8B�	'��:";�Tx<)���.��˼��z���ѣ�tV�صS(�dH�c���l��ނ��Vp�Fu0Q��bM��ui��+����~��Z��l���=eâS]�]�u�w*
HJٽ�YEe��y��^�@/������%ɟ��5k;�!0�5ZƐ�HX��e�W��k�( �����f�������Y��D��R���Z�*;���"��O�e��I���2������-i����a7�LrVi��e5�H2P{�{�V'��Y��%�k�c�����٣�f4��i'�����c�0����K���TEK�u~W��i���mJ��M>�G���h��9F�|���/��\�����0YlFZ($q͡��:��<�i�r^-�����6���Tڨ�/���D��Ƣ"�"t[���&F5wd�RUh����;�G[8������]�k.>����Y�~/j�>�ˊ5I\����_�/<,�Q��$0�[B�e@[x"�E
ćI�����v���vNa�0r~�N�B��a�q/�	#���B=)��`Bċ�R���1�l�[�g�Y4�7M��d���* 6D�Q���
p��9Ӊ�O]\gl�RJ�Q?�`[6'�L1��R��H�a<yr�j��H%c��k�PΥ�j��ľ�@9�.��h$��K&ƅ�<�0dt�/8l�p'���Ň�Aձ$$�l��t�_�R\���"i�\.o�";��Y;�lt� ߆b�O�ҳ���Γ.�=T�~�r��1�/B�T��JP0��5t��@E���)(�ٯ K�z3!�F����༠Ms�鑕�����)g>~�,+#���4�����.�:��b����_��ݐ��b�c&ԍq�0����d��Q/N�M9���4mՅ
t(���ۏB�uek��tA��E Br�fHk	._�u������bhP�a��l�[/���-�|���ҟ�m�}��:��jH��,%�ڜAj��Q9�ʂϱeS������% �ȵ��o!�?&[ ��� 4}cݱ��Nv���*�s��W7��1��Gy*�R�Puu��j�xT8�d��:�Sn�wI6�^Q�H]��۩���Y�Oz�k0�=A���ˊ�<B�z�v���_i�tjy *�[��*&1�A��|�R�C����!��ˬ��YQ�p3XI��Dw�褵�A)se�K4n�"tv��(�|+�¤��E�*�1]��4�>Ӳ!v"���K���>�BMJ��ݸ�#�	�r|�����J�?�	��Z34�G���xA����ϯ0on��#q���q������O[Х$��L*L�Od��	�go��+�/ '�F\��v�C���d����U����~�W)��j�A�Q��'F�����*�A ���,�`�5��>/��M�Ş��r�mu�2�1ѪR��a��&��� ��3/f	�����z��g��AM�����\5�y>k�{��kf@�uҾ�����B�����	�i������a[�f聮}���y=�Q\V?I��;�'ݐ�tɺ��y@��Lj�c��	�����P�L�]�v�E�[�Dh�������+E�����_19����g�����;�M^e�⏻�$�-��#��4��o��
hj����{��nE^����j�9�E��[�Pp��O�Bw�w����(G]��,��D��PHl}P��l���Gߪ�ChM�Hb��br��a��G7�q�8s/�B��C��<s�o�sz�Br
X�&kpɰu;UP}���l}��|�U��b�o���|gXQ���{s��m���O���5C0�HE�/�<*��z
[��i��*���7V�J�n���
�4#*��ɝ@#= ����~�1�օ�������?-�
^ �(�@��̓�b6��r6}g�W��Ǘ��(��۞� ���.�ӛJ6�����S���M�mK���UL��Dn�����#*��}x:9#'�O����דh�?���Іb��s,� �o�Y)!�"$�� ��y��:ͷ)��c̡s����ɼ�ΩX�"��Z4+�6t¢筜'�����V�' �b�*�)4z��M�~��b��J}-SJZi3c]Pn��[�)�>��-�)Ԯ$_���>_QD�p5���W�n~.9A&ҵ�Z�^#��&��T��M�qe�XO��`�t��� ����R}5eԭ��4�#�K6�_�箯	�3��%hp#��^�K�`E𪦯�E<��I6��^tR��x\2�#DI�ph�oPA��f��<*	��0�5�4�Ǌ,'�uOw�HG�r��ء������u?fn�C"*�M��J��s}ጯ�.Zgak	��0I+&�f/�&�O�Uy@&��G���u���{0����%���&�x��>�Xځ�O��5~�M��L�<�:�0��{K2�W��B�C�@��q�@n�������Յ�!mL�,'��u�c�<�����?ր��k��&vx_t�\B��R@nz8�}���EA���s�s=1}s�WN�S�1�)���<�
�t�}-�)a�{�/0��x@A�o_o����W~���{�5�E�E>g����T�����zG	N{�QQ�i����ޕl:��f���f�������x�Sz���H0t˲N-�q�����x��8����4\Yj��]����T�R
��Ҫe
Z<�.�b�/wdoBv:��ݼ]	M}�Z0����8=�53G�Q�����ܨ��%o�%Bm4�z���?���Xіz��ۼ����8���r$��[��&�P�*��9��X�#�Bhg+�GmHm� ���xdE"~SL�W�Adi���a��z;X[:��ܿA�嘥��("&NTTa�רc��c��������쯰�m�����)���7����U�&\��粓nK�Ȉ�Z��n��e2�p �Fв��p���mE�Mo���U��>X0}�� h|��l�e�8e���c�Gs���(%;�
�`��{�Rf���i�,ןB��(`E=�/��>�&+�½Vq՗"���_ �����3�ve�M��O_�8��3Y	�gsN��Vc3�Pܮ�����n8!
�Y?!�����V$�]��c����ۜM��	���4λ6m}�H��C�lI7�E��,��V>��["�c��<Z�7�����`�-O5/��hZ����y�����KM��ݳ\�]7xU(�u�:��$�����s�]�Uu'��"�0!є�T�<�+�����n���\���e�M��]��Z��Ų�t������R�ӑ��xdCZ���,n`�#��(��Y�v7�Pn�-2QU�ud��_��lУ�S��<���ڻ����TE J�נ���|Ds./rô������ֶD���h�������}���c	�j*�o���
٬����g5��y�"kmy=�ҏ��`Kmu��|�����>�nE!:}�^�KЊ?EB����t�Y��[�x&={���1(�6�k��
����_�CN��2��� ⩝lq�)��G�q�*��R�r�*lI����nl\M��-:���	�{l����� E�?���6z���{=�Q�n�o
�]b#�t�w�
�Zɱw<sz�C� ֠�2?��\x����)�C�M��1�|�:���()��ݐ��u{Nx���~u�L�V��[���ThD)���E�9���6A_���5%�aDkܙ���?~�^sR�] 	a��r#�'qi�M�M�=VCrC:����,l���[�l��_���C[�iw��>������,�)��o�5�@g��`s���X�E��pT�#���xP��/�n�䨆Ӈ������s��
*�R3i@�wm����/Y`R{=��f6:�������$���"K�s�ܟho`��ӂ��*E<���`A��:��6�73��[�<����S5�OۨA6�x6���g���Ci���k��/и2�)q�2a*�ILH�6���қo���[�Q����ޓ0�J1��jj	-� �M����������)~��h ژ��1!���܇�����\���gg:�ׂ K��#���|KU����o_��5&���	� @��^�
�N|d�d�� -� ���9�V�0�{w�2N.�Gani��4�B��%"P�_�ʪ�4R��H�U���%����t�
t�tK�,f�D,b"�����H�d�/* ^�F��8=1��p΄����,����;��)���[�HTGx�*:�݉����q�6���@��iK�]�`u�z�Y�ρJb)8n��2y8���^��iR�^�7��d���/�Ǜt��˯pzsh�ƚ"�!���XO๴<z��GJ��`����'�`߳��F~_qt�|�J�db��<�q�[9A��A�	���u�}E�vM.�E1t�Δ�������6�3$,�t)c���;�h�oZE^�kg|m+���X�&a�͕SO���9�R�T�a�������@�����Y��nv5cw	�GX����U�J|���2���ُ6'J+��+��z}� ��x������u�����#q[L�t=9�9��h�����^�lQl=�����C�<���Wo^m�@+����5d��PS�oU���(|�t�\���lr���P!'7��+Ձ�h�:v|'��{e�1�����/Q�L�wgV	��5�_=��c�bl�fnu��2D12��h�G���V#�o��_��Wh���xO��7��ۇ�T�0ּ�:�g�z�bqH(H���(f����g�A'�Ƈĩ��ps�36	���|�哣Qe���a�!Wvi���q�$���8���V!�ml�>\B6|2'�5z���8S1|X���ܑ*��%��9%"$u}������	:x;�t
�Hk�P�+]���B�1�@�)^֘W<Ŭ �H~�P����f
~7.'Ӆ��Mcc̟����:F=��,�
�uH��He���0�#dn��N/6��t4n�M.#��z�g�ELd`f�77#v�ڀv�^F���ʈ`��RS6�/�D�݋@P|�͂*6�:���k��O6�eR��5| �!u͌M���a�������[�h+�ʰ���� A��y�����!�Y�0�s���tL���'��ć��K@�*�l�y~"&S���j���|���/�;s�KH���t.���>�/� ��eP*����N���AEb���=+�ԩ�^-Џ�f�^��e�3@(��_��L�y���IHm�CZd��==���["�Q|���9,��j+�m����e�k���j5��C)��;[(���Wnc"7�ʷ]�X�´!�$��\��\��y6�|�ް�jz4z��d��˿Q��e�cI�&;���u�Y	'>�V�[W1�6^y��i���}x��4�'����X=E�SpJ|�ڈz�k�b���JW�G��o~�t�k0�86�^b���J�! �=�$"��tl?����JvZ��LAz���/(��*݀N��u�"�|����̲�3��X����tSD�!m�=]�¦aW|<���Sq��j-���v�k�E�ٵ`d@*5v�IŖ�Z�x��
�T�m�x{D�+)�áS �:t�"��O$��2\;�`��'����'Nl:wтU,`�N��C��\h�C�7'Y����	��K7; �AW`Z�!5F����|z� "+���xt8��m��+�1�YĀ�����U��d��NU�/��PHe �H��ɵ}�ҙ�IH	��:�����{'�7�.�$�T����y���Í��i�D*>��g�k񅥘�|�`;�h��&2�&Ԧ��.����C"�ԶJa�A�[,G� �9�-r�iz��:�:L�]JZ���oM_�,����zۖ$ҋUfXN��قc���y����LI�z��p�"aԲ���d5�u�5p�"�`fD�!
7�o8]�pA����<kV�=U���QU�x2W����1��۱�����}u�R�q��h-�i��]L���fh�伌�T؞N��������I�4��@�"uaZ���c\��vpGɮ��,/�U�DT0��v<+ z�ƗI�tў�D�t� 7\C��Z{�%�N�}�e��1��(�P"S���ef!<�ZX����X���jW^��eh]r��ptS}��"��?�3�#�}p���T{ݜI��+���(��������9XC%���_���P�e�(SP�E�PqM���1��5H�.f5�i�	�Oj�+��-.iK˕刧Q��ގ��ne,f]Jx���;䵲0�ƒL;l�&#Ăi�w�}|���ɳ�E �t�����ҫ� �D�皛�&���h9
y�-ݖ���$�TSD,CV���ϻ˸Q��"�sMX��֕�i�k0��dS���ݷ2K���V���������?� S�8k�n��S�{�H.��=���S��N������6��,�n�O,u�̺���B�{���/'�Ե�HG�~�?�=l����Hi�h0��4�+d�|M5~o��]<�Zʤ�^�F�+֮g��ø���\�"�����L�=&����'��.T�0�]8��ʰ����A��m�t��&�{Z�˾������(�P�@�����%`���g~��4��S}]������,��t4p#�<Kk���I��f?��	P��8�P���'	��}K�F�6a+��'-B����Ad��4�@��1� �Wlf����w!d�)�n+b�a�.�&J� ��$S����KK?���A�׉Z����T�O�
CA��������u�k��6���X���b^?�i��h���>��I}���W�2b �����9����N�j���#�x}�L=�_z� ����o�V���.D��5���&i�h?2�����R^t���Y�bN�i�C��
�E`d�����D)��{c�3OQ�w���^��(ε�G��Ej��eثm���~�č���pI+F'�����Dt@u�	y�W�L��{1�Db�?�0UZ�v��;z�Nو�ܱ�=<�tn6`��O��pw7 �VS��`!2�ݼ� ��z"^�c��<r`�z��l������ �M�2@O���]�����|��
�C����q�U/�iذ񗯭[ ������_'Ǎd�5����ڜ<��GtQ�h���Y`4��̆��{X�f�:�j�9W#�h�>��Ob9��	?��?}3z��m�����a��c����;��3��b.��6( ��O�zl��/]��z��[/R�W��%�'�v2d#�8���=��kl�����0�����ub�xm�֌�.��9*�����>�SU��?A��<8$�Ofr�R t��v����үC�^W�M ��c��p�)���4�^�Y�.D�7����+0qa7pm���d��t�9\X�*B)��.+�"���z���
�zT��+���vn���l�y�ż���B>��k�<���_�rW*O�a4�*��$͑��
G�D]���l8�jvQqdi�=kf>�c��	��2�c�p�U4�m~job���%@}����4��S2�����=�a����Yi���W�`�;{ܖiY��T�F�Bx�@�_ݘԁ!A��\�2V���H����Ͼl	e�L�>������'b��9z�j��BFuk�px��$�c����wj���" tŪ�f�,�R7�R�ڽ�鈼���&x�H���]lg��5ҏY4��R٫wܮc��d�oB��᫃B��q~��$9!#HȒ2`6a�ĵ�!��8�T�D������yB�r�H2��$��t[�@��&���~����v�'�K��6�*�K�O�v�d�����s���ЍzQ��(d� �PJ)u%m ��a�k*N�*;�� ��Б��R��,��Fn6TQʨq�%Ri��񍎩�ѳ`�T�&ѴhT��&q��%�X�n�D�ZIyr��	E-�Y'�j�_#�p��$	�v?��rG@ٵ2��Zxg{�b����
j=���p��}f���Z��R��.����öq>L,�] �waS>�F�d7�!Z�)�7��" �m�'a�+�1�'�=�g義wv�F��DEv���k�U�k �\{�Ng�j�2*7 f���SD{zV����i�V�\,cC�x�6HBpXq!ʂ���L�гE�X�{���(V�X�NMs�h�h�0� $!���Q�
Z.:0����ը�SS�TOE0�(r��>&q"�ȏ�ѣk%&!@Yժ�}}Ol�t��F��g*[íH�ƒ���4
8Z�K��}q3�)�l���Є珫 p�-�oP�;� F���$}����a���<�>�`���Z	�꼉�L��.�Q��I����G��g?��R��]��I�����>��4������a��?�T���3 �����L�06�*���.��2��3y��3����Z��Ǘ�+L�F"�+M?�@��aQ���s1�@����\U�D/���z6���t�-i��z��sW�jإF1)~7��G=���I˯Mz��ȳM|���'A�?�-S��f�|tk�Q.�v���yT� �`wx-?�f��w1㚣���#�Z�h�e�
�?q��˂+X��) e3
�5e0JW�/�Ċ��*��Oƺ�^6eU�"�JX��?꨿�YQ��q�q�N5���*9����j38�8�j���uy��n�j���A��E��G@�"'����]�{ҹp��Z���Z��ƚ��T��tzM�y�8q=�P� �I&��XՄ���e�k�.� �a�+�a���ҍ�O���Ӽ�P:$�*xr�������Z$:*%/5jӟ'�F����_P�3��b-�b
j;�%���ū_*~�D���S��01�3v����#�X����-��W)E8���/�2D�r�Ud�C����g6&W�^<����W�JvX���E�L!r��	��2=J+Ųr*}�����|�/���f�Ԉ�o_��sW�s���9T�h���ś:���+&���P6�KoH@�EAcFԺ��mJ�:mcMQ��V��%���i��[UQ��21>"�����w1hSU���E��So��t�涱�K��FN�Q�Tw9~��� �~�3ݘc�1�R�":m0r�+U
�&�|��C=�v���t���6�J+k���k5q�Y�6{�x�Y(��t�`���L�E
��Ux��� T�ĘSCf�����rJ�A�W?��v�?�T'��m�+�얶\��q�͙�3�N��x}*0��B��X�eߘP�d���#!%ȟ��H�Um�?p3��b���w3h<���-o��+��lQ�j�XH����N�(6��|.6A.�z�q�{d���t)Kn+��=d6�欓?�H�����a�h�?z�j��mWV}�0˷���3�\�}ٛV��8`3��m�PX�i��^���~6�e���۟2hju��)���Z�����rǐJƃ,v�l/�hGJ��2��M��;q��L�\�\�hE�}sL���S%��n	����S��#��"��w�tH�r�L)��S��g\ꭂ�Hkŗ�.Jc�����È��$�>:և�a��i,�+auN3Njė���~�d�
j�W�
�4=?c�&jf�x2LIû|��1��U�	��S��"� ����nBo�?6�1�]�riލܽ�\�T��Y7���P[������X�sT苓!H��']��;~��n9���U�*�ur=��z҂ա`�ok�v��`��� ^�{eڱO{�F����v+o�l��V�(O5��G.1�d{���O�K^I�I���������e&gɇÏ;����5��g���I���Ԃ�b �v��V�-�m�Yz(RctT)�1��2�M��[D�ͿQ���/��$,>|n�)���H�)��"E�[4Rq	h��~[VFj��z�Ѵ> pi�Xwg�aO�<i��k"��S�ޒ3�%�cSS���M���C�Ux6���i@("c�$�tOj�>y�5��o�3�Y
�ю1vc!�`HIb�еG�w<a��L�8��<?���ن�.�#]��O=p��]�}Y���HYZ�	P����',r>���XR~��,V�����t&���6Cަ�d�����T狪�?��$�N�L�)En�$����J�	���_UG�;�w�/q��k	�����B���	�����bgF�;��o���]��Z,��ÒbQ@`�_[52�^)r��o����ɦ�����~>JԐ�Lׇ+�T��j��� �ϥ?z��u.�����o�%d�&"[1�3\$Y}�^��Ĥ�DB/CE�pKi��$�F��������G��Վ�kt�@���N����p+�[G����ł������K�U��,��0%΃)0ʴ.)����]��� �J��v#[T�I$�I'�O"��4H4��"ο8	�������#w��9NR�S���n
�>��R ����rQ@ϰbY�pN�U���I�!�Ɉ��7z^D���ĕ7���>��B�6�!b��_j��p�0����U�'����@��\����a2�[���k��^FPg���N��7�><����yQ��l�� iﮰ%%R/0v�������J���o�Pl0+���A���0����M���ت~��8�,����<i�s���$k&*���>�!�8��{��4��
oi��%\�F��Rn�J�`?}Ȝ���:A��mQ�T�ϟc'�Z��G���h��{�3B�""Ց)�+�G���Z��������J'�'�m8=P��u�Y��1f����JS�G9�%��^g����l���k��-9�Ʈ���HH����O�/�5�=�G�r}��̱�Qg(�NA��`�A������,����7}��v�E�Fzѡ:�3�kf&��AX
k2fOOh��������P�n~��{�}ޫ�c(��}��T���^�'"������������Z�����VH���V�f�20ih����ƈ�s�̏(��ф�?�i�)��k£Ё �W�lo��s�7`��e��`�����T�Y�v�\��R]����L���)>�T�~
��8��3#(Ӳ	[�v-���+�����b&<��h,��=s�v��B[n����(d�j��p��ln�yB!U�?uM)+�e�ޥE/��e�0�V.Ե��$N?`D�����;}�Y;G���
r�	�1�IsK�IJF�lmFj�C�P����~�
)�������X ����Q�.�jE�=�ɢ����딚֟��_��d�LiQ;��/�X���a�C�LJ�5��]��S�G�8rWy��\�?K�\c;�����^"�0W?5�U�z��D�U��&��&0D��u(*>�s5����o��'ȥ�T�P�x�E]�
���f��m� '�+9D���V��kr�s� �k#��F���I=t��������P��K�l���S�f��B߿�gW@�ɏ��U��Y�q���kO����r��E���q�o�L�b�F�ى���g�K�?_x�]�|M��ם�#A�0�){���lǓP��b���>�p�r�����vD�[AX��4^������6��s��Og�
t]���H�m���:G��צ6��z��9J}Ǯ�XQӝ R�t�k�
���f22T���70��S)֬�O������J��&�4T�M�R*�w�ܼ�]��hq2���!���Xd~��vP�*�U7�+s�jJ#��s�X�4aɜD�be��z<�:S�}�c�T�O��u�MW�^Ծ������ ��a��ق�(�
{
�9�0�@��}瘻9��v�}kiS���dԏ�y�Oo�쾰���(lJ>L*��Y���Q>,A�P�`Q����� �wx���`)w#���|'{�M�� $�a�/� y�/H�m?���ԁH��H	�~�}�=���/*t9y\H{��$j�4c�+i���nRTKZl�:���N�qng�I1�������m;jT���L/6���ͺx)�N�w�p�vم]�ݳ���l� ��˥�$Hy�2�B7�ލ����C]0���Y��y�M��u���<��3�g0�Q��	���Ѝ���E�X�dp�&��*P�V��W@�.��dH�n=���RH���L6�$q������k�G7OU#/6�K��Dj��~[�9z���q/�~���_b�uvm�EH��|���p��@
o��k�,:&����ϩ f~�pV+^"昜&!*��\DF���8����=��1�܈er2��
�Cz�a�Yymfn<����v�`;d(�L�K��}#�U�%��"���l������P<��/��OJ}��������	�ɒ���X�  �`��R��������J�Q �Ŝ�8�Q��W4��e4P����.���!)�B�#N�tM%�9�����`���?�K�/ u�Llꎋ��4{���r�0j�Q@(�Jǁ�g5p�%��� � ��]�sb��CV�Myl)�����i"]��1�cb��$Z�ɑ2%,��%	?;R~*�Z�~�҉���U�	����@�<�bo�]e�s�/�
��j�5N�&M^n���*����&e�}��I�ӿ1]p���i�x������D���/><IL4��ok�m�hȲt�T�Z/��_��f�>g����ڪs��x�|@�ġ*������}�o�2k߯Y#ɶפn�W��D\�!�hH�p�$����;d�,�T)�8�.`�_PLGŧ�;;�l{u��0��NS	�`�f_���+A#S��,33XO+����Sv~�W.�=�4�ͤ����Bu����l�=�=� ���C��D(����c#��"W	1䏷��o�&��t|�V�MO���v}P�ִV� �$Ģ�B�P }�斏X�]o"KH~ܷ�7�h�h0�3����1(�Պ�\F�I�,U���+׽1 ��_hk���)`�N>T�1]����p4�zM���;"
}�����ek7� S=@#s\�BC|��H���x�Va��}��w�*0��tPY�����3�V�A�Z1��o��g���)X��"[<y�:(
I�q-r��;g��Ϸ;α7��x
���$�M3'y֦A]�i LO�Ն��y��w�
sw�ͬ��jf@7�KZi��?C�����n�%л�:�X���S����2���U���41uF�#d����zn_�C=# L@1Lh)�T����js�U��n�N7����T��[�S#6�Ut���xh-�/7�*�S	�h�&O�x���>절�Q��N_��I��BD
�A$y>pG��hc�/ˌ�鲄&��!(�Q��E?�����EJ���+�8�8�Z�yR;пֳ�IZ��b�����䒂q$�I�4�|���i�Zr�nx4vɛ�u�^��dOi�W�(c��9�8CU�{�y��I�,� �O��"��Ր��=����ިi-o_0�vm�14?d���W�g�]��7��=�<���=�b�R�-��������8���eN>��-*�W���o	,Z��nFZ�#�H�,gE@�uXQ	Ȁ�x{��ĥ�Q-P�Fftuj��Ǳhw�y*p(�r�i�-]��������K�B ��5GyƂ�ń��
V�����&	���P7��v�y5���F�c����$��\JɥqI5:z�n �T��D&3�u"�(�Ꮞ����W��FJ�Uk�v=��	�61�k�倢��&sy0�*�������T#]�5����:Z,�h�qK{��W�?���#ۘ���O|�2��Y�2�̨E�1U��l��T`ߍ{��:���X�i�˥u_	�ԁ��9fM'�\@"��gw9�T���	��1�1��=���%�`F�tbg���K���w;�s]avیz:o�=���;�o���)��X�_6�v{�G�WnI�@y2�D�M��o���f�đ��,��X�
�#wǋ �P�q�앫U�!u��Ẩ��d�_�+Q�z�RG���G0��&�^	����M/�R���p�-�
���(g��ֆ�]1�=�%Ʞ#�Uٙ�]���(8������A,Ř�,��]O�I��d������W����aQ�_¾���c�+�de���\��d\�q�!�����3��f/�j�҇����N��V^����uhD����J4K��-�3P�P���w��	V�}��0�����1����vB�S{�j~�>+��h¾y�X����J�
"�8v@�����a��Č:�p����dM�p'}55f'G��8����[<h�f�7�
���h���+��M��Sx"�PF@��"�Ȉ뤑���P�+QO�»J��*a�s���3$ƣ~��=��C��[����U�齃�Q8�۶����04�cuPlB{!����&�[�i:�8���߽��O��P��f�>��j��h4+������F�1��RfI��I���ok|����C�Ԛ����H�"�Q+����+X!��l縃�i8:.Qew�����N���j���H��<0Lh���|�뾂�@���s�{��<1v�EkX�3��F��z 8���ْ�3�Ӂo[��YLȬA�s%���І��K�&{X{�W�4�h�gˬ���*:<H.6�òP�CU�y��&�
����%/n�?9��kN�F����靋zP� �tr�ԧ��Jig�u�p����$\�{���C�p-�/�X3��sʉ�<Z'ifۏ?���6T�(e������3��[;}����h���,��M0��<Ut9zN��}f����B&��O���?fx����u8����Ʋ��j���D��}<��Y��G"�d*�J�Z�'��	��� �YI��,��T>�\;�hS99ۢ�fHX+ܚ�)y�}��ް�6QO��9�{�:�E�n�`;�N7��(�#0��=>�^����z9d5G�iɝ9���� �<�n�פG��������|V��Q�b�BCК�$�J��i��Ǳ	�%��y�Z�%��f�w��P�-8{l���*�VA3�^��@*V�2�6��ˈ�	��󏘤�_9�N��W�9'��l��1\��6p��n��+E��;|��#�a���r�w��?�-]�"��F���'��WDD�n�H��$�I�4�ⳛ�4,',�.E��9�4���IU�-��Q�Vx[n�zW��{����B:��D�v֐x��Zݾ���CY��h�,ݲ���Dɣ�F���e��ۋ����eq\,���b�p�킅�	m���H���ߏٯ��ZG$��.����V&P+�ãL��t��h���Q���<�$nX��3�T{`��
i�4����r�kn���Š��2s��ׇ�p|%����1
�\W���æ�s�9��A_�ъ�k)����O�)Oj�F�W�ҋ�����C�YY3�b�ԅ������R��y�|Ʋթ�Q�M����Ön4��CI�;�{ъ��?�p�0p$^6���AJ���1�_��[d��/�`�Ә���
�	?C��=d���75�<�:J	��'�'��&�3e7
�ʗ��m��!������Ï(\�N�#�0u�u�ɑ���(L���H��X��N�̹�u����f�;ä4[cZ.Y�'�]�)�/f�_T�d�5�rm��L�sb��Ec}�K�����i�'0�XI���
ƿ�S�C?�J�Kз�&|B}�X�/hL9kS6V$���(p��c�m0��y�L%��m��ף�S�9�/#�G��n�8�]?��� ci@XT^���3<���S�_<�����L!X�ڒn��P�����	"?�hH���%W��z��p�:]�'5@0m�J:է�r�'`eg1�δa������&T�h�R�^ZT1r�����̀i�:�~J��Q Rf=L�ݽwX�B�$��[�;$� .��K�wf���PG����p����Ɇ֊3����N��D/�b��kAE[���N���v���~	��Լ�
��/��H��h�A���yB$�	�ē'��v�����Xq�I���������a�<���kfñ� �c5)n�x-{V:��(������,�E��_�P�����+�d(_�z�[6�*���Н�=tݸ�sAx�\e1��D�҃�y�E�����r�I��`���B!��E�n��!����4u���җyH<C�b�V%&�uO9�`� �F��(�{l����.��^�%8o� �$s��RRCG'���J��J���'i�2�W�	G����H�<30���>�3nG`=-:9�0o}��[זi�����CzH$�ڛ9[ܺc�F>��_��b����T� �+�p}N��n��4���e�)eEƃgȧ�	�}��C����P���gG�#ށ���v�3��i�V;���\�@'����(x�1k��cL�E�����Ĭ�����䌠����:��;�1���d������E�`�����v�{��-9�����{Q�՜q�f���Bƾv&��P��-u�"��-҅f��s�R�
�^Ga��p������p�;ipy	i�fW�c�� ��O���h�w˵����Yi�~~��;.�%F��Ƃ�f@�	�4%���
�G��bdb��1���44Dc�76��塍��Ҿ�؇��x�am��R�P�ֵrPn3�/�W��^�khٖX��YeQ������F�Y�I��LB)6p�~�*��?�����?�C���/����t�܁i^�n�#
<K߀`�Ħi�?���f��H��,d*Ŵ�:�{�)v;C8�2�\k��ŋP��}V!������k� ěD�#����3����KT�)7��R�nV�Dܨ�o��G�G��s<h��l)�eꁌ��:��P	x���U����;�co����y	ƭS�PR���A��G�p\R�������z��ۼ$&FR�9����v�<�;<��'`�G�$���U��-�0~����;OFJ�5�#.��|��n���v�uUc�>��S����B���rU�Uʵ�ߒ�j���:�_#nm�o�v�oy9
<�3��{,��ǜ��A��X��3�i�>F��[Q��w����JSŸnKaQF��U(#=��p�IjD&F��V"oV��JU�y�$�QE�^P�Tm�E���?�7u�|l�=���V��iU�Z�Y,{0j��zx�]��J�t����lc�4���G/4D������:L�	��p�u�
<������Y���@�fkn�i@�����g�fC�%����S��5�_�aiY^gX��v��ku�ħo��͋
����[�6x�*	�3�x�j���H�|�F �j@C����/��}��r�XI*�o*�$0ɍ��Bk���.�K�VXߑc��iClh��9�s�+w�??M�4���_�J���
��Ǡ%%������Pq^���έ\��\��  2�O��Џ�ex�1,��ӊ�j�l_��s��:���<>^��ѝ탺M�m]��Ƀ:���J����6�P����"�T�+P\o{j�鈶S�#��a��~��6I��^��l�T��?���䦄�YK�:/:�*�{�y��M�`�ۼIYJto��U>��a�
�eZ6��ʻ�R�����y*:�h����x�{h����~4 �$h`Sx/EGQi���=���Xr˽�݃�/��ϐ�$�ׂ�S�N]8p,�,}}�]#`��n�;CL�8#���j�n��5k|T�Ž,C�V㚂��k�HUb/�a����3����B��(��C0uՉO��3�i��Dv(�����q��K5�S�١Q�;F����lp�HBi�gQ���<e�*�e��G���V���i�P*��!��#9i�K!�d�	��y4��m ��Qf�R�<�"=xjF�o%��Ū��U�t���T����;丒]�MT5G ����.	z�a��na������D��h��	sᔼHouG��D"��91M/����Y���#%Bc����B�+R�#��:���nYo j-�K�e��/��8x�������nehy�q_�^� d�BNH���
�r��D>7r��×D�����������l�OD���Z�^�<��
�Ϗ�ň��9��H5�4�����ѳ7"|;��A�M�`=�A���k��� _�*^A���%
]@�4}��\��*����jb�@�Ih��ʺ	 �VZ���Kp��Xo�[�"�vѝW��Ӆ+�`!�J��L�*���a��#�F�Z�!�����飘ٍ�v���\IV�u�)�n�`�84	�ţXgӤ�^#J���]\򂊦E�Heб���G|���@��'�l���-EY�6�U{�0�b3�����T��d��j�����J���<;�!4,B��3}ů���L�H�E^�L���\m�b�;�80�˔�gI6�a?�^����#��.mI�r� 5���s��pREB�)���)8Z��CmԆ��[�iT��Ҙ��o�o���9�wuR��U���1�P�׺��Lp0�5{�ڃ6/M-i�a��V��~�3Ğ[B���#̑��;� ��<Z��s�w�-Jд��K�8N&s�uH%'&`7���'	I#2�p77�ZY�	H���o�p%w ه�7�Bʀ�Pͧ��V��5h�t"�fQȋWʶS�SD~=3�§-����t�b�<���X,M��Z���)�5C�~�����8$*�o�0����G�C�Tr	��j�k�1�X�T�=��#CC��^;�xY��~`o�b_�!mc���ٮO��-���h��X*-�8.�~C�x�#�GY�Y��c!��\*��r<���0��<��/q�%�[�a�I!��ֻ��֫� M����%ҨK�?LM�a�Q'V�Q��@B�.`����r��v��������&V��\��j���B�x>�F�%���_e]6S�d�D_�w~cS-���L�����Q9������E�W���*�fr{�U�����Zn������4 F�KJ ����X��7d �x��LJC���W�=~���*b�7�����R�c�C��389�㣅N����b�vUn_$a�/3�
�<vS<K'g�5���A�%�(mD�����i�^ qH 
<@��ѧ�ÂX�0x�>����D�B����P��s�Z��:��q9����Ւ�"���K�1���kvo*����sb��z�\�S����؅�
���Ÿ��g��d2¿ ���#n���5%���q�:Y.��9�vn�@Q�#ʷ�-'�^��$�-�ze��e��d��q���#5.�����(���k�	1��޷�O��c�/������3<�R5h#u�eH�H����T�8qOY��
33�낒݈�9AmcJ /�KP z.�����>Ui|<Y��<�2ⴽ�QG?:Bf�������P�y����#���}�%�j=̭�;(�ӕ���-�x+w�
Ҕ���=�ެ��mg��<r�~�g��4P�����_��!���J��r�ܘ��\K/�SMl���B2V_G��@z9�����q��uw W�e.|LD��+<�+nߝa+}����� }���y |��>��]/>�|OF�i�k~���[��1��8wt�A��%6b��>���5���ȪA��ݏ��� /���u���I�Y":�ƙ4[|�_]�����Ƨ�t��	�Z�(s��e�2ijT�}I���$oit�,��6��u-߼�'8s�H���#���e;��Z*����@�k\����#F��M6ԿᣑG���p �TK��XI.9���P:��� ��G�C�̒���5��D{��X�a�FG���ťz�ͽB������vO�,����{��c��&C��C�}����㨰�7� $�'f.#p|̈�Y��A(���_A����v)�|2��7�<Q:�F����J���\恏X�t��?aE����X8~ݜ���[|�r-�|�Un��l	�O� �"� �x4��%'b^�%�S�7r��P�!�����)�I��N��W>�Y_�pDj�f��In2$H����=��������z���9�#��"D�;���N���E�]��ʚwuy��';�b1U�L?z��.\��^����b�HlY�����r���6��p�� �&/����LRZ�ED�n(�
������cA�:�D�7]M��:�N���^������S���1-�V�3j��'���gy�%��ߜ��ɨ\x*�_.X�_�O�-�E¡FM�A�
�a������l�<xkR��D�������8�I�^�y��3�� �8��k:��P=�/��H��ò��J�y�8�^\��/�8�/���+��'jjt���y������@�mK+�I���pI�^��>)��k�A�UL
�AQ�lh�zڏ�WpT��B)=F��'�җ�����5�������~ضq�g�`�f�p0���q�2�E�W5�K{��h2F#���?y�}�*a!���p#BO�p������H������d5���h�[YŰJDO�ru����ʞy}�V�j�BN��s���㤕�E��L�7$���J��E5c=?��F�u׵�=��rJ�)�~e������ţ�P.�5y�pO�ɹx�l�Xv,���ǚ��# }ӷ� s�6���#~pi�D��+E$Y0F�t��+M>�ܵJ�ȳ͕�C"��RiӜ���E�G(d(���2:9�=�+�ne��$P�!<�!oQѠ��mW=)J���$����[-�1y�.8^�]d�l�h�r�ٿ�UG���cLvn�k}&*�ں6��Sb=T��B�]��Rɽ�0���:���߬��O����*�>�g���]��vEzD LѴ����N�9���>�9}��EH,�U(S7+.�W�$D	/�.�+���u�tu�;�K�d:���鋮��W<�C��zu�x�dn`W�I�)�)������0\h�F����.c�&��JV_<{L84A �Q��˗yS�꼯��u�G���uDѶ�ۿ�*b�3u �r&�����B�O봒)b �d,|�h������:�ɹ[��F��EQ�[n�>iPD���h���W��9VQL��k�j�O:�y�Q��k[�dB�k�c/${n�S�Nk�"/��ɐ��~#StX��R;!#�M�cC���X���w�xr>�Y��@�ʩ ܎�I[�n��C9ݔ�I�.���wr�Lv$.��֨��7�=<6/���J�ߛH�PM�����Ҭ�j�����j�M����1Y�s�b:b�4ɧEi����
��{�Q�u�I�nr�+��h����=�L��9q�����������GA$�Uw8�%�W�5(��:��p�A{��1���w�!��̟x����������>��py�HE��	��V�~��؃0'��U��ah����Ĵ�[�?�a8t���"z�}��e��{�h���c	�Q���1`h��h�*�?�q�^�#�4u���e�;�����%\���_�yUz�u�B��U9��� )(
�͈��(/���s��@��ǿ�r�D3H�d{)ssR!L���1�4|:ǁ}9n��F�-��ж
�+N��-���|�`\�x'jT�Ϩ�-�s{1��Q��[�))q�Yn�N�����.	K�Vs-%����Opfp��v^<*6�'l'��l}�ռɑ��*h�{�
��ڭ�P-�ɞ�-8^�ӓ�\V,p���E����;��7[�m�.�Q�RfXJ��4k�\�+��i@'WMLN
��žگ�HX�D h���T++���fs��BI��7��I�I�_%$<2N4���B�$���Z��˘��s2�����V{tU
��P�N^&D�넳����`1����9`�I�ɘ�5|=H�h�=jSNIN����$O�a6��0&��(^��0)*�z�H|{�c%��6gˁR����MJ���ٚ��<�p�����m-�s	���%a.(&�͢"�����Ks��j����-�ƛ+N�����m���jL^������@��5�J�g9��k@����HF~����o:Q�ඩJB��,j9B�3�X�b&�h\�y��CI�n2�$T��]���꣡<����UçMc��ݝ��4^��2�nK�N�<�T�뒥p�º��r�	_qGnZ�T�W����v�3��⾱
%��P��z@(Y%K�@JKi��N 8�W�!�fd�~�D{v�K��������%x�;\����#XQ!���̯J���v"��.3��91�[U��G]C�q�S��*���#����ZH�z}e���Q��m�5Y/6j�4�(��&J��
)-�)���oDTX.�+E:�*_l������t�"�N`k��Ϻ�E�*jI����oO���i�|l`0Z��C�1`bʀ�0���?������nz��P���I��3D� �Ӭ���,z#7v�o�`LMǁ�V0��lT5����G�K��ƒ�9T��L��� ����,oG>��0M }]���`��p����<Z�E��t�郚�O�o���^����A���D�����5�א�@�Ϲt��Pz��df���]`nS��#�G�&�����\f�.2�o	=��H��M����j\b�]����M��grI�;}�ײ�B�Tq����k��v�L���.I�W�U\p�^����#�5�y��o�u�1�K��g�Cu�	8A~/�,�k�#���*u���q_^dn#`)��
D���Yn	�DŖ�7h<��z?��dK��Z�������ȶ@,"6�+���rQ~�P�� �ɸc7�qr�φ5��J;�o!i���|Z�㋧!�BQ��w{����k��&	w,"�b�w0�	�T���'��j\ˊ�t8[Pv~����uv�צ�RǞ ���b�Ө��y�^�?��o*'�QNO_�o�N 3A��������k@��N�>�����:�f�uE9�VG�x_����K<IS*S���C���W�,g�	������u�p}�D.�Z�c�S�I@��V��ݰ�C�=~h�6�����$J-��L�O:��WI?*����ՠ��^�>��c��{�o;�'�����Ҧ\�*��CP� 2�R2޷���61_�C��e���K<,Ф�e�hT�6��_�|�9�c��.��W�ro��:9d	�[=�}���	J�V�h�6��R��.5��o��t�����_�L9Kp_v���Ϛ���+��C�1��%Ԥ2Ȋ����'L����u�@0���������+q	�5?a�I9��6Z�F��>�G�#����ЇfC{\%[��g�:�fy~�6���")�`Q�����|��k0�"N���Y[�����L��m�/4s	�N��ϗ9wy.΋:�.-��h� ^��eת�seY�9�O�[c���S�oT)7/
?���Ff���α=?��wK���P>8vl+k�^8�9D�< �Æ��W�X��b�'���F���7}JT�K�����bq�^�|�Ә�������x����AiP�Q�-65��ֵb��*�*������q���H�� ��{��a���F8��N�"\��R4����N��ڴ�w<Sh*�RxM-���+=Tꜽ��$��ӎ��V�F,(~B�E"`p�C��_��jD6�u��AV;S�J����N���$ZD{k�}�C5�����Y��[����BW��CK��/ū������-�.C��!i�S9�Y2�ӊ96��>�¼^��m��[n������9|��-'2�T>Ԣ�����*�0d�I�5�<�I�	�wR���o����`7n{X��ÓE{�5a��v�v�L��t	�m�4`}
ėQ��;"��I���𹙫Dt�U�9���M|w�_��^��XF��ym��kA>� ��g�1��9�]���Ą���F^2��o��EV�{�������e�"T��&��2�_"�d��?�u�3����e�K���ܷ��k��i��o~��m��>�yU'g��X׮ʇ�y�><�������[�W�����B�P��L/�+w��m�u������!�o>�"hw"�:&(1�����w ��������dc�J��G�#��0�O'�VU��s�d�1�5��ݿ9�)��u��f�}�#_����?\�WU"&Ѝb\�5Ѱo�7x��R$��P�$!q�ٛ �f����$	�bؼekБ�󗏓qk8�Bj��7�Y�������3:�PP=ߤ�*5Gvj���=|JHK<5��а���9	�iY���:XpQw���_��޶�`k@Dv�*t�ϑ����kmZ�ZJ1r�{;>]���H������|��v�`���k��OY�y<a�W=+���Ft�Q]4�E��U��_;��C���L�I^������^�!�^յ3���uhf�,*�N�tl� ���w�����I��]��L/S�mj{����YM�~�V��6�r�7G
�G���|2�mÜ}�\Ԏ���MD�~�����z֐_&�]T������� ���9�A�;8����|B>`55#������) A�~-��5hx�t�n7���s�cf�m�t��>l&`:Ug���j�l]�l�ci!U8�9�$�=�^,k�?�D5���c�V����3h��	ݏ:����P�$o��憔���X��� �)	�)�FR��kUZ5��R��H���5R�ퟴ����L��m*O�1�6�-om�?�w��JX��Nό�p*d��;����:{���!vCV[�� 1y�p�R$�t�V��� MZ=�cZ�15%l��νsQ�' N1�j�H ��7K�c�Z�BE���}x�=�-ߞv�1�*,�ѡz��>�4�����]nea�~\�ƥS�T0{�Ϫ�@�0[_B�� ��+ĕ����B�x��XQ�TP�HmD�$�ݫ�����d	b�ǏJ�W�õј�{�?hܣE�ڄ�ש���:�?�؜P�t��
m���s�|24�t�*5M�͒��!J�[6V+K]�N��D�8���RS&��9���`�U{��.�͔�($ rY]1�*�]T+�S6���FF�2��YU�*�ڇQ��h[��ۯ�;��.F�9Ǘf�_g����$�6�]^���}�d`+�@�MW����g�����q$��Rz��I�aP�K�#8�,�J+�ߔ����6���$n����[0��n��%C�p����'G��H�3���X3�p�t`�.z�ⱀ���!/��_�}^J$���Ã��u>bQL3�v��{}1'��9:{��5@|�LN4������(�����o��+/����vˑ ZKx;��#�;�9!�t�ѐ�����ƿaf���%�����=�B��z 1��ٴ<6��UR����m�ٝ��ϸ�����ex�bFH(=��H��F(�/'���B����ܷ�O���T�>��ر��v<.0d[�����y�w~�97�3�p��5�t{�M@�].<^֡A�_���;#c#�}1m�	^2O��v^���*[T_�^�CP�ޕ���M}�ز(S��=)��	�)��a��ԣ\�C�� �9��A�SR�� x����$��{�!¨\$��~�b���H��x$���e�g���X�
�xO\1lk�8smL�6?Ԥpa�6�O����Mf�;}Y=j���<-M��∆�^@2��p+�qp*�I��R�^M�d���>SP���4����6����K�b�ni��s�X�z^L��#s��	p�^���*�{6<�3�zq����[+���$�py��_�sFɵ��$,���HV��Ҥy/l͖#�*�lH��N����xr��K���޶��~�7	SQdct���QT��R��8��i̡�)yҢ1�_�g��5��YA�s&�_@@xu����b墌���9n7?�/��)���n/����d6��I)��.�!���Y�gc����[���6� �{�p�2Pm��0���}vl1��g��'lR%R7I����>�H��9��!o���n�s����8�t�\<S�6�$���C����}wl��h4���`���Ծh7^bd��N�1.=���Њlp�{X��j��� 4��� !̏���>���E8�n�.�̳�L���z	�*��T���k�u�;�/Z�huZ�jC��|P]�S��̪�<���얆���m��"d;Zp��D���6�G@����fH�Q̞.l�9�q�6�7b� ���Z����@a��Y)}cr�I�N��	��oQ�m-�]4+S"����To���|:� ��Sn1��A,�$���bc@Tj�օ'�:}�Ҭ��b䀋g� (����t��������U$[��u�� HV���X~֘��d'��l��+�HU�Eff38��t_�5��&�$�.2��w�7Q�1f��Y�d�J~p9vA�Ix�����/�ad�b�a���^��˟|}�QB���PW{���!A�K4�L͂}�=�ꋰ.�p��^�$+���cr#�̜)"ċ��?y��<%���E�����~���V
�u��A��;�-�uO���	�9b<@eQAe�o��,�l9����%�����Z����oH��4|�kN�,����g^j���L>B�?MFLe�_Ӟ���xv׿�	F�b3�'KH����O�b�CK��̚����N��O&�
[n6��I<c� �yw��+j����R�e��s����
��'��M�s?;��� w0��/�y�d�#= ��ɱ)�~��>Ԡ7s9�F�z9?U`%񓞧�TH`��+2��h��i���7�y�d4?j ��-@k:%/���u<�n�2�f���`Ƞ�)ПH��tJTK�/,]�rB#�#��+�׶&�Zl.i/�c��Z��L���(���N�"u�fEݳa�-C�9����bF�h��r�H�=�ݬ�|&R�s�y�_�����o8&��3����e��\���ji|���ڗ��dJ?�s��BO���BE�r<������j�*}�%Q
~����KH�Bv������0Y���^�_����xrDa>(��w: E�E�i�]����z�fոz"�Ǻ΋;�=�*�Q4�־4J�z�����u ��I�1P^��錿�l�O�4$�E~lb�@0h��y���$���]�6T|M��;�p��
X'.D6u�_]�?F!��+��ό�h����	 +�WY�0%��.���\2�ˮ���Q3���i@��kB�"�(j�7�qA*n�Mq(�W�B����b).yԽ��M����{���������$�����MP��p���jjBe�8�ko�T,��/Y]���gѿ��{��z%F	�>��\�Q��*�Edc��R��Q<�TF�D��lj��^mXT�4�ǯ��3���5?���܁Wg#N~�c�GU����q5�:A.W�;<)N�Z�b��|��Vb�{?Ϭy�[�L�/����"'����f{+tb�@�0V�X^��Bh�v�l��f��$�'��d0�툐n�"9xu'�$V�.��=U'Jl��t���w�njK��F@^�^�uA!���T����s���
J�1
#̵k���G�$�Z�s(G��I����g��Ƭ`�l�z�qZ�(����v�J�>�R�6�b���[#�3{f/�o�I���=��b� �|�۬^����&��X�$8��-K��� �b���!�KdT&�o��7u��Q�_�����1����2��6'�gd[?(�D�M�j��YJ0`h	v��8�;mi��/��S�h����9�R�c���C�x]?�4fFZ�O�]B(�,�/dUl1�k���J�������m.���%�#r܇�N���H��L�1y_h�����^�wXv�1��kDgg��=и�V�k�����\� �O��b����� 'hZۓ��:��́�)m>�z���OL�����>������7E��^\��#M���hlφ�Xqu��W9�WǴ��p�H!YQ�WR#tnu�?Cꞽf�^��RM�
��J��W�g���I�/��x����@����a�vRW����5CG�٥|�>�R���E�\�Ű<�/��5h�������Y��Eeu�J�lx	lk�Xo3�v����o𯙊�3m�z#m,��xX��s��� �+=/������b�����Ӥ�pm�ѳ�T4g?�%��;6�&�<�BOr�2��]��@���)T�����Ӊ��Y/�  m	��?Wg�h���"<�Y�֎���#�t�<���+�#��|�+/SnQ"ԝT�v� =����[��(���E�7���������I��dU�V��h��퍺ȫ�3���?�Sܘeܽ�l:-2���Vq�Cs��$`@�X��Q����FmM��	�/�)�d�u��ҏ�����+�o����b�ō�����o|�WL/l��[S�+t�hg��`���.���2�gu�D�����^	�H�D�En\lKQ��^9}Z��S��TPV����d����!HJ���8�(�"J`f��<��*�њ!B�5��o����$�� �,���� �Ж�K�сe/C�6Ϧ�k��e4;���=Z���s���I�W�I���!�џ=�P����W�xi�ʼp��,�>\�:��e�
�rY�z|w��bSu�@��R�N���\�01��eޣ�����_�N&�x6��}�x����qI��08ſ?sO.w\Qx.�L��HBu[���(ه��#�H3�l�hEV&+��v�l�x2!���`��p����36=���H��B��p*�W�}�Sc��j�X�:T#���G]��}���
T ,�9/�e�A�!gJ�K&��uV��Mo���_�評jAg�I�%�R*�ɕ�Ҳq4�;c�C�hm��Cp�]@|8��ǩ��Y1 �0&�$���^��s�J�O�
`C��>3�Y��t��pa�u�?�'�#�TY+����K����A�" j��ZG��6����5U"�9�6£�R��'�7�5�;xr���\~�~�h*��*̆�K���i���Z��Bs�ǡz
,�N�=��H2=��OZ���x��S��L*[p�gɮ<ͥ}�J,k�EK�]�L�1�f�|g�$���p2Kv���N��Q3�Uz��+����8%���6��G����/et�nm�T2��H7v�� �;�|#_J�oj�0{Wd����+���lE���A-N���{�9g����V���I�m�V"��u��ʫ�6�d�0B!X���|A
�V6�:�a'�*q(Hzz��q��̺�h�T��v*�-�뱩X��u�B���� �Df����?"bN����+���8��/Ĕ�g�ߒ2N���e���	U�^#�%����m�Ώ�s���JNJ ��e+��J��B�K�Z=�J\O$����I�s��|;��D��d�˥��{�0�Z�>�����h" 2�V�EQF*��my�fBND.���F�]<���/#�?�i7��	t������l!Ijo|ߖa�ꙖT�ւ~��Q�=U�Gvd��8�9��˔�z"1Ȗ����o��]i�V>MU4�m��� �'��*j���b��L��fN��qj�K��22}�R������~��z�)cb)Ѡ���<��y�`�9u�,L'��.�цB�>Xΐr{I���Q��6g���'%"�;�%���h�~>���6�!��1��c�'������Z��3c�����w8-�E��c'�e�g�,��=b�Yl�����M|���Ҥ�hYv,�^t�t�H���$�Ԅg�䋕��	7U`]M�,�I��n��]{p[���6y�G�p�I>�O/VC
� f��Ny�jM11���q0�i��z�̿Ϙ����$��Tv�[���G�z��9��Z��X�e�xwh`컍=:@�-�m��$G+��܌�3�^YsI�u�Z��W�f���'zɶ����/�A�m�"�J�	|f"��ёh���EE�:�m5�%
O�2�U`��w�Ҫl�o�W�br�w=�h���;��O��|3u��V�D��w@��[{����g�z�b���Ɛ�7��M4�����_0e�ٵ�1���d�L��CL���\0���p�xe�o;*���R�w� e��J���c��]+3�JS�&��c��1l��f �q�%��N����Y<���~-�����Ti9�R8Z��zgI��R� �Pn�(��P�h��C��iA��	�=DQsڽ;ai
�"���j��1��K����?�\	%�5�U� �]2j�/S�z����yp��6�p�@�'�uk2����H�2.I�m���`�c��<�(��I�5�Fϖu�������,�0���<�����f_�#���>g��_��b�p�)����}�Aͥ��Wrℇ�����D�뛶'n�WP�ו$Vݾ֒E�;�J�ꗐ��P�fU�!B!D�E�N��I�tmʽ�LuYE菅����n*�"L�P��\�y�¨�=�[���Vsu���uC��n���s����v�!A���=�M�D<�ut���|F���i�C��e����ՉR L���w#�6 �X�t&���a<�/�  #Kx6��+#s8�:-@�}%�n�l6�/O���N�7@6#�i���>�
�yEN���n�?������73�]3h��t�oWً���U�F�L�
��}��S(N}�N�v�© G�b0j1g��T`C-�N��.�=���E�}�?6�}�[��]�66�J)M{��N��-F҈d��`Q>Ђv�!��^H�o��LA�m�OuM��qW
쏎�[7��񤞠߾�<����W��0��:���s��Җ:��3G1���ݠn��v3��l"¨zE ��j\b|�����6�o{
M��2zN��8�p�W �a�n�V�>�Ii�K�a0P�»*����Q�.�ǜ�-O���$Ʉ+�j[��0ލf��\>��[;� ���'�:�|�J��V4�d�U�,TUj�������׏��8J«I}��+$�#X�c��'�F�paў�-��-�~����n+�m�r��.Rx;�/�w�ݚ�V���M�a�p�׮��+*�L��RI+
�:��!t���{Ƽv�.`��k
2y��=V��"��=��g��"����p���<t�S.Zz���,@
R.����N�~�&�	��~���zl솘&����7Yh�,r2aC�O׿�������h��0S���y��~k���I����Y6�.wF`��.u��֬飀����][�^홮O�F
�[�'��tӴ�)��u��uTĞ��uʒ���YI�����4��+���`�99>вA}���rQ�\�Җ�0��6���֗R0	2׫����gf��V>�`��Q<�e5�q��F��#"8T��d�B�E1�썷��6�$&��N@6�B䉮�;�����=%�u~9B�J����{*�^�$[��|�������D�'�<ca���=�\�w2���"&�g$�xr��"zX���5��!�g^�!�RܹTxc�N�0�5��t2?|��*r�h��ǝ���IPA䴢����i7�?�������l��ኻ|�t*�r*���h[�MG!��F	ȑC�;L�\��Pl`��[�ݬ���C��E?�q�ǒL�C�G��,E�f9�����yh鏁O0����-D� �]���͍N���V��tZ���8���\sr�9O�n�R*���d�G�\�kuf��ں�;w�, �v�l��Gme�g�WQٹ���t�!Rw����e���s��&�>z�fS1�#��;��i�����v�RBY���@��|n{�o�]�)�GtmX�0�[��兟��0����̣ 3)�ɳKҖ�2�2�KZ��2ٞ�{̬p^����Ɔ>I̩"���k�R��Y��d����h�D�rK8����=��}���v��`�� ��8Gkp�ǅ�/��i�����D�v9��O}!d��p �`B!�w6Y�xm�n]f6�FrwP?8�������7t� w`�{��Ք�B�s�Z��˼���0����1H�ь��Ì�D>�Ͷ"G�\���ХZ{	��F)4,�r�J-6?ܡ�����T>��A�R��p��p)0�p�t��z�u5�<�!�Yd��Et�����]Լƨ3�-�>��t9� ,y�25�T.��}�8\�<��	};�A+�b����Ż)n��43�w*rSFoˮ�7��Y��I��v��#���Kv��} -�����Kz�H���~�տϪ�@W�=y<'���>C�}85u�L1Q>�c��dЉ�)O�LS05�ϡ�xy����=X�Ɯ=�J��83	�l�q��?��H�����
��(:���~���?@ #�M��M#�%�EOu�1=���T���+�-���'����ڰD�p$�S�ܬ�nS58����Ņ��ܐ��QOv�{��x���5� e-0����/]�XV2�|����_K��~��)KAͤX��b�p\W�w�I�P��Е����=�-�oq ����г��r��=�k[g�S��^�R):Rj��ՙ�j��f��
P/QL���1'��o���'v�G�A$7a��hWH'�.3��C�xx[�6�-���,Ue7��K���B0���ܦ>UwN,��K�֯ =g����,ɳex^�N�Tk�
�U��|g�j_h��H2ncҫ�0q����K�؝�5N����2�]xb��6���y\�魛y�맶��_~*�iE�:���T��>��	Z�p4��ٙi��I�I���*`aߒ�L�x14#�Y�f��pon���CѲ�	c��>����B-���c�m-�� i>{}�+��c2�>OؖK�;�;A�q���h$��D�DOȕH�n�(����.MgI�C�%��[Ο+��CR�f�"�qW0�m4>���C�3
�2Lq�����&$W�KB>��6�%��?XQ�?��l���Jwojw���lҪo�=*dխ�j���V����V߬�[�2˧!]7�%��;`� e��t`lU�F L��y��7RNCM�*�cP���4�"J��n��2��ۑ#�4�&����~< C�βԳ3I-�������=v��U�Ԝ�E������W��@�]'0�$IJ՚Gw���mL�t����g>�� �l�	�)�R~� ?�d��~e8xg��-��0?DR�<����k��C�ҽBȰ���^ 0�}/l  :u�{� �{9o���ِ̀���8(�����{������wU��x�nzr�u�D����2w�)QFc;����'�Z�!�~Zם5�Ќ���21��ט��r��x��4�YDCB��3���7F��Xu|_Hs�vu^���7��w��"k0��ЍY)��
�>��l��ɛ�z� �P�t������d��|dh�-!��q�#�_pk/G�8e�v	\��C&䕼��@�"��[ϧ�F�#�\>���G��>j(�1	��]���H����z�up����2W/�����ew�mR��$����0E_�~�����mbCx�� ��ڧ��/���u!����Bql)�/��>��0@5\�c��q+6W����K��|��*?���h� Uy�@��:�C9;���E�����:���:��,eƁE��w~n�}t>���^:�, �U��R�9��_b
7�PD�B�n��&�<I��ɣF%��p6��<��:�v~,��ųk�6����H#�qU��Ԁ<e]l� N����"*d� S���5>�-R��*=$�z'�}�����z��/������I^��JʲyY���hiƀS���d����m�����I�INi#`vny�C�$���f���Tn�5�8�� ��4��\vm�8�#"+m:����r&��9��{��4�Z��З�ת8�ؠ'�61��.���h����lAX�� �Ps�gX����e��Y�юf ��J
�UNq�g�U\m��8���6��i�ʻ��n�Y־�?&����s�e�4�/Uq����fdZc;&����?�����RPQ�^=м��|H�3$�V�����O,��ZXq�X"��1�,�إw��n{��'re�݂�D4��?}��}���)(sM��)�\�'S�F)Ǐ�|���3��	���5�,r/�[�
�p�P�H���G�]�gu܌�u�-����?NMޫF���R3#b_q�t������֗�ϋy)o`)��zEOס"N�����i�[4���9i����ˢ��qq�NK)ԅ���%j��u;�Jv�����d�ݤ���!)^w`�1�����!]6�F�:�8@�5��C(�����Uv���P�����O�I�gu��P{b3ft�Q}����|�1�V<V�!n�z.9�u�Ǘx�Ý� ��to(σ<2Z���s'IbY�x鏵f߿q�J�G�S�P�R���+1���ܺO��×.g���M�ī`T�����ij:~P2���t�M�{Uj��6����Y�$Q�j�{�e o����'�պ<��26j.F�@b�9$��S�$��O��^��9��&�/����YċH��ف$�^P6��M�s��"ݻ�Q� ��{d�y/<r���v�eQ9�I�#}ƿ������\�Ǵ��zk���DjiYs��QO`w㪇il�A��q�N�&a��Ț�cM���+�~��ݹ�g����90q�G��}�ĭ�,%�{�б4��P���ٙ5�}d��rF�ý`��#n���2/�~�&�
��5h��s(tq�m�K
	L��%@-KG9��M�֮r�O��_Bw�r�z?F�[��ι����Ӄ�){��[��`a���P,3��#�H5=F��g2B��}��)Г�/�êB�����RJ�45��Kˎ��ȸX٪*�
��I����ܩ���*KJ��v�zx!��A��٨�Q��b�%Ep��8qC(1���4c@�>HY,v 7E�2�̋�,�	���h&�BF��b�����8<�LKZ{����G�3�����(�PD�V���#�D*R�E�a.���)~��W�/scg��_ߢm����5�	���af��~}M5��|Ke��`�|z��6�P��'�0RB�׻cZ#��DCl�br8W���SIk*����k��^�K��u������Jx���CFi۰i��rY~�"|13�S��^�{*���s���ʐ��s�U�z$Ժ&0nv��s�r���>NN�1}����6G��;�ݬ�YQ�H��\\�P�Rj0x�÷Ñ�[2:jb�ˤ^��� ~���8*\��u��F?��mG�{�ԥ���Fu��~��/�C�q�;C�H��G�Dd���9",;�gSh�
�V��oX2�Ȉ��HP���:���W��l�? :2V�0���~mݟI��zjq����ۿ�ލP���kh��!H�F4��0\���5}����a�_�����D�3�^����s���h��28�&���a�`?�# �x�b�>�?ڒ '�JbΆテ,�m���_*OU�0Y�Ze�@
q3��TKO�b��F�������m���tΉ96�k�R���sP����/#��r[����H`��wI��x@��|l*��[����Sm����B�s�pK0�Dz���&���#ND���j�~��+�E=�$ˣ*�~%P���:-1�}=Ɏ&$�]|�c�:��㑼��D����B���;�LS����A�)��g��R�ns�z�x��`����/ٞ����0D�&n<'���4FX�]�
�T��h���p�$[�a�W����ꚂD�Vb'gG��Ƒ���D�����\�d��Z���@ X\���'7�������`����Xie(w��u�XCF��X����^�d���*�w��>P�<P*D=��|����ٿNq9*�4?'֮7�����奥����M�
b'�����RP��­���7���H��*$�L~7)���‱G������|G@� y�B��`��yð���p�瞈�:Al��V�(ʜ`�l���u(_���Ҩ��K�����:���7C���,C�����L�`����D�7�%�8�W�qgBw��vU�pVKb�ҋ�rl���D�б��BE�����^Nx_=�2�͑�N*}��>�aJ ����IH�^=�D����`@��h(]�V!mc0�;�lHW![/�q6{���'Ь���8�|aD���&��7��'b1f���ui�H�`��&N!������~�ֹ�6���N�BG;�TR" s����[�K[C�R`J��#w^�������@�?,���Yb�ĉ�%l&�)�m��og���ǂq���֑�Y��<�yGѽ�7}6{�jF��� ��K�A�E.X�7����mu��C_��_ k6�9���e��H�cL>��K=�z���*��6s!FԤ���jΈ�����c�D��U"�<�؄D��5�,�׏�T�=����O���G~�Z
�,{��B{�%
���\�iR�%ko���=��s��Z�1sbz�&�-eO "<�k7���j�e��ե�w�Ȟ�;�:J1�.C�ڳ�5[vM�f��t����,6:� �%����ڒ��B�쩶�o��,���v�S��.;l��Ia����t^�)�2(2��'D����-3��T���o-��+K3�԰fy�1Y����ǀ� �A-������*�!��=���mX���K��{����rC�5������.�Am�Ŗ�7)��g[�q��xW��I�(c���w󿯬,�Ӫ-�8�&���F�[�Ґo\�6�5�7�t�7%�u �ߔ��˔Q��^�ݗ��pyO��=���H��K�	Tܛ�S��S���\�z�>f���N$�.7�����>N������\����}� ���d���!k@��� �|�@���W$��O�.΢-�X/m��e:�M<�vW>	hA�ض��M̶���!�{z)\$��߃�*i�^e�1+O���0�(n�#�=�c�*��=R�����b�6O�3�O
uVE��*�[��G�}F;8�e�J*q��f�$�^����Z��4��}��N���=u�bVy��Z>aWP�#����y[�t��q~��������~���=G��r�s�c�&lI�t<��Y���py�, ,�G�;G36�47.#����g7���f<QU@�Z�$$��e��b} i�M�g>zj�'+�����(2qU6������m��S�sT�>?�p���"�����	����i��7�nPhF�Vp�s��!�jCގu��=o��6U�@j�}M���6�_��v>0�x���.�
�)�ۺz�T4���觷�.i�Dx0t%�z�����/�p��2�zt��_� 5���ݮ����Id6���6��S�-_�'ժȉ�ʌG͎��G �����a�f��,�ڌn�1��s.Y���!Z�|F�����ծCu�W+C+^�	���}�a.7�"їT,�j��G{�����Є1{��G�o��PS܂�N�<����������[�3���}~�`�]���&-ڹ�" }�f�[��t�]ģ�����!'��9�pjL�pԬֆ�S����Q��;�g�c��acc}��Z���8��
�Dݚ{�\��4�}��`=-М�K��:�1_8Ѕޠ@�>��"c��p~Q��+9)�ߺE2$� r�d�ǬS�>��ݞ	"�k
U��4!�z�^�D��٫Y����n2 3,��C`)��yW�,�{�W�EUH�B��p��l��o5�:�{��l��i����|�I�D���zcae���azau�@+����lA�{t���o�j*7��F��Y�m�u���GG��A��J0��~p~�#)��e:��@��~��ٴ�k�ۡM���,�y@R�Wb�~���?�L��s��7����P�:~*/�1r�����K��>Wl��P�p���wf���B�<��@�+]���m�3#4����䩃^0��5�r�����6�e�P>�4 |$��?Q� >�шٵv�M@�ye�߽-��~G7��G��a�j)�S��ilke+�� �u�㨅���G+hOM+�.��9�@��	������n&!��I�}�Dʚ�F�g���j�m���y�����FG�2ڔ��Fp�M���x�ura�g��$d�o�ӑ%ժ��ā��1l5�4Q��IDY��zL|��ٲ�9�p��&Qk}���j!�h�`M"�������kr�~O��0Ҕ�'V�Z��Q�?������c���Ŭ[(ӵ�́�p�ChVu����TR��R�O�G�Mc�h��^����	f\�谔h@-�������4���-�ye+M�[���&�%��@��A�_�i]�� _���Øb;�7����`���L�{k�i�װ)ȴ�v�E
���~�ΖJ�ߗ�'N�AHh���xl%G��p�T$��3�:�^%����L�������\-w.SU�߂�g���>��e�?���T�b�����"��Z�,�����fh@�FJg˲��;���z�Bj9�O�YM���aL���4x��a�Φ��<I�\p)��xܱ�M��L���A�!QSڿ\���?��w��-�G�d�i%1��^/�w�y��C��%J�
�*�ɱ�3<��o�,^�c ��]��Џ�}.t�Y�����J��5��x!�
��t}�.��B�$���V;��3�P�_���7���(�s�[N�~���!�ۨ��[9f\�v6�CO�\�����.������L��
�O� ��)�M��X0���Ӝ��E\V�Ǵ�@t1�mu){�]�B	��
�fe���E_���
P�#���\ׇ�u��)�#�Wd�&«��A�����g����N�X���E����#���OD�F2-Ovh'��e`np}vI�88��*�ܯbK-F��@*k��ܥ�R��r��cGE8��-.C��3��
�ծ)�~�~淁B�U~Y�q\���=�Tw�q�~����n���=���c�@y�]�H����G ����� !��1�<�L��t�"(�>x���{��5SF;����W�s	�a��?�IDb���G��K�
"�C�9`�d��嬡���'i���gh?c1S�uy�[�~�U��|}I�SpȐ��7��-�<uډg��m>'m�9(��T_/�vٚ�0����2R�O�4D!��h���F�̍��3�ɑ�F��?�,�Ek�A�[|d��\�B1�~��4�^xF��}���8�t�My7f��z�^g7
�|=46�2�ࣉ��tj�����7��/�����e�<8a��
�Ҧ���e�9�QВ�4����/B�H��&�L�gx��I�W�L��3��اv��s9�0���E�	%�$h��]�j���b�� �iiN�w� ����Ec���Gw[�h���_y��
�G"�g�2Ӆo���v�ĭw���ަ��rj��Hk����q�xTuG2�J��W8C��mD	���I�JEz�vy$�F�yZ6�7��<H	 
q�n�D����:j�ڬt�8:-���9��%w;�Å�"Nԯ�G �/ٱ?v�K�rvj0�G3�C�5Bx"�H��l�nAvz�����%_���g@���8^0"�ݮI[�hNR@�����!PK�|!�}�6ҷe�����\�h���+��;�抅��t��r�зq|���>�w����k���0�L���r��E/Kpu�S�|Au�E�x]��a����9��3wc=�+&����2���y�C�b?�n�PŦ^��(� ≮�.�}X⣩�86«=V��#J�	wI��8->nk�0��lV���X�������zFSK
zP��%�8v)�B��V�7�<���~U�ŕ�ǡ���WX-���:�)�Q�)?+�7����5�MQv��x{Z��R��9ˬ[oe}��p3Ċ�n��l���D	�uj�=d�*ŭY�#c���U��E���#�K��s_�L�=�hl=m<R{� �	ɬ����qq�:�i��ο��SB~��3d��Zݔ����y��V@E�^4v_P)��Ehɨ톭�7��5�b�<WuP��C,1�������� ��h�}-���A��ZD����'�vn��pӊ�LI�lv{V�L�(�Q��,lbSZx|�Z�w��0r���9=�	T�A��O�y�'߫>>����TM�/T�k"pbXNSj��X�HnѢ
�%�c�y)K�����b��M$;��ٖ����rXc���~U�@�3�������Z���W{QÍ��wC1k'��Cw����S;]K�@�V;�����L�p�P;���} %��*��{3�wO �]�C��1�m�w@7�Ek���[I������P� 	Ak�,��z�!S>}
�D�@���]���hc�� �W6�,i/�k8y���ۄ�0���g�?�0{E�Գ�K-�l9u	������m��$�m5��QhoK�����w��D�˶k��~�s�����H3;
+NyI��!��\bkZ5i̤ՌK�o(�-��/�u cF�B!��M���Nϒ;�	�2G�#U����b�|�úk���%y�vz��CiZ�3�-�#��b��u턇��yS�Cu��l&�H���O�? �/��5 ���8������L.B4�x�'l.���J��*n7�ބ�L��x.��Pd�YT^L�lp?�Γ�TfP�y�SJ�\�KC(�W�/�o �-��� O��gs/o>��\�)4C|��GF��v<V�!]�|�\'��Y4��*�X���f>�d���qt��sVixl��U4�ͩ�ƔK7����.�jĎSE�6b�q���奤/4�b�[��~�H�ah�1|(�x}+w=Θ�(�U ��7�Z�Bu�U����=
J-Ir����P�]�u��B�i�~pAN\���I�G��I�:q>ZbH��f$���;��o��L!c�O�y��3U/�3J�_0ĂIc=�LV<���>�&�vL��s�s�쳋�
J�O���`��y=�G��R�A�σ'|q��A����ׯ����)!�^������Q�s�b�T7��'��<H��~�և��67� �AHq�jy�|5�Ȍ3a���yQS�J���Q��$���:��V=A�9c��*�.@1K晪	���!E��OR��0%CP�$ϗ�ڿfro�pl�r�q|8�4����8J�����ѳ`�	������!P�$���)�ܭ,��r������,1v�=y���_�W�W?��z�M�)��O��K����r�(҄��Z��X� ]Y�ωU���?ԃ#��c�;%��h�Z�T���b丱z���}��SSPc�@OL�`/w�Mic��N��([�>�j��9L�%��	��T��A�$ �[��S�>�#	�H���#�E�H�..��\��&l�wF?�h�*��q�d>����"eomw\R<g�(#E 1s�7֛Fx׹��N{�k)9C�����Kϕ �Aݬx
=��Ԕ@ב����J_�����(yμ�"�=֏�x��n�G��	Ae�,�W�X�g��:��Vka������a�ׅs�iz�����kK��x9˰��Nak�jo3+����+�ɄJ��ЎqU��hO�r��l��hy�Q 7Q�R��f�&�o��Ki��.�Iy�;|���t�!�7�3Q9+hE��o�6�l�%z��z4�4�T�[�Fk��fob�4n6]��i��.�y�\<a��b�ZX���
n�?��_��P���F��V���>�L�3FA�,����ɏ�x�!x
��s4\��q����& ����6t����k����8묐�b�Ϩ�Vw[M��u
c� �>��^~)m��O��z���'?�i��0�s
���z�Ċ�	����{�ĉ���1���Zs���o�54�o{H�~լB�76��;ґ�k�ZM)f���ky΁�)^"F<���CZ�����{�_��B�#���n7�8���p��'�[TDy�^JH�eol_@	� 6-:p��Ԥ$WA8j��z�Ea��i�Y��#����KW9d��ڎ���}�ZD�^�[#� �J:޹����(�,R��b��i;�s̞=����������A/t�<uX3�& �f�N�W7\ۚ��)��ٚ%�lo�&�Ȝ�9���vT50�.�Af���a.H�T��_"x2}<^�eن�o����\���Κ�ri�`�!O�V�F��f~�����ʩ5.�G� �b��3K�`�Qi���C�3�7J�! ���q�?;e�R䲒_�y����,���"0�>@��T"��{0u���Ҝ�=+ܺ+U�;y���˲W/�/ctAjH��{�^l%eȫ��!��2�>��-�2�-}�$ޒ�H��������b�G$�E�z�v��������'���8p'�ގ=ҋ�Z>�`�"V-��b[��JR�ט�7R�ý&~|��I���u�5GwA@tϩu:~�`גjJ톊�50�z�����;l�Ԕu��tsm�`)
S������}�[�'g�G����5it^j�ݯ�V���"/�~)�=���O�u��T��B��͎y�\{3�H�s_�N�r�t�c� B|��38:KyY���B����	���h���#���m���X���d�QH��C��,�w��`�~W�
{�BrWAJx�5r���DLg��2��
)�x�֋ƙ���_T{�Y�)�o����^5H9��Ԯj%��B#E^���Y�y8��h�qx_��42��Z���QC���g�d�T��`�˽��]�1�-�i�-�*��\5,���(�҂~�C��a��TkyJd��)�a���a?�N�%L%'�0�r�?˛���4�LM�kb��)�Ci��=�C��z;����E��&0�s�w�H����EFv(�^P�ދ��~��j�π��6�ӝ[m���^MNra��6�6l���g�^5t�}�j�&W���3�N���9�.��� �h�:g�N��r��K����k
�����-���P�U1��谕��I	�m��烳��]%����ac`T��Ġ�{�"n����y��5��l�2�9&��[�zisG��
��|f��举#����Re����L����� ć���v�[*듈ZGĺ�Th�0����fh�ԣ�5�姁f�%�zX�9x� )��_��10u�:آJ=��yT�Y_'�:8�\��[@��C(�<��';g�G����x���*�-��Xg��C��l����Um��N�-����,b�§S�x�?���'�̝^��i-@zct`I��zb�ܕ�'���s��qTV����$�zL'hɐ�x�=N���Z����� ~�������cn��i�`�n�>Z�a�S*0����cK��]@��'V^<��uC���T ��/|N"��0+J������_��b�<J}�����g�qK�`,7��Z(Zk����6����r'o9K��4��{��S�v�V0Օ����S�t������ɾcp�����zvQ[�ǡ���f�?&u~_M�mO<ur������EE�*l�9�HR�2�N��A��?D�|�~0*�Zf&|�˳��q����� {K��t,�Q��l�1Jdh�}�x�����8���0碼#�纐i�P>�>�e�h��r�tq���o�����d�P�$��d�$�{�S�qv��)Og	:�ud���T���[��0,���{��O���.�\0F>�R�@:j��P6��G�>;�j�ʱQ��|ZUQg�'K%$|A6�C�>�s��B�,��#��-)�g@'��[�;�����Q}���Yw�̘Ht�@�`Vf(��	��y��>*hiփ���s�k��_ډ=:����[u�������ȡ�
6�>��nN��^����ΔM���H�Y���s�2э-ܶ-,����Y8��)U���G�W]ò��[�ayY����}�x��&tP�$H���b�t	'�ܳ�`�!�	����������L������-�S*uI�\���qld
�3��˞����7\�}ǭQkZ��"S헞1__1����J����qG@�	���ID�M�qѻ�}�Vj
?\��%1ق���O�1s�Z��}����q���сnIG	�/���R����1�	")��H�eK ����z�x?���Cnm�İ��^j�-8�'!Hv�B��G��y�`�s��K�B�p�ĭU�M��~_�v�hOj�����\ý�3�����Xc���zu/��k�����C �D7M�'�!��XVǽ_��To����S ��)�٭��=�[�0�t�&)�[��.aH�-�>�v��2$�7�������Q����Ca���$:F���p�|��4�j:R�TW���.s��C�U��l��r{�8�:]^[�����Qk��5���ή9+_Pk�z끎�m����u�0����T�z���������!_R��&@y�H�c�V�u���v�:�b��.E�-��ۼ���Qbz_�����1��\�?���ۯ����bk4Ex��Y@Pϡ���<,�kOzq#��l�sju�ې�Z�XՒP���XS��ڕN��C�^2�2��g���e�1ԉ-��O|��ޔ ?t�La~���Br,j�c�l:{P�7+����X3%����z-�Hk�|ī����лJ�MWy��9���pz��DT �=�R��V6\dS���%�iW�%i�8U���m����͟�\�Z�����˰G@s�,��<s�Ɏn�h��Y赲��8�*}�d
~�6��b+�����s�[��DF2�R��l�u�4^��7 ��t1�?�n��xI/���sG������c�������S�ĳP�r8�]�p���3���EAg]E�6��v�^c:5 	ރ�`�CϷ���O�Np�}f��i�`c��)�h��r�̤�ofA����XL!ޮJ�[:�oB"�
���5G��N�|�k���,+�}�%P(npw��1�g��U�l���V�WҌB���#KI��e����z`S0
�a4~t�/��7C�Y�� (�,���Q�\���uJ�(-�j�T�^�А��ۆA=K9��yW=1y�'�.^� ��0�MC2�ǹ/:._g�X7⻞{i�t@���FŹv�5�k��[��;���2�lK���V��-E�La�"��Ob�߽�O�c��q�	r���i�}�e���b�4�$�����;�6ƴ 3�K�;�xg��rD�D	�n����|:b�c#�Ly��Ƞ4��ȗ[�n�d6߇Ņ�J]�>m�Utc #iU�Or���t���a��ir�E�i�]yrGEqW�j޼�C�h����#�C�i��������P��N_�{���^u�d��!�������$��	�]�F5ax�o����/cj����Ų�,���RL��E�9Ҧ�6r��ɺ������?�:�m�r�҆�<M՗>I���b��ⸯ��5.�Q0!Y���WCzm��Z����^c��99�������n�W5����}m�K�U�}���NsV���y�(﮽�!AS#5<�`>�G���_H�vk�h�#n:b��2=�� -*o^7��I�Ӕ�}���3��b��x�Ψ!B;(>������+��o���Ga��Fyy#��X�}n�Ɲ)� %�o5��b� �<��y�Ce!4��V�PCpyMp�+���vM����4�ӷ�Ĺ��bFo��:������m��p،�2�]$��[qq��߃��%�P;q�Z����U��OWQt,]����%�k���f���<Mk~������ֶ�.�P���������@5\�U�r���M&�g9�� 9*��s*��z����Z�!�����/Ŵ'��H����n�+����>|\�l_�&aR(
�b�i��Hiw���J$�`�n��	k�8���V~n�|[̦�r;E�CA��t��;�l&���T�����؜��7��dEj�`X���թh�Y����g=i׫�vǡ+w�V��Y����lc��!����7�R�T���(�P�����6�)�V�����㹡�}N5��>O���	?����괧��MvRD|�ƃ�J�����O��[�Ѿ�G�\B_FLg�n��V����ޙ�m�TZ�P������J$��k�Zm�־��"/�����ҍ%��*���>x�B��r��1���䆢 ����БF���E&kb_#���� &��V���׃ҨEK�Fv�J�����P��C�B�>��n�a�-�c��n�߽����PVa�P�rÇT8h��U�:���2��`h�ێ^��
:�����(��ZE���	AT(�Ym�;'�'H�5a�C- �']*J�3L�ƶ�J�|��N9l۹��a5]��.;�m�Ca[ ��lT�A ����D@�D�:7Y,���S�v��r�	I}1��t�U��۷�7�<u�"�$s�d	���KH�ubɲ�b��K��`�@�Q����փ����R��;O��%~�Wz����45�d��I�m)���`{P��d/h�kQ�X_�Z�>}����{���꠬f϶1�Z����Z�o��D�?؂o@�� ��YPg�ʙ��	Y�Ǹ[/��Wǹ`� ��cl�4T��s�Ϥ,�9Ӳ=�9���������C�rƖ����o�B��ް�
/)��� H@Ya��߰��a�V��͇@*��u�w<��o=�^N4b�ȹ���V�#,t��
N���1�I��۶`��t"C�,��Y�D��Q�5�zdfW]z�y�瓚s5&A�N���T��Й�4f5�byz���L-�|�W&���&��L܆p�!�I����u/ �~���1Dq`�D��XL笧+�h�'~���_�m�F*�&e��v�L�1�?�3�����2KX��.��tx�(�&���E� O�<�����]X���% .��ăj�a��L�;�d�<i��4��I����՜�s��:���DE������[!7�vjaN���W7(�6�N�,:܉f��V���ѶBLC5��S���Y�*B~ G����~(g������ۥ�P�
���6rQ���C�
?��ysG{z,�<�#Yc}W�Ӏ쩔 آ�ޖ}Y2�Z�駘��I<珻���mƸ��f�#$)x�xr+�M��
��L�	X%���I��O6�[ތ�2�F޳Fߎ��d_��c�������v��xɄ]K͈�AӖeKf�~�eIB�@$��=f��#@QYү����w���68?w9<�o{���y��=���H��S&R.����]�,L�W���p��1���%���݈g�Hj_l޿��
|�⬛¿{�qx8q�U��[R;�#�a�$�A��K7�YJ�gN����|X��1��7��������� 5��-����B�Q����3��0�<��9I��aC�ȿJh�Xʳ�qM��&B����6��,�WG4NN嫰� lŅ��so`����jK%D����"=Y��b֒�r���oKͧ�c�
TҢ�Fp�Yp�h��Zg=�@���g�Ɲ _^�U2�� �,��^`s(�(4�?,�t����ĵ"c�&bI���i��^�~���t��`}�)����
��~��;�oƐ��L T,���؏���X���2z>��+P\ʺ",�&ɸT^�R5<��;1n\�$�=m^�\R��\qj�o���2{�}1,�P��N>�?H
��8G�
���_T�1ɬ��0�����Lo@�Z�|��_֬ݳ��w�b�?�g�5�Q^�/�ޏ�=�,��
^&�v�q�iP�c�4`��V�N��.w��(#1�5�y�[�Z�_����n�q�p̓r�~����)��(
�'���5:B'��ύi0�U�?AY�� ۸�vԭ������ډ��N�$wT�˗����5JǬ�B��?z�<@��Ԋ�����l��J��NI��+������q�y���>����7d	kw ��9��Lx�T/��,��mn��m�?���<Z���ߖ��I�&k������f���N�3ԩ���ԁ�"�|h w1�����bw�'��8��t �J*x�H�W����K9��3ɕ���on��í��I�0���J��wO�r���6T>ZH��L�+75� �W�g�J$�&�����Jl ��A�M�n�]\/�J��	�S(O�h��E�ᓫ��O�3��}a��]��������_%5M/�h~��[�ބ/cEs��傼)���G��d��ڐ��\i�RR!g�B��_�� z�`����3�G��F�j&�{���]�oIJ�mJ�K��]���W	��= �J�%B*���T�Ic �n]'�������2�BB�#�m�aE�C�\�;�l�u�i���sE4�}Ή��cab�/�W��Y��56���?���}
;��(�Ş�ğ:U��e����pP˳�Ğ�8`8jgkX^>��lN�h��3�w��ѣ���$j3	�ٙ�]�F�����S�@�w}�V��A^�"��h�Q*�ǰt�R(�­t��XV��`�Oa/�3>\yݾT Q�_�0O��$�~@1�W�ƴ�I���,z�.d�id�(��q�� ]d+g��u����}����e��+E�	��r�� �RVQ�_lY�<�5�q������Cq�Em0mk�䯜Gnk'��Y�bG�SW�7&�դvk�X��k��& }�~�ְRE@�{A�-�Y�}�0g�_���1�f�{��eѡ�E|��Qu��[�@T���3�;�1%0KM�1�0��P���yKX߲o��_��1"l���	����=-���jBj�_��w�\��-|	!�
���B�-��h�&Uƙ��\ݲ�����|H�?
嗩D��5��LYe^K�˯63� {���ZBH�86��G�FpK��%��M</�� �A'AA%���h��;29r�S���=t&T�k�}!ܝ�`�Ԡ'ʘ[��ͺS4~r�kq�M�.J%R�+3���_��i�+n��ʀ:|��+)��Oy��/P�ډ/
A����g���w��%�E�}�����
����w�X�����d0��D@7J
C��S�$Jh��.�j�S�ʱ����z ���c�� Q�&%��/�G3x6��ᮅs�J�|4��h��O46�&�(���r*��ۼ����c[�%�itEϾX���E.�6l�4�ja@z#"Ƥ~���웖��|�xJ��#�*W+psEE4ߍ��@T_���zo��fAdƌ��u=f�ɉ�}T�֧�����+��&*�	�s���g_|D�.؄vTI�:2E�G�H_�7Zz��^��h7^��UbNO<?��T[-��H�� ����?�W�}��~�Kc�����r�ě��6� ,F+��a-��G� �u������{>9T�D$ϱz2qT�@���5N�Vt�5B�:[��w@���K��|�xE��m��|��|��\W�ã��W�"s�Ǣ��8TC#S�;^8>�Ͱ�W!#n�B�,yv��z�D��Ƅ?CZ��p%�dd����H��gg�Zr��5