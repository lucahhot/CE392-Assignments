// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
N45DbHs+Zys+eg277DltFoCiGHRNtcirszfQLgzXj2pZ1GH8GDVSRbNgPn6KPnM9G3GyUmjF/9/e
sA89lEvAL/u5B/x2VA38ZHi7dncL2eEJeD58PQUpVSokehcNa+X/NM5hzKYsLTG3+YGUzlLulSRP
30YaN3eW3DAKZbu21hQ+x6cpMxl04ChF+UV3tz0vdQiRIG7XxfivXmXtbgfwpqLvDiQCEouLJURF
Faimvg9F6fYi03q/U8lbEuyhbMS+esSgWnryTcmyOG6QlIYUfNolN7SRYmkDopeEKvK/rcLbwoUI
6fOCCeGEDBPReH9zLa2UN13c3I+jypOqFD2NVA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 27888)
u7lBdaUJdRqhocgffqvOyFpCSeuqhmWMyCY8Ks3w5yfh92Qas93HBFki174KC3W3Jbo/X/GIP+df
s78tJLwLOloMRhBqBycyYB40pdZ5TjOfykckNPfjwCmmmhoIx37twqr19Q2BX9gZe1aWowrxVfVa
N9JRvy02x8ryoqAEoiCfJKHIaVOq7XfnM5rAtcBQMp1Ruie1Nt+zmTvQt1kfyDdcWwjZOKMi/QAz
u93vNAxX3FvqaRGdFwboFNjjs/5HBEOshRPX/ZEt3CQu/XP5IihMNS09NzPZW7id4w9oFcU2IhTR
UV9ywyjXDnGMD41QxotkEnDTeejtqO6lubVWZTxSp5Y+Zc0JfhiQo8iKVcYnBzlSvPVwx1QtCFgf
vadUThmvzYcaA5m+V8Vf1yUdFT/l3gP8h1hXfIJrl8v994WTWjVBTQ5UXDBGAHNDdl5mFdtCScEd
sLs9nAjNJ1BgTkINgNFmrn6hxbBQrcah8lGRwu+1cJIHf2ckf1hATfaw2uXkP2hmkapbCUMmPsnn
cG4HyVMaotwSqVK/XNTQt6iZPx1zqdzHLIJzqDF34WrUJIrDUBaSj54T5dbVkcOS+mnEK/RyAqtU
5wu/w3Dj1/4tjRJHFt7hVYtBciIJprLPSXb4mLCr1dMA/+QRC/WGk8gBhKBI7jFmiC8SgGy3SBBw
yDS9VNY8zjfFSF8eKpbVKGbJfOdqpT3OGZ96fgbdzo+a+hWTN4POdi/l1iFrKlKqsQN8hB+iUYAY
BDwDhwwcBtscWYe3xU25Jvnj5sY4NMom+eW3u3unP3KT1Cpb6d88++uVO1E1goVA+luSg+ILkili
tf3c8QVn/nuE0HMaTFzorqb7A2BW7A7MrYLfFGH0FKdRTAggqwquNYaGVNmxj3TzVT1HTfZ5wMVH
CW8rmCyy1LTPkUYYWMAvPNDJjPMmIMLQFUPejIBHH3RgdocoJ4YCwr0Iqi4e8YpMWgXhqetp5XAj
cZT1Sw8PHuPaj5VsevnPK+Vpo4jIWNSZUYBj1cSHBjnxtSv9Uq7oioJiwyKD+0jh+I/ziVVTacN6
LWfyrNfFnxC2KkwTCl9UjMEVepaYqxW08qf9ikCbOA+tavrT/FsaIqnXZjervCT95v3nq4++cavi
/mc0dHAVDOF++NAhf6WgcmpKcTFj3AUntgQdGx49NenjAppKioxKHQlwYxOnVUWKnEhN9JBsXgET
fhYSjUzQlSw4aDXnX2uOn1VjwVSRKGhOuwxrskZk4vS/IKNvVUeDgUZHYCPv1x+mpGki64aVvIJ+
CrrX2tMNpkYg+CzvC0uteTwpG1Dd5pK4+kFx/jvXNwycnNZXlcxRu7nLxAuW4y2UdbikkUSwmZbL
Sq58V6yR5DfyM32svJocI/gU8LWoWYTZ1GVkAAXypi2WMbFsudxj4yzP2p5I0FKL2vWPaZaNS8s1
XAvraDwnYeKv2hhq+IMuN27Z92PBVXp3nBmAJV/a8mKF9pWldpU8yBp5qMBZxOMXsm8e9TSR7pw2
ODBgTWid4n0B7V2tvndPNKHA4/DCm9V+kcN2rVOX7Na3VEaPwv8T4JfIUbNEIbG0cyVai8wMBIq0
4xigIKeH13hQTVa5kTdTBP3m/oZ12oj0fsrpqS2MYTeKFlbHSi6XGALh/LjsQfg9XlxWNkzq6Myq
H+zdFktlKrfpQKfclxFOcotfGoPZd8dxL57jduJIErchaODptQds8O5dFuCgolj1UreCKtB2pYh5
fZ/92+d7Y2G0a8ND1Ns6MF6peRIguPZemURRVRZiuGVso9GBHzBeDNAujNexG86fOybxoGE28fuF
/8Zx26TovQ4hlZrm3Wzx7U3tyD9OcYMHNK68LZ7IYQjU8OXpYR2wzhoOlNPcO4dmWd0Jm9YPcm/N
6BKCR12CcBLkzQheY0J+W5UgqzwJ9IZGOAwD/zljKrhBir0Uy/b/kp4oJVjh5SEvU4UdRSFXYuEi
woJZP8JyFxNT8l5b47lfmmvj7oVew3Hg8epZ7mnKzsknIKMBKmwQhDEC0nuArfTBXZe8cEE+wDa3
HpeYnw7u5zf9KJlfkBVG8+C7Xv36OD1Y+6kV6EyzUVT4rOKF4gfFEb3X4+Sstg8g2g5ZKDlB6Z5Z
kHX7Ag7chxOUrzILuVQt2mMpsx+YKt6erEq9amiYDU56HKYAVjVOk4YO46cZ3Xk8SsIr5fkZNfvX
rA23Px0hMw+TE+j+By1KXbbwAKGkeht8HBG5Imm0Ye/egSRyQUH6nWReSE8T+n9Qqif9nVOMzPhN
PFWIeuEh2L5tyteaGX18W5TWR3H5wZpwYk1EWXNi7Lj67iX1yW7Ejmi1R2gtjFGYXYSe9ArQxs2i
zRJHraTod4FsdShT4p98HP5rNTYFvCFCX6axtmvOtjqe9gONS7hNV5+OuVIoHaiocxvW6GO5l2f+
U3oxqel5qHm7gb4LLAk/H6axNvvymhVxDB1K/bDIwfpqJOWeZf6j91ImRgVjHEVJIGuUp5OKEsxS
Bl7V+gOMSV3YhFSnrQVnkpiaM0m4o9umqjnHsABNexShKG4ZI80VSZ6CQXT2Q62cGjckEtDFgN9C
o1Kyx/xHHdMbicyYVQGfou3jJ9SxhItaT10d5l56c/NC/5SOkhhWJuYEuxj8Hk23QV/a2ejBdF7L
h8o9zLZsXAP0TNuAWXJvg+yNQk3fXX8qH9ac69xlLyuwwdoE1wd0oQSTVp5LvsMTggGONxIxIP5F
SlBReac4vcPhVPlKGqx3zxtXRypmOTtv2PRIMlHdpiiD5jBhe8zgIVXCUP0iwaxyfejJDAqhyWmr
PWh1k9+EGn6Ffj+hAOAmQKPFjhQ//pWLtFRjZCzA/wUnWslZavU6mbIHL/psMR07IE0GhXto7Xjv
9lGUyXl+bOCuCiR84e8hCTvMISTg983lPq/nqFYOYtFQUjLJnMhqshs+IRTmPGi/Ssr+wOnNDUBB
XxsO/s3qbGaUxzBBmSEvYHUCLRy5f0TjFIK5PNwRmWySoYjAnmNn4TnkExRoct+t21pvRs75GRwd
2fYruHhLqVcgmc3As7JTp52zQ449q4y5/uGK0uEmwIbpA0Q0SFQyt4RQ27HfetW3Iwgd8AgjjGfZ
q7RwEmavwIRjBkJAMy7dn4fVACr7KTeOhNLVuAa0nzwQIlsTj2aFnWieZRw8O51VrsCivx3URokL
unJSRERYTq6AitPAd7OtAjfkTeeDNjE43RSUt7j7QyR4MLAEnc79gTFDJmTlfEADWGqK63ormJWu
c1E8js6uxgwl+0FC6ti5fPtRjv58bRtYF1NvLqGgLBUfvfMtXxERSFDZt2zuSpI1ieChDLf2UP2I
Vmou/NW3U2PoL47dF1vagmSG29GnSOfNHsHymo1gYVFz762bVogY/5bIKneaoLNFPpz2kapMuTsL
kjYPT4KF4Rmg2wIZL9idxH+yaEWI1YjPWtOMEI1M3DIjFPmJg12ozZ7g8Hn6/v5giGJKguiYMZ94
Y8liTGvJKmCmqQYADClSTh5E0YTXA+++qnK026mp5v/KMO2CGcDpS2d29U4k3Dvu4Lcl9NJoirLP
Qj/IlUL1Zc3vuPWQVR6NaVIYRnoK8E3jSvhXbEPxLsGHONR/WzUYUB2UuKs9AmJIkkNOhzT6jf+L
pCZsrkm10On8fDwzTu9UzyWv0mfFAGxsbpW1hPYewHMV94M0LyhjA4gamg+zmGU6tNvBhX39bBFY
VWG/xOcqg1chfDWKNyAA93qMLpVcFJ4yKKtBbQ5enlaqWABXG4Gpqilli4tKktaxUW/1wmTKgl0U
wEoMot5X4tha5ZeC44M8m0xum26luJn4o2xN8omXEOk8rkGvRUWAMY9XeMjoT3ng7qapnhBL5jsd
1yBsZeWIEsExdEm1W4ddXusrbwlGcw9L0Ix/VZ3duzNtjwMtQP8JgusnDpnnnTOSfdFkYVgWCVuH
G9dE2zUAmxAs6vXEyQG/bg0TMtkjda5x0TExck7cO3zB1rl68lvllsHXPyaFaQt0J3TDz96ZEi07
1TkjdE45aeWXyenZEX0e9FUHYxcSOtGLki0xDu0wIiraFiN0hc5qwLYs6JJDi5QxGDecf+q8i6ef
jR10e3uIJ25CDp1Bdmycz2MIdYeEX+BAydL4KkEI2MRSMYhLZO0nw7zgnYWckHPg4YWeVo97qb3f
YpwJdjjMJN/k3J7Vw6PIQ525wPAYIMmug+HJMMk4x7vVo6k1UrhIf4f+NbvrTrUmvGoRBq4AF68q
0GqfDOWBgjZh/AZ+xpZlmOglikJvGqI0g6YN/g6DxhKjt/H5xZtUxP3QeEYgiWZTbikAHTdqLEFu
nDDbxqGw7UJ7Htv1IuGlkF2gwh5IUGkoRJmSGcfDVO2AjFMfb1oxlc4xosp+Vo3nnv5B89aWMPEr
bZ8jF/sL7UX/5QVLYoGKwQZPXtJoot66QISJfJwGC+2phaOrWMMrOPbTD+Ypw0Lh/QgCuAWd4TUV
yY834kJZZxwYevC5XfUEIBNIsJ1mba8Mmo+WrgUNN1PeYP0zbR203+icbdqn07SEGjWUCQweRLVH
9WbZoKiw/14wb5EMSdx4gFcXSuYUA4eEkadWUHxkEkH/8CHDd2sQzm+FgyD3HGNSJ8SqKyVhGaSG
itEMAWiwVMM0MykTo7RZ5lEMQy35ipqPSoR7jJJPdMo9qNK7Nwbirj4zigQ+QdxlPS1CPL4ep9Zg
GY2acY25l3gSUd/dsIFdQgDOb0fY4RGaUO/G6UOgjYc91CEkCp0+l4zGCO5Yni881gEfQXsYwdrz
IFjPvRX5aIVP2l8r5msKnWOgiH+3Y5n5XpzHRzn/tjcLn9KhHmQudzoWUPeP0SSoIsmwa5/5xnFe
KmBF53JBQkMv620ub6mUOKjRhnp6pyledLlCBDfzm2ETZMjKpZaIQo2xtl38Up7jxFRtmJqOZyYC
8xeJe8RWpIWjSkPMrtKuTUInLQYS1TmUKpdqtgYYJxdZC809/bvqlzdtu0fTxrHYdtwZpat/Z5V3
SDKorgwOfbpt5nPi1FLslBrbeAX4K+LUdfdyhlShOzOBT3kUEJE5g9g5/DYtHENQ6+xB3bKTRg+Q
ybDo6C4yqrIEX2SEsAQnD3ZiI5RQgmuAW6ERScXqn4FJZ9ycXijAXVONnaH7aauIvxa+I7hGrrXT
5YoK6KLxzX7BTfP6vmgV58iALTtcthLg4IuFqrR/KU07prTSsXILJAXk5Msym2Q/67vB/sF8fxN/
lrRJaZe5hiVqjkgsWmFsqwPWvQk/YT2sxAX+IUEsYzZU1Zn88CtbJY0JfovvXDtYBJyL7O3KYCEy
DIo+HCkKR16ghcZS4LjnB4Z+3sKye31psauNDcqtCDhOzhQwNcngwKwtuTYbnCy12DU354R0cQLa
n6hbwwqI95qdl4aRLCX44a+mbHzXk3L/IGXpIVIlBBd3WG1U4VuTqnNatjHUECb9lENUr/W2LcoP
5ODHscPHvz2+jcrLNAuBQxaIrM1Qre/MJ5bJW/csKFKgU5yceJeiP8kvk/tKrYzh/DxdMUoXEMAd
AIUfb+fBrSweV82uXaTL8E8LuxaJLADQ6tWQQgLSqKyF/obo0B+GJ9w+sd1RG+aQ8WoKaI/8bcE3
hckkqRdipKCaDUHsqdlLNuIZWoBzVPxIsLrQQf+jYDgz9CQMfMZ37Rt6G5ztyx/eRnMFY7W8sYAO
+u+RFGNmjdHNBuz5E1iYVZ/BQPztA4ZBrxY83kiwW0zLDqsI6NsW8LI4XGuvex/O40mOtERmlheU
fGdu77psOxDx/TxCxuSE42K0PUQyvkdA9hqDWzRk0SEo5zHnEnbXAY2GHi7kpaAJlgoVqlX72mHv
XIpJ4EI1QhxB8TkI1AwmrgYHXcBh6CZams9n1Gbjhpxe6/NjVVzBVvU0cdzrBLVTcsNEKPMpI8+U
KkpvReD4UJOo3iDGrjXoCpD5e2q1/CXisM8gtqc3YUjz+ZEYrCJQlPbqTpct6I8D38cMDK8lX/LL
WzozOflk43gTtxGJrpEHSYvcj9yUpdYS8v+ZW/BIov2/fYiStGqBv+gVGC5sOOuYswAU2Ttv+PMx
RTPTCcu1kgTVeRJeWhYMDgY9CuplU7/MCXjLmzpklWO5V+Kpo9eC1rg9IUBrn5sfeZ/aDmVwvK2j
dZDytA0JAJMKsIv3GN8aosEFv6uGpcFYdusvJmAwAWvv9Vf3LlSST7ZVk5A7l+vk2H9yumLH2/E1
YgXFUXpGx10slbOAOU7allxiRf3foCeP82/SbTO+x9m5bvAXaiwhCXPFIwoqFi7L95zVbFK6X4Fp
g7Zoz45simnFLSz27RjdGQ2Zd1gtcF8MFKZquAfEIXLYSu2uyQ9GfobxlAxpXwrz1BbMB5ew5Oe5
Adt/vSk8fAt9WOU7lY85aColFZkQWQgYka9JsHTJy1ZaroX2PBfT0auSua7CBX7lW8HvVvLa3Xgo
JAqHJgpiqZ+s6U11M7w30bYhknCI7oDMj3TG79in14PzLhQDovZqanQsNJoKBDpVQcrbXafNAQdr
rerOoRfVe243Tx6CPs82dusnW21JPsdK0OWQhWYj1xEBUKJ62YswPJ+TzOKEhvHETi6OazYzPvdX
aVNY4UW13YQEmp8boOR/FJn42WGvbidFiPrCnMrcICnj/i4GTw5TJc0vUsZq9YC+wOYoapxE4fyn
MiWWCI4Y8cDQ0ILUWNUZl1n322i/d1jfBXlqmCd6quqE0FSpfc2rr2wLgIZTHyBu/vnnuGCmR4hM
203LgkF0ZkV2xDgE74FyaLGxaSlKtgDeQ/rwk1wf6MwDFmVU8HfPZHHccqP4x9nu0ufYkiiYGxC/
SCJY+JxW1ETTzPK5cQQ2vHBjhZLjxpyxWZFPdQ0lCocKp84r/hiUDXJqIQ1arBdayw+wqdsm3QoR
lN8kPOEq/UU7Z3K+E4U240CHkxCr68RM6uIJ1kT5InHpBZwwrGBxBWpknChHvXFItDOVMNYs+eHq
m98bRyqvWcbzyc3ncYby1UJOAToHKGA0Qn48iCrcJChmdimfVIRwsq9Tc77fXJ/0eBmdKT8pl2DI
3lK3h62xIWMPA8ibOxQg2nYqtrxUrkANkdlDZiKm/hTZWAzAKTbSMknG5ssdqve064KtvEXiTz6I
EINmb08nB1BQM+CNg+jRnfzSSQ2q+2u65vEtHkqsS8VRUiH3xUDGOSPfG32m3oSISc02aT5kKPeP
rly4u+v4tZ/CPC0pDbGvEzLeDY+XJoxFGcM2SeObkZopCNRMmReZA2d/myPgfzoPMzlJ48DMbLIh
QbfvivuvpRoJ7i3TZvEqSQpZVCAGGTZDFGOKPC4hidKCi7N+e4MtDq+AbSLyzxI8mk+dkJ75280j
KQ+1Cwfxb3IXS6dQRNtttv0X3ddCUgDdP8R7tTJrBLyGjXrTE5w7bek/T8yBX9kWTETU9CD3bs1B
eLQSeL9GBMZwYfMQWnqSKVFqJCpnQL5ecK72D7tJ2xwiT0TBzF2QZQPoiAF0sDRWdGT19Bc7mmWi
zXtHoCiZaB/pN4KP1pS+h5NExkAphYcC+cJNMWx+H0wNP3J9mF53Bc/Z/4NG9epU3FmGRXbvDqIX
C3EURfHpCM8VUDHepsDXaQgtVSflR9NvtAlWRFHiryNCeJ9zo4GT5GnuPL3mvtxFk8gQ7VsjTQ/o
+I4ibEcdzl4c8wWN7zUNTNnoAZopmXG9cDHPs5HchuDfvrCSypdFMpniYUWHAWPZ4bv4Vs3SjmA4
MuM8Roe7BwW6ZhcoPypKwADY1DWyahf8eUjADNHupLMSmielGlZtsBCPyl0cEsVeaQQggKxLC2Qd
wVtGgGh8JEa3akRu3yumUGxc9XuURaPEXVMM+VuBi8hDGihiz1Nd4l0w9zrc5JW271zBLEbE1Gmc
ImOLn/yTngvwAaBc7bBBAKLLoYrsvhPx3Z+YV7HpGlwdOp/VscHuumhkrTeZBBF/pDheXa8MzHho
907YrWQdhBnaVZiLAPBI63+924ovQ8UH7/sVG9Jq8qzhOAGq8HW4eRoeNADEMm95jNW3OIRBbKTD
iUUEd7H0gaMur72JqRB1IXDvh6sRuA9aFh/qsb9PzmKsWBuMe9/enNRz97w6D/6hwSGVUMMch+aZ
OmjObzQJgMuFiYvHYFVHTwPy2pB+ez0mUVZz0TupREXdUK8FGrOH+GZpE7whkj4irlntG0fLsj89
oS0/AWZPflVx2pcvJ4fp5xikQiwWbl02xkfpAuBey8QxSepUyBKbs0TupFKZVAY2hNNwtb1EfMw8
4q4M4yvsOdJw3VbcIWWsuw9dv2QvnVtn8AD1Opi/FQ6Mjf8bWXyQrZ30KuTwzA38YsCfORQsgBdm
Bk5LlzkRHTU4P2QXIoowTTn2rkVb7YyV3F3DVvqDKKub05qBOwzC/PfsU4FtkW/gKI+C8tX2elHA
EvbN2J5zlP1Ra39U2AqokwpRgflpkuPW+fqQnoHjQF5moYtfcgHslAVPESee56nLkHs6msQxA5mE
+eucliFlNgOOL9x+/d8e22beU01/syfeVpVpQB0BQTZx4T3uSnyEn39iJptXz9vw4InlFO+vmInA
WXK2FhcVzvgkyt96BNCHXrLO95fglOzz6EG/nF6e554LJppNVs0NNbQM3JREEb/syzHsHrHj6i8o
P79tuwvt0/MshBASMwvQMpo4MCERshInXsy98yjjZhsr18T1/TJKW12v/ZuRqEyPjLY93cRrQS7i
lfTxDTzkUkFWAN02/uRxBbsG+Cc9aUvEH/by9Jetwgd6TXkViDtfE1r+SOMBMgpp/09gNemH4KUp
Fc+mqmAftc1Sd8GQlK5Q/dy1ACXZe5fDF22GeZz7LzQzzOdSyNCQvUHvYGUooG05j6Kx5H9bLrdC
JKQfeRWTXMaNDRWyYMiVXni30K2qJsX2YuStWUfvh8rVRQeOLTgFR0M/msrbdOCx3RyaVmSksZvg
GdNUTd1ZgKkr8H7eEy8u3ksh2JTjLFqjsxNRGei0a9ly616Css1JS6pvu50gU1ZeSAdhztz1RQ3b
Rx7xtoms8v5WhpuReAgWn0Kwl2QhTm+Cxum8BdspqlxKw8lo5r9LtDp9HubcYZEIzsQbwFtE5I1K
UEKi56bEuu7xjcrPPevKlpS2tHSqvK2yVr3y6lq4DR2YQnGvqly7JtDDuNLEMjEmcl6MWBI1apAM
th41T4Asw6DJUT8FLips46rAubQ1r79RV4ObFleY6f0+R7of6YN6+PL0UJHWI6yaum5ipYoTmYcZ
xGfLA3kKrsjSPa0mbco4RsGLUsjKGBz9IvhPVcL8e8XM/7zPA91KIvIq61RCpaqebuI61KeWDnal
dN7Bc9x+wUnaaVo9oTEk16WDWdM72Qvo6Y86kV/ADxBDs/Pwr019hmlZfijANkwonMOD9YX3G82/
wfy1adh924Cq2AC1zSd24jIgst3q8sIPS3PdLWdzB+7V7cBcOy882bKeVC2V3PJhDhCRuiUU0ZBH
48JsqViwDlnwpHKD/ATGSLknvnaXB9PvWaR9YeykJTCLecZE1r6y3q8XsN8EyMM6R2wrhyFSAPg0
+LEj0TgsfEzYgMuKwKVw+MWTtE9etMWvg60kx6CundYvaSAsX65ISa96mn6v/vAs0fa9ti6f7iMU
S+RRZ1hw9nQhQSTlmCHjieghsipSQNJdIU+TZv2n2XF8pnNySc89yIbTxvw8Bk1XVCerF4R2OlFU
D6s77d4E5GxtzljLPkm+rRW9MtF9pqwjSxBLaHpeAuLcHSqR6jEDZujXVyhzbk42xGRHKorlqX0F
crqpT4nwy0lXfbBlM7sVNLRjbORJZFjFcGyEeGpxz6DNWJtXSFE0JP64eNy6sgRpWI7k8TSwR/A/
WL9lemMbJIVDrG5hRz7bJT/4yKB3/BZ9fwln6GeYKuu66iH5GA1JQI6LcpNzYu2EFuw8w0QNk2lo
eC0FhwO7JshA60MgesOuoipEoUUj7F5fmNXY6DGEfoq2TFfAGcUVcIv2hTOemv36gCVwnDoKL0HF
r7bUJqOdCXLi6VebW/onCc8bYs+E91c7Ao/NrF5sIAyL+yKyQFPcwUD1Yo95dqCLJgBKXWgNtTo4
LzJy4g4tTXAdZsUpucJ895fpzcGQ2M9YKxlo4hKz7t2GuYrVK0mIvAmF28sA7d3bRNRq4n81M9rp
K+qaO18HMqgQTcr9wvATP3kS/nSy75dUBz29BZYmOEjwCzXtqwY9U1qjd/xtQs9Nyc5JHhgJp7sh
pVVtNetzbzPw4xq/+Edu3RJX47oH6DAs6tulTJ8sBwabpQ6ffoh0BakTGWaoClZed3QfL7q9qDas
JdlEC/FcWsdRWHyF32IMzB2V+TYlgfqZwWzFaZe5uSNKQoQJUH4tjztu0SqpSCHud84S+JYIvBCt
9a+YQDSXCAZZpRuDBcFWys2j7p+ZFCJOMUNBW3DablZ6I0yvYx9whpWjGG11uXNolrydZQ+eH7WT
3kEZxmQnxmvKws6PfpJKP0zmfF9Sb2tJPYJaFicotouhTxJqCQ/wcDVOi6wotGDl3cP+sX1o5FKX
pBf6U/Ij5dpIMN9+24ZwWpwVLkfjSU+x+BkrXlo5u+HH8gSQhsifnD+HyuxRAQEL30TBu/HxfTjf
YNhPKG183G5XApRNUty8urJG/5FCZ4hqI9SLXYCIn8LS9ujRB9OJ1/YmObX/uYvz2DKTVuz72ZGg
BVkvXiYFegH+Fu2PMpoSGsiP29IRT1PdkLn1BgGw767bbel7NJ387osY5WMODOAu7oEvYscBWFfm
DZ0PMA5aASHHdhOA8Go76JU5y5TVppuckMRwpRxJ06s4SXf2Mr5SSQPbg+avccQTGvq4/T1GbCuA
koiBPm0psyC60OlJ8ZL13VXF3/OpTqO/zzWg1Y5mvui00xORwCBY85BJ5W/cbOAtAx+owfN4Jo9Z
nnciswrPp8MmFRbRiTxgtrEQbJ6ZNoJR5Fdwhs9rtho7u5VUp6MVrBzqmjbUPCnsUpeQ6eZwjmm7
27w/YsBgLi9WMQd6Bw2srO4HNfI8y78r2G6eGJK4oRQAT3n4EQJQfzYK+wQlWuFiAuisCVbZ/rfI
ruTxLSXOxBFW3WVTnUGWRD2U4340lhp5YSmpj5/rqBuFTkKgtPiv6qs0s/UrcC6PYeSeWnV5bnHj
pTHVEXX8e+COzFwm2l2rAD3ycK5j20EMhlBdcaNAi01FfbdxbVE3gaKJzCR7QedwNG+j8jhO7TeP
sE8d3afsYuAuhfqRWz3oEa2pkYDqULFu/s7uR2KV4Br5RtfbTAgBxs0DYvM7MDIovQGO0fRXK61I
zgyuy6vS62SjRRpVI52bLpXyclJLG6y0MackTK+/0Y/iP695cIR0d+MjCEmPQDY/Dyp7oj0OOK8P
anDNUAajujJocp5UBrKTD8I+WW7Ay6KaJq0A+inLpHp1TCkghN/hexi4FnA1b1eLGyGyol61VNY4
QDOWquSHGzO+MbKcmqW/cfyiqQOK/ctsuHRTCWd6MOuWxJP+Fu3GV8NzyZCsjAW6b0ywpckxPblj
L8B/upd15FMSsQ5xqdD/F6w1cpDFG7NJVUrFcVu/uIAgL1TCtQ9ELGQxApoRHXK8REXyh//qROZi
FPYbuksCM68J3hj6nuhUYpZXS3jzT62MIl5j2oxhWZLsmygtjtMZZUfBZpzuhG5lPa9ZGLMgT9yR
IEwKXNiIh1cTnia8EhaIaU6BdLPc49yw7gnpgLwWbtktyye3o3+YxFx9IIG2Xn2uOmdrpQXIDFmO
Cit3RaTC8urnNdMvw+ikgDbIlOrGZKBmjf9xkWhGc9ubUYkN1BZpKB6ICDT0hOJ2fTiUmaUSMr3r
LbRe/ArnjI+FfPiO0f5flS+He+mWrIV6vboAd8rQci7dtKHrIr0UgwQSyrWYbZUc66eAm+cVJpB8
0yhPaUz98ms+4DKeDGlemYzykMI3ArpQeDbJR6M4u9M2tKjEWx2tUQxuUSTchOuP6H74iNPsgPrc
AnH6YlCVWU73zIzG8lx/saIYiZduKLzOSJraEf2f988ixzgzDz8wYMIuebEmgsygFSgNvCxW15Ur
m9nznolNEUrlLLDC4MBJAcSBNGGHvFlwyLENq+bk6Ca2yFW8RapCE8jtG/E1r+u2VZBtJZuq7Dy0
NQMBtmn9lqoHCmTggXgWUFEs2AeG5sFTO19/uSbPh8Pww9Bjamum+W0iUnrOZCkYBZfFNQfpXsL0
eYkbuWOfaH2LU0sTcvYDnMWrjhB898PzhsdykzIo3YmPijXPkBaXmCy4CHPNIZt+kkiJqOaf6YyU
JxvvMLFGjclGvZgHRgSEVy16i4Zcyx+9wOutbEfxIiuvh0Ig0zt7FCR+hLN9zIB+81SWSLKLvCcH
dzEQjvO9zba9xChZN/b487LTs5XwYWjWDv/uqJ9ErhB4mmZldsiF1TiL0/xuOFF7KmwGxdfp8RZS
VSgNHXSwCS81urG55Ewk23tFI8HS2qDuLkYulxxVs32RNwt3L+141Vac9W+WsE5954UWa6WB0Yx5
zIlvFpI07HqP3p5deCj2gJHVid2EKQHfqNUgxekwCSVhzB+WdLvlDjVJrFTmCv+1oEMqanacTi0V
1T8BsjboPPNC4/QEjbo0EmWla92CHcyeJIfgrmH/MNpZmG9E7IHJpYItwp1ykwHlghOizv/pC0xJ
36nUcjFncpVUZKdeMh8A10m4ejYu9FiUIY1bd4HfZKY1B3A9SLgkUGP1Pg0eZrACF5lrx+erfCLE
KBPd7UCrAaMazk1w/DsDTvk3A6q0gB4dvw8hkaJRWrjG7xDPh9ZiktkZb4BhT7kde6GBQHRzr2co
kDKGPjOE3apltCcZXtpX13HWH00VrozZl8oXCn6riFgmX+QGIY/s1tjFxp1vqmuZf9987lf8yW1N
dtJ+i3IsZ7bXGitrlZyoF0X7ld7slxl0dBb++hNismRkUzv/+SXc1snoos6evPZ+kVel/MbrD5Vb
i9hi98YAhU7xN2S3J+SYFoZ6BsLg3z1SdlpQlY+/L/f+bZBUiXmS/fRs7BE9/FSV4TFLRnfTRLKD
b9Q4dQx9Rfj9ppo+NK0UJBhEiJj6ta0rMJ+aCYANi1MalPdp9wxK2V9F4505N9+EGxkCfQ0BcXAk
yiV3wVeh+SVaT80Zpcy0WbqzV3OhdkCjSuYfw4SeiHqVpmgIPmVtSTkLffLN3oLSYXZhFpPLEL2K
49Tyaib7dBU4KU/orxO+kjwi4rwhjkf8BqYT4953u0qVmMhuPjc3dTo6B7dKOQrW5uiWGEEKNmoK
ARtc5lFsUan0RnIMBzhxoubzxQ61GrfgyrkufER5EUEo3GFqaMRc7yoPfAjlOmW8E8+jx5wrKlO4
1pmAbxtTs173L2Cnu4LIaRBx4p/PM87QpT9gMtZ4nvCPBXqzLYHtZryEA5ZnYLqAeYuI7JchVskn
TVPyNzJxF/Z0agwHp/Rar55EebSfo2Pctv+iPXvbzoS7gZ9m5u3fzrxRkxvoCcgy4FebcYT6gkC8
I/e8UoWw0HVECdIZSxuGbBOYgt3FyiC/Vv51XmsPZdOqNzkFXXiZKY/m8Dw6HLih3KjKBZg7NEPd
SmHX7bVFR7dyNehcm7YwlRJWqZuAa28HKw2RpwY/dSSD1xbMfmWbCVKSNGm42yWDHfVasM9rmkv5
pazxBlNL1a/tpYP1EnON0NDi33ySRrO1mbxBcdkU7jvUQo4u7iN2QlII5s0EOo4AOcHi/0Yua1Xc
lpw5vFzaxc+Iy4UvOPumURSd1DZnRptGn7l8xMGivAzFkteGgyOkYtOtoq69AdClN4Jsggl02p1P
y5uzM5CoCPBBM6bbZwLytuWsAwQZXcRGYEsE2jkJnXFI5n1okLFdnDxwoOHhyFAnk182wCwrJUn4
UixhREHVKmFgMBavrI/SskrLczVTdx8HAQe9fkQHxkN6+RzlsTIExRNDV0cn6ksGlUJ43oj9eWA/
2Xhp7JV93nWuzuCQ7T259h6KXwFnaslY0kLupvqENXG5p+Gp6jjk0yuOZDUMEYFfmMpCLP3n+QOS
07hGBfyeAiiUd8rRiaZlPbE1ZklX/VzMg4FkAaaO5bd3SQFvehrMlxzWLDVATpBjAsZdQdV1FfeZ
v4ZWmsfaXyGj0fTGgxSyIaBzX1UqnWWkBP7k0Lyw2iXXTvalQThW0LwmoO9jr5Q53UxdqnxoUX8h
VZ/HL+lB3oOM8A3/MkuDeW48QgT+ECcF4GwKIE2DN0Ii5+ZFTlyVIDCiOdxfgrJfvHR4e606ssx9
9Eu1GDPw3riXenaHXlSSMHKJT5n49NXQCdof8TQ4ErKO5TEbFPJHA3/dMdXPQ94qJOJ/hGioPBI0
CnhgKed01AhtY8Cju2j7eR2aTLyDVDQVx0feesi6k7Mi/t8T/fcCm4FiOvrEG7aRxfevjmZ+lpId
AOlQVj9o8ZKsYSpONsVtY6XV+DTCV8hBDHRYWjsSClzFFxwjyxoKhVt/hyAINX7gItqzZizT85hY
rOTKbqWL11j7ejeEG/Xi6H3MsjOKOn+2YkGJM8OP+ASgXA8/zkGmB0bLBw2QRatu2nh4ej8MsCJl
R+X82JtJ8ePuZszv0PIRDvEH3pzJCSIZaZuTFJzBV17elJ39TN4/vZLm8RvMVcICDU1He8vc5W4N
QMX+5Q4eFTHhuTsVxDgkhDhV56hS5k0Bfs/XLc42k2XKSglHrEDjYo/kiUY9YOk+9vBcxXQlaj4Y
plimn/d/l0iTcym4yOoksrDgp7c95Uujv0xj1DUjvA2+SgslLAWA+iFJJ5d+88YoQEB7d7byJi8b
ppo2vxeLtwgTaIrjjtIq6y1Tchk11/BS3Evxh2MAToFMqhJJ/9/nhODZcoEYRs0qpxzMyoxVS8Pr
CyCC4mAPsw4ZzFNuw0fLL2rPIz+VuaHGWgDZOC0QcDYAhNTJx/YVMfVX9SJstlSlQIZBFCGHW+iM
UPixHbpPwuM1jRnWG+TfiG9PaUPJCS1lvG3uQnvsdxDnuIOdk4OeGAMWMaKG1nzD5rchu1A1Pycl
nQKJ2EVBUwfGvxejEw9UkSvN7spdEtk30t5AfWRewwHZ28VXOQkzLS1o81anHPFyTX41chCcQmwY
HjLXURVRWFPOkxxrEQ01DW/+dy9tjZ9/1m+pOOpv5nSIsbiekGWBoWzNtnsCp9YoO1UE2JOtRBS3
BTNGERXiuEZf60bb6UOq89n5Bj3eR3yqbxGyKpYZ4Ts6VgM8khUs+Q7Ah+uqq+zHN/tQDvPUJjqH
zBR2WYJ7dnmVYZ+KlWRVk0EivrWDvm3pyVBf+BA/C53xrbYmcvhQxCjAtPS4d3aFPiRm6BWRcyDa
ENpuKIDqF7mzRQ5K4S8XQ0C7dS51RkODl+dI49fvqJwrWN7NkSa1no2eowTZjsqpp9OrwKki42b/
Eq3jrn/qAl7rCKFeeSOv/Mcan+6YsYbHB3zIcGdKdLPJ++s3NoDrYUg920Y0lwYa0TkKVEfBQk9L
t4ip5vKaQj2ZhOWm3yEq0mRFANd5/rVa6faJcmQ4+rmF921+l/9W0ESslyolPfwEroFpDMUK9/pd
DG17L1iCdHBsiDYH+DXauaPvqSUNHXqAqkX9/Pi75Bu0hezeozGNKVFlFv2y2+P7fNitJTkTTp7n
Mefks7KdqUgrWMSMALkwi4c5OShVGlHYPt94QNdmBSf8dov/iBPFhPn047ZibTO1u4Ma2wUJ2tMF
eBzS27EhETbb9yPUrLKol1wRp8QWyxkMqXTWtXYlorT8hWtSsDgKytjCmSldnpUTtpKkNrtG+3Dx
hEhLcofmhM5gDMEw1x3uvTheLfaEV83Yv35/bnpMZN4ryiIw+6SSKShHol415gLf9o3jjpNf+5k5
zRuWVlNAv9/witSjWsToV3ybtWnbusjv44iDQ5naUaHrRESU/7UXeq50bxE2z7ihp9rARaYtBaMR
mA/No1I1/QZCrtKrV1GIv1JXbHi8/Xc34OYfPlw/sQyvZGMYpWFImPAZcN9WcqyLYXUSjhHM6JTu
LYBPWw0aL2eZdkv56hVTT3DxktqlolfOaUAPtRj4unoe7KsVMOF6Y1R9RON4Cx+VIR+c6866ni+B
Hw9fglGcWOOFkdKXOgDUR0pHcP/EswLz7hnrrPjpJX53hJTMZYkNRyl2gD0yhz/6W+5WNX7n8RgK
L6+5LIlCQVEEtvJWGQ/Rt0UrkPd+Val0FX/ZOlQZTD7JJ+gMRpc73P9lEkGMMnxlpqANm0FYRlxz
1Pr24zqIkYUOc88BQswSOvwjlbuSZ+fSnDjF+Qyq/X18hGapGF/bxc8P72oOodZl/cL8CrKcKLZY
PcEM0HMkZ0nhUUfV+Cm6kpG4xhJHtcGZfwPkr3EEeaRiYSmATS3cQE1SzhYt09nfj9fRa/MJa/YB
EWGJfZTuIPSWzg2WZifVo6xynQDF8oFMowPjMkL61k2lGC/UlTmM3XvBbrd7VRcNsw47EBxkbgUw
qmDdnRrRE5Xk8S2xd4y2JOc04d+3B9ksIQCrU3fpBpD3T3A1X/lbC65i0rrJ1U8XFZpGzllK8VMn
BqZtmd0GRD5I93/vHdKjntjNikyIl7vYei79NpzHQUYj/g+FR9Rj4hJNE+zSplIBojMv0uJQIhPo
TqicbNr3Wbd/rN5JVw2opi0XUdx9c9+/8BO3Txs9rppX01vs044wIsCmsxsvDm7c4oJmIMVHSuwv
ZanHR3kRimTBCFtIoN32gew7po0W6ySWohEYcvtjetCZ7VVTVR+YiaO3uJ6R/G7j7sy7S4X7jfAr
3c3kCGM9nX66bq8E9alLkbBgz/FhmifLG1OqlrvYOG12jtdDMmhUQk5Fd81wP2nmTj6bhvP0WCUh
olOM5yW2+TIcU8owLhMCLCGz/oxf98er6/iXQZcFQSt+mtuiyKO44LgrcbttZ9vxWJShns9ihFov
caOocu4AfA8qZwRelRHBIV017GAcAjCApWcTJPVVqMkydyNqLUBihQTltDz8ziNO7o7Mlh0u1Tx5
d/fRWe9bV4pHvzt/iDEEnqvtGRfYihI7JbJ3qSq7+j1UTg/8sOntRM+4eBvuXtTWT6GCsQfnqiGR
M8wuBjhZSSS1xH5poZtVd0Xd8KXfGxRMdXHoT3fRUzK4hiOKFUbwrZ7kz/4CQYJ4yov27JLFEtBO
vqHA5dus+RrlpcZZ1m5oLScEYMuffZrlfy+P8AXFODdgp+k1uIMwMA3Yf1eQR8Xd3QYFBW15RIcy
V9HAndtmUl9i0OQcnVgSAS0nA1/OPhsT24fQkLrwjXI3iFwHbqxhlRjqksCz0wiiCpEzyHdwBbIS
nr/Ipp91ZWSU7BvlpCaFxJg2fgcfxgBNY8ee3vIsDy1Tq2k+F2jhy00Dg3EDdRbCbdsJyZf3cNbl
kfH1lBh8zi4L6Lo6QOo5iQto7CsQOEcES9GRjMI22itXFLjXFwIZTwN48T+egmiHRyKveUB9fVXD
6ujmYbV1h7L3BxUThT1Kz314zPHEdaHBdL3JnJQ0UQ0azaN5MVTO/sSBVX4ktuKG5zLPHm3VKepm
nrkcEWs2J0SPxKcpTuIsuoefrEt8AyQE3sGIy9z5VL/74gV4bnzQE0EGCxxX3q2EpOjl3PVk1wCS
DT2yuz81hdX1slB5lZDmfv9jCE+YpSKkKZTUu5k7bbKsMgg/V5Hx+yJuhD/WjxL5xDMteDoxrowo
COJT/5/vhGzCKlKyZmwLF6N1K1A3LEY327e1g2Biod+xr0kYvprMLdh9xK0sWHH5+opjNaA3s/aa
FcZHvjh+udtHqbifeurZzv+xcZV7fYuiIMI/0hPhOu9mlsWfOkGx0dJVdlF29TP+9y6GFoa9rJah
Buk6uv7tLHK6me7qhyHcZF5XOqDdkxyl8ijYHNBwaat5u+NTPoTV4QSKUNj3vxJO0l2t/P1gjkh+
YjtIorXLySXhjASKfEUzs8IcMgnZ4wgQxzhg4w6TC1Acj8La02fczAxTimhYDi1yOr0rYZywOGKO
j+klTr3JxcEz3i4QnL3NEX3oq15cmMO50XODCFpz91G02wfb4fkbm+itKf97WJB0vwUU3+hwHl3A
Y2Janka9rnX1PPHosckIda4UJla4dCh4o0DkFVeAv4U+AEdIyw29Q9benCM72d9Aegq2p1h1V8Hv
WnVv+kUGji+H3dPyG82TvjTPjgPoLg3Q4ayRWw8NDBDHT8woZBWpuiFgl+NlE7uXp8QUp91jvCoM
ZMr7pzU0BatmWB4Tl7LW/NRHfUE8IFAmlNpx6cNhb1Ur3BkeUIWb+BWNDjHF5hGrq4Wt1LvPs6Iq
Re4Lh8rOlAwAF5OHlk3w1qbPhq89BA6Aw05QDIrv2M/7/P1sX36uTtsiK205qnOowpyCDLPz3wUn
QMxjTmbJJhrFxOhpHfl6vAvzllH7WJiJidBH9nFNKOKMfFUosNqfMB7A/nfoweUO9gZn9sttIARY
5z3LZx1h4lFUqTwvHRN9ptbG3NUbOHA+UPCck91BBVLVDkhgQ3f3DaOY4DB/qEVt91IvLVZmt3UO
Szx5WH3sNbVLyOflycH3Es0m/ircfWy+FX+K/l719Ov0LBGt94xmrNZJlCjTgQerjcz4OCpUvJdp
0z9Z92QsGxECJa6DE47iRR9hrKwhgQssHRgM3Qrqm0i87W2akleJ9ye4gArYMpmebSwOLMaGDEAB
wZ1Don9hGjauzqOpWe1kzTJz/2RFuMoxOp4f2S0rZ8nikvp3RiUUWOjifwqvSrFpU15n9fw/Vo7S
KiRSa9qD3Ngv4yVnxWjjh6bMZCpFODwkwSyvZ5EayumuOwOd32o9GslWkU112Nb9s2dSD+sEVKXO
Xg9nJBYNVXL9du/jL75cf6z3FrTEpPCnnckxTngFRtLPrCAygOSRqNcmcHA9Sl92XVbwGBcBAZA6
x3+WH87NJAQFvUYXISt0qCOoJNFP51Pv/gqkqjW0aWt6mCnxUC0BWv1tHAs978EQjkkcvSeqDVQT
M8hs4dGe83Ewsk7vH4C1makYM0NsDOWfYwflUs67py1Rw4ufA/V9E0ek++m1FtTmbwxAgx54siUI
T/uks7qa1XCzq8PK4m8q2gCVhHBekoGETN0zxM8osHnmy29eR6cuLWpDSYJ8TbF80BG032U8v2xk
AtiaezoEb3QdAIe8BjMxxESPyG/1t8/A5grhCD2O6+GfByL0oJ+uPrqopUx54n1e86OWOLUjeQuO
Gf9Uq7d68zlGiJd6TWc4JChc4tOAQw4uaD51P2J/UTVLl6LfVJYMrgR1eA9X3sa3ixyBfeLUn/eh
MD6agBJmQAE3qQVAZr780X64huzHi+NDjQHJt5FkcUULn+zk47FAyI13QCXb3jsenlxSmVX4MMJ/
MPPBcDudb4M31yn7q87h8hllORTuLjas8I+HCvksz8tgjlgdfYtFMK2q6sJgxzM0GuH2Fq1aPJEC
gztyT79kDdUMZvf+Qq8rE5L7kucVTYiVbYYoH02gQqHD1fo9amzJ3uFR6AJA6y9wjNykW1Zavh1z
IRvIV9nNP0b+vu5tZZni//dwQwCcUPNp2CQX/mqIkfFFDW9VgOE+JHVF0Lz/yR1QgaS2b1IRQh5D
1ZC8fTlM8ICz5hE7Xo7kPidf0Gen8CrENqzIGPARFf1Q2q+CvlMvddXom34J+qYY13UIJ3gIsKcv
ezLWIJlBVmnbnNWX7gRYHdienlpABOH3bRx8kaT/WtNpo1uRS7kQs4224yQcpT9pBUHRpsAgqt0g
taCTe1saZ/1sLLoHWrE/RoSJC9dFAoQ+ehkOyjk0uRESUEIdRv5e16YP9LbDVtQkNqsDIz+K2oSy
8d7STY8OR7s71KjFNq7Hq7hE5xzEUfHZXoLDp8XNVnUpv5TOxoCrg65DxbngdHMELfxnEIr5Luyj
0+70AUT026C+EvQd8dEHkCm4wETaQGhEpbO6LdFqyk/cgno5U7o3DyEupiAq171Dvw2b/cy/DddL
fP9ICJmzhSdl+mtdekS4N5OaRV5CoLrcrUgp/+/3fKpndTHLzNYAx4FIbXx8aBxHmXCIOcK4NRU2
WcEte+UyeuLT3emtxTljoynlP31VXLTEuXkRmL+VuPbwRdq2RzRNInx2VlYJATmpTM/o1yqFrWE+
awQ6juUt8b7dQ2qlIkCKOhqKvdkd37Dr4zE1qDfHXdDBrYIawUe8hKQ8vHaAJ8dpb2MHPaM1xKS2
2VlcDvDt423uMbCy49ZdPznLf2/c/cgiomC/BGBTcacUIk/KvPmPdgMVZJuIsKvmWbnxddfok9sc
Of43JnyyVqogvRATB6BrXt2s9kHp7WdkPZRna1OIfixKRMn3t+oOj/X8QC0WhW41kI/PTGkbIC7S
bvfUeIF4dOUeiz1zd4uoNa9Zc1zd53bmox4+DyOBz7llps9T3smRqZJZ/HffC0EB4DBPWjuqetDu
q5VSsmBhnW1QeQSoROo486wBYgsb6PdPV4ZK1N/zZOdOqseeN1GZhw6oVUZ/YOZWOsZhUhN+W2ei
JoQJfqmF8EhinWQsCnZ9nzFaagDKnb/Dg/50vwuJvgITfo/66YyXQL0LLMBJ95GEnbay++gWsK7O
Ib9TbNxJ3iYpIEZdcpTOJzmtmCgZH1bYQt/jGnn+57Bqxqzf4sp5pkvhsaismoOs8xwGC5WlfqNr
rfnTICEYXeeLXZeoD2SFePqmJd2y7sZqPGyiYT2ZgFpZAg7NjncPkWTSxTXdyvagP+Csa/MHm4VY
NhoQuHz85WqgCU5Vuv2SArorwuY8jjt+iqZ/rvJBl6uKndcWr03R9STsZnb07k/f6ziYZJHPUOEU
bmw3cnegtIRL/zFNmCOvULQteBYVFgr7WnjqQJKkbwAMFIqD4spTXi6RIf1YVjhWY5cmMiNF3ZBi
pio784BfRP+zsxfAuD97kRBgaxu3qZBIy6DfOhUIdn1v8WCl/JGw7J2sY94KldsJ4vY8soheOK9/
3mAF4YNpjSZlIbA5gkz0ldt1kg5v7MsVAND4On2W5kXF9B39Rrm7a30+ijq/+zB2tScUsrYap8BB
9Kn6bx0RrwKKV+EXM16xRx2vSA8LKbs6bgzc9Gj3HZhOjDnWcZ+LPQ42pqs9izOCpm19M3UKv24X
JxWzJ3KkDO4kgx3Fk0L0HtpCPk59XD8T7KliJnaFGWz5HWP7EXGNeayITrL4eMlXtmPP3L9lLZfT
uykV4Oq1fqIQe3dzNiu4l11rtGXSdziX9fUkdJQYTOj7UDF7I+BDVjHaJUnHGyMYd2h1jzJp1keC
JX4EjcE7dz015KQMhVXwZW5bkWqqgAcOwFxct1f/kjXi5O5mso9ifMX0SoTT20FEIgH60htQJ2KN
yk5Ljea2b9kMb/QT4KbqwS5+gfB/3wwqft40fWBQ0uqIyPrqWIzxspadXfsPTLbkLj04/xyGDiRd
X0aAsjsQDlwtTyLJOEQ8c9P3jaCTo+dGF3JXOhk98VvW32Mt+N6cV7Gf/+DjnNlc4T/RpmKsxBk4
TfctPVH2ENbZDvw0j4xivongDA8/UikkV1LsGyJqU3UAAK0OYZ1G0Goejj1neZq/pnDB5tMltAq2
oGqgmJRk1dJSF6ToiP+g4nBWu3sR7n2/NtAOK/7EYZmlrPxmbZmycjNHwqGLaKx1pQ+gLPtZa4Eu
BcInZ7hpFCltphJVTnqCR/0ZTKZ5LpfWCvGfXWaJOQspCRX6ajVsPE5zwsLDDMxC5HsZM4f53VaN
SnAL86fI0fKT3WFG3S9a9U6ojgqrkRnAUh2CgpItrW0J1W9zTWQ/y2EUCpfxnkf7xfksUCk1tP5j
lHcrc6JszgyDTYSU0Mhv5lR+GPMCNrF9HSG3xhCTpCw1tfbXfF7WJnbECeRaYhjTr6IFzIjzPYMQ
UDi/iuqQHo7AsMhHkB5IpNjOb/w6utK9y2/OYJwfewTVYWSd/qR4uN4P5wND4dV48CQc/qAPTTcp
xoOWp9kqlhNN0ardgPSfwovjM10K2h4UySMPvUAdNmL1dyH9j0srFAaPCLU+AgbPIP7zpQDkW9JU
cViSyOW9VIl193bcd+7D4rR/sFDqz7Ez2WP7Eosq09cvZPRR39QzX8Su8GxD+lngHVz6nIW2nqX6
GrI7Z4xM8bm4qVpUi7dG8cOeh4KqZDPnGh4PYN8MpHuXN8rUV4FcEZNelSpV16spoBen5JYLtFBl
FKU8ZlAhTtNsxkpAUcYLwBk0Ry4AealCTPNPj2Wz5WTPsxVH3eCAPTDqo9idNiNufRxzWq4dvlLq
v4f9ndcD8oCqKSZqx74qpk08so6MFQNpyfVgf2lKY3+x4zJG1Q0d/fVpBVidJzWwYqp7uFfWAesV
lMlT6KCrM+wYd4OV74zDHhbdu0z4K4jPWJcDra24dKVYlL29yxxUhBvkDJrUQuhWGYxTWLUw/omX
tegbVcc7Q75YuJPmwWXrWZvPkKwVuQ71uNJWY2BNpByNS87IGZEaoQKuwkgdRPX/NsRZSMXLL/ox
0messCNhOUwp7nGx1u52MRpRQHxZA2PGAoJkqFTxtuBzC1lj5/Yml6/OKrreQDMfxPT1VO2yZVRE
Uk41JnGBmAwOxIR3KfA6iaP0Ry5WuE2eS/uLXsLTMaksV6dytGxnv7FMZ89FGcIAZkEB+9aEKuIa
/e5xy6erixHFWnL9uLUaKWne2pXaq+sw6ZV78arqg6gH3eg9CQwnMIvwxEDX5/FmkJHbE7YsQV2q
k0/4T3X4cVCaqf10bn7gF+diCNLV8SxN/H3UXDymyTKCaHkcEAxk+E3Jl3KdS3Vdrf/aD43J9XKo
xQXp8Jr5v6LUQ89Fs8C+d+igDNpPnDSf+oUZztEIy0ijtSX73JOJTC8bFG4lOFkVsl9zsQ/iKglC
Y/7qYp8VM1HYohvz1mQncwLlJzWInbb5374pvuQFpMpjjLsPDT1ClE3gK1QFpLtJ08TR6oyGbF1G
Wf1VGEK2LSAty3fWuwg0EGe6AsE2Zf4r1mCWfL5Yj5Amo2OcBBUxsJHKj+h0n3QENTZHd1gFyELA
J0RpLQv69t8/GxrcjDwmygawV+5YOlzpOViPXpDbM26oXzAZ7F9o5T8qoM54k9Pm5CXuBzmQftQd
g6peLUr9HE+IfdSlCZ6VurUbEklaWC0WY7hYFsh3hxJJkVlUq+9OZbB/3HWGLwbgoL+r1eKYWxKV
qHYSYHoPRna3bGPCBS8RlQTsHmw9Y2JS6Fwnl2EAyxAk5JSfoQK1gENqOcqXtPP5BU/v5RO+Q5Ox
S9fPeMPtvoiGnsLe+TaBiZklbpsQ94PA6O/FRah8DPSGkVntzQBgPGebp3S7iIsnoYiNfv0h+aiX
RYsxqE3oZNhKTh4RT46h2BD3RKkdaBMFbPaBZhKxCHZSr7jZ7qWGuGjSwIbdhenem0St7UpZ/bhI
SVjhyBftPhQoy7rr6DLYb892/K2O1pngbEAQMHBtalbVHgSUoCFKaaWQXSfozD1S2QaQcTFgN3Hu
9V/hInKqo+VXc5QvFcxaMcLJQGZsX3Y4WWy8Htz8PwaC/M/9lGZWOrYkhOptDy6gq9uh7+g8PLRI
TsG9b4oTE92uPMJaxZWXhSk3DBYK7PkufUzT0WkzUuhhwEpREu8SSzrb8enu6pwRpf7kTSiRW4J3
83MZV1dSrbJSXe7dLkEsTf7+PNRrUTu6bxiZcXV6zFcTYbRN0tFT+KJAx9oC5TL6KdPkGfDNorQY
lYP2WcPbzr2KcYbbGXH2sp4qzJuLaHFZFu+s614EuH5hkqXNbnlfPxk3JQ5wS9CH95ccTjkz/m5V
7LDykoQDS8HYs6dW+kpsifSOKwHICG7GFRV+fQ6aDq0JVU/CYf+bqHNLnZHj2Lhd7b8Fqu+dgqwz
ZLbCpwm2JvbUVFWO/eUsRWg/1QXR8iorMGTRZaMDiI0qnvWCrnwD7G0jFnqQY313CRmoi0qXeciq
JwNac4dZvLDbZ0RVeI/9HxiKlV1UeL183y/MjJ9mAkhupS4anSOA2MbEp9ePO7kwNXGUqOCCVA1P
5UIfqh2lCjwswpBJ/aYay85hw4dLaN5TOqqpyVmPuNyEdS0C7MuIjoN2vzDlPTW/LKej0qJL9RwA
jGIGWQdZlNpj3GVzwjQiyNSH9GPcb70tmDMtlKW+ROaGb974kHgxbbLUQ3V3TtWCY7lIcb8RoEVk
1IllzDr8N1JjFugUTgZdXVu6KVI6vvlUVu4Xr/qwwj5z0UHbvEUl6/cuPjm9TSO2rOus+TSQtHAH
41opmXQdq3tq615F4maL6MHqJaNxCdrurXF66oz9sB6278gVpjMU/TfemHIvYl8nprU9ofpvqQgs
pd4m1nVnYgcMSnVBojk5dE/YRnlJA1SG5zKH+gwQKqGp3iuAWi9osUJs4l/fVjTLodVl1+dolG3Y
BwGiqA3ZSm7Us127+vzc+KGnaWZAOmgEph+u+ANMVNiiiWtkJ2aSWG5KNzSe6IAHx88GOPlwVN+P
aNfMBNPPsQ7cn8YFxInEVgktgnH8tO7gWswAHJvCnhYzonp+g78SkH2ptiTcOsFn0+/Out8xKzt5
hUOEIzjEFyxpwLoFWuUMn6DiMgdCA8WBCdCag6KaZLvndzlq1r4p7fzW5pJ7Y9CzUpuhm00d3Kv1
xzap87zvhh/mo15aR2W91Qz+2FgBBbBi3z+ut/q5mhsSggC/jaAGWxQT1iP+y2+mF3OuGyrlsuIj
7gSJJey4lij6MEtbpu+TC8Q1bJekAjA3Wz9etEDvoVTgoJn5xvbUe/Qzue+nhoMUjZ9/Rll4zALE
Na3E701hf1Z5iGgrC1DCN+OUf+4rSZIu2+403Ukpk7YPTKFkPOY1tce6FeHmLi2IbrSb9TMnWQX5
kL4TKWk+iV41SeUuiN9PQAXpKYypjTHAh8mhtQ5Dm/QlgHhgvicC6SVMCEvfRIz/3HWSlPLloLpr
/Czdd1VaoFRoq7eeppK3qqr0iX0lFRjHdqQCENQLjjkKP6EsNGfQ/wnkU4asxYpL9dlZ6lRObCGd
K73su8Ze2M5zN/GQ+xtz87wSq32pZ3f9m1+qNDmYAxpttev5L0dKBW1XOGpFinwuECNuR4ZOqiux
SZWgo+FOLBLkKtsthNYH0lLtwqJqOuqMNTwk/y6euMcmmPd08bO8nJhj6Q0QP+t/NNcrsOCuSPaj
5D8NVcL3B7wymJ6mcsc7J58Io78cSFOAyYQ2CQZa1igUuvzY/6VutEnaL7RhHmybvPXHbZtKRl00
eTXxGJRCbvQavXMSzIpYG4IZkFopZpy0q0YQ1J2GAOkDV3UYmzYZ3wvsCvDViZiGSa+nc5H8u8xK
Vw+vJj2QjWgqXvhpfG6IstqsEYMnPiqupZywBD2dtAffLG0gmdj8wGdfwIiFbvCDP2iWL9uwW6e1
55xbFLmts7D+tgllB60OndS4zSl2owjWPJ6je1oQPzzhYF3JgbA9Z2tJ2xScNKW8G0FUMem9Ghuv
f+hgK7ftvfYd8vDcOYmP1kJvduTLaPFsLi2rM/Upq5FxKCNlB3Ln8aUxesZogAYvv0X6Zl/wnWf6
mrObxyJU6tUzp6Gp41Po7ItnRIaiLJF/rYVKT6caCko/+qD/5xklB1HQyEMfwMRtntrk/0GabGrr
SttHdC1Yl0aSZdlgS9sbWxIH20XOyfIpKkuUEbpfDQQTZ8eWtvOHEl7Q7cJn/ArjmZlERe36HAJ9
hPKsbRe7Kds463VWE77yX6QBa8L7+3IPCk6CiuWEK6O00WeEpJOKBOf/x8xrNt+wtm3/6V1R1rtP
Ng74WyqAB5f42lkpc4VbjNT/LY9AlwJvicEr+YgjKyzzv0Tn6oTX+vn8VFXh3QvbZAYeauCQ6Ys7
OvjcA6BGsHrTyPPomNfSFSiMP6ucvjDEfFwuuapozgirzbxTS52sAcM8aVG5WcwKGUWbEXXQzqRs
Cl9r99iYUDta1dp2vE6b80k8A2ZIsfiEj12Hd4FkplgYPnSC4FwskbV5S4A3nYwcWQ1TnQBYSt2+
HaaO7aGXbYIgt7004nWjjlBIDDSzEbVuJYVKBbSYf5tXMHdGm+tyAIxyNAxgoEac0kHQ5icz0Rvn
T7T5yAhAzMP/WK4P7eQn1bQe9kW0e2XS4sRzDgaUz5Idip71Ea7/mnxB5qfr3dRPhr6MVi/9gAVJ
1lWYyQ43KhnHLgDtpYGfjmO3p7e0Qp6ppJ2NOPf02BGVDKiyIqIsIakM8AQizbFgkG23KkI40sWc
OfBlHfE5up03cHoOwLydBplVBZIOmNzJJCJroVoezHFGF3/VxHD7G/bZx29R21zRNYW273oKQvbh
L6MOrh0Hwbxw06NTyKuYZZ8u5TYDS558JHbJnPuQR6PKYYHPNPl0tw+CiesDxhHs94p2iRBo5d5I
cJrGkAZjtHGhNxjvmBrU5wA3m76atZ/o+rS6Ib0tVgjAQ8MJfyY0/D08VW9h2yLLzFO408sNAZ4J
40ETN7Sh7LIG3zfLM/t9IhZ0V2QnJzrNcUmybyHkdtBER9Wx9qBqV0J+R+CL19eDvI8W6tWP/dek
l1bV3OsL0F7LTauLZkvgyIv6d5MKR8+0U+r4EW4c0/iersth1u4v8i5SMI6cnXlyKHvb14QAPVeO
F6Qa/0dd+kNTig8qtQpw8HoNa7g4Roo1ilGLp1u0swy8S58+rFV/pjkaonU35yECW5WOIN2i6Ew3
ggjlcjzJsn1i6pNc+qqEHxQLvz2uU2oKo+7DvOK0/z9cr8mp/qlslrFFIVxnUmupJ2ooSG77aLML
gBmFFq6JvcWv5lJRyE30HKPBbaeZdT7dpVqpQgbs4nxq9X8KPfSeBDV5XboQuTJgFPwQtQWqfHNb
PJ35RiDvXNvNaDb4uqHEmRWdqqJdmGPizJ+CLPCBwFI+OONKNbs6lFYlCiihGaBDY2U/VULOFhUk
MrHxqrL76C12G1xi4eDSeXU1O1xAJtDOTDJk/pMsbwbqNqb4W+4086+rms+ITkqSrETCkmDCnvQT
pijhnIxQz/k51u8T+cPJy7na2AU98K/eDiCQ5fhDSgKfqkQun2QXPdOeMulcsA2pu56rwoGqlNVB
sEStTTM70BgCbvQMG02qNgJ3PZEvX4bvgohucyt14HwXWzwBK/v0x044sFwlKlstyc+Xe7LDi5l4
RwCoKlGeS5hklHZRhz6OhQ+sEq6vUSLT45VDNYPTfCIS33Ug4s3+N2Onu9mv/aRT7Qnd1FODKQRT
oOynQ6+bxAFlDjPsoM8iXIRPwdp+0QdH4+3Qcved81edI+TNey4jT+m0avzon4w2UL+MzPX81MhU
Y7l5XAjENmSkhU1VOHjV+omIyfBPsTjkaFLWPu3E/ACjpnwaVivZeJRy+yteNnz7vqUYTjgUAyjB
eYMCR9NSFc9XTfITwwyXqzTMqJavKk+7J+xhnsJtbIayN56GTNgr+xN6i9WAzeVTfMMA+OyBVAd0
JxR1kx2epx2rH2J02AyuzbJEJ/oLpr2+GBL1+YzdSoI7EBg2FXph5BFeG8KScX8joaZ/Qp1Xs+dz
/avn0AbxBS2xcA32zy61dnEKzZa/saoQai+r1tSiFq7E4kVZ9EceSO9Dpx/Zu02lgfWZqPkL1hh9
ZOfK346JME5xLL2ZCm66mtp9hrTBea8PTggOY9VeYUb/PEyLZQQTd2Jq/7M3GP0PQ3kBVy+fFyFo
gA/8uZFjazIFRiSWHzyPjSWrTSoipKIF+hNdl1NmfqvDRhlY76VjBoSbq7hiQDbq/ckJym3/h+wZ
yI2FQ92k242iw3sTgxn7J+xOuA3Wsjr4laQCvF+sc+mh4P7KGfUFCTnjfg6e6+lPmcuccBg3OFmG
GwvU7+Cq8AztgeDiIkZfpf4b+qrltqdS2ZmeYEfNDy4WAi61pqpUqgAflvTULkXxTUDUFmJ2R/bR
qd3jx4ZZAbgDwQLdd54Bl7uPy9NbIUQSMyqjGnVNwM9PjYu0JcKbHmx2te4PDLWMIbttP38RvhXX
v2CmfPc1nsIfW0/BGm+QEbKAJTuvXbxEklQ+hLIsiEvXJDcSP9vBak6583xTftaKMuw4G4q648Of
lDf5WMSwrxk3nfISErMUvNIQEN735SDzHu8V7mPvLgbrHsN3hmgU3GdgsO7et0uoiXNw2N8B2r4E
/gmBSieG9E6JYGKyATb1BsXVS7pdys/yPyia29fB51E4OC6MEjmkQmBz0Wnah/bL0FBNNuuyGDlE
V0AbNG85+HE3jNeu4+javaUefkQ5yfOibYO7cPzXkj9UPXV9lPpvi4spLzBC+qVOHkp7HW3i2Syj
Ai/Vt8jGte0z7ryjajHQobAGOscluWQ3HZ0jqr+OXvn+Ve12vMEAvhAIkpKz+y48c2w6Wk5O5ONZ
ejFwfTDuFU45qo3KT9NnKrrfp7ARIgQBqFCSvMWrjifPygwMW33XU1I7BXGr9fcWnzjsupMGz6QR
W8diyeKm5PMmJXXv3WJYJUMtdTq/+oEIgItnTpF5QuYqLbAXkX+J4wrVQT5t6E2DCIZzTv5gEf9/
PcxChQP8WEa8kvpzkDZMiPa6U3jaGCKj6SslygbnpShZYvgAJQrl3RjEHLHJBRuZ2p4bVdp7EC4s
B8+oC3FFlHdGB+sAlCEGPWygVavzIgTgtMzhvwhtWNF+qf2w/b9Y+6dtG9v0faUtoG9g4oSi/A17
r04rCiaoQMI0MYtCKZQIfAVaWofiVZGBLjnwUXFv4imTnFn51lkhyf4XlmBc02gDGwS/O79Zz68u
w5VepEtYJ101NG02aIB7W5jjSAXePNbrZANBR7EeZjG/KRjLbf7F1A7GxgZWYQN7Dgl148dO433x
PDnDzAOyhMuZF2jhjcNYusaVo0JegAiqIidUakP9QzlTO3DmXoo1zgM7uaYFqHQPtn+31ztnZjJT
Ft+swSwGWjNyBXNpKX9fLKxs4MyZjLgfWZ2LexTDUnXwJtPL5lBh/geWlDniPXBKJQuiol3w/7+n
ysnaMaGLkzgt0df9KhloP218HFDUjgX+az5pnio0SWYAakxU6uNI292vQd/9BtaMP6U8O7PcINbZ
A/UBZVdDI/BLjHzITDuWln4I2LDNkz3ojTknUYLdh0sZTUoP8LWrKUQvZpThlKOZeMG3a6ty3SgQ
PVpJWkpGXeHJCAgzqSPqqHPxEHfDpk98ImVHJkoImbFpwS6yn1FIx4NYf6hKrUdBQgF1tyVKEluY
S0brmvUzNWMnWC+LkLQEZ8DoOAT4KDECKmnmxwRTbGZVfWWI7Mf+3LN1tn0uJolvdsWG+DF9C3g8
QrdcpuPylgdXsxSGvNAeiSs6CZLb2xjhhEjzLJs0ABbdJMq/QXbKG+dvawo78EmCmVpSsxy/vDT+
xPoOoXjAlr54d1+4ZVrz0KhiaSo0RyK9Z0TaeglsSCDFbLZVgBVsZv5xt8/v8KEktBgG+VW4N81k
P4BsV7Gqn2SLtZ+eDCqAyY/D82axYUFCdIde5I9Om5irHpzr3skSPSwfjiRtx5Q+1JrjWox28xup
ieZILFKOePHNVfYDOLK/YQhiK3aDO2vPwnaCeLS/4mVr+s99ETTY6BWJMVyQw79rXwLKCkn/IY/w
Cb+/JDUSJsMg+5EBd712IFHlr/wSV1jvf0BMd8fUoSgLw5i0XODflupT7k0v3OuASh19VhosicLG
kKMx88ZruKeaxZHA6bRSDeHO/DDaYuPM5Je5+mVl2HzSL+ZgeVLZ3IkjnZYpC7iFprisHqu+/RTW
YqkhTD65s/u3fg+ywMtDuPhKHYsbkmcmhIzUiBS6K5S1O9dRfFxJpkwEWenIhIlgvXlXLe8mvYIJ
s41X4t4//h4uJqeaDoERmRYczop1BOwVNkI4+orcC0Wwk+9yzThLf6iXxOQIGUpi4j4Q4FAAeeH/
i2L4mjhMfcfXjYsrBk4wHSikYuYJ/K4ch8/6dGnaGTBdFKHMdGpjpLCf4HIUlwd0U7e9i3UlwdyH
SHuJBh9LFmE6zeZkDlClUtI0RJTsSP52JYCSxdA1aMAO+rgvdS9Mm5eSpzQfYQF5NI/YjinA7ZSv
pqGtkfGDL6Qsj7+HHd7RkNmPqXDbwzXgFnxHPmjOmFkgovKf9hJmXJi2GqQ12brT/Rmwb3e8laUA
KysR9UboQzmKLbH5KXfoUJH4rvPVvvuI9yClMOxhdz9LbIB3d3mDn+9U6bRsLm7fueW3gILCeVd9
3jvhXQwRn4VhgXZIDlw9HWJUipBMn/jSdwWhh0WEyRQ0MYioNo4H2FZwwMMSQJlQsEyQGvrXzkcD
tiz8ULj8ENjslqIVG6oLTpagdfRrLQArxp79kB6TImkipezGuz83w9GeWokxbri85d4MLf2tTPFg
tuRILnaoAxWUNQgyxDK1dyuq6IsNBVOliUZQ80Z6oAnluLr4AlaZILRHRwgDIcSWnLqt9HCA7YfV
41e1H7MYOlAThtpPWIj2Ze5BQYkFOFMDvzUhFcAaDiljz6Me8ZCAUFYC6rK+bwf9sRMRvBwhY5L4
EQkrTqUFqX2G9CPcqkWN+Nna8HqD0RdlVBCOE+Ambp85qxfZOBUJ1L0H7mzdulDF4KHCLnnlLDbr
GF7IuLILXUwRQ6Bc//VUliKXle40mFCNT+eOgeUpNTX0eL3ad+XKEmCOtXBU+AJY/vzfpFDg3ID6
shlf8kznCBEA6f7H0786++Br5WaKx6v8coKXlLPfxfTuzLp/6wW1uH45YCi4b71/53F4bqDbu/cA
uzHL0qYu0frVRWdP1s6veyDgr8AuM1adcCeFzRlb3gDUBNBPnUnJNPiGfTCvQD5wCK2r1rIBo5FJ
+JTtTo4htP7/0yb5JfCNMDa2LrQzDJ50e4wqkNzPqFg9q3Z8dZMPdEYg+MwzxV81s1TreeYsrDkb
/kf1HgU2VScOfDxFLBSmx9X4n4WgxYKyQo5vMlVMhDYyDSDEEw9OEJuEOVjR16zgSKYSgA12k6Ye
udrQtT+f5kEL4SuvsNKWEKn8VNI/sokw7GD8wyLZ0FL/+OHaiHbxQB4oQ11EKunVxfKHSj6WvqCZ
yASXCGsFwEn2E8ap8FpAtppmhcahOCZFu+nbNpgDU4xm5O4YLLCsIexRl9KYMMaD1pLfdneCGHpt
qNkh9FCkzKi5vVtUGGEDxyXgh0Fn3AuOrvBz1YKV83u9VI4Qlo6uHzq7afUcgEXYbK2AbsJScWZO
43+4W7weQda4bzMsuO8WhlZ0UCxuUTm7PK4FF3M0SyRV+fPQ74KjXBwLRpUTXOTzBvaTeSPf3g2l
1DmEUAsMfMWdn1O9oCzTqeHDrUBUri1/HWuV43uhs/pD/RUYE9aTSF2S4bRbfXzFhWq8/AgLM8ZP
8cN96FydO3TwWhl3zhknThKy5NV6a75xD8lUXgNePYW6qYQ4bYZaILFSBpTj2pvoTXE9M33wUWC3
18TFBVsTUPsyP8qETxIYmBNgic/cemMuRef1+Oe49rl3el5AzKGEWn/byfT90zRKvUQF0GhqWNtM
4ddLZLltUntkzDFoQlvLoDRyVc71oYYjPkV45dKhbJUJ6TjM7p8UWk8eoU0JuAq2zslHZAKZXwyz
3tR2bqL+6HN69c73jcLR55JHhdU03IV6tHgfK/RZPjZ1OcslOk10ZDH8dFtfOEDzrm4wfxYPTEVu
TBNKh533s3n0lVwAk0DN57+jjiZ2La+gt6DQXnsWRAQEcjScC3irXFFoBeRiDztQof834vFvojrq
YvDmlXe/wjVMr872QeiGB9doFZ5l93r7GqBuTBSgru/MAxttZiCzzq+UXpHhw+scOznbRcSxUKz9
0RE5IHA6+fUcZLbguXoUVUqArdpQSGxADVc0LNhPuEy2IYMKQ0otuvqTyWmq7PRoQLd1WSxs878f
1P9xoSujUWvF3UgyOpq51SAoeynVpKsoiDoQqtewx8vgxD3cNOtjY7KEKyFtb1etlpWb0XgiRat5
YinGCB25X3IQvHRiDunDBzmEdhWRzeYta332ONYQVTTosW7xjIfDSVi+CI9hyb/I5S4uWwAoPuya
55u6xxOLUTetvPCtgMoI/80Q8xAFepELDfz5EJdm24ekfF3FiTmm3dt9ef5eE0EFUMLWcM/XaLbp
MlZYricwC4HurKtd1ZEQzULgjJfMtOyN9UDqrTxRQrhYEFbQIbGJLJXn0FMIEKWYA2EmQcsFfZFz
3BvstupYwVKEGDsy5E1yUIx26mWpsgH33o9xsfP9R1dMLRz6qRonsczpeUZi2qfO4Yfkk32Xdkkz
p/A7rW5CfQDUG61VSSgRkx0muSoZXGk7Kg582+F/nMtzGIk1UIvvLmKYYlKgNDXqel3mb79hjLHZ
oBq8gHls8O8ZDqiF/Ee3EjohCi2iEXWHRpsWymU/U2vwuAjRDt9L3jm6wvvy+XxbvLwIwiL0fOsk
bsolUoYa3ceSET5bd3QFU9Sg0Os1yZkWAt2bgP9OgKxgx+A411lJ2BoIk3LlxaT51rZFYsxMTAo4
3jZxech94HX41GnUghPneO+xgp3Uaaxk4LbqjBOfkRj0WdTfm4voAqYvE6FmiGUG5T9xLGBR5hNv
PGTq0u5qmYJwaE+DvzBiO4X0jeGykK8qQf+/dIv4bzeKBCq1wYwc9pUvdnFX0PANOjomfsqCDbZE
mTh2OVfcAF160dOuteO8DukRo7D3lqFpTBGTgwOuZp2cKM9lq1N8plpMWFFc+lzpwpF2WvtfYeig
EqLUyjN50Hy82V3o/xxSiD3xsYuOYOyUs2cJTlWRW/RFJf5WwjQIz4VBBM2vzEkyry74Y74Esukh
F0Yk8pLSAvcGVXTHFcrEKGtGovOVr22u3M7ehsp7aFqiQ906yJTN9f820mtMw+3oQybrsLTlTwUD
WgBdT3HBlJfs7b8bg525DS4o4J6SOIWzmFF5du+Vml4ZzcUBYx+IT4S1Dr7H+p3gJ2TOSmr+zjMA
l1Y2WRsPl7OXOQoqFtSlGC/H/cLGoigbQTxUqEpG6LRUzNRejOxV5MvRBeUQAmUWydNL0ZR+vSXX
08mRURxMjxQox7wv259qTgueBIppZOFnVyADx70iywbL25OxSLi4fDevUHkmJjotZo9ct1HYh9fp
EfGYYm/b+vfsXcWgaZa/1EyWyEauRuntrR3aoPNPViHivoFlsPOw5lY31mCiHPBNtc+esIVC3O7B
PWE0oDnSnjEZ+EGcAdhuMQYCAFlcy9JbsHnHjjtg73Ez/HZUT8F8Q9W4wOuJjjG7dTmCgqXfmf70
68QMqZB00kuX0n4See2PVRHL96HDlF5GSQRnl7nym6W07LfRR3/Wrt4kZud97iAw31i9w1p7qBUZ
t9JFSRay+gsgxvhXmC7ktF7f2W0MTpe957JjN2JzET0mUd/vyLObxAAn/UBNQm6YCPwftskT+ZCi
lKzKAwC8IkrkQmU+nKh4RWh1b7avQq1w/yW/rfSHaKsFwAc4WsBpxpmgvEq/HRr9qvt1sX0vsvrt
EChwNRUKZj/viAzFj2s91+nP4sPTH8OyUXCD+CCw//kZVsK9N80A8cgt8f4axQATQvTrMPZ8EkJh
4gogwewDxNElZacokYIOK3PoyGO4Slh6D7YQbtcnKKGYJncxrI66sJDsDTZZXKoLTIjQ4dmLb+0Q
aQ2VRwYZQ4SsnT7jjzMAQpmNxYJBEp3BfSY1sk4yEXsLuZjId6NoTVJwIhFL7osZVNYvraxxfUFY
RGfWalbBQEx77/yDuVFGA1sec246t3hY2bGVxu1JE3slPChsKW6bXmeI85Fpe7HgBq+CPoXB2dXy
qp6UII+ycJoYFbsKM1EqrElTkGpf61Il+86h6F74nEcPSUXe2zP3Z9VPMNwBHtqxSRh1CThW6jcY
sU4KY2N+iWblWrh9aF0q7dzpN/AVnf7h8ahApbzcBLOV3295tO1cLLTRMFxIBmNAbTf0KRv46i3t
CLBW/Zfo9UHaEY9d4ekFZJUJCG/hLs+pRRdHi90PtScGfDrNUWswN0kB8+mWESGbhkb5LFBYGCAq
+ZAuV6mpZU29AqiHnGMgkJnG1aZct59DQNAd5mup2RPsvfFl8d4tgfynBUtIBogg4o59yFbWmDSn
LuNGlTy7FEixDnllYkWgG01Dpp1DX/6+yjOX12c/fk9s7RsPnc5YSgbs9ianiIL8Y9EeDNmUaw5Q
YPz09wu51mUNxuErrFM6ZfnO+gXvRFSdort5mj3DSyRenCRHo2NoTVc4wk5Vlru60PkpiiprO4mc
AOsACkTbO+qTesdgQBDxztdaMdGk5oA/ijAVF0mLc304Vap8Lz/fOU6xaDvc25YwL+OPaJ+XiwMC
mnJ+PsX02VDy2YLr128VbiNqns79xz87ZGFjOsGFtmO9lIcMfqedjLfnPYYf6YwiPe9JO5DYC9de
smC/qpHFJZzi+iKYlUrPhaWXsTcgN2w7vicr5u2XvVnIoC0c1oDMrQ1TDM7mE38sUupm9tuIdN/e
cJL8VE8Csm91oZH1I24ah9I8nP/TrgXG+b2xfzh3yzAAOsDzrrnfVajK7AqHmd28cHNdh8el16eh
VkDOVY/5orIOYjFI9ktu79PjOKcAuBMl8OSptwgiJxMgAazkQz9qIAyAW76b8SChjsw81oZinNOp
HLxWyP9ZKsQY7MAXAje6OoiVettxMYrJLu6j3sXNLqs40wlmfAMKIWHCpe/74OLzeUbutzByvtIF
XpLETN0RSmBion1agxxXm7ZNq5sPKIRkemO0eesgV4QgshUsqDfUFK1ABDN6iaZOCnIHCP6mxwsS
A/jbTQJpT7Y1zyiHM/e6GzSiD+ke8J1oj3TAiyZA823SbKShXJEruNb9HHLcPi4ALXydt0267ASr
sVa+scEEtxs8N0nrqs2sTzHjGbQ5urSeFxjiBUf/9PL6Ra4/3aNTe3ta4s8XaYpbCnniiHsE8diE
6y0+4goxtob6kmTSRsrGmMbVrbN/nuGoCDCPUtTN5UP6kcCMH8YqXT5kimyfkqcWR5K6IEVKgBQi
Re0o8hTfxUOMA1LAm87RDoQojjGp1bYMP/Cj8KksjGn21N8uxu0ZBC1S0x1WtsOOVO3lHdhM7ocf
QtljIzc3/qdstndwc/MbacdIRiR3vxBJvgyasWY/kgSQ5ePboNF+6/4vC7cck7LE6LpLy8Qqa2dn
CYMtmlaE9+1NMdgukwpcxEHsq5ju8TjYDr1GVXynwCwHygrBP5y24BGhLmedNS1PmB0+UOF54tmc
Ywy0hzIpqvoWFBTrhhB+D5hQ8GXzKLNZlBw3heYB1NDGlXaIdG/j4UhN48NByKyogA/IELHO0PHz
0qR9n/xucZDH8zaFgETYy3VYsFaj9Xxoot/QYj7ENuOXtDXGDnTk6FuvIXf+Z753R/3uVkcPCxae
7RSwHWNAlXSE20oB+0b3gp3LVC8YHnEQubOW3UaRv20EQzLpNdVKa6DAdXtSDolRscQDwGaYtw0k
hv046Q/4D6Z6RPI0jPe3JLMyA/oUldfwhBIcw5OPTVYczKLz/1nA4yyktIWt/81xPxipz/4xDiln
/CEsjdXC8EPmPKS8pMhBWO9dG8bCQs/ckwglU1ZW5GIlEH7xMXfodoho1cuvC2gk83pnTmaesTnQ
hGraE6ug73ZkoksUpBLAH7x5cvpnbMWbc0V2CakkQ3xKTNXt5OkXAidlLOOoY84DwilZ3QSPBzfn
EizgUod0N4jvTgX5GQFkmdWInQY4pkYJ+Xr2jJsYwWdiO7CrdhCCwvFXXjpGjVYMO+HiPA7G+pQk
pEz0fMH8CzGRrRHFQ7TnNGdX3BmU0r3FborCngpT/+TSVRQvnABnb5HComeTI/EZTespukO/PCEM
LbJnm6ZWQjTLhJwHrAW7y0emdJkHbB7n9koXWqQVDa1PT4tGS7FZ2a73Np9moLmjTNdrhLs6TNLw
6nyIXGEsNnuxGql02/xBV1AQK0SCTu9u2E+axDCXHwhTKGlehMmU0HFPmkg56fm5unCqF31A6GqZ
uSTqwNSxA9tW4BqiZSkp5T9nGAP7eNKfNHtvRpMgVpc+R6GsoQugf+0yM35heQo6A+Fynle/svJC
44Om3iivKcfjLgbwEJ7FBNLwExHp2bDanqGdTU+cX7V9s3opnsD9EPsFkRYw6o5LwxigUx27GR+J
WkPFGofF99DufKbC34sX32wJHm1bPmHpKpjdC5a74DFikQYI3QVl0e8gi7qzkC2KPyNsNou3L5uZ
yGDzkS6lOh+bfwoeli0sQ8BHwGOhlKRuiRrPQ0mv2/OjXy5I+5deOg3JujfdGb4V3jZOwK3uaCie
TbAZJVdu0gLBPTuH/ZSOBKvo2yl7ZU2XOPIfPyITwtAJf+DqH5Hf0gZgNQeRFMD3gjxkK5WvCFfp
IjhZxz5OwWcaBI64OEtpxM0kMfYJp/NPICI73szTzzjP8V1nKLxL5seDSBGYJssiyyMr/Vgj5f6U
Pz9OblwxgYPUNtbkLI8yRNHy5c+FEAt2n81gIzMzdfmZX/4q15AXGD716xvCbttZdTLNJWNzav3P
MbptDL+gdDaCyhBDUTJ8++GuJaSZN4EztpQ6OlP0GkckzjiEvcnIVJJN3XqT99YMKmxRiuaN2gMt
7aJjpLvc5PCQ5K7iDDknUbLcOfNwMjlUvAwaJ7QWe+zfKSN2SHycz1ACO6h1C+IzNfxr3GtvyWAo
Sxjv8kHcNX5lZjcPdktAPyBH4T1aEYoL7q1l9phHNZ5aSMDhzjMJG6HSD/ymhPk53SZzpUgGUfxw
x8kbnVmK0Qcl+XtL6qHM5730RoJUv1AlGs4L1hUifwh01m9zAqF+/XTATGq74MFuN8UwFjgBBnut
sbTIqIk+oFe/Sw/Y3MbIiHwNTWUo3lFJuz4UDm/YyNQD04s2RbEeXM6kd55DTV+OQnTckeXfhviy
yEMPqLL1mFKvbYkBUN15smxKCiAZpc/Wp4AQKM0qULY/JKm4vxL1vrL67mTXZP/1QNNKQUbZDBT5
xWtr3dXP7tBk8K4pAjPG6ihbZeoEfp7g99h98faUJEw4QWZrotpx9llmA3Jo9sn8zqAo4PxVW/yG
mzA8/76F25KkLROXkdYw6oa+V/dOJTO0qAbiTWgQYFaNpbHRWnpemIhKlMftgaCp/0vjQzCB2/N2
s9XCD+0T7iuA5sm0JYvGHlns6xYdO3/81Moc5duUMDdRTazSPKtQuLJVpuHDDwRKoIyjazc+h1v+
Nr09GnqPP9qbQvrXRC28
`pragma protect end_protected
