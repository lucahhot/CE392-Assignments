// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
JVlflkw8gt/dd75PEhoqkHFkOO1Azkkw3GMvsfgzO8sZX7ZU6NT2bzQDa0Elt6F4V8MTu0onfEi3
mOX+L8NAEunEUiZxuGpxat0c2RVRYvjgyVaWYBSN/vsihjtKK0LbrC3makCfox2XJrVtTlUkhQyx
7HlK5PBbrFSEMwSvWFK9jS9X4SSKqCDS7zcSxq19Y7FI7PmjsgKdy5xqQbLvIlPak2DwQHCu9ktR
7QlK9bz84qDT29Zz8IPnaLG5ZW6pOmQKR3EwSRN10TYDmCrdZFrFexoSCgVYjYQ54BPTA0GuixTr
C2Wqe8kij4Kf98PZ9lRtiD3DkgD6wliZssfeKQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 29776)
13Zmn4P3xepJEEHSaU5EaKjuZzgOllfdhx5PNbvdfcqnLTt0+CJ7NCkYG/v2+aFHm9VkeIEhE6ZE
Hgdd8mpXck7yW3Ms+14ZZJgxSe4PyvNqZc6+HlgXGgLYs6W75d31HKGvCCvZbjA8Ko2QySoKxUP7
a83k1WEJu7fKb/ShIXpW5Nnfr96NvbnTulN8alP6+JRWmzBc1u+Vkc4X8+KpzOSUEe2VrmqhKPBl
tTXMoN87c77bJMF6kX+glU/JHg9WwwI+eLfGOSiRmP/g1cDEX1uKJ52ofKjM2TNTUyB6GMnj0Yow
CK/b76zBtlHznMAucRWkgr5q0GgxBaEf295ZT2StWE1WLHxLEivYoc66bXbCY7XAVFfJC8y2IDuo
oeL7lOnvlFQUAvsKdwh50bh9fqOzPtbGDW1fToFicND6O8G3tYDo5Kuw9s+kCoE8m9CNe9UQ7UIH
f9yDLdVU86jC4VW6DZlwzJCI5ft7kW/fomU4jaXqaiIFEYM3I0KBYJFV6WB/TyhHptGyaxSDB1WM
Q/h3Pifv5im7cvzS5kEhxQqXrH5jcL5PtQ8Ix71iNTJTbaTj8HY0NSIkcHIyPPTwkM0rmQg+CVfG
rfU7ttaRsIlHYb8mbXVYz9lTbs9qPOzaTMq/65APdVO4jpTzgFMwVilLMZyG9pysqdTUcgm9FBmX
OQXz/GR+j+SMqzMow+CjK3kS/3u7ZpBRPsefIJGeKCHXPHAT7o0qa5iSb4ZFs0ComWEp1GxeAVnT
k8+pWAdIlQ3noqvs4IoQUZ9LQyq8HWoVohFdzBC4jpsv7xWdegnwtV14E2t+2+HllWD9fo6bN7sa
O829ClEZhiS9R1RYt344g/nTTGx6eikxhR6uXnk06E3pssv46PpY9W7/KZyqbrf08wRcyBI0W9Mn
x0Y10DS02ZFo0G+Wn0ANDG2tYFSH8Hnvt/QI+A2fSQ7CjkJOwFsWJXWJFutVGZFQ+7lr10X5Avu6
eF6bQUIXuwcrx+JiXVYJJO/HJZKuV7cU0i9erDjPwiqGx58ub8Q1hAU2bg7PAM1gbOmCkfUr/PZq
jxdZuuaJ6ibfMuF60RXuh32rzEYaU2LoP7xSUpn9FkNzclAxgvmwHx9CZ2qyr+khyw8W77T6jjtQ
DsXxqQRn/WAS1p21z9jQYv1lYqXovdcyAhj3IjlrSVfjyDc50ZP9LRwB8Msmq+k16CxPKZKas4EM
Ugr2jA/Y0Z6uCmpkuU3dP3KPRW97ddnjtv8IL1u7MpotuyniFtZB+uYuCf/rkbJ2CJ9HdJ7xZTLV
GsVISCD8ZMzvM/+wqQSXfs2cRE75YaJQF4gMEb8pFoC3ZCi9eRbgLctkBh+aQiZnCOvBGdPJ2q7r
KSpNvwUr/m6s2snM/mN/KghGnxBa4U/ySxJxdFchRX0a5o5xUfI7TP5F7m8vUD7WOwTGpL6ETYJp
2NwerY83qpwXDfkQSDB62B/qk421bo/ZB/n4qr3zpdX9A4jm57YpzPov6BWDlhgA3Cy2YqbRf+UV
+BAmfkiAXoW0d0nLmY36Qofg25UOYeSW24pq/VHFMBan8MTMXwlqwSQoBLVnm0jveYSvslN4phjz
JqyQQDePrK67vjvZEMfcLlX9XpMq57UWjWT94VCT4cOSfzP1DiIhW6y5LpjcAHyEVvOenxhcEUn6
DbvNrsX0afS35x6RP913ob4CS6SpItKiv7vupfleEB2qmC+i9hZejlfwcHMUtIHPglwlSmwqhSBQ
afTtjOkJLEzOn8Sh/FalDJlEjP2SQjTfycIIlM9lltQ9rzubMHaG/ArFoxejRrvc7mPJ2IEkyls5
9MRuoHxVjPg9vH5GLQChhC+9/jt1BqGdhMRDB8UkElWEBP5sh5NRxEHiM2R3tkvLdzmCp+NXVYH6
zGceXdO6XmnDMLaXD1dUYu7nCyCMtayy1iYTjUYa8BBVdXZX6slQjZa7II34rJ2idvFljYh81+pe
jXCCRCOLGUbWu75l2yDho2Ta4G3o8mPLhKWzfryLm9VrTd5USz22MPJmqznbB+sBdhQzJNEul75y
xYMIQ8iBwnwS/sKzAb99AD3izSh7Umasjg9z76c3WCquKkINJ8lvXEal3nP0qeMmNovjhOHiW1oL
Qy+gW2Q9H9NeuqJJpjRlmDNt8gRN3ST4nbiUDFU8murlvfIwGJhBoOHlx/ZCSYtPAswZoKdV8CHT
FFkAf2g8jF6t42jc+z9jRpIjR7miUHvAgwdBHW/sIAVC2Ah3cP8h+UazRvKpIZkIXlhSnxj5SDg8
GxR9Ww3vEMVOBRsX1N4I2gvLRx0NoNxL91oPNBtHFLnCGBXMuZNm1ILYTY4ommHnq4rhoWfpf7Kh
i4WtYp8mN+EOFdQI4tGFWDRbfrsiyjBfJoDmGRXTAeH4GauGTviHAzW86RaqL1JTR+Yu5QmFN6et
shu7YOJerQq83i8PXYhC9+lTBB2/SoOQIhAQq8TzsUviOhDNnrwAZxHZNdiGEtDHIM8gfFRWYqO1
CKHjj8D9teaX0Dg1FY1Q8hnORuq6RphFCyoRihQpL7OIKeuXZNUmRCDlejKGOZuDXVhI6iJc9LcH
DyVgSMGol7txmyvuSLf4kBkdHp60ZfZ0Ti05384GPBklfrQHuxQT9USFXxSMzyHNGlfrWPFkbb5g
xOiAukwSmHEvFwkFF133vTQrbbwROy4lAKGQDwXkjSSsc9RtAd1Z8ZfoPbRZpYOeAe8KarS7kgPE
RfgBVGJzs1KfQY6qqfTwI5zc8tHzDq/wZSrxibFLvNrExanEKRkbQQpaIodaMu7OlHmjz2xscYH+
dsS/HLiSWy0W7t8eVYRyYJlrSr4epNZfQtbocA3629rwoupMbfneq7Rk20ImWkLn1w6pjGCjhjDl
DSy3p1aXXey+mEac7LXIS8sSig3SFVkxGQrzOzVlwM3wcOKgVy2O2yailggdXqD/BZzFeoqGlsQf
cBI8LZUiLsGFEIunN1FS3bfQS23f6AddKZYsxlVMNQmN1ASP0q/vZyT9ukjQM5v7oigKDdMm3aiv
BU8hUNDcq0PTUbBwBZKmHsi7k5Dcn04Oe7yvAsD1XWOmo2HGCoQcgPfivRXEnw8GcTmq6El4HwmM
ztvo3o5TazTOh3dI1iTmgIjhFT5zqv/Qv6o+fa/V4Vq4jZM4eGRM7DnbVTZ2/RSRURja/slBJ5aJ
W4C87RSQ9r5A5w/MYM91DTbyKdEv9tiXRv2X1RTfauaFdzD/tdK9rzt+OFA12tUWdNMk5zcgQnHt
6NeiWm0Dj+tvaA8sNH9kDgL4N3eZameIAuBxej74RQyi3+l8XSLoBvzWuU0YQ6lNAAMMHCax/+wP
8i0bg0uSgeChK0r2H0m7Tf1cULIUdJSREldcQi9nNELVbkZemOS1PBt/lxiWzyNzi8uzji/keYAM
K2THvYl4dUfhvxiSWae0lrKddTWUzBW9NlCJ/PX3eGmmyg5Hb91ddozr/wOpw/bwYsUUegvY/OUU
0yYgle7ybxTqTN9FLknchblpBAIEUakOOdU6oGg3qEh1OsR3btnv2XFlcYeABvQIpIAa5qJfmvdC
9YavDPI8apsYpM+D2e3ITyEkePeWuPtGZW9aHdpELIjw/wZ/otUCTzh+ysztw1GGTikPdPovsXLg
VRtpMfPvb83pZTrd1gs5kflEW3EXaq3tc+QHW1BUX4I3QChs7Yol6o8tSNYNdxFLPcahXgMim/rT
uV5Zd9JqDKofMvaEo8gBwgRBAlMbIyiSwlA/lcyLHhzQcaohRHM1N7/QCiNVKoAY624l8848zioa
OgAnG0kQCBMQ8oaRrZXOpbthLBai38uQA20pJBSsPH51ZJMW6/W85tKnYmSF3grg1Sy94mjcvbK3
SyhY1EuHYEL5SvfM62Hh5UP/hL/Oms0gX3fKSAvf6OHbffyiC8SfxeU4IaBlNiGV+MgN2l80tlQ8
tGeveZgOqXnZGyG2srA0JTKmZIzl5AkrF/WBv+ajW/kVihpPhuvQyScrbvlxJxKT5guHIEPDiyWM
kRxsj5wCFQO/Sk4fgsdF1Zxz4kkDPg+F/t3dFPlA5KcNTnpslLKVJc25kIQn4XN+i3cInuUt88iF
UqXtQPLWqU5QoSWgwCCKD/7++eMKP6MDKSwBLdDNoJO+7+29fFhUYHC2Z9jQ75Kozdu0X+HalFuu
LeoGN5VFrLnUf883KmjA5SdLCy2r27yWNOyRduc7lYPHdHqF/nT/eZ3bIbXg1GI93f/Re3svovPu
fA8eOro50n6zXkTQsHykpRD/Z7y1fYEWGoGkQs7A39ubdKbo0mi65jundlUZhX99jYZIcJpeD/JB
Q+TLdZ9f4FODiAD+CmQ6bj4QFOdfNv61spV8YIo3Csm1bgE32V+hIT4Zm3kf4Rv24JaneXGqp4aL
SeOr8NLSOei4FPlopcgBdWWJJbGCPv7oUTIuYpn7mi8GLCcMgDx+bRBGEgZyzGctVzR8B+3fyvlt
Jiv3u4bsjmJKTq/oxHFXCSzAlUJMUAy+LxTfKfj6Jou7ItuZQ3xoJoqrZRnh6dtF0W1zPcr/xTf0
OLx3LbAzZS2KvO2SzSH++NQlGw16D5r6msLHuMjMLMwfTZSu4YUvgSjmkuOeaNJW+cx1a49CA00H
9khjPsEeUpf63L0fdCarDDN8g9UE0W162lqKRVAk7cDNZarsEtSNKkMo+MnQ8Cc+Kx7YfTZMpTMV
Jl78V7TY3EDoT7g8VQPSrHBw2kxOfivbz9Uwrb+pWKhIqVlKTAskQ05Q5WZskdHvH1YUcSRG/TVx
MgMWM5iPvzr/EyvAJ2R+6tJt2lvt2riRmS6ot24L8UiBgYY908eGlJtJYYKxX1CRezuRqLNla1x5
aLSg+0Gp593p2ydhNaPJBLyXx9n15On9Qy2QYOyRS7AWECfxDQ07V4b2DhZAOCkCTwUHD3ng/rWQ
9HRwmduUMXNaLYfTHjW/NM9H01TlOUzYatp8go6DBjnjd8DW1EOFgydUvnvYvLj4CShiDb67m87p
6mCCZCTrs1X8Z4JKoRutTVCDX64XZQ6B6rr8dQJwodyQxtVxXYD52KSZ/TStnBJR4ye11JUiOD38
oUVqb8sZUOmf2nIcGCRMFDAwXz/a+hmunxFWTBAlGQI8OpGa7iZkak6dbsMeY1FSRubMJ60EWEZx
E3WobMqLp+b2kR4Eg68mB8JaxMQoj7rp2q1haSTpW1ebqGa4cCGTAw/V9niv9/YEo2FHRhn9xdMV
1F35GZN/A51RnK/beTj/9j57F+beG6pq3ICNcQqmfbN5l7LThFO+A9FqI9F3Lq6y7rmkht6xmHwD
iMNcv98bH0vxiK1TOzu6mx3NoMC6GOZKkVUN3ynsG/vJk7GQORj+o9vRJQUxGgeI2gUGnRU5d0FJ
fIdBxyuKpYxiJUyUWM7WlXEbLYzJV1aeeLJSy5eVSZNyOuVoSisjvxyUb6JGfD5/kRwgsAIReFII
vq0Ds6JzwLgbuEytV3/u3Lh6w2iU1+avH7/+6OG6fWlT6LfwTd029dJZ7nz842+dtPqUw136NIc1
QfNbbDlp5DD2hIy5cAHtbhM7AZPXpPNViaBolDN3VJcqFcgpKlSEcL1LiY2ixbzZr+TAdc4mJz1r
JjKt+7lvfn839VBScVtFODokA4a21/u0fiiArqEjSUG3PBVsiod+3Ww8QDzMpcRrNHmfsvAbGoqU
3GNFuMJVtCeFBuFngqFsf6fnXXI2XHn9KPn+MQHSMyjfKKkBDIN81fH5PluFp4YEwLEy5DUXhhNM
HNeulwWCQkp3KTGxfKCjTTvrO612VtjpEUrudap0m8FiR4os3GwQI5C1L3os+7Ic91/jRDwkR/S9
3xdRBf7Tsf2nRI1Z+BnxjbgnWOoKqdkjpqpXNE+xZSJnw53ThaHRljIzVsNNpLNyNdLLQVW/YQIi
i7OUMJKW8uNt3e5Zy5o0P/v7DGEKxKSPfGLruxg4jwMyNmaTctD+jdTDI5BeMBlde1BICefvWtYY
qQSmBOjYqqvEegGkgzbASQ/FunRcEppwxHzeYEsGest7hSsdQ9semEba5fZUJILFZjHQaSx4ijhl
5Npkp84pEodR4B7H5c+jRe626QcxHd/TbEhz02gzp3gg7yT2Lu4UuJJaGr1H9Bs/GNufbHpFncVy
mIj9+NlyhwarlmrVEnz0fSa8F34SZyTI7KB7IvKI5Sp6Jf8Ur2Nv0Sz3vZdh5TXenbpsnuUCM+3h
bi092nW43LLMAbvijqXgah06bu6Bfv7N/pt/7euIwSC0OTLInCtlBdOwVbz6/UUbDy0PA4lll6sQ
YOWVdD7d5GyEV0IV1LOMmHrrIp1xyBygWUBOoNWUi9m5OXRf5j4Mqww3lUCRnquv7SwNL5TP9oDn
Ab6zzcCjco0tDg/1WzQ+4UkR6e6ItT6EapU47FZgj41IBTw1ggMdniIY61VBVy5i3z2u5ln203V9
d/DNF4zIUbAT+rjFsaPPeqvkXtlmBQcb1DcPbJ/jmyODSYb9QPDhoYm1rIxs+jHXrrhIbLT1nclK
JEIBbsQrq7/wXo3Vod/1G0dOHGeI5K/blgWo4d7km9ECcclNFNLQ7v84tZosBy8WH9GbmwEh5KFG
dx+PbhPrp4qHA1iiCCveYpoWojxzx/LECWB1H8/VJRlgbdEtX5HvqD0yO64rAZUMKzNsQjXl6sX3
k3hiogBLd0ZBQZSiJ0H6o6jYFAJq6nhevAFdhlZBCFzIlYhS/8ErQ9tAJjgqL1sBJvF2mp8+vCME
/noh5L8UkGpEelNeqTmSP9Bh63bcPuPx2FOXITS68fUtAUb3efsX6AZ4xOV9FlQpTWkqbxaOwGyY
IRu7q/LxnQpRA3rJUsVFC2KiSGjtrTKgbi4havTwCckwM8H3j6+9JMisFmLpC1ihTKA2qMkKAthG
E4fKhIiGd9IXoGmgHRo08SfZACQxNWtHwhVusEsA1Kv3Vbov0re2vnhecRnamK49u5q62whzkADc
Yuf+ElR8JvZ/PUl37Z8BVqY3fesboJkXdqod1E9cQH6odNHVRlXnLzPzOaaccgPBWAU0fqJtu5g9
XXfhrm/lpVDYCRT/f4yMU/JO+DtX2/haibFXk4Q5UQGrvey8oLeoJe4RVf/pIdrS9DUyCS9v9GjM
qT+MaRkoa1Ktrpf9kwPsJTKbcRPh5PsX/gAAPS2nt4/RCHdLyMa3U884QsdZBAblka+GzYHIqRwY
2va+TN4sfLoVKdMEyAft+NHl0ccIKVEbROH5FIPppMr8FAzvEg/jOhy1iwrmlAAjSD1XP6wfJ9Jw
8DAOrIAIxUXYJl0bdTB6H+rfk+Zqy4d7JbZ8YaA6me/1BxTMtf0mImXnhlI1QFgpoATk5RQ9lAGX
RY5+thQO1/gO1dDMzh3sjLF0QBMzVfBrZVibPvx6ZSLQWf3bM07bgzrCk72PhUS8ROPuQAir1+HA
vI066AHC/t25qBm1jk1jGLTFJ5Kbr//qIQjEyUoidExMs+ZiD7cysXbV7QURgams3U1Reev6z2Mr
zNSzh+UPYF/EjFB40otBWkuRmg+oBHmRJ5cFLYqqLuTHVkGto1feL/uPyTIvyPRaGFloRKufHhsd
dp6AKK3lmrAqnNT8DnOzOdciyoD2OJWeYrRtDdMr9CXfqyE8fCqj4ps0/4w6VBSIwl/oJeoxgOiq
qi2neEkGokjka7jXCoFA+RNPpxfmqlN3ulAb3+WEWxjg0ICA09RTd+dZXm7k7G+0/sfm8SwlFToX
Wh/lYiW6IYD82Yop5O+/7KHwn5fE2grY8pTRhn4H7tAKW1LsLirWDwtVrrPR86Cnf14xhBp8k+qI
4z6RHZgRgE24c5fPudMMMJn3V3O7QG/QD8inXryvrlEIALDxxs87MOOEPzsmA8U9/SesZpHmx3cO
sQw2jKrG2BvknRzRjvOAat9dFjcsOfzNXRqsgF+iQPAxOfffb/Cgvn7WZSgV3d7rzs2EwtwxGKKt
dqTN91eknu9dB4ZFYMe9DnpkS+nmTfq5lgtZrEjQce1/zfz5GPGHtOkCthMDJ3lWMhIpJ/oL09Pw
BJUXosO2nvM1IFhbxisJqQ6b1l9W1KYJRSwrIPuSJ1IELGTF8mALQVdaXfH+L66pYkUK4hlmupz7
3Vb481fjabn9NUQYZyyLwoaIzoupRRf9Di65ZTZsRxMP4QOmCf8TLM8u5/f0J3iuTDlY6pWvQ8KC
iayxElvf5jnfskLJN4+GCMRJHFz2jef8UdFvsVxyGGpncCPeQxisZlNhW2tTEr0Z/R4VhlGUXGLI
pEhhdMaQcF4Gp/j/xGCXI4aCbTpm3NI0KcxqK9k8iUcBOUZIJU160dJg9H+3AHEhzu93jxtxiFm4
VxbCMDgktd35bTt+OoFnaHOHmcKJsFgxNL/2o6gP+VMawsFTn7aq4qgusb3buuCbqvJ1fBiSDfJS
dWHnH1ao3v1HyJCLfK82FelSRAykOow1NFstSWp5jHrKqNdvcJvz4tbfBD95ZEZFFqCLvDrAkgSu
d4tFBPsulw7L49IO5MkaarRpf6J6kJJM+wa7fst6F6xGIVlrDctr4iqgwnyq3rDGbYBtqOo+Ttsr
wp+Cj/BHnNbOrcK83FJpdPb+0UArcOf+WlODz2bhK0meaL7RFVa2D+oHHxkNksaCopxsRfIL4492
HhW3H2WjQ//7wFr7eDQOlCN9BCskmiKnf+d/M49YgiD8C5G0bset9pzoTreWeOQ/BT5lfgm6jQwj
1HB6um+O/h6o1IRxqcFH0GuQJ5P+5qx1VpHxw27LttTY+4JXr4FP6z08soGC7vjbjUbAC1q8IX0C
PX2tSV+RpWC8aFh29/WSUM6rzc5fVd2eOgvVqQmKTX5ZPuzbuqt0iTxLIoNHCeckALaibyvPu9OK
icHXRHggrPq4YjxZnTrof5siHCoWtRTUSUDE8YOkQbBySlbNS+QXLTwUrx/WiwWPDOaodihH183j
RagNqGWMIz21QBAJvBUcQj9Rr9NDr6HGQEv1DRhT8CmKdpZaePVHrGqpitjSDpS6mYotNct4dCdI
3y1ERV5CQb/H7Kq9PbKvYp8OiLWEagJcsymSVCkLaw1Dx8KL1Vd/RaH1CW2avDC33q7tgmGzbBaC
B8hKgrJ+jFgVLoIdSu2fOAbJ9wxh06jHqwLZm90WVq9bgMhYs3i1572mIe3cj9k3HA84qShFzhNf
oYByOyiOqB818g6IPmDLtL6IhE0YHoy7FWTHK3Y+ctEqZEUpAkwE4xQIdG1Gj4D07lf9BBgOjU3d
7/zpsmdGkCsJOpRPb/8lrISLlDHVwNPTvBmw4JeMhK7nvy3k6mw3AvZX09qyYm6KzRhl4tTtSNHT
6vZD24uSTqyrxT5J55y4H9nirsuAk9LlDqT9CPJdMA+bonSH0P+cflRqnaIRxgiAZksqFg/WwDKk
9fbCHqKqpu0W87Cb3oRx1bMRQYo6DoJNmQFtGXZa5HAKtBgAeqxj11LHw3BG+oC9KAzAptzM2hyw
Ozm8wOWX9iAHn/OC5uGtuI66PBdF4qkYhigq0w848RmTi0WojnBpE7VmROEAT7bd29Pi99x6nyo2
0vJF8yR05a0tOpQDsAxdB1MP3cO9YjzwngRiaEUP3QSz4eZFDkS8FyxxMkkY5zL4flIHSdEHfJdk
lJecbs3irAQi2kUCfYb9jvVOCl5f/eTv/PQ7NW3DM2VrK4MIcZCBWARPP4rEfkVhOwZ1hT6au00L
BHmRpEEukKpoBroKbiSDtgwNKy4obJEosrERKbqxzXD3YF6dQR2AD9Tuy6KDMBJH4roFtX9x+uzb
WdJAD/2MyWn4vsrpG/QCTfFhqn+DJ4AdbufGXztaj2pQJRxxMSde4hHoZGxDJGE1wBVH6l39YQtZ
8DlB8KcR0nhR+pGuOvfIgFyernFohXAQimrNaUPtVRyIdNECDywYoxqFsU+DUDwYI0NyeRy+pVRY
XBPxN0K+Gs9SFoPlXliiyHYMyT5DvTQNBE0ZZCJfno11jJk+wAIuFOTkNlGF0Flu4ptMMWg0lyFK
IrvK/gU/6Zp/aQNTk7fuJoTkOO4IdVybExtsJXYjGcoq3VWDQpQjkBYM09bchps7EXz/z/PnrtY8
Hfz8vWvqNlbc4/gwAhQou72K6l9THvIRRCIC87F7L4i1bfRx9bqaJ/01UoSy1BAJ90ZlBBeI6KBv
zTmT//1jNUYKLZ0oRCrnu+dxwg8Q46w2CxQzPpJJzJ0MfGp6TF5L1iHiT4b2/O3sjz0wdvAADfkl
xnmd6lWqtYfgUnUd217QzLJEfXbWQ+OVWiZmbTd4FUq7Pwrjc5pnG+G6EpNxlbcGScP7+q3CGejG
JJgbAIh9Q2W5nywrPU6A5y8mnVuMDUVtZeLHqwiqMMiZhsfu0wSfvw3el5IdDVrWziNC8h7JEBGU
CbSV15Jg04AQ9yT15uEZoOPIkjQvSLnOV47uLoUEDnKHkNwoimGj+hzAoLlHi09QPSpbvlcGqrdX
N+jQ29ieYyufNWmQJy0Hlw7mH9FcAPtMAEdK0R9o+8oUpYnXON3Y3On9KWChOzGydo8H5skAm0CG
kgYH2liFGsJLG18Uzor8tn0Z21v2Xp5t3Tkwi9F/XwQreBoUWi/au7zHVaBph39a4K1fZ8dLhl8t
80y/ZegIlISJoIhI3fm8POyprO35y2WLp05JhFtZV9q0fXvUG4PDtNd3CGr8+PWbN0C7rIKoXzNr
kdhMgVOnGE2zqgT/WHx65ltgFV+1fdDPLZPIuTuGOZriPFdJZ2LifOvnbcBkm+7SyTRPh3q4bREr
uea2UyCvI4I15H3m2WSfKkeeNB+zdUh5LvlBPk7pQ0qvh1rMqLpdfB+fUS/2t+5UnRiDpWX3hpB9
5u4ovLnN8Khyt3iIiCU5q6m64Iu4lrDn5bnXSv1jSNeOBUNQUHdSJ5jJF6RiWMUHpxPZA4LANugE
S6IS964EhIK+ztFBevnM0ZTGxoG1QYaWUqwa+nDjKqMkVVkGsMU3kH8cOqjj5kec5VI6Jw3V35dS
cdVU2i3I9SWumJmCxy65CjpERsD4DosfVHInAoyDs94OXvrYUuRd5exsbOAydJwaklbFaJ27nZRG
Wq/B51R8F1aKGW7hPNs5+sJr+on+CD226ooEoBipebALLAxuJnEO0wV/nHwQ5KB0I32raU65Y07p
mzPRPK2VXf8gDyG7epGgAbkW7YxWblTzdZ4PaQfVvsbxhSKYbdLXljWsJuXZ1D9BMQmlqA2U1mWB
NsIFEG5TMkr3DLLLnU6hVwMosQy57oGmjEiXHUxzvkVvbLQMVzcw3hiRmtD2eOA60BIInlwA7rP6
EdEedC551+TZJk6BWkBd+I4if5nppPzRk+52M5MncX3Am9px3P3qMM72L3SF7czq61vjdt6tI/ox
+Mv7ol3PukL+9wdY/6tB4Y5KZftgkO+O5Ec86VX0lSTGd2n2C4Lad+LMxt1NTrx4tlYDXrTmghn9
/OB320TXELapV3Y0WIqthzSmjCmO/XIpZEVj7TurhQAPqmljhj8rINvTp9y7bGW1iF5vn/fNmNtJ
EN2iCf9Txe0Frt+1auoX17d5wOxREctyseghpFfHZmjvWJujDFY1C2AC2mKP3POJyBpOlcivet33
R7IDei+usa4853HKCKs1LGdWv4+2bsTguRUmOaJYkcM8R7oKyySl102UUqj2ZI/uRFc1fbPHMkWM
jdG530oaXjRLS7rbvGU0jHqR1RTztTIDaXCROdEKLoiZu6sEQCklQBbjKnY0OGizTDMZJbOx++Oh
iZueCPreAe72CZqIivnEM+kCLgGBxopnkcU3sG1zVUSsfSgUjXUUEmFBWdqSfkbaztYYavsxY65o
rXHXEQ3/R+dn2bU3aJOab730L1NCTLC7gy6ljUD/rJsIX1L+9+7FeQ4ceNSGtR1ufz/Tq5HPGjj0
ufAbXRAHYn9BIWxBv2nhWGhHOpMlG5145yfcYtt/JTyKUp9Ov60zuOkR65IKXhiD2CvQBrOENj6Y
LFjHuHXl3KvFGwAongMIsAS4LaPY5i+jVmuQFYrs+cr76eUJzbetiJgExeaFW5qnfaXPbWklaFUV
Fqj3yXqYkbJw7N1DdbI3uhymSQy3iJGQQIy4JCKgcSTcMK2tXB1qqNbSUUWLzhHupT5TqJHJGb++
+/o4qWIwXVoD7QvvaUj9Ls/It5TfbIie3N3NIncDzP2vVQjyNBRR4ksZEhndfPZx+5jZemG90Q2k
teeSWm7TM+Lpm2KM/8Wcs0sgOe2fh0dp38iesRPNfFPg8DDUV30nU3qhPdJGLowEoghcib0lvjRV
1dV5oMQ7A96Xt4XjAKPu3dMAGvuq/xn/BBll2QxxR9as4JDUsRMeYrJhSVdO6pyHI6e0D+2jmDlx
VlAw+f1JZu6vp7tHZuaumKaQPvpufpus+SSt6Y9Py7ibfoG+1PFFP3p4qFuCeolYHWEkX5DdaeeP
PlluCvXOO1ShNk6zyjNMTF6jdNadUDMfN8MBDWBqznQQPf9sReFr/dPLdkW/oEcohjIpPz+/1bin
UIY6yVBJZoF0WthgzLIvbHQcnKRFJGUi+b02oTJmhIFNFJtk931mebk/O8SY3JWvXuCF2k4OHoEG
tdAup8D83SCDmPijXe1DLMHDMk9lSNRQIYXfcrcIL4YG4DNItq+/H5Y2iioAZ+5mFDKM3R73wSMU
yCQQhnlYImj8BGN+DzcKEbNRONqcUqQHlr4fOZrgpduxyfvVU6zpXr0tQOYOwtZnIN9Lu4UivBOA
E3HOVq5iiEnvSfdRI/zqtWqasK22yzb0tdFSN4C05QuL+kt6Sxj3ZnhwU6i9ZOwkJMcQKWl7fKpZ
JL3O1Ja02d8VNaCbNoHCkqiaPgCoP0Fqj+aIpkIGfHS1ktqtNhUmyaV9PI5MRG7sTbRjemWtDZtA
zGmBugMymQcAHnoLgu8QmoUfmIcx9am4tevEqlbNufBSNYzWfs6ytq1ioURW9zSLNRAwdmvB4C8d
rE14hZEL9BhdPTiF80HyLfHJGe/g/wRe0Zu7diRE+33fw8BJ3t4VqJlgPXl+y47lueqUPYNY5uQQ
YgTj3YFsng/Q8OOIAKu+gfl+JkemjoUlbh3lyjNM2EmthHmPObOl7oMZpe76GxXYW9xIsaPb8h9C
il5qNKthGw9MbSqRLtqxU2T2gNzpB/UIQxm8xGYp3TDjFIwudja8R+CJ8Ey1Hi1fubrfp5zrANV0
UoOuo7IcXWjL+qVM7tvV1K+3ics5piTEr2Wi/BrnGTijcH+geYj4y/8ltJTH+jwPUHT3m6iEY5vv
kUiUQbDJuvA2zlwx9gKZqIwUE5PLVK1unaPVil7w/R0h3A8Zv+NtsghfkekueeqgYA0UoH9wp+au
042iDCyZKRUysnanU7mklO274T0cw6yBmlq5Y7SaehXBBOo4/xsZHaX/gdrjs/PVrEak5Nn49PVT
0zRWJVXxbaR3stZa5vKI6ge2u6k85qW1JIGxq980tOGwKYd/Ai5qqx4/aqQlZc7lYfeBp7qMTVf7
di251gGwMIo/K42lNWxrPHr4CWQ9qq9C1daPU1t/gnO0p3VRbktvLDadkDhyGeBo1Ni3zE+lC0WE
FGN2/cQ9EVX7Sh72y8iw24/hFB/lyNvnSzfeVhnIst2VzLQIjQreJCNbmvbiPmNpJDDyWdKFaDdq
c/L+3IeQSPR620omfoxksmCnf+etx+Ciduze+YCee+as5G3wUsZORLfIw1wQYE1gqj7o4mJ4sVnP
rLRExyVByAFKM7KPHEWLp+s12tO4y/RtiKMyn/03CjoKRQekLRFe77iunOoPFBfXh9/m35wa/UZA
kg2+hsbws1GEXsfw1H1T9FsBdBs8GFvzGWuw9e4DrE4wibIjEpwi/BrwhHZf0+I/M8NyRr3S/o1o
hOtH4LNQX44uroWMG+A1iigCQhpILLUsQUcM/wt7idKINrU4RqUDQOTlAXJ8kR6qqzDHmgfWNZbw
5GK2aWrEbx19lFFZJy5fTXqv8Jod+DZMh+z0+VOrIJSwa+DBP9gGETVf3VrXEO0jA4a5Ozqsl5CT
ojDFvFupWHvchnLocF4Ol3iTJ3wmu4WwmrZMxKKQWmvYY2ZKwOv/RXTWqP8Kc0LK2aEdZwlN4AAR
jwCVeTUckwMlP7bxmuGNDY2HR4gVGMZcNL1kES82+jB3xq7a4vtzAiAQ/LizJv8jz+74NQ93yDAg
Fepjq4mKADxI05XWbQg96CoWGwCAvlKYACWQg9pNjFX2E6Df9CGPSgm402lr0VVxTF+03XaBEj2X
NjhNP6j0JIe5vMzuNzRVms6DQmFIA3Qq4VpAnaGOweUPOL/AppvbkzlPI1D6sf3DhkWWqhTM7uNd
9TdB2tAXEXd2RpCM3rNKmVLQUi9KWeKrM67tAR2jwmv/piv8l2EjfphIIxdNilTLlcXEosKGo5zr
vcAr+GrlpHkUbr7ziqzRVRonzNo/BOFFmwUo4pEQeuzOizhUqPPMxnj2FF1XWBXNwyUKedMFZpJN
/RtMljrVsq2Amm4gvdgTUzittZXWUqjZkNpBZbgG3OXtaA/PJax9QKSaDrohrRIEtqPaWit17o3M
bMSO92y1SQdWxFWGivmSYElWoDuxebg79uvPkU4z23jcYjD3cIPOmMBRQp8zFcNeyPZhWpuT05oV
jLGUfTgzVOTfutF7gqol0ztNWt1LEVPAheXRynJfkPxKWLsz4DQ9Yl6IlqSTlKJ/8qBnuU+9NKaY
Dlre+Q+FOUZoxsf8AV5wQ+g+U4rx0GUVpVr/HMlCi6XzBajZlS3+XKV0OPHM6eWUtAKVQXbzuWy8
yEL3cQVAGXz9fh/L0C6Pb4fSddadoXjIqLPizdAQyWTs/kZ932J8H54N5Es4REFHZa705mt0DzOA
0T7wGHe1k2s2tP/XPT7Yr0mAuqbgm59eyQ13bFnicqKGVOTBcwwIN5RZmcvX+T4l00oM7RZXb0y3
ykLFTooUFQnzePhYhqC5sfPuaTsCDmy785l0VCaLTSOTKae1o4hKjVVDwqAE3bYsANJGRJ/GbQHx
wUc/4yHOab+l1oMJCNAMO3SAtaKkGso1/765vrNV5Wvv68biHdPCIaBHmebc+7DKHfJb65etFiRx
0v+7hBkycyQyfGvmDCFFnduB+O499yRHuUH6ymGpTQAxJ+GtayafqTy1NgssQjc2tv7DNQ2dlgih
sRbZhXlpIod+gELV7ZxewXE6zFCPCk9rX2dvqLZdSMxGlrfO1RhvMvyexvl9LErZwzs7m1v9DljQ
nzaiAgn4eIr3Urg2Ma6iJnKut5GsNVoLi3pT5kNZTOVKESDnp31z8DNfSCLi1Tktm+8KG5ceKblk
O5OYti8D10Xvuz4hP8mBIRyM6ifTNCGXvspkfhbiqqeofKxjQ9vAn8q2WoG2CD24rg3o/K9q+3T2
+/jtg1YC4H4cpe3dGZgNRGPJtRmfBND8yiu6V3680wjaxPkAeGP5+GHByTQLxaQbdOwalpHF81WJ
qZ7qrSmCIBNK1Sq2EdJ5afhWfjOWVcpFsIePoYiak4ZTh8/czMhIFYLACagvA7Ie/KxBAzi04Pik
wIxG4iwqfgcWOv4dG3xjjFNxkEm/ZumKYm2Mku/bZP+LnkGzf1cO+zhLm70KKEfa0jTYOWYrGsEk
2B3LmvQSQAc1JRpHNUKvaUBOla8yxltjuTjq76y+nKg6+Ri/LflyK2V9ADXgl7HErH1PxXh0qcdW
DBiBB+jn+PpJOZIGlbxtl0meR4CsX9W5oz+05o4PjvB+TcmrT+nlRMZQQXiT1qAMWRXVekqIILWz
nnSpWJO8ldhH9V/SOjFmJIUEDwJnhfT7mRB2xsm1cQyqe2HhTvtTach64p/pQnJlQTPq1ILE2Jg2
I4O7HL5Kh+baZ4v9fv5JKOcPTpdA9vOVx/zMMXtRfAnN9jnCH6H/MquAJlIxmI0/DHdt9OORm6Qr
zL7DzZoMyGgubTvtg0+6oz1feRu1N4ytIiUfSisnqqNzB4ctdBqPSxF/5j7I5xda/Ki2IKi5WP0R
+BFZeJ5JaQNCiJP4US8/zorrzOdk3aqIeAONJSt+LatoQ8pElYVYNETZ/Fy29n5JpCFXATuwd6LA
75O9CwupUXM/FGNyLDa/k1blmU46x/O+SBPYkkoZIRyU5ziBm0NZ0Ri3pybsZkv3WdA+OPhrmvJy
TMSTsPAogsFNkAW+9sOXPf9QURyoZtzG9h647ewsr0xpqPeeQpJxb4OsTFScoJaQY0AWOZWm06MG
UFy2/e1ZTDzzVTA4xnqMPMRoYVsley+rIuEKzPTBxy5h+OrrBGnRs1g1Cl2zORJgDnzjMDtD2sje
uKRFlvMxR4JzDgxq3JIw5/eH5xpxjlnivDwzSjzSPEr77ESzNs1VbawrYLwG2Vni7OWCVnI26pBK
y9wejG3XglsBZkQa4fnBbW9M3fFloC2euTK+T/FwoTwSvdmbS1XltbtrWR0BhY/nj8B8Dv6emxCq
koDdgzBx/jy0L/kX7zLpE0c/dCb73T/x/CYWAdlNYT0fE3feHRUVhLPe0CypNTna3JZ/28ZmUL4j
ql7WCfNzS+dPObp09KJAmVHR1DFIddbx7CAOQ1AN06ysK8is7RFUfB9GM/KAysVStJvMC7K1Tq6c
8z+wa5/ovqxQGKnYpNlETrHFTnd8tqxZ/iSOTV/yvQXLpJ2Zps0VCTw17L3UOVZwbVdMgeVU7kLc
f2zSav6aQ/PuZIY4zy1dNLnIVBaGTwAcfgVbD3/3mXkoVEqcJQXnXRCPZpBTuwuP6NJiq9qR0fyA
3OwvfndF393dW0jbRgvIWHxs2Syci46GCaZqJUz1Lm3QFMXQSshr+ltoaLTw7g89dkdaJFrTADqC
yU+YX0qt0AB9FCqrBUfJ10iHWF+stLLPadujtkPSdQK5O5SHKXHgUq/YIxdWq7/v9Tm50pSMn+dV
jI82Rxc5YDQ1AA+7rch7KOC9n7v2X/I0WcAzT2SD4+k3a7qKHpOtxuhghyFMTbM/y6GlEXjfmVTF
qsCf0a90lxx+eD+oqB+nbu+44KxHNKDljB4IPyl558busoG6sqFrd0nptZssWRiA7NBAkK9FUHBu
XSH+ROckTp7KqjcI7Qv2V/Pxw3VH3mFVmoNsyTz+DlVVkyk1URLyfNnTcuoa4agpxBKdeGo1j1dl
XM7G00Hdy7EU44nEhCOXUsedwf6WXAjvS5nAdmQoPjdo0T2hDB7t4UvLbZd37cXae92oSadi6ipW
iCK0SwaQLjdyNFIjpodVgdoVEVZa9aIX4tiVoB/dw8E7rzj24PMHs62y8eXRg1FLRPUX/tUaz1Zz
u5Mc/IChZshKoW6qTYbhRzTGyDdnG7IN3cxF4atPx6BNToUF0sNO5ZJHwbtRFgH+wTpfRqfFCUmL
gCuxOiHdDMWp49+vc/gRhEKVIooYjzKKGci9HGF3xtKZvUN7U23UDJUtAn2gtcZ8Rc9UaR6X/sT0
+vM15nAxUIIst6YvCuVA5BAxarjHTZJGNJXsvt2ttzMXItAn/7NfmiQJmibYO/ysQHzGEqSUB5ke
PZ3GE9siPl8++hd3tqUgwrNu1bXrbT9o0yR729rWGMF3asXhflacGC+djoUzObdMbwPiIr1fbGh5
9vQMWWQFFthAjZ/zbWdRfkG1zWd3tfQUorHmunzmThTmwLo2k7Yq7POgeXbTp1KXWiOLMMctGYq3
TJDh+qoKXwR8V6f/74jylnI8PDn4QQ7g8rWf1PKfSziLJo8fo1kVpGIrnLy3Ek3i6tWIDSO2pu8R
KEV/Cka3SjjMPm4f5nm2E1o3bzCkhh9d2WR0CXGiRpfEddUmbrhBVkwYbE/CM1jw7V9dAsosTpQD
ujnoHJkwWTluobTQ3iNC3ZKLZ6sl4I3M9FqAHoN2V1H4eNJ3BOG0pRTzqoFa08I7X+Xoua0SlGw+
WbT0p/EEQNSKwrzVnAxFEzeOSJQSguRfw3FFGJ0poB9moLZ6Lewn0ofmGV9RaYXoo1pjQWRKrxQd
FIx7URWxEcxcdYdqx6gmBSQ7CFaicApDiYOcTc/Cihveev1pEgo1rUAZnMKYwRvdGA6f76kZljNc
opkkBcD1C5A/x+cWctqE0tMLdqNtk/FaqkGwGsgEZlXu9gniWVgwr3ndNlXmZxUT21obI7H/5/sL
tGkPGEt/74nZBfKNXQ+VPf8L/AQoK5sL7C3BApizRXFa9cqEg3/kLs7ZkLHxtbxfL332m87RUztz
MjPa2a34Rs220VYHfmMErDgsRyz3DrIRqVz4qfgRwVkmYPWyhK0tuXoZGKA6hVZ8GdnRsxLrR2Mt
kDoHEbXnwRh4ndL2IC27CiPruq47au0yGjR9FnzjqOPiuuhkQiuviIrwTxFspoj4laZtN2mFRAbe
RzHPTU8bwy7WoxNmDw1bigrz5i6AYRIq3GpMmicAy1IGw0Yz9QL6jGCDZIMWXylzDtFHxIC74OIh
R6HXMBUj6q9pOkD85Esux8qCLJ1RNJp5VVnfHcsVfhDCN0TUEfN6VuTZDbUrqxULVkz0Uz6JFNBB
2Td9+cjF0UiEbNKeStJsO6VbkmXeNnlDOamBmsKpceIxEul5pUAICLC+RhYMzHVNNW8iqGreCQrX
5HSYQfVrr+B1GQ8KD6gqcJ5RKpBAdkZ1vGWmPQkHK0xLoL1UgIYesYRnttRfoisCTSKk45AwoPeU
FxLQnTohR7Z1npB2WRzat2bbrQnuC/oWVvIMyCAFS3biJ7p0ZyTKb66YwexsSciXe8wockX4JR6k
D3Lk+D5R+w4G99qoyculH4C3deOEE6eASgwaX23SqqS+RQNql62v6hdagFLqF+RVltzuNUp9aJYs
kfJW/BIiKIbehOJotSNfLGX2DPR8qimtOdTPrbpf4d+Jz7PLKFp19Ajk7OgvzL6qsuZDQsfhuVEV
A2oTfY6n6JsJVsWJ0L9X9mnhims100T01zn9qFlQKGrxSOzxHht/PpGa9r+J8syGUM6WTToUy1Xc
YUDMN5ifCN8oMuXBMp2y1dp+xwQzlxderQjvGB+ibYvdMyMiHck6GCsSMlVZocx9n0YcmWYeRnLz
kBPR62PPLEJQtLEF7lsdSVYHMzkHcQMDnpuD27c+Cs/j43ysSBRByiCkUAchhx/UGAxEHusqgwUn
tKGJ+UpRD3Tj1ADKADPFQjQ4Q+vWP5d3kn8LYEOU5q8yj0KO3S+Ihw5mmb98yQVrzk9QjBqRlO9E
LxW4NiVnPP5eHjWQvPKhUVmXAs5rXGpHXUh0MOO9lggjIHdHEtkKy/ITk2O/j21meqFTq6JsUacB
nk31sUUnY213doCJGPJrLL9vHJ18oaq6SiR+rGAerUJAr0w9utV/hBQady8DG1x1Fd0ndrQU9gv8
CrOAI7cuQAvBSO39eof8dEgv650mFAPiS7njqLkqXFbve9pF5JH5SXSGmgiRc+priRx9PhTRtaO/
Kgwobzu9fznDTuUvWC8BijUEEYyLgZtvE+qf9+U+qmeX3S1EQDZEtTK3XIiBLRUwwho+ZrOkWvoe
dKoKyhFJyNAZvgd7uRVzCeK3w6qd7Ro/1NpxzfYb+jjZxA0SE3JwC3sS6ksYSUHaCd3OhMhbOVkj
HWx0UyLOTqQ35VmCEP5Q/npO4jGaQYov4Bx1KYaN8wlQTxnyexAkOOEsXZ3u4DOfNQaXXOz28yjW
E8MxFKrWISg6x/Mr039tjmRBOx65ld90VONvFZfRsTSJYOzmHa82XnR8U9VThv4YZ7cO4fOvbagd
pPk+VdsBXI1IZ8xulP7YD3JJUpAtkoWBs5yVstvpu0RL1/IhGHXR1abxH52xPIaQtvrPOKsg4C/k
Jvjy+Bnor4F6KGuABsFoTSbdO1g2sT63kq7PnmI0uf7uCtqEzzOz51tGivJh3CK26lZFjlfe3uMx
I3ppZds026Y2nnGX8L418yVw5onkIasxXcAdNslYIkAYdMfQx8wryYEvUKZUcAeuMeeWBtGFYCSN
PbCBIn6/rA0ES1g0+IaGgFpJ5ACuQMYTdFmhfh+mnFKt9jQVP/XuteL+Ce+oFS3MEPErXWAdTOCL
vFqkXhzelaiC/GCmWGsrp8wnMoxhHjx44ef8B3p3w3qZU9X5DjTKYwkHHznSBBQtYLYoaoxTKCR/
qUClS/a01O39uKLn60TIBTA2cAs9FI9xlYNJ/XVFiKzFo1TE5o/sItxEzJGK6y9QMw/Gu5QT6CL0
8qpO5pQHLaXBq+jrAKvTAUhFwcs492IeTqoB5y+fBAxTf2qLuFSbqoefL2t+0tEcsTwfObN+d+HE
Ch0nM1fL30qhJbiRN6CUngdG/WeEkaoGiHvso/3vDZrIDB0zHrbpjUJBxsKeTbbb6Ge0cQnp4q0C
GQhXm6UlYGNOuX8xgur+4NUXnnX7G96XbT4yKvRyAy9mL62IwvQXplvGOQU9PsdBqOIu6IQIpBLT
KONiyWFusQIEaqfULgFdTSNaOfohHG5Fl4+LNcxvA/g72StGevcf2O/r1vKjT+TOBAu4Ett9aWqz
MvYyxpdvscNsIPh/Rho0GEA2LtdKItiUbY0uLr/pEfd4Z+L76/5N6GdE+aw7zoun1n1ZuCgI1mYJ
lz8+kph9A0Bk3SZ4sLfIOrGfYDuzeiR32lFFp/bsfKtFswaIaaeUOD6/JZShPJpqIi2pDQqk0t4a
PpLnaVFgD6Rd0BXX3jbhvpax8syvcMFhcPhbBb295Ok1Kw/zJVrRsqBhqW3CElruyTjc0LyXMQBt
IBj7V3JJRJDbYP71P1FKnd71G38DJGnxl0kKdQfmnb7hEKSUyC2S8QyRZJrw/SHpcju046XJJNXh
yfHCRbRLyTKso0ur9Thj7P/QE9mnr88iGuVywJqzo1lhp+fcqc2XiwxQCMoexJejje2H1s4wSnMc
n3xCzUgIEUEdzET3wLJ3nblgrVDZbzxrjFW9fWHuW5EwkxpIwMN0KCFKnVTCixscm7DNHtjexbgh
CbVk77KcXUyDGGQE1fckhsEWlOs1P/0filt/dSRYakcsI2pKAqQ34cI8d7c3k4Zya428BSa9Uxff
MvgvFeyw9F7Z1SXbGB+l8ypfcYZtE61tf/6meGjTSPjwYQgvQYqfEPGQG+R2W46oss9v8R0YPWHi
z+8lXBEYXFfzQdHlmkhobzEi4zIwxKUK5LqGp59yMTQ+/kiZqiwtzlfcWm2/Eqc39U7M+grcl4t9
bsuY7QYBK8K1CbiBiORYbh5gJIoo3EM4MEj6W2jvJISn8YpBm6h03lc7pt2cPnfmq8U/scBhT05K
XeFUDBmuIOVnepWVz3AIma82+F4T7aibYuaGh5t/PXlZXLxcxNyr1jAwG6jnXXsxPC2mmCG3gl9n
X9ZeFDvBYrvNtWP1985U1k3jqScBohR7L3ogHrbmiska+0sJempJYTakpkMXGpd+mSy+cZqrbL5F
DCaETX60tMyjlPNrfudQ06N/0HpRnj1WuMVrczc+asfAoFBg3zuvqfkvF8XcV1YaYKm8aEthGSFu
DQeVmcSYkmkwO0fOm6ft43XDX7MrdFxP8aOSey1ESbE8pWYgCM7GcKf1NKa7oWiPAJov8ehHKlD2
oX/kpq3G0VhjugRSr2JYQefFFV6Tk8Q+sOV+sVFUC0hrLqMXZP8y1QFjHMt4e6jEMv660JSeaQqR
9NheIPea5mTzp9tBlevXhjMgrk9VmBsS3s3bh85K27qpd3k4tlcRrPZUp1dqicqNE6a4WMXHD+Um
BsXOwlUzVld6J+lpfuezfEyBcLmSZc+lkLX9qOwATbFt8uoUOdR4djQlrvkKg5Ap1hZveImlaPyP
XsHwH0hDoKfGjMVyzDrBU6VOefMCCMhjMObRCC+prkR/LulharNCS4XVvUFCS//GQ4ah3ioloW6M
xaXkryGuW7gbsPWvA7E3LqqYNE9jJhP2FKVxO2C35Wqla0/Z19zCvyIGQVEBPl0HItHEvtrVBzh7
emts88J7XQ4KWfFTbaNDZ1TW6rwdqXh0iisBwxHeRp5ECAFxCTqM+L5/dico3hkovHP6xGQYIO3P
Yq5wwZXbbLzJselJIS+JbYrhmLV3+8ULwTCUADoAfbKeTDOLfKi8wtDHmRM/zpYqt5fpHLxZl7RU
vswNHBvqG4V4JnwCoStitoY0hZEgAdvwpWayqdYED/WnIskgp8+sVz1l92rtn1y9MBAbCm6u+sJX
+1+LrJYeKANEs0tmpqzVGTzkUp2jnxjMfzfcnrPA/ajXEnG+/1zpmtCwb3aKe+qC1VvfRqBEtVQp
kSkHHKybnmJRvZ0x08UvY1D07EJ0iM/jgYvibfMopyGcn1RsVycJTc7nHfIDpcw5BoOtrpBwBkXf
FJvf9fLH0meRIMqhuRiNn+9ZAdq8fOf9oNUOmMpvQ0IGuav/HHXTCYk0imdxKuNfy7ax7cCk4dpN
+jBXV3uJqi7hjLqsBo5stHUVbtTImYzyYuucf3lQ/kYwQTvcbi+Witahmugdceen5J4FTROfVzSk
8s6waBNowzbvPBMXx1VW6MHIBcb+NBTh1fMJ//EQaYH/Fh3uqVaJdmng55+ZXP95bGko78xmSB7H
/1yjMonr/1X4ONAXmzh5iCFSZO8XfR5ToG20pO6+Jxrz6LjInI/NUn+kmCY/7sOhQ8ZDRxqzJWGv
7ZAs2abY+Dhhn0EV0z0P5SbYX4n0z3sfHejFzInJYriSyxX2Flo9CX6cEhhpE+kvP+OqQOTJOxLM
xIGqfjLjQwjiOBx5bdvaaBS8HXFOFDYNe1t4/7NZ9uCJ64kenaxadT0IQJ2YWx5hT0dUFH4KSaqd
k5J07NfECv9TDQdpe4mMpW+20x7bs7aBtnl1XLsrqyinMejVNQ94EY/uAIX2KcxRkhhNHfl9FJec
AwQmiRx31/ztcA8mRwc12LH5NYeP2eAmg2VKx2T8ROoZ6vkzO7vnJ+8SOqzFiqnbrIk01TcmAcv2
QLh26lmI+id4ycr8xa032cZkdxR40L3nOSh1iaWsaydZ72NtHJiMCEwIJP2Sl9P5fkj1f3Uprtrr
Hfz2aCMIgCAlhq657rzAaxhl0Q+O50KPZyZz1y5/sPxQMHQ2MIVNA4oThrFXPrrbgCbGXsCbx8Yd
lzcFim1BQ5ZC5rou2CL7FUct41As9kSheOg/qLjlizxhhpaZX1DeJO6mY0p/qXA0q1u/pGQZtKeW
hvAnJIhAHCcR8WY7TuDKQ4wfwWWvq2Pr5j+XcVAmKYD071ZEfJojMNiSzo9arhMkTI/W6JLdFYU7
57T+BbQvyTwSl0EO0zOAPk/Wz688XTtZ1qxeQRRu/3aGF1XzRBveqeeRj+P1NeBURgVetQctQYhz
KmJS6SphxuAg9J6cWsB2FNeU839Aqhto0Lle3RBiqTO92IUt2tixe4KEcQgg/77EbRbUq0y4gIw7
x95ivuf6cFOFVk3Qcht6LNPpU3fxC19k8OD9UAYTi7eXO14vKKy5ORrHHgzaDY7iD/LguWMlSZl/
ShIvCpwa6GrzavdWr5Cnj0quhrnzNqSg1E/mP+Y5uq0V7cbKUDASHpCezmRCyJ4uALxRfBS3UjmJ
UyaaB33+0OFHYk4Xt8hzd1Chp7xUA+r+zzoANtcNPZY1RTGcEdy5MLfu9xNU0QyUM+0ycYDJEToV
Y3iw+wv5ht5dEno7SAuR30/6nlgMjkJmYhj0fkgSOHLFimAFbIBUn22o3jeZ8Zprp/D4XloGfNiI
gu/x7fmKxMhVvzEVgdxDLbPGSgzZYhs54H2jQgP5z+TJqRHZdBru4nCpnwyrRD1nyhnHl5SZsHKH
7/gQC4OjyoLWoKV7dw8Q7uuhVnI4g2vDoCBICjdp4QLqnerDwf5GAu5mK2Pb0iKXhmQq4PM9sCPd
smdZGY2+rOPPpzOGzQk61xkG5zftC+np0jVYyhq2kmylNcfo1MXzrdj67zswBIfwgWgXGOmaoq8j
pbKG/nJZKWWnye7/QPjwYbgASdalRXLib29LHu+QybVETqy7zaOdUyHUXgVjW6n87Wap8ahjGxNJ
T5hbo6zH/MEn0CEQlRZSXj3LQ1H7+LDi9VPtJsVU/JGvobgJ0WHQS2QAFbB1RmkuHE5Lmzs1knQA
BG9tbTCZOhX6t1nEtoCPfImEJ7it/8hsVGEzkay9fRb8rboj7MEuKpoa8hcdZPmvViMeGNAxTHv3
oPOc+xOoKsKDEJCL+Xhl/C1Dtj258rF9XJ8l0ptofmHincHjIwaaaO+2aGOwGqDSEHLobWTlacjY
JUAc77viYXSnowEw7nScbddXky1wNuxrELNjLj84jh+Ld/N/qzR75PQ657YL1pj2v6s9xXpy4MS1
rHDfVazXf3iUNVVz9TKctKXR3P4X7YaZdRtyPehxcMhsygZDKdomJd0jtGlYXCUFzA8Mg3jVgIcn
Zt6fQUjSIcBYP2qDi8HVqukoBz7o/PWBYS7K5DsnZ0cLfyamIPk/ceFS817M1EOrfI9ESBjUKQcc
NzYuYBvznx1GKKyLIFCxvtwNz33iyuiTH7gdv0nZZC6EIb86AOrqpvwWvkq4fZ9WZJRWq+kIx6aY
Es7qssaAVJ8Fwakdebg7P8m0nraltin33OVKaNOOgXrZFbqtt4EdUaygD0StH6miqXyzlPO4zZT3
0Pd3ZZ8l0TcmMxCRUQJKhqtsgWyWdYKbhQwSZimJZK1RpvkhSRq9p9auyCs5eFvnyiYjOXhvkCrV
FbHEmypPIBtIrOnkXY2xFl1jZJILrxO4zGOQPgxj/x+aQn75h8OP4oIiZO03FGk9Ks5JX7l+JcDg
FeQEa8ITW55imSdjnvZkWs4LkXgsFrKSXHfnSW4eCu6kEpljW3KqA739l4ereTblWrxqyewL2FOF
ncboa/QEo3hzUY7+jZNyNPSOwvS6VlB30s4Qb/DPBbJZjVHsIP4xjlGPJ0GdAn90VhrqALAa0pg5
EDlZG3r3tXAtf2dxMdbBfi036hx7ZQLRjf8hWD3wdEV+hevIr4OAvqJ0ERbKEwmyaLOy8ofRkALo
dv4y0Cg2VCeYI/c6ktmD5WBHCQe0PGh2G7oJ0UCIjITj4gDj4plxjkadehRU5t4btEXmaVf+bvgq
o2u65t1/BMBfcMbsCaUrDkLXJHaFc+kMgiXvGAT4B7VbwzeFW6b/D6GXijEx/RbWcMiX9m3hV6RH
MI5x9BZguL25FWwCInk9S5yhySb+NMUEbOtl6zOgwXcvGEDfdD61NgqL26uPHhAro+D3uB0yCJNP
I8UA1FKgR2O+QMChhd6GDQYn8LHlbejmNaRUTMyrCnA0/z9FTIlazp665MnbWrO9nKZWcN7A0ZOm
8xcssHfaivxnDEIMHUs5VTOcrRwFFqwWJ/5dmtETl51PJMZSeYNvwksMT5wXo/oRrr44HEh8FflY
S+MTd6BmWSLSW00+L6BG2sD0X3NvhqDT2dejgp1gvpK0wHoxJresanDfi8esAENBSVj5IemMaBBr
wY4j4gKMQ69mMs+1EK3cUn6DYbcoMPC4OXKN3BfkQOi+5VEWS96nkGf5MbY7ZOgfQCo0QIHG8kCy
2CO0hJ2j8i5AfwCxkEX9rgDON4hgSmdGvp/AsCtJizTPxPBJGmFRqYeG18cSdFJZTJiGEAGrSS7S
ERZdAaiL1DblUg5A3089OroVlsOt67EXHL0o3k7xgnlC/l5hY7NyDKsONOi3wLiKGlQWAusRWO7a
b5wgR/exJp/B5qAGHG2Zq3+j5FLSApjTBaUwn+THuZAQh4a6Pa903oE3vBxZFPmuLwuT9d/4zVqk
g0n0cOWDhjQvBUJ+D37W+7ct2baPfkXQCvxM+YpsnZVQaRNiJVE8zApNikr7E7Do3T6/9Yav00xT
G+N1JRdCeSLuxqW7YRdXpsj8Iwd35vvTATvcxrnqn3SBK3clbqbqWqndHno0l8fBLqKimjRAMeIV
iUzyMtmwlYFYZV+CyaUQTFBT+8kc8x6zldt3gIdMkskMJI5pSUbEg0EQBgHwmatJwkUhKKcFUO8q
1Mj+vN2LFaTsfBX5Sq6oYctrKHQlcasKc2m/howCJdKcAF79ttBCHmAdiT3Qu8UdKY16bnkZkUhd
dopWb1q3/+kYzhMLrZC3c5MkB4WF//DpVzFR+ITIJNVeEVNKdn6DNYqQlJEjliIpOQ5fi7DV39LF
WQiyER9b23ax7M/1Yh9neSB3mreqwoSulMcRNuS+hH/I3Vakw+pYMc5PBqcubn2+DBwFeDrXxuvM
Kco3cuh8XUCmfN69UVZGiOA949jJXAw2KP3xFzlSvdr4T1aKJNfGv9Tf5PbfohRABzgGITf4lwuj
QfMfG0iUVnz7FnKvfulPpSgRTDwwtyvubMP1OjT9W45d0u9VfxJ5tkAzT4nJF+uQP3coeIpUZ2To
JALv9Ii1tJ1BpN7C5xMBFi4STBlUnFQhBh3WKxsmk+PXB+SuSUufCozqEo8g8IEsIQSgzWdcaik2
w3t6WyipUcZP6Zi8qWBnwpJbiWDJln7ImtC3DmpOGoP5WHYQXH7tE4/XN5xoTC8P4j7x830+yifk
LqJFVF9ZqhH+ORKAWA8Ywy+etwZ3eqDwKB3we5lH3a7Q2YhB76rxkki/pbTiMX6vtMP5rdqOlrjx
dCX0EcScZPlO0uByuPa9ygnJxTwGf4FXGMRlSFN14ESdm3zKVdZ7aXCbdXY2mP6cymlUP/BCXfjJ
W+ZY2gDEjeKBBkYnp/jU+RoWoZWZ3LlIc+NqRzZffl1VkCsJx5ez/Fv+goO6n/hlCGqZfF3ZP/L0
OmYxi4itNhN6uLhjvDPhFkReqo1lPf26tqiCddK1vnOB1wgPPVA6TKCV0+Yt8WNbpHGWPhuFrLf9
fLAPuxvxO7yb6ko2d0fw9mZ5rvBnsVv1fIPDPnE8tX2HdaQP7xTsFIgbvk9oWkqTafz+EehtDLKL
f39gCtBvMO4cGICcYMypZngQq6UQEI9Mao+sf8fZiClEEUSayF8M572JMcR5tX15H/QhmLHkCq9l
gssoj2RD5urm2MlVvIqr0FlD0ffgOt74eAk5RXOkwqRJj+35zrzVupvtWAUa88wWeLDz/WYTqA6Z
EPnkOpgftHll8jk55syXXevr9EB9qqfT0OqDkRxVOWahqZuuCmrIOYUiiqd/2G8WHgEF5GsVTWU+
V9cRCPQDpaS3S9JmtbKkMC6JjCXW7cBx6puNpr92gJHR0FdhDCpprXod+cGrwhscHr+iGUhFbxQJ
tMDaRIjt9l3YFk4AeuxgHltWIDxMdF2zfDmdr5hkXgZwkNEV0ppBrhQIHIBmOVBr27+Zjfi9vobO
G65miu5kmaqLO3ryStK1oPfNAw5d+6lxyi5z+SKgTulJHH1nA8tkQ50CNe+6dWyzvCX7IxUCToP7
6MmatbCmc/IlwSP8taueMANazfzrvi2ngN4DQaXUPUvwRQp9TWFxJX3rEy8Npnww9eDf4pI5PvvX
qO7y/6amvYfgR9L7Pjei5KxHIfaZFTF2SxYA5TpgZgGd0rluPTi+SRfrNrMo0PfxRwd+i+dWQ0Br
bdDe3MQyEpvP7MdeC4KMWqZldzhFa/eGXYfDHiWO6qThS7oa/m4mu6qDmkjsrc8U/Zz2j4tP+1ii
EAQH5R1qYc34uZ+UGfHLH0XcKahXbyLK08i7mCRepxYOSatTCCho8mbwXmfOF9LbwooUZGQYS0/y
r4USA1E70kNxthVlgm5R53kCWWhH4itUESjqlklWW7+S05+SmtjBBQe4s+5K9WTuC1rxJ6GXbwxn
qvImINF9BCsWzooj7Dnveb7+bBy4IkXC6+svf63RC0+bVn8cwXctuzblw6NA69OxXy6qj3vRUVK9
ZgIOsWPhd+EC+wY80ifXoZofMLItvCfq3CpW0VdFair3hixZ/O4w7PL5jljO/XMhSGjAYszKIe6J
Pa9043pqs0GEzK7TjXs4IxFwsZGyUH+FbPglIR9zytEvVNxkT6DB2i1jRH6wkcL1YkfPjiOp2S5b
PbA4BCXqZylF/dOHJYCxSeRwXvzkwj86kEtV7/oBEG2WPbI/9zinGrRnw1fnbBdkmdVQLDNdk+cX
ARse9XKgp8EiWFr8mXJn90D+0LYdKBTo4PwRHI+s2pTqQD2LtV7Eg3jvt+jqagLyhMqhns4SntYK
4t6sTc0AOs5d3mgMmO8lwCbVx2S7Zv6O4mmWBJoXqNhiOcnV5jmiobwvHT7ilBec361riaOWt/rt
u3LjI+ZohKnNFaPK/RqFz6jCBeNHJRrwJa0y6QRijqAaOQ61AN6Lfx6Wk03qJRDT3BGML/u9/5qT
mzhgL30/GWF46cBBwN0mXFCxjbNh5vUJATehuLhh5U/eR/H7t8Ms906hGbukVyYonaenyhss6pPB
rLPH6tUwqczAQudaPiZXvVNVeJROV9ehig2nS8C3hgFYPc2WThMaeKxrfmpTeQ6LeCFMIdT9N3Kh
XQAW3PKwTAgJ//voj6khgy1Yph1iBnbxrC8HD4Owrg392c+RKqIHcq41bA9Oh/dXOso7fbUz3jEG
CUn9KHBgDygHzOWW3QDgaI1NXoDJ1BqZEzuDu/TJ/6pkfaWTv9zxgCUepy+IFpn/a/+ONR5i/67G
KjvHX0f9fkrQyKN6u3wghI1xvZ2wxYwqSRqqzQe9JMFeaXedRc4DdR183LcpYX0h4Xdgi7WH3JeQ
EAP1J5D7nwAXdu7IpqJ/0o6m41ukx9D1EAwVGNQVnhgTUa7N1h4ZyCk/nCqlddR9yHOOMs+Ph7L2
yDG2wB9PQW1SuuVAplIIVovgs8vcGLKNS/6lg7GbpRXOg3ULSFbUbcRKsBxxYbQsRSuiNGdUH6io
cXgLg12/pHOLAz4XNlMP8yIHhYkm+WcIzxAijPaLRmT1eGbbsP3SYpiLMio/O4c6SVhK1HIwiS+j
GRD5XygvTiTwAymE3/qKmBVbPon5Wnt7DOGDIjrE3uNHLaE88fPvylBo2mNdJZw2x96P9Gn36fVP
rpfld/kbVz26wy+UqHyDszBgc5L+3BEUX+V8WciLheQ5dRGJDi4FOhrrsBqJSU1694s/0ZEcwEbn
o9XgJOBbSLbhzqDCkiJR5aobA79D+HcegNVG+byXgkPVmbDtRmmb9O8lTBdVM9cKcHZx7pEQXwLM
AdJ4vgo0Ge9s7Bac2fz1ZQUROBHj3vGbQW4JcZLf5vCfL1Gl1vn/f9IMHdMl1sPH37ECQvkE0ajg
tsX16e3er44mdPoxamPOJeMqMGUFcwltQ53LOhHygwholjU2eFwZMm3Ta2C4hzZ64hhOIjZFevkw
lAz4YTpx4ayYksd1W6169EQURH0xFEaV5HjSgZWiesOY92Shu9HSZUIGNrBxvs4cuDJDWnJWgY3x
2rQ8t0UrTcQHPOE+t9i2sgmihrE91rj3kRnyjMG9PRylGQkzR/NBrC5N1MzKB88Gum1rhimXx8Hz
09uDo2cJyVFLsqXzZQp9idx3dLCmIvbKO/gpiXemOR8w9TADQBrTv0FMzpJIruOBmTbhg1CQ1spP
BU/U5AfQF93BtDHHbHq/Tz/ftl53ZrLQOHHnCbL2lV1KB+8eVZHt9adpKQPupXTYogY69Eg5BMEv
x6hT2bpe5HXlCfkjaaWYOMq3L6r2+3hcnlEE9L8UKkc+tf6LST7oqgXYzO9b9+MfxLlTtLqb8+4p
mu1LvmlXq+VC+AwY7UYFSQFfgfyBZYqdIDL8W/Rjq+1HVCJH1OR2zwjMDG5LfS510v7QT9z7FVRx
1nN3b0aRp7kN9cfEwp0h6VAGT72mhxwio1yiz5bioWGgGdrNofQ3WCcooO5OnqPzmlDNcoKPyiAW
AcdJNzQ8kckUDKvZGh4MVJthJoOGUZ3BsMvJk5aAxCp1TRFtJ7I4dOjRE4LDV5Hd1tl47McWh/SB
fvqBwP4X9SSwvEkl8fbq3DnvuXEHwYxLahiVUJTM5H9nY0rwXmS+RdfAiEZIYhW7cFkd8wTwJfX2
NDCXNdjjF9acYbcaB3UrekbonIm2zi2N646nj6FLl+zhMmBqPuXZBGiHAgOSH3mnl0zFJq8IOOz1
OyFXl9fIjaJdeXjc17yIX55PfVwN3CKFBXSM1KDJ1CDxww+cbWg0SeWYJwAUlL4tzyTYnokAM/uo
hmT6wXCgzFH4WOn2N9jFb2cab/CkTcmZt0KMjaEwvpwH35bw4/hNp4qIJoCPLLUWDRnLhIlMEuRo
hOhbh2j+7tiGIyf8ZeYzPY25G9xFxihQSYhauayv6WaE56Twk4C0jCtp62oB++GJYu9rJlWefYNv
YnH+wJ+KQWj0iEHNB0JDMWERRb2QCA4dzZ5RGUMifDga8Ayu+3mOMWL2Lya+BK0iC6L2qdgPv9sc
zPU//J8KYMCOzEAv346JbkS1q/FC9dFsYhoTb1ynysMcGnhbBBNy43uR5Jq+cAqfZvPkPTe8L44q
1mEBM53dLJc1otY11zi1qSSzyDDoGLLONB1z5LgP8GV1A6iJe0zOOW0irTjdgWPLMdI/28lbaNzG
EtJn5/pwVzSvl6OZYjERmrj5cQJNUtRcQmFAlmIQB4hVKBaf2jAcFqiEWzzXu3g1RduMUIW+n+1/
dn1Dh4cbf2mGXovOHLJ4vv4z2NCHk3ipC7tlZqFF2N6ZJKDW0Q+UT0Ua2HtqR53YsEn4CwS3JYRH
qZFKGVaZbUQ1WfJa6ILaEfzvx0aMHbHkRBxlWaFSdxUz7uTFrGLcyZVCmvixpwBi2xd9G9zSzuCe
RdckIlNvGbKNXZS5GeFi3NTg3ModUU2l1m6iC0WuRvM+2/jVtcFxYO2P1PHqP9MVCDzKFHjned4w
r2Mnot+WlgYsrOj9QhyXTo+QATnp7hvddkt2SPnDcqai4ybps9RxRMLnQg1eowB4z2V0m8+3DFk4
uSCP2wLVS8RUjXJoPQzlj2iK/VfFTPAUQlu4CY8j9k6nxgwQvJy+4v58jx42pKleGb1lOluWLVNf
orlrbz4Ur//TboeGhrtp1chSxmVoLxDe1E/ViM2+Mt72n8t7dNsYPA9hQExtHegKX5nu2b0TLWe1
UJLfeYZUG+iJeP2reK45ch1x7NyrJNLYX02yZRMQexL/ZxPv2zSRtmW8vCF7MI5TvzcVwKSFnAyt
pwUAMTm65/AaE6t0gOyJ3txmJvRlfPKLF9KqcM74R5xXMB/XFekJW0QIBt8Q1mXz8Aajrp5AlmZs
ippzVFVvlnJEKwDSh1dCtt95CDhpSjUvUIlGQaCag4MGHotexEyLffgthasYnGQKPwr5ELpwPZpS
/ZmSJWBoZorAssKz0JsrsyNiFjrWXkeHtWvzs9T4Tp6APS9156TuYzwwk93dXEYIzIexpA9wpNak
c/RykvbW2l8C+LimytrtilvfN+k99Ma3j7er18XAKkZFEaYq6tuS9ay2HAT6rUl3iuf7aqhw0Bst
/yXw2savP2Fhy2chz88n3N8tb+4YB/r7zCwWI8jPe+FAzLLzqpXgwRIbK/osaoFgPc/u3Qft2qy9
0+oawXqaDNF3aEsvM0nrLs7Xj+J3onLHGeSYb2gmIp449ODZaaejWNHM8THnFjgSR3tSITAooC6T
PuIW+0gXHyp+V4O4/M8aujpxoliLkhba7ILfu7bES0dcfwty03wHaRoVX1IQmtAVBXhr02NjODuF
gZlYWf2hV494eLCT/1v8XCqo39WLRJLWZ4jl2W3MeWvSUP2TAW5yHACeUms1okUf+lE8Ttq4uFgj
6ld+N5Ifo39rHsqY+/R3CsJMWgyXG+AINb4Av07uh6XoJOnIHL49nUZ61wg8Nu/p7Lq4D+omrfOM
9GMlo0ZhTisa3PL3hogkQSPYp6b0CZwCrwv/lhMiG/MQ3+FJGomq6c9UQWXUrPtZz22NH2wk06Qv
4DOi+lR/ZTwkielgTwdzbtTex122CznuXINMpuAQC142DyNiMbwrLoJm+ec9Fnc0jBLu2Ndp5YjI
CFak+TkZlF6y5KQYSJzcq4LUMkDKE2wLSf/wcFaz+RsHc53erne4kN/RvCGndfl7FKwtvVonxON1
Px4rP8GQ+lWclBkT9tOdaZgSsSw10iQUNXHlTWl7Q7T9KIfhxurmpegtPk73VbdoU8dZKrOgwyuW
RLR8QHey0yoGE4Y96miYRfpsG1HJAzoVTN2Nk8MzmHMaGqSU2kK2X3FM7XoCravIIQlE0Cshudhr
2JmvHzvVlw3HsVxAFa9l0mUfQs4x+m5fkbcEqiy0+5MQxK7zBFOeZV2pjsySl4xPnDnPq50S34Vc
E1UlDgP/f+HuscpaTaZjgTXDGs4/N59fiWzM9I/Q23QKwSRo8HWqNR0pd4HeNSVjmcn1WVm3+cdb
ybx/wSHZs5AccT6WYKnw0kx5tjRRjBEVGy4WXbsloD23bAVdTlil9fG3mdrw/zPNfMPuf6kpDqli
YRoukT4h8o/zSrdjDCBlDp/O8EIOcppTLTbtB7BmSMk7B3Tf92V4zYZ77dunI9QSWZSuZb43GLJL
N0CZTJoq3fo4fjKd00OcFHbaJWi12JYBcWDUsz60edMbFfUQQbjy/L1gHfTnHjIu+H0GyWsVrZF3
whN7+sbrqnYOXC6F9LU0Hf9PUUdFkndu521lBXhaZhveymJF14Q1UjyE1aSC97FxBbieKbL32VPx
//tcTpoDEYnldt4JkCTm9oXXlYxINXLMwT9xjgqfqlHvRcR64X2DW/2Lf7/jttAFPvGxZ4KLLcZA
JVENOSOyHNjHcWPx/IayxAlQNvxCqijp9Pf9R6boglm+IjyYpXyf1R4XJL9La4xeRtpyxeOUqlvP
Bu8mcO6w+54pDkKxxQvX3MqG3yzTfIVQoUM9dDPYYw324JH/7yk+vUM++AKcWHEN20ni1qd3hBbx
xMP6lwPWp1f2Lx0jku+ZglfRIriecOEGxLnmTrNIBDkXwVm28bEVPrqhYiY/0RdPAcBLKS9Magyf
zf5OFr+o7IG4yx4sqCR7//m3/0PwlmM30kmeYqPXtRn4QSd9HoIONVV9w2F/1qQFhfAq4DgLcRR1
VvIxG7BPNFI+usAxQNhtwwMekuja2haJzsLdwur/fn0GMY75pOTzYwZjp/ycExEy7ibJBPvKaZPm
1Ls/atjUpxWrxT4OBT/CiQRd3W5yAYkGS8UV5q4wAGVMD32EAvrpnPZUVTI0XfqmDyAih5Hgel5F
9X9BYdnl+pOcuvCxbRY04O+FHhRR2orVkY2oI7XIFcMV7EtHj7W6TxdxdKOYwGk2brHIMfXjuazR
acilUYX262VHe/SGQhI9r4KcCgsKWktYFSe3ORe0KE7DS/IdzXRFZgcSJRAk7nU7aypXtR6be373
4ldMES6mudvS41DFm10uWGdT6LNpKBUY0TowbjKRp3eNfFH/wewSG7Y9SDNGPUjfun4lzBbwC2ax
HsGXvQB/kp32YwPenJZN4TSjsHXr+0B7F/5mrKtEGPz0/JivzbLEwyospNNbl/O/drgrtIf/elnY
y9wcEpXoQjyCu7bzwbkajCy21jdU9DxFy6aJMKE99gfQqctA5HhgYPKndBjjapJ+VIoFKP2iEzMH
JwrtuAfKr6IUkRYxkk3UKvorj9HMoi7gF2F38sTVm8qbssfIH99aTn336DMXRmYtun6M/oOtcyCY
iwpCgL8uYn+ckEindYj5H37IKs6iQFUOBwsApjm9VCb4j3VqOEkIEjXN2+FFeH+osetyHIOPubfh
W7sRKKOrTPS9SsaYAc7NC0QKevKgbeK60HkqHvvygiVBz8PjS6agBad1Xd4iNLkN6YkcwwrA9qFg
qrYuPm5eqQKE8/oqpf+BjWSlenuAiHDOkvqEHVKn2TycYpfYdlgaCG1qN1yRKo5/1s4q/9q7tbzf
77ZmB9NqMf37QmwGDzrv6kVLZaeYbQWt7BaczdLV/5NFP7kreHSQcPgmKezICieTWJ1oZ9QcWuOE
mRX2LkkYR8Lby61spIvsjUNyZXLrxCFPULjjdcIs7khJj7cBW/9zrf28pSvOV3rlE0cMGRjlPtc0
tSrTHjNQGiV+JfBKimWk28ZMIaL0GPG6zZR5AX7sECaearP628S71BSoaEEnJKnkmTZ+LI7FyEYb
DiUVR3K4SUFxobIRflCPNohIG+rxzYfj2heI2lWVB/btQR6eVWdSn0vW90akOD7DV/b4LFV9kxzz
MXE6bb2Tai4bg4kINF+X3SgKFnRH8FBnAbwz7Xnq6rYXhSjyQCcaDbMKHjWYCn17W8BxpZzRSWOv
yAal83hBxBbCACEaRA6tHYKUTTV+0oJuUqmqPi2oUhyimbBuE56cSU5bM9X+zieb8HGILKgLqICU
gYxQkG6U6reLu0xfxFxuuR1Eh7Ct/KJpfqIDWo7KZyo2d/a704j9TNy1oTqL28qdfwHXr0C5VORz
C0gPPu7D6Ap9vNTgHq1bEK3+bOzt3GviHBjdzBhj+bFUaJuVT4Cp3D9Y0kQaCwjYLYVCwjtuZmBs
rnlgNcGgWYUUugjt3x7UuQW8lBd69Nl65hpYjS6V3IQeifhR6066R7aJ6CksbYyfj9X5jwKNmvnF
vWdYrVuL6yXcDDsvGX1yx2mB2HG9B3wfdEEylsxzyUc4tIeaDvHiVcEpQ/EzcvDIObcL1w7Dddxn
Vl52pSBGPGVD9sowpV5WJExHpSTlO0OLSKkpiXkT6P3fWVY42r7ODiXtd2vRqjmPeBLFE+R3LQo8
TCKid9l83S7idVF0qWPWnpRvNF1mWZ67/nWoIR1d23gPJb1OMdUICRAcFOLGJmK1p6HFeZLv+MOY
4y6H3wMuzOsYXUyS59ho7W/cfjoW2cwaKYB97izHM/KtF8N05ChPUAKFMgiwKgSa4CCZC4s/xFVi
Ak1TYtqK3SxQa0WMMhYijUtngtbLohGkHYMlntxPf4GuLWFJEiw/GA3sBXKrhOiRIm3M8wQEyRYF
A8b3GJ37FD6b6RvYjDh8JH9wBdIvgVrtAI2Jy4lovpFGE6Q0yGkWlF11bUzYaTNJ0DYF9EtImWvk
b+0e+GE4WAzAF8JErPaxXRmHFM7vGEXpcgbFZC8FoGW7X7ND/i/QhSQG8ERbuFRclO/jstDWs3Ez
l0Xzq3emOBFCDa8Ag0tdpFDeECe09Zgutqoh4AlXPSxW53slTO5kpRtgi2h82dLTaAa9uq5jrGS/
zQD6lU5ywpcfAQc0FwzVU5Qb5i2h+2IYvviCsgMdHhPOiBQ+iOh7o4wVuEfB6VcCGWn7XiiejRWF
UCsZjdrdAOhs6TDqJPeFQYmtE315y8cwbNS2cZwt7HGLYWWJwmKjqYNku2rNJQTxdj2VqpW145vq
rWGNSwLvoYBQoNHNyRXdGTmCALftuo9zytXBkYcpsgWl3hwfw8b7pbSXhtohOpOYJQzEyZwQ3Eeu
8nP/wk71/YpX2g0tPE3wI7EOz0Fhtzuqg3+VqovQH9xsg8bKYzv2Sstr6As7ez84tOk+LJg1G0vQ
Drouq2jI11mu9O6fpp7jeIQ9trM0rfSsyrrYohInL8hTkGaArNre9AJOWDws8a9DWKFtjio8vmBk
7Mi7NrU2csJ23xQsOdu0mb7ky3er5cQKQU43JTUR5oP60FLxCycLwBQJk5MRlWx+qbjMSn3gkZom
mDvYjPOiJaFx0cDuhlSVh0hLgEGT95wC1CiZZFfUacfoeJbteVS2ZT4f3bw9XJZeSQDAkb5MPgUh
PQGqHb2tJmgF9uJZZqTyp4nx0UesLcnrLleVWKkeSaPIdNcl7RhxzwmpapXjJo1snVZJKP/v6pxR
9UEnHSlY8ErDeqAlhbZa8jB/pK02z8u2nedVnARS0aa3pJAYMeK7tMbDxVSXJPskK24yitxZp8Xx
BnhH8bjdY8qOz5VLEJTMCH0v55er7wGa6F0CPEGre20dr/hEmKl2tlxO7COj4mZZfR8eENUSVkvS
hlodSZ5zWOUgQTCRfRbbzZK5h34oY1niII/enaIzYNLadDNvLJM97SVbmv1sGv3RslqL2cxKydQ9
Ve1NJUCjy1zNy1gTANDxPVLWRGBxnaRd8TKx6y2l9UhZO1TZSinD7i5q7qlGi8798VDJfV1cj8ss
fkUFvQjeqT3LfJ29aiSCl96b9plo0TjU1QZxLbnXR4+Y1fi4NrwRJPSOtm333YA8CztzGKey3GYB
dRLAYrvW38p7bFFxmWK6R7j1sV6sjlZem+GFlh14CL55sOVRJ1aYC+wHEn/0NsaMlgrVV75ibFY8
keqSJtV4zpzkrip3r7PFMgfohrUhmEaWijJGZ84VuFMbPWBoZqPFRnjXVYR7iqdc8aZA6DuPw4Sn
fr6O5rUQBXnrzrAdVgm2RJ82JTcbDxQhvEYgcwhiNU0pqhS9BzLX56VM5C7EQ7IknPpbEVNxBHAA
IHmDRnE0Ymucnrv9yZ0KvaOv/43bG8J/a68kYVqAyK8sFPPXluPiyvWDKCDevW9MtKUzola6/BiO
96CxJUxVAoaZyXtpzFuQy+bywvXQJvZP63olbctIpyXqh8P0/rVL+gBcV31VekSDcXGjDpan+ddw
/U9xYgHzEOEezoKtF9qblfZI3wKWc2guMsL/GzdwInjdljLoLYTr7Nsdd200LYWa3yb/40v//KNW
nYnH9qLWReq26VzYiCZ3br7aGTOfJrh81rN6p7I5QFUqMPYT0cz20t7EVYpEM48RbAjmYGdQdwl3
t9kDh64tjYYckD8wrXAcUbJlJe9Zs/2X4MBiDn8ZazD7FCXnblbllqJBv4chQcPhF4Za3KTTvC+U
hI3DPFNoTJJp1icWmTnn7bHI7HBL+Q1ct+r4B2GUhZJGuo8uLZp3SY2wmOpfu/SRYQuE0PzlOWRx
y66fAFq57zTQ/jdIygNl2C1/MmrbwwadMjhN7JxKhxDTUZH91k1DUx7tEGrcm/PSrUBpDqhqehvb
ACHEgTZEthNKYloXoGDP3zszmVzf0LwS1MxEEIGX0DT3X3DwNreXcKkvJIeRSi3m6m/9bCDSjyht
h9ZBIxdeXJXZazwz3BK/Du3hP4ag2mfsQr6UteouaEBUD0v7vEDabFKw+ZaxjQ4PYYegYIjrvUJm
XXz63pkoJio3tXFMkTQnviEUPJ1T6Wy4lfyKsTFnN0hBp/C2azZ/wgkYCIqPNqqL5UOBAawKo/Ik
Cnzp+G4GLe+7lGisl6qvXOQnIGyxO+qmc+/zh8SMy21NQrca5TA3aFhg/YNDnhxQB1HrPzMwY+kT
v4BeI0xwKfSyE1TcWqs4UahlKlJxtKZrS6N8kyMm+MCy1dzMUjBDiUIHnLkH4m37KIf4os9W5lYR
Vti9/M4Uprorkhz4jBk8XO6jnNuhqm1ZHbEwu/x73B2dRAJ/uL8UYh2fbH+1dOD963dp2AvuRFqk
mAbT4nernf2OOnt1J4u8s1Kn8FzH8oyeWOKr2jKu13eT5LSN1WeeXDRyzMlyYBs863GjMBCI8lYQ
yh9fAiz45umPPD9Ig5gBpd/0ok60Dl71Q7zFMn0TmJbe86BVyi930kzdLPzhz9f2mPDYOIhkX8ek
zShxRZzAhu7WNxXwpD/nnE1caeMRypOxxIL21eETrQCGgwuwvLF7q8R3M9uyewmNdi0k1v83Vqyb
FeSttFZ8z365MuUarQEm526ajMErko10EZOHZ1qP9pJeVQsF7L36mmsGQ7FEUFwBaEzzk7AoMGtq
A54oArgAlEaT91wk1Z55PEJOdKvjWl27NGQ0KbwwCY4J38dBuGhYOVkAWGdUbhpQ2YwyBN7n+S4B
IKlRpRkWvel2MmPdvrbOALoRpJMUc1Iatvow5sTnwnRgKHyi5a0uK21h8q8/g/J8aSIVpnU6pFOb
ctx4Lh8D7lOUdpbi17SwTy685dHQuqcoF/EzzPPpEzDHdWmn1kbZA0ussFy8s8d5EsJtXAD7QyM4
xWGxZKb1ShAMbgWkYBTWx+DGq6o45thn2CCFzL9pZHvPf/8s7i+ta6+IqHAGsQ/wigZa584B6RJS
lSsTv9jbg5PCxOnC3sJGrtu4BnwGm/diAnYs1MWsGCWKKwLiIjOUXk2epo9zQN7VnwV9a1qwi/aL
QkhJUiMdnFDQgdaaDIOsxg/850NZn/FRXpp71L4N4HYO2U1sP3la4+CTSat+GUHNL7bFnj3zMKqv
5PvNeb7xp44iKUjZrgWIMobtgJS9zeV3tln20fGV6KAzb4zWp1MguMOpEsn/yIJ9gVYCKwH35MgX
2xI90hFoi8VM+GWcig564kbDNMqXcZef/VZGvJEWcY9bhRCHJTShG25ShxHzSQpKeQQrJmamCvoZ
abwi3bYRgtqbuPu5xq2Zes1piMwDyY67gPy2qk+HIVuNGbE2vxWEHFq+0Z+0Tsva8rhN53t3l+yN
6JNg2JMaVroTU1IDwTe35m5wJOEX1WsHwCA1/AmSHLx2n2kq6vq5q/DS2Yxaocb1gkUYjtMZUVPy
Evb3QZtTlzjFYvFiUeABDowJzCg5xAK0zBmET0h65+zndThEdzkqk4IHEtiDfm7PWYhqFgYzvO1R
uqPmzJ+V63rF4x5GaV4udrOazJwhpn3thU20HQOzV9LDKSZPvx0MablcQCKgj+XJ34vE8wNxWERg
kVkwS3RqZDAgP8rwmWW34Qux5iLXTw7mYHs/JsCIfMTFiey3dBdzI9m5VU85lobYwaX/Bj3Xh7tQ
ha4kQxfrNeEIPq3txN5/RcnlhRwMxlPuvKdfYCzdzUIhXqeoUfV+hnzPioh6pQsTsTcU/qdMq2al
x7jVanoDYLJGRXDQ/J9V66wuuursdAqm3VALAFbSu+5UB15HUg82R3GyNT/FsnokeHaRdYGMfCFe
3fL4d7Xjr1Fbf3B5lp6cMDrNhHriyvfo5YOANooqOjqARx9lHJIYM6uRimuuwi8uX6d1P7NftHy2
fvKBOzM4aTIrnjBzKZsxzuJ7ilZTXRPPCRBxFgF9RIyWwnaYluR5TR0d5x/bF7143yGO0qrGpMBq
Jni6w2NNr7A49ZE1zcfMuT5c/9chXHASa7U16JIEVpUku5jJqwN05MsZ766P8bSmY+3+vJDU5DgP
BD+UBAvFE9uFtciWWH78Ac6rRBWJp1vg+3F5ko1fHkooRZG3N6DT3KQb+Do6WpRaEJKMStX+5GAr
+E05VMEfQ8KYuDEx7P/BFYi4iidqcwvNDkwnZYi/M43XHZoWsTa4hr6ERJlAa5KHQKf7XONAN4Qm
cSMm8/Sy2V1LlpjADWz7TG1SvXuUmchvDzkjYd42GeVgy4dLqBxe95EVEOgjsTKRjirETR3q0EXa
wvBVLcSaAN2kJ+sXCdG973Z8vU94dTGYQ432v/aaUdXHpOtCBhIfbDJodGjxp+KEVH9UKc76hcvR
fteaq+SR2Z/GTq9d3fdVaPITySx7dlbCp+QADX/m+qCetruJsuOMKsOpfr0XMR8MneVHrdt8xz6z
41cue7uN+OLQhlaS8bFTl1Z6OVgfc5fJo50m9AIvPJH/pG27f817CUqR0VkWntcEXxi61S1rc1u1
SMyj9zrA+WZsQPiEzRmu8jXopzKJFT4dcdG3bTNA0gpqx5GAi9pOc6JhhymIYDZCAHs7Bt1n8fhN
RyETfNcPU+2twL61P1W30ENXcadGBd4waEUbHdAEn1nsxk+WTR/yZ8YDrIp6ndtUcSijVpsQLhJX
kEgM9ZZvPE69PeBX9iz5CVsSg/nbP+0luDsitRprlxrGIiDZIlBKNeXL3/0TAiFslzIO1Kn+DCFX
ZFZQ0k/5aT2+Y5pFaBk6Un6QrJHI7A==
`pragma protect end_protected
