��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�a�ȝ��M�(�A@�=u�R�%���O0��FW4��y����1�;�g?jT������T�0.���3]�1���h+����s�v�E�|&�3A^״�h�<����;!�^���wiD�n6�&�v#c��*��i{8�T�Np3>2�r������"�I��[�?ϭz8\�v���I#��+بP�̾;�}s��2ѩ�٫��*y������id� �3T�縤��[��Y����ڊ9�ؿsT�Bc=��E����4,WA�P:�l(��Sy2}��G�\Ӫ��ͧP�-�*�$:���fu.M�ay<�I��@VM�`+J�z��k�`��}Pk�r�?ul^A3N�Ð�'��θu�eEZ�ݒ�����"��W���t���>_2��lՙ^idd������Nň/�8��rz��$�n����3Y�Sd����0�/S�D����x,7����lR�h�vj�.�Z�]��#9gd�7X�
��X�UJ]ƛh�`���K�I�-\������:��ʀuFi%�+^6�o �rmi��F�W%������B��nV�p]F_��_=��&f�����ys��eW"fT
��L<�_�sHB����u�3,b��8~�?���쏪*�u�wd���s�eK�J{AG�j�Ly ��g�_V4R|��Ŕ<����B0-��,{E�y��sa��c�����R/��EF��iqq�΅L�% ���܈��+�r帋5m�V���V���{PK����R�fa����u_t��5'���ç,><�ݗ���k�i'�t5�n���Δ�	@Ě����֥�^г	�#�j��y��p��EO�E/ḧ�G�o�U5��U�A��)a4�9�tK_O�>��(�eEl��m
K�"78�߻{�0��C#J�xө��j�e��$���k�I���Hk���2XzO��^��'}��E_,��a��L�Z�}D��!z�\s���0T�O׼c�Ǯj��۟'�9R�z�Tsw���)��1n�Y��09)܌����5��1��"���y ���K����/Zz�8"����);/�)Đ�}{���>�u#� �����V���bª�L�%W���)Y7��nboF���}�B	��X���8����4N烽{�ov�!�.��VhE��JN������&��"������M��s�E�����115:�1nCnf�0%LL�)��|~����6	�ké��̡���H<�XLv0������X��[m��2�P��Y>��M�\�9�f;%�S����]��F��y��)���F�0�6�IOW������:MG�(M�Fd�C���ҌT{�x2k���A����l�
�]�?'��M���!K�y��/�p:�>p��!������l��ie�H8M����I�8���������2ÖH8V	�{8�P8�D����+VϾ�۝Sm���r������;����-��5��Y�=�K⊁�T��ee)��Dy����i~�bO_�!��s�����Y��
�-��>�	�?���~1���4C�5Upv�5_' z��I ��E��Ĳe�A�Ǡ+�����yk~27u@�}a����;����|�x��^ϝ�z���Jq��5CPf�I����MW�y�ϖҦ��׭�ܱD�D9Q��	���\y�%Nf"�o��j��k*ffz�U��ӊ�W֥Ga�����#��yv��l��R�����I]����J������1������a�S�7����F/t
��0p�=�[3ˇ�T}�/Hĩ���L(�յJ��|2̪\-�>���t�>=�۔&������1h]������q��UP�ji��Euw����뀧b�DR�4W�J�Q��;V�o���X4���o�?�����/:������ >[@VrdK��!�՗�E���W��k����_,� ~���|I�=8���n湮�B�I^Ռ�G,�D����{f[�N��b
'�\�l�$�Hl���[�Ԡ �1̅K"�{��I�M_��j(�I,�o�b�l!E�%q
��7V 8=���b�Z%^|nEv䊜�y��9:lDx��z�[�8�i��I<Q�N>~|��D;�/�q�0�]�K �C��A����2��e�Vm;,��ıP��zg �O�FT�ʄ���#�}޾J�א�7EV
%��7�څ�6O$,*6��'����m,ȹFt^?�*�/ٯS�T��kP	ñ�{�)'F�[cy����ʂjZI ���z8|�r)D�ރ��Z�M`����2Ժ�{�x�l%�QXJw�t�߭U�ǂ����BݨE�?+uP����R]�hs$̙}S�9~��b*Dp=��[�{D��O2+��r�X��B.��{p�}.R�#�g����9;��Z��[���u�af�C�ާ�L��E�V�{Z6y�&�Z�Hy%@�4=����F~�����P�-���B�kR��)�V��(�ǀ|B폌Z�a���XH�O�L��I�������v���IB�s�#�E��8�63ͱ���`���r�㧔2�`�$K�dтȏ�!��ψH%VM?����I����$�p	�)*�+�	+�9Nõ^U+Vv�k���C=��y4��T|���t���|� ��f���3��ln����  �POT�?hw��p9'�j<��)�I.�
�ͼq͚�
w?�)49�H�
2�xO�����>k
�;W����;3?�|G(����m�W���#��r)�־��wZ�^�vgk
@��,�	�s�R����S�^i�F����UQ���.��+����X/J��<��`p�L���y~�i���ᓼM2���r����I+��社���eIO�!��\(+�&�>��5T��S���:��`�\����H�� ��`����S-� ��τR�ԋ?FGC��#+���Ȯp�6K�����yV����_���j�q&]��"RN=��b�?�DE��%���`�>�A�k00��h�8���!3<D�R��2��c�[~xz�C��W���0�����&8{勗%��H�m��j�]�"콿��22�q7A�E�X{�����܎6��Z �gMN�&����K7���F@3*�^A�wS�l���v�hav�?��.�f�}����:�e�bg��1ݪA�Y�r�5�_�L�3�]��������V�BR`�
K��47.)�L{����bl�0�H�����z��թ��j�I�a~�M���aD�k�gl�Q�gح_�nL�\�������#�1��A腫Y�^�r�B�`&��v�������C�\5"?�����H5���	m(��"�8K�n�$���C��q����b�pb�Z�Y����ʋ���F�xy�&�����%T���:�G	m��O����?]�h�w������8Jz[��1���z���{�w�:����Q��5����ԑ耬��d���S�l�H���gG�@eW�3/�$��n$��x7V�r��я邜ʰ�U�� ��������>;i�pn!��N/��F����q��ڬ�NB������3u�*����)+��p\l�1����Ϩd��Ɠu��}�Y	�69�3uZ�nw���P�Y�<�2�Μ� Nàa���.Nt����e�}ul�s<2E���V��KZ�?�	�)c���ŵ�������8�W��u��T�G�d����g=�I�v�_"�I�`��S�=���~誨�Ɖ;�з�T��%9�F|`���,R*�Ӏ&ȅ���Mѭ<إ�����&Ρ�7�b|>g��p�o�w���X�/��YBo��1���mH�w��!+��̰��=� ߑ�y�4�y�����e��6��d�/��ѴL[G�jwe*=�=;�]�x:�4�������G�l�5ߔ=j����p�@���ɥp��/���4	w��̅�إHm�|Ѹy�H����U��5�U�|��x������.�5����g�m:I2�,�R��~B�����&�����N�Q�ޖ��ئ���fa��c�?��)K����^����dtK,�O�����!���"�-�W�Fv9����rNW��Yq:�{�<��_��/9�BgY������ז����o���*I{~^�����i��>��	hx��{~@c��~��� cKu����C�F���0�~&�/P���_)t� (��B�pȚ�� ����x~טO�fW�o�|�	*!�wu�Ӝ��g���m~O.�]���_�2�{̫��"�h���TX���&f�O��VNf9�O�Fv������<'�{ԋ�nr�(吋g���i&�'ˡ���sD�\dw6�Ǜ@d�*�=�-�������NtM\�`�JݰŰ �7���� �$Q'�i�R�kݽg�J[�N̔6����y����� �F�+-_�K���r��S����&�ae`�m���s�C����P����.��7RIx�E7� YmS|<A�'ϋ�������c��L\��K�y��$+��N��9�,��'��<T�!���6zR�k̉m��.�!wh�La�h�s+d �8�9ג:� ��s�v�-�9'�:�@��N]�z�)p�k0-^��Ċi��5�����S�>fد��K�?���T��Իl��l�qn�ɢ���~v�7Csˣ�-Us�Cv�4�d�L�8!C1��KHc]����MM�������VUD@v�'*9(�l1�[z$��^Ȫ�>����0��Ϥ/�;�̻Y�H5f��$-k�qc���'��*-Ϥ�7 $�A��2��LI�jG��7����|���,]5�i��Ym�m���ꛖܨ�?�< hȻ/�O��P���XXX�/���deT�U��b�n�sѩ��n2��t��&u�#T��� ���^Jj����ȋ�b�8׳�VR2ǎΟ_� ����F!L�V�X�A��;��E� �qf�0+�����Ww0b[��I�SK�S�l����K�u(�;���Uг<�i��|����n�ޜt�}7�����Dk��kЁ��y���&��܅�'����ʗ�&� �3��E(.��������"G��d�%&z�+��o5��f�Z_
��1��"B�m>K�n�
��������A��3�s��~3Z 2q�´B�M�ƞ�2��_�0IR�c�Ѓ�8]>��I���:$�R�/1��5�퓞b�뭳^5�a�O�XzK"N䡖1��~MD���c�ۭ��������͚ �թ۾A�FK�t׉����F}y����D=�J�2:.�k�yW>��2P�2*�H��=;�+�ho�yr���i�")?3� ��7Vػ��28pƃ�s!��)@Y��<������ϕq��ڢ�S�'4�.9��4`�7���1��t�W/s0����-���5�iĺ{c� '����m�+8��g�ia3�B�JWm�Y�k�֎8�� jsB*��U���;8�,�"�%�jR�= ����l���X7a�����d��aǏ�����aE#����u�{��HE���Z�6}h�e�LN���K|���H�4�M��G��U����gb�Ь�5�)p��P�zJo�!V9Hf!��HZ�#X�諯)�t�t	/@n]��b�*#��aM4}���X��h�#���":š�먍Qv��mP�\���v�F�<�j�вE���i��9�2`�i��W�ٿ�.��Η^��p��D��s{���Nc�!K�(�Z�����5Zuw�%�%}_g�'�J�/��M�KLx�	�+���9��6"��wKv����1��c������ݵ���U�cIIj��W\����1��\rp������G�}?����N��vG	:c<����Nt��V���î٩Z�`Z�~�� FY/M[f~Ņ7����\�zp\.I\�f�(!������d �r�]N��J�F��*���de+���õ���'B�x�j�BN<$I��R��t���k�KN��#���	�p�%�0�؅����Kgן��%-�"�;��\�Ҙql�o��{3+/d�yEA"RG�T���P�e{���v#��ȑw�}tr���=Q��B5o40}g
*)��ԅ����fBڊ��"�O��G��r���.��|e��)2�/����\u���`�Vq��K�����I�=�q*�k�]��(��� G@Ʈxܷ����0h�ܗWQħ�cp#�]�j�`hD�"dh��Ka1�i=Ҝ.?�w��|o�_�����c�d��8�Tq��L ��wʻ��|�/�6�A�Z�^pՏ�]��6���#}�\���!��V�, �\�*�V�׸*c0fEޥ��]�I�qA<�n8��Z�x�]|(���@�ul襳Ա!M�MRi$dfl|�o��k�e���0<���t�����I�ҍ��*ȶ��ta������O
��:�ώܒ&φ��<�J?7��C�M��Z+�/�_ܔո���1BJ���^�[�s�3�QO����E_�j%r�ؒɱ/�C�G�ط%���4n~����LSbɆ��y��W��1����2A����0�HX���!��_�X�i/�܅;rJL����ڡt��?hCߞǧh,��s�j������/KE�V�Q�h��g|�}Y��R@� .W'���u_�q��������
�����������y�ˍ�l���3���21Yh���{���=>q�y�
�g3$lx3�%u\�f�s�IU��?|E�C��7�f�a�g��<VM_�!��:�y��F7��_���ڵ�:�`�pO��

�m?x���z/R�l�����ǲEe'�%fWr�|�$|t�Jv�57�L�9^�6��#���ͽ�)魆��k�Jܞ�׭�2�������[ٗD뼽A/�b-�����O�� Y�6�,���GQ�|O5nt�-�_nن��ÈXh�4 �ib�$� ���F��@_�a��8Е�H����!l��i�%uU�;�j�*qs��ȭ��l!6�FC�6c"p�&l*t�Af�b��HJ�@��|�h�@�+

H�D���㙰�w/��0^>LP���O�3N�Y�▫,���w���̐��-�������w�AjJ��,U���{�*C'��e�����(��n�wNT����i5��$�a���âGO�������a�7�ߤ����Bh�L��$��?��&z�H�(�o�HO��3��y�o�f���oRJ)�j��S�N;vN˳�J�
� ^���J�[��>�+hA���t��?A��[b����C�516!;�!�E5�멿��$�\���Pр?�$i-����I��%M��[:0��߻ݥ�8���7� ��~}�� ���|�@]a
�6�Ti螷 DWDn_O#�f�(϶�o$�y�̠jB�Rܢ�� hdI(�%�/���z�f��(`J��5��v�L�
����aP���/�F�������U ��jDK�8�]��G���O��A��W�o�6��d�m�-���2��B%����>>�����.�FTo���]+��C�T���T�-�; �	��@��A��Z�W��$ɽ����T���M�^�v��<�KIt������(?�WC��[%�_�(�C�MV�Ih:O9o�+�U����%�r���z���s�i�ß �3��C	/Z�f�x<1���D������c�x �K×P�ΈB>}�cP��0nrNj�'҅�j�B?���F�<ΥS�`��~���y�N?P�܆�Zʲ��\�ʵ����w���(��AP�Q([H�c��O5��ߤL��XnS������)��[��z,	
Ӳ��.�d'��}y!S��3w�.����������8��ف".�����/-|��3���M4���\������}�� �f���EZ9}f�`e�"Zz&P����@���t;{�B�H\�uGi?uF�o.~�&M���1,q����&F�U��z�)~�Y��H�k���j�ۑ���8���o�4��yi�ߑ&D�SC47)�15�l�.����<����-�98kmC��G.k����9���K�FԢ�6��2�d�B�vp�G�+G�u~	#xXe������<�{O��)�}��r#��������%�Brg���[=E��Nug�T��7���^���p��۩�� |�lST䳻�;��5�C�y�40K�U}W]�W����X	>n�\����Yz�w�b�Gi�ZS�nW���^�Ta$�N���Ry�\��dQ!&�y��t�\��aa�_ysέ�3_���&+���e~E�4�Ҁ�T�;���Kw��w��h_�RuE.E���Ř�9��W��6�'}����u���\���~� �"��6EZ+������vXN��@Y��*�!(-*#L�O=����[����B4R-��]2xbv']˛��� w�NdHK�F�Dg����!�9)��$N	�Eʮ�9N:��Ϫ��~=��o�*z�3�쫺��~RY܌Z&Hƾ;�A��k	h���Y��N�+Y�Ł�w" �8����_�;Q�;>D�-;�������zq��0iD��"/���q��A�?�� ���I��m��Q>��v
I<zr��ni�.���I�fQuS2�W�$g�K�O���u-�pO0�s�Z���רm��!�ڿn�I�?�Yʘ�HO��,ޮϙ��k���#6 �ú�io��C�<���H���)qed�_$��.��U� 3���%�+8��c�/,g����ݬ�aM.�{�Sr����<&�'Yv�����
���+Wy�H�s���b'i<�4���?Q��AWȌ�.)F5��bp�a Қ� �����D	��;"/�0ZG͈����-��O�"�e���(o
��8ƷJk���S�Z��>�Z}Qs����)�^��?��,ם�y0:Z��c�����s�º�q� �n�j�"�nL�;�a����S��G�] Gj߿*��8������)��%��Y��%�ێf�>#:*�9����Q�����>~Z����b�	ѡ��M�c'�f��`�Y����	B~���{B`�-�0��m�Y��e2�:tx��k�N_D��htss�	��E1�ǃ�~FC�
s�U�Lsu)I�T�=���2��8����D��N̟�G�'Im���>@~�0���B�bmJsTX�j��!�#6j���x�7i��b"kN�f�FGx�|4˘���&�c��Uad����1�����q�����O��R,�(R�Ծ�	����8gh2Q΅)A���/�O�f�\q�p�T|6�.�p�#b�B�h�xYX�x�=tLx?���v�Lp�(��@rv?�żOp��������Le���m��4�%�z�"�
�y�%�ma:�L};��BFJqп� ���nFxe�zC�<��4	|��Q�m�>�}�q�˩�}�q�'������_��6C׀��.��aH-W�[��k`��{\���K/2��s�����$���V+�Je�5�)��x�,���9A�6z.�}�~g���z��5�C�s�mj�c��V�����<4�{'�5�EI|/�ѝq�n�m��"`F6�f�M�F���1�I<t���Tm��D�׼$`l5L!P8Q�M��{�*��V��V�u�;y��>O�]ζ᧥D�g��������uS9�3&�{9�ՍuN�6ŷ��Ϊ1��rC�e�@��+&9�`/��	n{,��J�<�1e�!�jS0c֚b�����>Έ��ag��Ԭ=O�5*���D��`���S%��Qi9Xآ�ш�e�;ܽ���E�����fF���O�A�"�؋���.��|��)�rhg��C��M삦 �̣��@�1-C�	��i�@���u]Yc݈N��a���O���A���s,���l�b��~k������?������Q��S�,.�BK��� ��И� .D!er;[1<)F�p�tp7��Q�.�.)5���p�I~�\fq��������. �lf��QԦ�����kB{�!��PR���e|��9�o���]ot
�h����n#Cj�5r�G<Y̑�zr{,�?<F�>�A���/��$���9��$:Q��`�?����߂̙�~�B�˾]`H1(d+��U/��LeY��^ �Z�}���6z8�l��]q���`(U�W�������.p�h�XJ�朼`�
=�,j����Y��Rql��ī�t���|�Ҡ� �d�lZ2)�`S��Gi�-���H�����I!�g�ԌRy���-��R���Tw`wy
�NH�f�h��az��HǫsW�!��@]���=��/���X�q�L�L�>J�pe�O�3D���QSź��?�@Sa�,�8��'�ޗ�	�$��M_y��:��i�"x
�\�b��Rz��Ic�D[�ύ����(��<{ ��8S���+�ԥ��-����V���<5U0uVp۳x��1DZ���T�
���m7eƂ��F�xA�Gd�8AMc;v�+�sb�H^��q�Q��ǥ8=L,�O�ʧ_���i+�-9Q̢zZ��<���~�%�� ���qY9V��w�ۍ��0��K9Tw��Ig�d/��,A��X�P�$ ��F7yz�4�:�a��7�����j.���1L��G1�9U�GZFy���ì���fO3�ƘT��|䷋g�e)t�:)�AV� L˨���Oz������#�X)�^ٴd8+� ��GY4�G�L��o<]P;��2.���Ջ�"���&��qq/���������9��wUmI�T)7c�V�h�;Z,�DDĬ~��E��m��_B��b�;�(�����"Ă]�m���\�����V�� ���)�|�*��$j��ʂI/����j���d�f��[���ds$a����~��$�&�u�����Ό7���ᗄ�J}vX��s5��ލ��eE��Z�5�$�����7<^��K������Ȫ3-m�1���Mv��s�#z8P~�3�"Sk\3 ���w�}�.q��G�	���-��$)�7��n�H.H%�Iﶦ��R&��d�q�\
� �`�25&�"em �߂����;�d}=�X����f:�)$������]���J焍��ھ��$��0m�\�>-r� ����Wwt��?d�?�Ls��ɪK��|)�g�����>G���T}{�dtE ؁H��<�5'�}�� T��C1˔�� yNY{�b��%|<���b���C��]]�T��p-����,2��$�����.E��0s �_�G�g���>
��[�0`B���aM�M�����J��q�B:H�;��X�2*��`azg<��Sق����}����[rk�c������m��C� �$ä���p��dΡ�ny��L�ו���7N:5���Ľ���/S/�����N�ZA7c�V#U��f�{nr���_�?|�BB܀0�p��0v��O=z;��^+��»��P�(6ߘ��"�@zㇼ���Gy��w?�L���X"���f>�:�G&Һ=��-�u�Dm%�h��zb8^7��C>��g�&g��g"ϒ↶�Ŏ�;��౑��9��Oׄ�!�����@�	���0�����ʕ�'�s��m���͓��Ih����~׳�?\zV����-I��U(���%Y��|Wy�&��[��\����PdV|C�2໼��������Ѹ�B/;�v6j̷��:��8tѯ*�E� ^�"�g!�A�n�
u�W��K�舽.�R�\��]Oנ%HI���]�
c[/ia&f��/�����C�K������
�rN/rhy�W�j�4�H_�͹�&���
g��_=L�o��@�o���K��A4d�
ڷ[�54�]��*�zu2��-V8F,�Ug/���!g�eȕ�%;�<[UM�/%�c��O���B�JE(X10{�5e3<�8������&L�>9[ �*�8������h�g��@(��V��*�( g2��sÝGY��f���"Ŀň���.�=|�nla����3�5b"��'ũ��re�:|N���r�.zFf���gl�.sEUw��왿��>!=��,��@�'� 2�S� �?"��s��"�=(^���{5aD3�|�Bʻҕ�qX%�@K����!Q~wQ���`!z�P�%���l�풸gZ.#�V�œ����U�[�E��u�D���hM
!�p�f>�h��e���tOp�#�������c�� ]�b]��x+����K��-0/8n3f��Z��;^g��!��B���x~��Jy��L����Ġ��c�L9�3�r�"��+�(d��w��B�H⛰��%iҜ�W�{�&\���N-A3�!��g�����@�DGLU⾦#3o5ܳ'7]�y�ml�$ͼ��%���!%�:`/7�i����!�����Z11"�Lmn���0#��Y��S#�'��j��2�� �Oh����S�'���ssH��Ş�\r��	�q!W�k�@K�D��s;.�lx��&yϒ<M�d�����k֟1�cV�nkI�`Y����-���t�d���e�'^���F�E��5V�����|V�E�g�LPx��>����zuk���Y�VL�dt�j�4��iN���>4y��@D�)�l�s�tD��9LcO�5*�� 6M�M��3Ɏ0"���.������of}�T<�_�ܥ�o��
�K2���$!oڮs���|a*z+�ޏ�?仳m����2Y(���q��5�%(�.CH0��FοRp7�Y6��C��(��?5����[bj �\�?V�P�iIG�0���@��tok�����*���.�YEW�����r�2��e%h���.�x����!�x��Fs�!�9��@>���^����Oǝ��qF�5�<�u:9Sȋ>�U�@��\q%1���@H�� p�c8�/�d�:�_�ar;
8��έB#���S�1��UQL/�X�b��ymA��<tcViu��S��b^�-��Eᘆ�Y�θ�z���|���uB��w���N�m��q�*�J�yT�Eä��!F����7Ic�b��c�g�`7�%���Kt�5* =&�`�q���oڷ$H6�ԯGףMn�O�˜����V\>��C��6SJ x�4n�|Z�U���R�e��D�ɤ>)�j\:K^�u�=��*v��ZWmAl@K2a���2��5+���s�6_��ᄥ(<�Z)���@E���x^�j����a��`��i�'�J�C������.���(r���O���@�b�~h�����F�ޔ	u��w.�1����=��*�#���d,m"���C;u��Rn�K��YBm��p���i#�`���>�s��R�x>�V=U?}�E�9��?Ԩ�i�wߵ�r�΄bZI�|�����fh���Mh�]���܁�UaI�C?'l�l��5���TaT���>��JX��g>$F��Ɂ�2�~��V;�ֽB�&�u��^nI�l�b�Ҥ�\Z��X�0f��o�]?�I�����x*0�$ZQ̂lU�<ɴ�;ϙUz���<����:Iщ�Q�gZyaYp�"�!�h��@�\��k���(9#�y8nޜKL#F+g�	��k���j���:�☞p��Z�,i���hs�k�^[ӵLK����C�S�CBiG�j���|�0�v߯q��ߍ��7��<�*�/{��ZƤ��[A�IU�}�b�_��њ��]LW-oa}�����2SD��W��2��=�o����]��[p�;&)&�>g���h+�۠f��Xt5ٶZ��dl>�d'�碀�U���;���MO4� ᆩj�!
!(�_�gC�m�qx�Kf=f���X;�����R�h�tYcq^<j_��~Вl�����O8f���*1&~P�<f�o���.�_d=�|����o{���_�VڳwB��o��
�uhg��Ԭ���������ʶ���T�Xn�Z���x��c-�_���޿9j�_*��w�]�\�̔���ӭ�N���|�N����4wb۫���ZX��	��j������Bg.q��/�n�����AF!F�-{��0��WNv�[*��nW�mN������DZݻ�uÌ�!��a�����r������#�Gܗ�%���Ăt�Q�Z6�>XT_m��o��l�pkMm�n� K�q�)O���h+q�ba��x]`���J����ϟ}[v>ʶ��੆u�^m�������A��������h:0L1uMR�26q�i�`��۲08�Q��'��%E��͛t��LMY�}fc��>���/��*�a���v�?,��4I���gD|Rtn1ǩ�o�L'�*m�ȯ�1�!yL�r����S�И\���}"�PgZ>�����-�~��DFrFĵa�����u��kN����ִ��JBKƞ��
Y]9\����TT� 'U�[�� /ldViֺ1�"rvvڶKw�Lq��܏7�h�dӃ�ե�D���a�Y{���10ԇu�ڍ
?�]g��Q�.5��<���� ��c�쏿;t���f|,���p7u�l�m<��@t�I~àtQyKҺ�V��Ue��ҪB'3^9YK�q��z�Oc`7�*S�Ni�h�&�
U.�g��F�� �s`���Gdqf�]����q	���s"W�	ͧ5��a�~��h^�x�s�M5U}�h[�SXV�K�-�^O!y,���/�^y��&�G�G�+��Q�u`ש$ [=omd`5��I������h1DP��@!����v�[�I/~��n=�!��T�����T�vN=b|&��.8�]Q(`� �d���W�Q��� ���n�֑Ĉ�3Ċ���<��G�t��x��1��υ `��x�1�;+z��2��[�,�`2�='�VN�A��\*a�$(���R�����^�Z���w���i����6Z`a���=a��뵕�ݢ2JL����fQl[-��k��L@+��ɭ��ztJ?�r�&T`�g	�7f+��l�y���`��o��l�=B�4�1����4��mY�L`�*E���Y����-�������?(#��w�oL�JJU�aFa{E���;5֡. ��H6�l�㋱�b��pn��V��9%���"��<ڂ�Ҽ"�#�ۡ� ��s\����
�}���p��� �w�
b^^�KdlwD%�]X���!��)q��\��W;_��iu�O�ޣ~�5�h����4	l�!]