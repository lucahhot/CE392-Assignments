��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{j�X.;߅ţ3n��}�K�����in
n�=�߯���[�ѩ�$.�}B$LSH��P�|�Gp�L]�߭A�n��_�KBG�UӁ@�mْ0	���2/��%�&��Ʊ����� zH��@�A��"hܞ��dT*Э���v�0�s)�0o�s3�@fzTa��jw�/�.�Qs5A!��l���D��>�g+#+�4֪_�&�Ϲ<#��vMh���{��~�;P6�M�㺚b�/Y���LLJ-�LM�Sk��8󢳠a���߲�<>ln)� D��|�6�д�H=�w��I˕=g�a�TL��1�˲�?]�	qI�~5�ePL{�]�|���/-(���>��(�ՈD����ԥ���W�UĈ�+7�{t0�_����B zX���w�?��E�����$A�sE�j�h���6$��{�j3y�pX��C�G>W�Y%���O#��8O��ɻE���{�d.䙲��ù>	���ⷌ֬�����1�c�L?��A�&܀�Ə��P��=I�Ksq��ͭ�CD=Ȭq����"	���k`�*��{s;>���Z�3���E���l�amc(Y���#�Eǅ�J���c$\�M�-�.����yi7M8f�_�*�����^!��%��W�t������1�kv��[�L����>{�צ�2���3���h�Q9WղPwK�����F�H-�A���n,��.+�����A��0d@eG
��^bmb��2%������O:w�ߑ���a�':���O9�F���K��P�|d�i�I��ȀǤuH�aܨ�W�>#��9|*$�qL��E/����VL��N�˺�WΫ`.���U*��	1כ��v���_���_�i�DH��2J`����ɫ�����G������tl00�܇ 4x��j��M!��/����~^�VI5Q��,m'z��c�HH���VHԝ6=;=��z�RZ.��~�P�ed�m�c)�n�r�5����֞[_�q�M�}BEV��6b��X8?��(M��b��"���v= �c䢣ܩt��_vC�L����<F��9 *�/,����0d���/@���q���/R�ӥ��_�Y�X��ޥb&j!��.��V�Pޗ����L�YL��>J,?�4�;*�J�C��#�߼L	��\_NL#���������?�P�5V���=�c��h6b���h{?[��<^*���>C'V����g!SXE�ߒ�t���I�+�[�҇��e�m�|�@6>����s�Ƥ�Ǹc-!-V�$��Ȅ2�%H�)����C!致t7�2���r�Tof�'��9gZc�S�8=�25E�(r¦��c�6�[3��uu�G11/h��
�$�6�ٗ�^l��+�0f-����r�"��)a��wm;�y�4��t_��{�H����*}e��Mϒre��3* ���~;帠:��n٢���F�ς60tvE���`l�^�`�U�����do�UR���#�"��U jٯy�h�1e�8���D.ܛH�i
�:ǌ��|��n�3K�hm�I���h���[8�;�ZW+��rjhg��.�a���}����zhf�B�|�"P9�C�������f?(n�"�qV�k= �k_�^�����z�MH0�,���2P��n�G!��4+YQ%���Ȃ����2����	��=%਩#��*�w0���[�� R�9�V��v%Ŧb�#;��W�t�����G�`�b�oa����-{��Σh�A��]����l)Q+m�AՍ�+rkO)�(�b"���k�F�o!����S#>d%�� �o�m�5�p��jΔ$�MXE�Q�w�k� �p���JYBi�<����;�䤭�Bݍ�y&��^z�.�;��\U_]���\nzQ�I!_S[�V��Xj��k��7?�Ӈ�o�+Mm�q��D�g*�+�^Do+x0��`F��c`8b��z�����R��� .�$*-�D�r�6<� ����W�Gm�DB+5��"B���Er#Q *��Ï.�??��6^�BN��6Z�I�\�nn��#@��j��L�(����&�b�M_+�֍U���R^J�3>�I��>����PI� �z٪t����g� PXB���┙\����((��X��R��536w^\�u]��g�A���L��0��� ��[�8@��=Ͷo/�q�v����3v�w�Z��y2�SV� �-&D�����L��%s)��{,�p;�x2��:�m��r����
!n����p$(քJ�<�F�G�9ī �~�[?�̘��a�zrm��h�xu=�5i P��a�"�`��Ҫ�7*��e�Z,�l�X�KԇB������ Aۅ7�p��taH&fH�Y�d�ج��t��Xq��vc9�VH{�W=��ݞy]^/�0U��K�x��\�x5��'#~[����_��N�~��*��y��Vw���M�y�~�d��h�7)��I�K_��M�I��~��:|Y�K��Q�'L`�tt�W�7Y�O
%�� �5ݬl3-^z"qnVO!���n星����i�\d�X���z�Uګ�U�|�H)v,�x��<���� �M�!:W�R1l��k�x�=���!h�W\%o��ǜ�X��)<�I�l<�}^��_ח=�Bf��瀸���[K�5�^ܞ�����P�N$6�N���f�l���4���ݸ�� �2���\9�p����I޺�@q�{j���ښB|��w�k4c��H�y(���X���O�Z�/�Վg!N��v$�A��f�8�����Y�':���+�f��(]�k�A'�B��u3�N��/��\+d�5�(vlf�U�nM�����'S��yH��wlW��b�4pʧ�˾^+���(����Q�Ɗ�Ȩ���M(��O����8n��p���dS���sσ(J+��&�_ͻ.�C}��%zp��&�Aq��n:�dO/�y0��z׌iu!lzFt�G>svB6R��2W��s	G�$u+���,�~�*UMZ�_i�^��9U��[[���@���������
j���I�,�#��"�k?��է0b�x߮P�N�������ބ�V���I�:U��\<"%zTI�.��,h�A����>�<ܸ�X��+F��Ӂ�
Q4_����ĞYVtS� �|��+�9�hFÞ
���S+0���6�e�%�\�+�
rF���t���ש�<5Y,W����y (��;��<�@�6`��B�y���L�lF��%���`m��O!2jy3��LB���}�ǩ���	 �D;�$�}!��/t�c�R�?�S�?������;���d���;b�ަ�� �g��Î�+_A_,F����on�q?p`w]�e`~��m�����G{��80����[-��� �0�f��<�n���|x!��٣m�x�d@@��!���j��M� nL���Q�&��$�-7�٧&����54l�G#��m�i;ګ��[Q�ނO�f;�%Õ*���p���*��0p��.��
���@��-�~�K;�X7.���6~U���i=�&���Gf am�C���T��]�]
�_5�[���^CK+H���RS'o������`�E�6˃��ζ��R�-�{�(�׬oN6���u�4N2�M�K9�-��9ͱ�'��te��~6
_�̒y�$����O�㞟\���HRq^��4��Q�"VI�=�w�&j�{�>�nWBo��^� 3��C�s�Ӄ:|�Nf��~�[���b֑�$y��l̲�Bew����K3��žΤ��1<�t����o�!���{���UA}s�b��Bg��M�-TUδ�O�b�]�v�Z>���D����H��.'ڛ�y��c�r�'@��8�.��AO�2�j^�(�������i�q ��QyNab�i�op����exOaА��s�L��v��x�2���=j�՚�k�xkl����l ��[�/�Ҋ����SB�ݦ���
EZu�����ς�ɸ]:q �/q�!&��#�&2R3/��@&D�~;���R�L�vM
P����f���z���k�����"�u�#]�R�/�u�(+�������;�;:�<��w*
;�N��-NP4d�gt]M��m���̓Jn�Hm�j���sv���Z��80J|�<��L^�%P5\��PMW�E�v�찭�Mڊ��#��G��S��=����Pz�i`b6������� S�>��a�]`�z��L��b�?��a��<��W��/�	/���(�&"@^�С�����d)��=�Yj��A�v�z5ʖ������'
�!�p8Ǵ��6��U���NT�f�����]M׋!�	�S|G����Q>�pOw�/(t�ƜE�{����q �$W��3��3�'�ݮgex��� ��5p�W�ep��36�9����nf|:�J���o� wk��L� ��+��\8��M>n�(ɪ�]P�`9�S�k.��.�1�����7pՊ�G��\�V�訡p)8��Օ��?�Su	7�=���müIq�vG������L@���I��CtkC�-�@�sk��'���<�f�^��v!�_�n�9JU��O��M���Bl�B��=v.��[jl)t��6E�������xyҙ���,�3J�s�1ta<�5a\�"I���6�ɱ!��N�����<NX�W`�
�<oH !����"�+=�����S�?�rڿK-!�;�W��;�kP�A�
�2�p,��SD$����[w�}`�q>�	<��!C�S0�вNׂ`�0���SJ0gg�YL7	�%�lZ�:��W��]m9�e1<��2C.�ە�a�v�ј�O��8��YJM�@~D�+�Z5����3r����/��E��F��r�o�����V����Vges�h��&�M,Y�⺝M)��٨�����A\5��U�i.�@W�F�F .�JK&���=<*��@���һ*�D�.������$oW�䐛�+���eA���4.���Vr��hX����˲�/JLHPy"_D�O��>˔�M#��C�^�U��#.H�-�N�z�h��_�G��C��\ h�i��� ��?�%��[iG��Gc��;��U��r;����x I���g��k�	��$'���Oc�~m7��\��22�����.�NV�4�`��Q-����(��<X�?>��of�L_��uR�.�� ��
G1�[���a��%8��@�ᮁ�6ƞ��oD�m��/UU�Nd�H���/�iv�%4ۨR�Bu�-��	�oZN"���;f�L����!�ĺ�O�:��~J�Pl�.OCީ������q��M��Z���8��G��n�ҪE�I���A�]�6V�Z�m�.^�9Z���9ڿ���`�nR�'�+�R=z���y#��?b4���+`��(!y��ƀ�owc�z,)�22�6d� ?�D���� 2����\S�m�8:&����G��̳\�?����;#�zM�'����wd�~��G)Э��k�|
�*�%AA���,����[V2al�<.$]�e��G�ɫd���������&=�k��.�h2:�E������0�&&�Aea+���Eб�F&������@R<WƢ�(6�z���?z/cJ��;Ɯ�����#��؟�PP��n+'�$� �VK.l�����lT��M�#�"����U�<�^���u�s/ȯJ��=������s~�v����@G|�]�����Tq?��!��!E�6/8rp��"���41�
�d��q8D0/v�0�#l���- |����6	F����Zfl�����&f�9�S ���U��0��s�'_���(�+v���_�E���Nw�=�x�4���,`�(��A8�q�J�a裞�Q&�Ӕ��;d� '���Z���Ƨw��u�q�۟����IM<*�J���e��ְ��ODfǼX<!�
�x"�[���	�&��'A±,Nq�7;�6Y#kZ��I6 �ixة"��b&�k;��$��;�b�C���%.̦AA���V"���ţS��ˆ5A�xZ�^/4�l�>�����h�+_�9ª̠9�G*>�G=p��=iZp/i�~)H��ʊ��� �/�< �Y��[�L��$jw�.�m�t<�Z.1 ��7���v� *i�[qM��&���2�Q4	!0K���{vw�`�P1{�$��٠V��]33�fCJ��4KNUR�j�{}�#�L��YyR&��Np���׻q�PR~�+�;#��b�*��F��|*�^�-#L�� ���2#���9�B�$��Hc�-� 1"v���@+P������3�0| ���4�Z��I�Kp��qf��3\b~7"���Vx�
�en�<Y8�Їq1�х�0�0"5�����2�+�\tD7�m5�O@��C��˷��j��W1��5������F$���{���*l򙵘�(Վ��%z.tJ�6����2"R�ƴ�J���4r�I����6���5A����7��s��-%��՚�9�sb3c.IV�����n��)w(}����������6�y�s��0�A=���i=���"�Y��R�1e51Σ�n�>*�ih���FZ�ɝe��V�a��Z�����t�H�V�'ٽ���@��k�щ����XgF�e��2D7\��4�l�e�!t�j8��)��Ln
�.3b9��x��[c�2g��T�R��5�.V���<�]SAη���g�8�����mű�z�(:�롦�9*Id���mI�g��k�?�^�7�7���Ϩ���Z;����_H�jF	_��>H�|�N~6؁�b�1s%��.9n�V�*�
׵)�'��2fU���_I�<���@]�:��p��m����e���3$*<z�E�0v�(W��yVNk��3��,ִ��	�Q��,`z���|z+5�(��j�1�� R�WP�mܹ�x}j�� H�T��.M���u,3�����D�b���]ޣ��^9;���K���	�Ul�+5�.|+�R�^'����̶������;�+���4���+��h��|��ԋ�(@�C��-���k���8ٗ�����?J��Y�:k����RF���2l��|A^b-��;Zː]UA�R�]j8Χ���� ၜ���I�<p=� W��_�mt��^��Am��:k�`����5��PD���"7�t'mQ�"n w��ӟmEO��)�D����1��A_b�9`Y���<�>
r�Z��/1g��e���9`���yB���&a	��-��Z:���|�j�S3�$J�相L&�%�d�d� ��������Z��h��_g����-�Nd9�i0Ū�˘����Hk/��F\����P��ޅ�	�n�ݔU_�@7���4�DB�|"�q�\$��Ҩ�A�il�O%H��b\���;�
��oɎvh8I��"���iB#���i2��n�����Z� �x�/�"�V����Q��-�+���e��9���Լ�y柄H��{��ם�P �*�F�ʓ�u v�WR�#_��B���������AR���5�B���
�CT���*��'�D�Onҧ��K��1����:8��_b���"�<B��y�C�%Xi!l�^>�2[| 9r���M��#ݖ���̬�+I�د��Z�?���<�&"�hs���Ʊ��?*�2�[o	���L����Z[
�o�j\�w���"_��p�|t�N�)���}��T%F�6��	`!��;���������qx��i�v�j���N>*[삶�V
	lCu�V�𦠥�
�N�S��-����������M��� ̔;9�&qh�癿�G{����ׁa���V�Y|��e���ֻ�I^���R&�|C���QH��%ǗGrC�A�42)BJG�_R(�1m�_�tM�9���hҠW=�����Sf��	~��̾h����Y�F���DLs��)���hU"�����h�Iۥ�8W7d	s�06ŝ�&~�H�Y��Y-ĺ��KE��B�~{|�O}�������^J`k�uN��{"ӱ�cnܙ n����$)s�v(���:��r�gz�E@�a��i{j�L(T;Գ�k��C��U�Sl�C����Q"L5�q��*(�3%A�*4���QEU�RM�%O�k�����d��ND�õ��U@�������%�����6�dn��-o2�WF��>��m��_���@�=�ΪE�]ݮ>��;��a�%�%�:��j���Zd�����=��Yrv�m�>��Zꭖ��de�,R�}L��j3��	�zoV������C��m��Mt1o8�������IB
NS��>���>j0�5?Խ90���u�m�X'8)�:n�$�\v���;b������H=�@���:Fν�p���I�Pʸp��
~�(XN<?dO�Ⱦ��t�]W&4��1J�⸐eC��(6�#n�Q�c"�n,�"�ݼ[��E��i
WjI�����Z�o�O1�E%�<����(4�F�qY7h^�!d�&C������R�� �~�F>D4n��,c�ƶL�q ���d�T �QU�t��R���I�+t�~�N�Q�^6΀����N��[�W�W��T�ҧ�hҷ�]&�@λ�<�m�d��H��{�F���٢+��MU��T�ڣ	,�I�jgH͈��	�A5�#�p�B)9Q^��R���	K
_*ͺ��9��D��ϸ��_�����VO1u����y_�޻�v(CB��wnQ�e�e�����E\�;�l����ە/<�(��4�9���f�FZ�]ҦVn]�C�յbV$&�6�.�\%���'��G��Vl�tз�lS�uW�]����#��'KkH�Tu�T�Y�0�s�v��c�1�'6C�%��0�: ��}�En.ӎ�a1+��jj�*<Rr��Z\��ka��;�lo���y>�T$d�L�wE{���}�����M�6�)�k?�a�9��zZ��.�R��s<��WaA]���+*�HU��:?�U뿶����v����9}[E�d����WU��	�{8 ]�دRX}^��V�S���t���@ `V��pãv�w�ϢSa���MC����Z/�����E�C���Šޭ76q,�N��-	;�Y��ݾ�C�6;���_tY���8Ū������~%^@���ݥyRr���:z��ݺ�Ө���Z��""�N���E��/��s�Ґ�KF�<����=��Z�����Bl�d݂��ѓ���r�k�6z��ەE
���7Ň�G���<2��6θ)Ui�}�B0�pT�v�ֹz�ΉR�=�䰌zk\����a0�i���`rDu?�eFi��|�w�=.Bb)[&�F��u6֍e��y�f|?��s���#�ކVtQ$�ڔ�u�?��/eH Y����`�V�������Oy�W9|VH�RS!�K�&yi���	��MH��X=P]H�H>o���߲�!��h7��%��;7)��ya�ޝ���ٺ<hS�z��@�:G���-�
_5-��������r�j��G�tTŮrTzJ�����(4����B���(`ǿ������u��:�H��-�K�Ŕ%2��h |�O�~g$M��«��Hw}V.�uC��L�E����e���\-�kL��M� �in�����ŮODl�]���k��TR�b��=�>�	fZU4X���e��!4�n->J%�)r�$ᚗ~����~V�ߜ�G@x��3l��:`�~#iŶ9��b��4����s��a�Iq����Oh�1� �y</ZU��`�8zl��5�g[�����x��z��Ќ��q~�A�Y�F�4k/�Xɼ��qaDV��L�-�� nC;$���ڎI"�~������E�bh:��{�[7��:�̷�P	���?F6�Vd$D��8�N�5�u=&ƨ��x��V �����R����"��9,�cVs�(+v�A�28>B�n��-Y�-uI��,���ī����.a"w&J<M�wV/������(;5��a���j��a�o�S7�{���8����i�?%���a3+���*��&DX��%d�~DC�J��j$�G	l$郻��5&��1HX�e*��]��y�g_օj�&�ҭ�=Ё�t�_������|c?�a�),� ɉ��h��\���f� �$`��*��m
d�)}>���4�Su*#ċ��� ���jv�Q���ɏ}5���a@�j(����,q��孾���W�us½<XA�'�x�$�&gV�I?�%y��
U�V��'��uVi_l�iԧ�T
-S�>�(''�/o���yAߟ΃���Z]�sbgj9�׮޴	�j�� ��Hi|c���z��Y�f�)I�L:�:�._�;&����JT�6��J�E���z�̲�rF�����tK�ڃ$H��������v �~��b��-t��r�c��mD�l����q0�C���F,���4c�Xdh~ú�Y��#�/;a����B�Q�x�����U(��1z	6R9/̇Cp�T��#[�ݒ���w&��V�d4�0���/�}Y76�O��~�U�.V�r@p���T��v��]�c�9ԙҮH-����QK���b��Y"֮dq,h(�B����n���;L��*����?\s�cJ�'���6m"(a�h�3��ޤfl��I
Q�Nd��^��R*�G+���F�I���ł��l=ǟ���U��a|�5_[~0W�6����<[������*:̓$���w����?&�����d�P�%]*��zf��8{�:�
�X��n$��h�Os��Ŕ� }��/�ZZ��1P�2|>ő���&�Vݻ��U��z������m_��K�Y�l<(�'�Uhjr�sK��]�i�R^*����*�3{0���e$h�j����ঙ ��'��s14�Js����)+�kXݒ�#ɾ �Tt�xG��h55��Ɗ�+}�z���Ԉ�%�ډy��O:+	:�a��	��D�r@��5�z�T7\�|Z}�2�ɉ�GQ�������K��`�̺�i�4g�e��u�����k[oqd��Jٌ%�N#3��^�Jy�׎�R��,|�a������=ي�-;����JF^����~�l��Z�@�L��G��Q㵖B�%��@BN6�|xW��p�~ϻ;�2F��m��O�[$���Q�tM]r2�DE���l�0)D�w�$7C�[�S�P ��NR��B$ʲ�fw4�����Ԯ�UξKJמê僝1L����7�BQs�H@�P(3�U�Ƈ���t{�I��X���H Y�n��.�����;ji�Ȩ{� �s��n]�'Ԁ�ї N�_H��D@ݡ�V�$�Wli]��6�Df��V����o澵iY"����BB����#������v�N��Fp]b��}􉼼�G/.��cI*T��B}C,)ǹd��Q�H���{�q���e�����q�?��g3.��BO?U��Ɉ�H���E�h��.�Y�k�,!��m��I]7��6~X�u��|d�� ����7<�Jrp��w�//����7\jb�������opㅞ� U�t��q�"��4\��d��Ql��9_"vY�P�\$�i�P��H��}7H�p��"���ƎXQ�T��cz$�tr��i p�d�:�T�ld� 
:��Pm���d�&�B na���������Lr��IN\�	��X^�ݢ�ܔ�!���x��<C���_�78H���㜓�R� /(��.%Fۍ��������e�"��_�v�9Y�����	QIa�	4Sw�����Q��d꧍���U���(
��-�	6�dG<�? ���,��ʊoՌ,�9�~��2�Uﯘ��)7,rG��.�ڰ�h�#��ޙj�![����7���a{��Z>��/��꙼�MW�1;���J�}	�җ��͊�0��W"-��l�T$:٭��K?���	82�ɋo�f$���#�I�M��Ah��Z]�=@��w�~F&�@x�଱�<冪11����VKx���6L��$.������.:eĢ�0�{V��O���+qcԾ+-���o��h���1}f��0 1"�Д YyGd+���2�	E�ksya�J���!�*!���<�/z�.�G�6`�y�M��O�g�r5ß��t����!&� �F���o}aJtW�!O������n.�9����_|����~����\���_��K�B��FֶCӈy(0���&���(!Zz�4~�����:m2K�l��ζ$��,��Ĺ�iorJ8� �W����j]V�nU��d�zPl���sy�J}K��rYS�&H���D�1@����Bʸ3[�����Ǫ&�=�c%=�Wq��d�#N��C�������χ	����r=�P��"'����K$�άN�(װ�35��Sq� ���?<V/��Z���m�A�fT�{���?���TJ���E-�[����)kSBcg
g�Ύ�/1�8<�X��xC`����2<�Nӂ ���}S�p@%k�6?t\X�h%vQ��"�6�M�\�o�=�%۶��y�=��2���2Qmx�*����qe�\5���g(=�$���P1�o�ă��d�� �̀{�Kh����>�b��-�����$�*�h���뗧}��EF�<fF���9\j����:�IU�����r�n�������X7SOk���S�Fud� . ����c��ǖ�
 �I���S��FUX�r�e�`Fx�T/u�3�Fs)64_2�d�hV�ed��o;�	�\�]���Q��sB��C/����2�EVp����^���
@����pՕ��k����0l�X��=q3�;�(�fIv��W��	�k4
븢-����H=�����Am��G��e%1�z&׹�8��7�(i�=�_��{�Y7�}�B��s��FF�1Y��v��_��1�+*��ˮ쪃 ��z��j��k����;ތ[�rxR�[]�f�ށ���]Wd���/2-���!�G����q�$1lW潥�'�5�^�
�M�s�L{{Ǽ��}�i\j��+�����J�\��.�՟%��]� �=�f�N�����q'pS�*���U%fl$Zv�:f�o'��jʩQ��.a6TC���W�n#��[f8,o/b��o�f�������7]�*[�V>�]�p��g$~~ h:�x��gE��&���`Y眞��n�n3�R}�A�Q���jr6�Pi4��S:�����F_ǐ�a�o�='�=���I�n\�Vsy�:���qw����ƩD'A�	��ܓ�
���>�=���N��D\}���ካ��j��N��=BWDU�(��L{�}�-C�ri�.����;��;�z��ŘLѵ��c�T`/v��jk#m�Ew D=j���}�u�2��
8M����W�5���u��	�g�p�Ar�CRB��J�H�;��~,F��"р?�����a2�e� 'ySn�λ�X�������)���c7)�V�ۦ}�W���d6��4��P�nK�G�/�F�m뀠�Vv)6ã�G�
�-.M��V7���%��xmI��U�F�S�ږʯ��n/��D8´�/��+���X�dA�O�'XA�!8����b���]��Ի�K~�8P�y�#c��>�;%������qmBx��� ����\7|�i(.�N���&E_c�MڬD4Kq�ň/05����)�,���HB7:{B�Jh�^za�_��(��ʌNJ�����-�.0Z�/�N�����Z?�$z��z�|,&`��(p���j��PQ�E.�#CѸ͉rmm�cn�a�"�+�����|_8o�0�̣��� ���~��l���l����D��w)K�z2	\��ՠ���+��<����N���Su>yױ/�i�YXP
���"��k�R=�7^�(��^�a�t���%�e�q�L_��%�eI�H�_��):$�NW��4A�ݓZG?��Db|_3�jqDL1�z��bY�P���p���YKͿ ��o�|k�w��x��FQX�hf���@�T>��Y�C�\ݗ!cM8p_����-��\Q��N9�\�K�.�wD��	4*j���ܒY�@|8�t3��s��/�8L��=ێ�`�=�������o��t�|����tm�^�:�d����C�fΰ5U�P�U~9'&Of2_n��}���5�1���ɪ.����|JY��^B��,g�d'�ݟ�_���k;��gP]�OՂ�g�(�_��A��� �!Ev��;g�v��>O��ί�]Ulh�ysZ]�-��2@3�E��	��it�u�ا����P�
5M��q�T)�zRs����:]k�����X� ���=�ݹ���^)�󯧊ntv�4$�5��L	\�{!Ġ�B���S�x���6A[K�h�\HMd����c.�g�=��y��DN~7�/Zk��KF�<��ȞU� ��/�E�����:��Ēv�8�䤪�8�l#��f����������4�"�&c�[J�a�}	d�*�'_*��/��>y�Ml9I���#�<tҨ��,�m�� �z�\���x3[�ڟGR/�ܲ܇;Hln��\�`;G�0��/s�GQ@rib�����V,��3SߧM�~��*4T��'�O�Iq��kā_P�p�C��	�Q��ɅU���=��4�7� ���V`�jj���� hb~m6	�Էsr��8�,w���Sz�KKK6�ʌt�^�����Ea�
�G��Y@!�{8t!By�p]E��OTrF���6$;��:�wA�8LR�;H->�b�8�Y���ǵ@��jq����b�4���k<oNA��2f��O�������"�7B��*9uWo�G���%6�����g�b/!��-o�SI�ϰ��p^9��Ga�+����~N����SE�%����i�{ex�P�����	d?��� t#�Q5��5y�#��Ș4�����ii8�ó�[�ùl��d��?�~Ew���Ϙ HC��E����L̜��J�}pI�r76Q�9fp9�CK���O��� D�<,)����c�Ι�[���a���x�G��0"��	Mz���ܮ�!Ët
/�� �Z5���D�JA�p���k:��b�?�� �4��d-=t�w��2!�����_��5��+�}�J�S�&�(��F��g'B�A�C	$�9>bj��\\*�niڇXXy�����jc�=?�0�������:p$��\)V��K^��� ��X�=W��D�W�Y���נW3�#=b
��t��N�ھ�A��[%��(�q$>Aȥ���\Hl3�����J� ^���I�� ��1z���{ �,�$��DHOϣ�� m��e*��`��\�{t��P�$\I#�0��fp��Lo%`����=����5�)��� �c��"O�C�O��>�I��j��v���l��"&!/�{�+F�D#L���D��}!�Μ�!KC C@�K(�ȱ��F�{��8�y�sʓ��r+}�E�Ǯ��W4�����
y
�q�y��������[lJ*UԽ��/��%����o�?�]�3y��x��$���� F�y���I�z=���0u�l<R���q�q�(�889
��]J4�`*CE4Pi�Ǧ���?]�z�E�x�E�2v ���1�t0�/�ij���$���@P'э�'�$$n��o���h �-�5��HCK�H!f�	�|u���7���	�����\�=�#�"di
��$�-G�m8�lQ��x������8%-V/���ru.Ѓ4q��x��n�:Sg�	튘O;�k!)-�b�I��Κ�"P�@����,j�P�V־��V�����͔|s��EF�hO�5W��2��y¶2���yKtӵu8�e���p1�ф=*�G��-`�3��6��~|2���>��0�q��M�;���(�Y/��m�<��J�Tjc+]�"��$:&wT'���L�r�P��/�Qhm�R:u�ԴӨ���^���ɬ�/�����n��P��g��`�/U(���qS��z���9 XC�㐛o��,���̫��2*��T�`$Y䨳�Cv��4;2,�|m�E�c��w�%�VC�������A@ٶ ���蹴���x��x~!ot� w�&�#�������U��)]�cBďk�ܡ�+�-ۯ�b^�:��i ��g���_!���=�7(ګG��Df��*�k��jy�j���="�?#ar(�4��7c�K��r�=�RH���Q����Q{����|oe��Z�����r�di�$�=T nY�P���x'�'6}�孅R��tu�(G�H�2���h���yY�܏����v-��s�/��:�����`���˳U��>�{� - � ��(��ա�������R�Ɩ�m��s���H}�7]D����т�+�5�| R��\�.q������|�c� N��hh�"����X1V�7%���ޤY�G��Lб%������I�C+���\O4�R�3���"���^���dk�D�� u�E�թ����D��gz'j݂"�T��<ـ�*�*��<~���
:ޚ9N��_�P��5��9�x��}A!�hX̪oS�����>�r���}�+��C��|D�����hh�5X9��ڦ]��n�����V�5�)tǢB>=�i�}Uk#�l��?�4e�
�:�#.1)VE�Kγ����7��|vwXI~XNT�����V������D�����- �DNa��:Aϲ4Mik�" �M��g���Xejr��5�)&��Ѯ4���B�x�����H�X��
�5�=�Vm{�8T�>�)Xe;��<Ri��t�bGz��:���V�{�@�2�=�6��nō��8[�Z��3l�Sx��3�|�VJc%2��(}�	�d_K	�>ٛ2�����x͊ݮ���[֕�U�O�c ����k�֙	����x�e��_��*k�@�D��hk��ժ���yX��QD���T�lKi�]��0�Ӫ2�GT!��V�?�B�*�=���8�nK���GV'�<���eP��\pu_H�JMV���n��ꥇ��ଏ��b���	H>UAݷ��Y_����;K��w���@���W�~Cj����2�J���7(}��Zp�9!iT��K�ǅ!v�K�Ea���l\IQ1�*|��r ���%�^\�A}� �6�vŠ@�b1�W~6Q�[�ѹf댣�R�@���� �+_��۱��2mXv�@δ�����Y��MNЂ
���)��*)s�Q��z������"�Q|�T�[7��o��*���r�\)�*F�f�p�0����g 8��֢O�a'�� �v�b�����L
�O7��1Uh���=Dё_}*��F�do�O�Hv�wWI���p���9�7Jv��z=l�ĸ���$�
�[�ɚ�����A�C'#h0��`K�լU2�r�g�7�l��h��̷tA��.�}�J|	���STؠ�u�W�����!�F8*�`���\��R����%�Y��(2km㰲��8p@u	A��d�
]��0��i��_븤>�Lj8�sJ�߰��M�w����t>��o75�v��@/k�h��*Tap�͉�( � %Z~��jD�E4�{>�q���cd���g6���\G���K����7�Yn����IQ�!���[�2(�5[ن��ƈ})/�Y��e��#�~��+���F(`��f���������_��Ob�����2������
ЃΘ��"h
�QN��[���{��w�������t�����ogǳ�>�peC����RDBo�p������} �%k{�:"5 �c��T�Ws���KX�V��y�?�WU	�ɀ�4�WqN4c]3��1|�y���/�j�۴D�P�z���=ҋ\�;o��R�a�������T�pg���b�����9sEL�"p�-?N��|��Zr��{G]Y�����N+CA*ᡔ��%����M�H��el��s��y"n�d��44�G>udHB��ƾ�y�\���:�� T��7����D��/���H�k����ɮk�	�.A�]��ʀ���(�AihRA�4 ��������η
���Mp�z5A&�׺���|X���(iD���>���K��V����W�#y[�l'�,(�;F$p�"}7�ί��9���O��ǧ][�kb�k9���=k�wQ�s��X�4�����q-ᑣoa�� <�����C ��m�$��5�)�<g���DcO�}�ϑ)�H�i�F�1)9�]˷��+D�C5�B}҄(�k[��~�"��50�Gy�ǻ��K|D>&��K��5X��:{Rg\� N`�z���7���,���S�(���D�MsUsdp�q��EY����ӼRj��ZG������b��~��yI�i)l s��In�J��R�w�;� �!��J����9�j�_���$�cI8�7 �~G��4ip�F77���T��VbZ��� ����,�l��x��4võvñ�;|�f�r���~:}7I�	�������n�P�Ϩä����S��3�P�dCcǗ�q>���EV�Ϝ4�F�=��cpۉ�Uw F���;r�{]-yT��ko�u����B�Y$c�2ڢ�#��":�d�9\�m�����GVV_����P-�S�mĽ�\����l�/�IT�`�}]�ל��UFM�?������3dS3�S�"s�jg@�]:������5�u�B`5�?�,��_�*�|���X`��1���,�Ɔ.��Qۃ�Z?ׁ����&P~Ch�H�*	���}��k>�VK�/C%�J㈃P_�����C�Į�m-�%��l� ���1�=�Il�ഹ��[��&�=�~6>h��<q�ܽ$�;��б���}��PI2��`�*���?&���`�#��E<<�/+TYx�����ț�}D��M)k-�?C'm�@�iN���HG�M�1(��4V4I���<��Toܩ��A���1���,k$u`����1܎;��!L�J)��9y�	��
�k}���m]�iL۶�
�P���x2]�0�P-��ύ	�#E������� q2�T�B���_�p�f�����q>#�0�������:X�R���a�J��>��T�E/KM� f~�x뙕�Zq���,��`R�R4�ݬ:�У�W?��恟7�7H�~ՐCR��g�O5 ��Fm+��������mp".Q�{�,f2�,�i���Q胴���V�n��X@C���V2TI,RRNdTq����37v����4�ujߒ�t�5��+�n����X�O�q� ����Sԇ��G��|'�7dJ7_|����~��w1	c���Uߎ�#�����(Q�H���^�WE�w#}qz�/ ��c��b�h��,4��V��4��'�$��k����H�.�����\5V���*�z��֥� ]�?��6֝y-s�Q��b �I�8�P�c��VJ`I��Pz�$�a�E�`���������V2D�<j�W0�A.w�����n�̊���,� :*E;�ns[p��Y�1��JX-Dɝ�n��%�>�	S��~"a����_��vJB�zsR�6���Q�1�UN*M��8���#ƒ�d?����U�WT�}٭����Z5�Nm䊦���t��a<��~L�Cj��6,�f��^��tT�<���~X4�	���#�����P�n�����$I�-*�-�.�cf�O\"��0�	(9�N��^�g9�eI(�[�%�BFӃ����MV�Pk�?55Q�q������eGF�@���k�!����Z�,a @ai�����ӈ r^��}@,	�>��ga�ӑ�rY _�󈌚��r�<z�&ܾS��ixJ@Κ��H9��I�Ś�:y��(���
��<��>� �(;��$������;L4:��ɾ���
Q���� �w��;X���4��Eb�l�xՌ��G�JL��_@�Xa�{:�z�͝�ӖDd��z|R�ү�d{���u������5��n��p�� $p��}�zqi�{����5��<P����!��P~�_�G�Y�x)q��K�Яn��g�M�`.�;CJl��g?�2
"���=%C��W/6ynr�JJ��Z�4J���Ȁ[���k%�D�ض#v 6G�WY.c����'�$��!%�����C� ܽ��Oâ�7�nī��b)��=(� <�)�k�����SE���x�N�L+T
3o.󚓟9�A\���Oe0�p]Q:��?�`An��n�m���s;�oI�9�fp/�7��G���F�y��߿��<(�N���u�/��2���dp���3KCaH�$�Go���L/9]�0�oC�����}��!�<�ޚ�ޯα�b�\�n<[:�Æ�k�S�C�H��YN�G�����Z_Zb���0b[��|c*c �EIEz
س�Rj����:�V�U�D�=ÏJ���k9=K(���ëq�"��l��i��S�ݵ3ّ���BP���BL����gϢ�>���lvcW+j��r�W
ƀw���">�&���hș�)���j]8�(�zd�%C����꤀�	��s�IM�߀�P������;:J-��yV]2*�%�\�	�*�QM08Vly���̶� �.�p��,J>�Y�3�r���6�>wАw)YC3��콈�M�8>������������3�~�m��DV&Ҡ#�����NK^f��Y����PM1F�(����ٖ��`�O�S���_�/��U�Lt��_�
ʖ�c?\�U� �<�!�t7"��K˯�]b�n� �x���g6�_���
;�֤` �e���@��N�����=k���Э��ֹ/��f��wz�oF�%Ei��@Z�JC#��˂���!wo�ئL~D�g��G++Ƃ?��H��o���z�����*E8s�C�M�V�Uf�j�X���9h\wx�lH�,�e6���0�L��Y5�.��e�j��S!�8��w?�j�Zѧt_	Q�h��I�������R%��cT�y��hރo�K��%����i��hd�``i����V�i�DP���qo��8�t�!�|��-�ʰ63Q%�+�ف�P�OP��{��!"�E�_r0�h)�TR'Z�/Tn)�v�wc5�=������αf�M��|�:9)�DU 7����T9�� ���Щ!���f�\\���m���Tec�tfE/��.�t-��/�������i���pi����	��꽮sg��$�)���Qt��)�s�h��T��8�U�E�s%i���R���6�@�P��Q�V����GY9�!���-&��p�=�RtЗM��r�4 �K�^n,�O�&*����\fBR��M���H挈���b�:�(p(���>u�n����K�\�3~�2V�M�%����9i!�SF&�>��Mmt-���J����A���~[3�f��h�Fl>�FJ%M�8��l��Ԗ��M�Q'e�AM���*J��_M�+�D^S�C����=�-?R�&i�nu�q��h�]	�<�"��kv���5#�p����^���Ϸ�m&��p�0��� �^�U)�{̟�2�3��I=;Ij�?�1�Aσ�
c� a��D��r]�a�����
� �̇��a�P(A���(��J�o�?F�j]I%�i�+fV.g]R�k���NG����p�7l�s◃h]5��'��N;�2��u���c5γ��xК�̡A(u��$�-٦�O��)�}�x��c�5C:]�,�9�&��Y�R?��L0쐚o��Kss��c3��˽p>��(|,�=5j<NӦm�h��R�'A|d|�^�	�0���m|�l/)�#*؋~q�>���a��C$�ha٨�3v؂�Y4�~��R��1Wz��=��q��(H��0���W/X$V��}�?LE����-V��$=��w���(C�K��T�2	@����C1���I�w��{���'w�5��D ������x�<q����x;�l�&o��j���n��|��9�X�@G���ճ�2Ge~��n�8��;1KL]Od�A�kҡ�ҥ�R��o@Q��X��+�|M�Y/����Q����)�Ǩ4uz<�l�����p�;k'{w"R��('Ҷ�Y���*HX��j.��ץ�c��SڹnɎ +Ŕ��B��w��22����������4������-n=�1_+�1稉ꁴ��gt�;�ȣ#��T^ũ؆^�B�'e!��mD��YYS����������N���mv���I������\����A[� qN���sS��	�*5w����YU��(0�(� /oYP��Gg�jYG�=)dc�i�b��-�C6�+b,��#�'q*��a�����t]k��4��-]k�'���Ϛە�cF��!c���t~�ըm�� q����]��B;���c�bY�߈����'�%UծNZ��z��y����Ͳ�(t��D��m�@��1=F���][8b�6��.dvn�� ih���+��R��"�g��r�ǭ���p�L	Z���ӎ�}��>^!��<3+�����:�r�;+���Oݍirφ��9�M���$�'B~�rgt�{k���䞵M��ـ���t̚'�o5��&$)�x���ǜg�Ao�E$������h������	�{ٸ�D3��w��f���I7�? ����U+�@�f�5��;��oe�FY�31�#�`{������&kř��ВqŜBhn��1��WC������Id�N��
��}��p���S��Wj�.�/��h�b2n^�%�^[����?��á�z�:�[SDE;^�S��%�w�SY*y-ϼ3,G=�?�Z�	�����U�!�VPk�ck�h���Du��}�yF#�Z)���E"�ۅ/J�3t����~��ȵ;���(�2�}*����`,ŧM{n'� Oo��%�n�.�v��	pg�N~���x�*�O��+��f�I�"����j��f?xY����JZ���eԆ?��\��O\�J.~t�<-�'�$��y�����w|<�����̚^���^�����u��;>�*	ջ-���m������X�a+��T�¾^S���)�!��m�a#`��1m߳gʸN�ߜ�8L��Ai r���~���G�;j���T>��U-�%6�@7��j���O�
�v0?��D80��M�'�t�v����X������4MG,l�(���f�@�1k�C�K|��,�H9�qI�oE���w��c&�8(��:��2�p���f�-��<#b�?'�Nl���C$�e*����%�Q���^�@dn�����D���󗿋�C�4������NQi��d�w㱳�<�M�'F���7k�=�i��5sF�\0R�]ۣ�((\Ǌcrt��M��ӜF*`�B� �g���U�64���
ځ4��F��(�}\w�:fn���-����0K�7V���g@���z���1`���(k������u�Ȼ���x?�q&�4w�I1B�r�LzT3�b����⭱��l� ��?.yÒ˘�Q�>���0�!�"����#d�2Y am�3��¦O\����w�*w{�f�������VA;��^WK���~_�u�4/,Bp�ԧm�^s�7��M��� Y~�ѧ;V �����Y�p	���8���m#���M(*��b�'-��}Э`���*�.Cݮ(�=l<|?�DAs��%cc��F�;-�&eFb�s@�q�sUECE����9���?s����t�+i�zwbؿ8Y���O��
2���'Q��C5.�h���� �GR�@�	��b�*�=V���0��$�/E�h�2�;�!鈆��+#~�0�dp�a�wo��1�,���|�ѽ�,z'T�eN��&��C�l�J�+0�k���&������x��x'�(�t_1�\�~R�#�ݹ��2' ��4K4�Yw�F�,aWo�HX�vė��#�Q-��
+U߁d1��j"��E;�uՃ)쪄��0<�kL�@j�b �!g"}����;�� }���/o���8G�i1����;�PX�`�	}��Xt'[�>��-e��x��cZ-�O<5�
��s�"���P��Er!����Pf՚B��^��-��nL��ݗ�{K�O.�u��}%2��4��3�a+�F%/D���=���P+���]<�P����}&�p�Q\F�����D ���m���V�v�ǳ��"�ݩ��Rt�I���6� ����7
0/ڈ�B��r��yz�Xm����}w���y��^Z�=/bv�ƽ��-K���`P-�����z��)��Y
u
�6/�����&�S�����RKCAڅU���,��'8�r6��sr�g�B��ӛ�Ib��&!��=�b��+cۈ�/w_��(%�!��#�����hz��mD�6�WU{���o���� "H��>PB[`�d��G���gE�]�����+��ρ�:m�.��AU����ھ��xv�c�"�}�����dL�Xߣz��Y&տ>�69�g��_	��o���&�D��K���q��:&�rL�Pq��?��H����Z�[��_�2G��Q*�jt��G�/�AqKt�ϓ�:���C~{�򠉘♟�'?O�����J9(�=�R	0�$�n���K]	��<g	��9ȁ�h�ʙ��,�G�6�����)EA���0֙�#��n�.e��<dQ�lb�����hB����=�
8���ܻ)5���U�O�/�_�����9F�����l��-U��qy悾��Y:i��WDd�үhn���z�߅ELt�ߠY'�b�����rOy��|�E'���$�D3�"��P��몣�N"��nY�ouJ��iu//
]ٽ]�!ĭ��E��D
G*ř�t�����GG�7��Z�'���b����`������茞⯦�N����Y���Т�����~���vT
;������o��?!1��@�eLz��Lz��t��J�qle]�0��������q���|=�M8��GQ3�L
gdq?��S�Aީ��ћ�F���2���e��p�"��;wV�9���7Ynt�/Z��U����M-)������RNa��s��`U���~5a�e�'�s��r[���:�g��s����{,�J�@�ف���8c���1�O-
e7����L�jq���%qx�Ծ0�x�M���1��xS��p�Э�mn?�"&��������}�o�e#*�t_)�^���M��ouA�qâ�v
#*���Ǫ�0��̤�Nf�"�x&7���C���*x�aXp�<��Vlh�3ann㾜��y���́�;���S�hF{-��<�����5��Wy���\�1waƼ����Eo������0cշ�(Uk�8#�\Sm���7�e �K
Fd]dYL��R�4/`g����K�����Nؔ �UxN�#/=4��a�K��x3�uT���ZnN��Yt������m��s�g6^O.�S{�H���,<x!D������������h�l�">)�����􀲹�3�
�"���Q?��o�j��'��/-�buZ�<�;�����+ ;�^R&3�C�iH�3�J�|$�ҿ�e�6>A�s���pe���2��q1�@��=��Bڗ�4�vW���E/٧1*���_B�-ި����S�i��,��Hl�[��t����r���z�$�IFZ��(���ZVfW����i�A����g4e�	R�H���
�j�7�6Mtg�͏U�%#��ƲU%��]�ڄ��.����u�5{�p�o1����Y�.�b�j��].@������V��B��LB�Zq��e���D�2�J`� D���W�?8�א��~2��Y8��e�>��+�	{�P�>�JD|���D<1F=#�6�KXB����3���n���V�>�bA�f��aE��{�U��4�L�+
�H�ʃ���S�}[�t�3`�E�y`�A��Q���#�:�G�Z������j��R3�tRk"��5�q�U���r�'��Na4�g�6����LD�� ���{,��#	�?qK������I� ��o���KC❽�6�(h��հ��ຒ��@�H��#?������եeVRv+��Yl�m�����H�����1Ǿw/��C��alv��)#�g`�-)������N�a��	��{� ���m��ZD�I��j
��7}���An�����9����\�� �!�
�`�7=[<Ff#�!����Dǎ����?��S�=~q���Q��;���$�<x�njˁO<���Q�������D>� i��)�>�$:�򥗧TFLqrOπs8��O���ҏ���<8A�G��Qι�Ma<����"��� "��!Z��Ǩ�+)c
H��V�)b:QU�>�"�.�.�����l�n[~Z<?�J��7Y�����V�<7��S&7�GeF���F����S��[>�?n"P�,�I��%�f��!�R�L#�&�,μ�o���� h�Β��]�MV����m}�iK^�����s4�Q	���Ԏ���o�:X����ͣF�x���L�7� p�-�ews-�����|��B��ctR=��h���}\�V�ӣ����":��W�L�XFp��~�(��ZF�Z `<B =|ib>�������_X���F�%a�P�A�������	Y�w,��&�6��a0�mN�WMY,爗z���,���@�ſ_��/vf��5)���J���C��qS�׊��U9��'��fN6j��ݼ��:�2w*��7�螗
$x�fE��]�@�:@3p麣 ���·M�=	�␔�O��G*p��YK����2F\�p�y����i`��60U2ϱ�s BO�:����K��BbL�����|�Z��(�f1a����w��W�z���(��{�'��V���6H����7�sua��2�?3(<�K�l������G1�nA��># '�Q_)Ɂ�k�fx�ǐ.��g�{h��	��z�V�V����] 눘=�n��ҕ��c���Ћ�;����ޡr�U#�Ԧ�/��<u��Y�c��^K�b-�{��a<9���ao�R��o�4��<S������5��I�ų��Y!�6�v�&�y�vt����H���, ��mŝ�4�}Z-�x��F���h|x՟�.4�Bk�9pxH���h�"*/�s�À���=3#b����B#���[������B�Z�$ �V`�L�Ӣ�6�� _����ț��i�FwO���d&C|�A���:�|0����s�{�K/U݃�R$��ӗ�(���@�[ݓ����*���O�.e9�%�5�&�9�� #6_��_أޚU��2FF��8�-^�.���V+1��{ȟ��u����L�sH��c��vɢ���n���!H�P�FO� �{*�C���d�o|=�q�6!��b��?64����]���YP�r�,̭b���ÝSCp�:����ǩFؙ�X٠���wMt��&������Z7����޵���E,f�0Uo���K�bܸ�;Q?A�k
��ѽS�V��@s��V��]�U`���^�6
a+g�yCB&%��qT�EY0h�k�3)%B���v�W��/��Q�~�
��& Wsa���<qi��VR�Ϳ�.�T�J߷�'�AG��F�E��U���W&K��WP�u�Z��.�^?o�Z�`ۺ���d��eɦ��F躞'Ľ�90:��w���9~ޓ��[q��D�of� )����o�grů�VCO���p��\�#E��<dp�4Pf����֨�b[aܤn�+����*\Aɑ�ix^N�ϯ��)	l���G\|�RC�Bˍ��t�l����k�95	J�8F�E� ����3��Yȹ`������&Z�-��gi��X�EY�-@�T����-ա\���="���#,{4O~�Q��BM��������@������p�μ��S�s���!<��(q�~+�+�O[P���	b���ӯ��)���lw	�6�K:���ְ��.q�GZw
~��ٶ�qd���vG�+t/`u0�轐�Q	ƣ�=��pj��㓚m\ȤN��As�'��
:�����V�tY���������B��,���-���d��D{L§�qr?
����i�"C/C:�x����y�Z�g���{�ܛ&�㨓�!94�k�afOnI�&>aV_�v���z����w���:B���*B�sk�9��jg����=��a�L���2�v
U���QB}�~R6��N��{1<�El���+�;�c%p���F�9^Fy�ҝ$����U"e�,�.e��
)�� �*����6؄2��1>��VVM���ڀkœ���:>�"yx������{�f_����	-�{�o&]��r���E]�����_	@F$��7	=_�p���������Wƚ�p��
�E�n�&L]*�`:ߕ�l��Q�~|d�䜒C:|��>��W���k�)
����E��c��[ӷ�lT!��&���a�_��a�B�!��]G���͎4��ʓ�L��`W�#�{�L �%h깓�IH�)I!"a�==+�a�㍾��/K��3��݉��U�	?�t{��yGj���J����Ktd�뛮�W�A�Ma�O���H ͟H�\�	
�}�@�j��.-�P*ޗ�!�|&����nN��D����t����(���e`9���/4q�S@X��O�ӵ6,%�0���>ڒ"K�]:��T.�:�r�ڱ�a<�>>�u�l%Z��$o~";wAs�6O�v��?��'�N�Ou�G%'4��̣� G����c�j��r���s4�8y���pS��|	&$��!��[@�#�%���|��M��jxŁi&,i(o�vl+ًnъ@�E�Q��zE�b��ĝF��f.�Ga�,�8���ˆNb"X�6x�-/����KPQH��o)���N14�nS�\���2�4fU���ڵ�|,�9�cB�%�h��@�In�h訧�&�e�$�w��t9���3c��s-%Y<�i~m]�<,�f�.�.�9��r��Շk��Ϗ\�� N@E�`L�α�dG��,o~
���%B@��,/;A懂��j�m��s������v��͆�:2�Ĕ��}��ahCD`��q��=���
^�r7ɣu=ѳ]-L���%԰(��Hj��H��ԅ-��oP+T"5f#ƈr�-:T��,B#lM���Fm�y����ke������`�-��ʽl_JR�M ǆA~�����p��P�oyO���H��̢Ě/ԛ��*E��\>����r�������W �a���㿎��%VQ��x���1�(� �$X�F��p!�"��<�*�i�%Z�3��I
BF'�Xi6�j��:�r �D��/���f��et��=2�����DL�,���Ġ���1K�!�x�/is��ŅCC,�	��i��~�|�0�pc��,���8��"������7�n��6��t`��Uq=O��3t�����5���3ìrz�:�ROUt���^�1���gV.��֡�k>�pH ���;0L[ћ���?9��EH����d���?�}��,���S��L3�sC����rs��=��YO�CwP�(����Ϸ�8�1k9V�����ߕ1�5�{W+�տ8��`�����Gę�)A�-٘���;J�[	�s#���nm�,��C�LB�}LU�H�Ɖ|�`�:��gU=�HuȖۼ�y��������)�p��z�Xw���Z�~�nj����T�	(�
�Ji�M���̗�u�@���#�Z���]E>�
BF�BG�m'�.�J��!�7_^k���x���ޅ�g�^��Q�X�3�m��[�<4Ez��~i:לH�%�[6�� hD�U�r�d�We؄��7R%w|��E�0O�p��$�I�ޑ�����^����Q��,��ɛÜ�y5��urY����S�r,�ᮛ�t��`�i��]�˞���!D�~��^��G�Ԟ�)����h��Z�;e�<�ŏ�V�$֜��	�l�L�b���g���v��
Mw���y$��S�sHvp�l.�n�֣2Z�-Y�@�:�o�HI�� ���zN�?�ɴ]���Q����n���M��mE�DbR���� ����D�q���*��]!b�Js�qa�F`fs�"�վ��˨^��?�t,ۍ~�����w�̀R��o�ͨ�Kc�������q�"��F�e��$� �Z��3����i���EQc�[B�"]�"���1�d��_�B�k��(���#2����̌�fa�ub7�\�0�4U�x �PH�>����$=�m��w��d�ɕ� xǐ�Fʽ�~��b*o���IM�u�(�9�XҎ*'j�m��6�(�V���rA?�LE�CHy�{�Q�P �����:d]H&�s� ��(�[��!�"�}����$<��/�AL��nJ��
&m�2'�3>8�&#2�T?�漬t ���`Yw�����+t~�r��FZ�yyPF��d<V� FǪޕQ#��x����Z�.���dp�1])��5�/y��Q�~(�f�ɿd����k\}��!'t �gW�"ˇ��ڡ��.K���V��u��5�M��`&�?s�|�2 ����-Tɬ�R�Y�]�;!o�<���@�J�������Gl<.J<9��1��7 N����C����
�Ց�,��cr@������SZu}�!9�R8�W�-��,2=.��C���ϐf#xg��p���3�Щڪ�E�t��0X��U�܍E��\�.pB���4st�w�w;�:S���-�
^l���O�H��r�I���0���4:��[�4̤JZL�e�.+K��az����XW9����|� �kAhd&rJ�nMS������V����Z��FpC|�n�S���t;4���<A
�^���@4�]����1=�,��r|E��TK�,S����˲�E�:�)H�����#iX�C��터
�����H��x��*�>� CG?�hyD*�s�)�QiO��û/�/P�ÿ�$��}Xn`�Ԓ��aU��0D�V2|9�ز���:�� ����������l��gf�E��_;a����&j@H��E��Ɗ@��ɛ�*��z��͂�,�f��>xS�c������f*�ܜ� ى�̼L�ڶCs�K�u-��F�� �O
87�p�]➈�5�w1�7>K$�9(?3+	��!�m��pbJ	Y�#K��T��N%%��r�yc�ʑ^ޕ0���c��6/�i' 㣪mcU�����]��"�	��F�9���07ڻ�	R��|�v;���T�.gM�D:�S6@`��u�v�H�8��pI�Q=yP��q4�Ӿ�K��M�Ȫ��\�T�d�:@PF���ٺ��'��K��k�A5��9G,w:n�=���@�uS���po�w�K�dW�	�T�+�;��}�I���X 6#4���ql0��i;�G�\�nW�AQ���w�g�W�X7��b���x$����,���z��^%�6����Y��;,P�X�p?m��*EP`@j�´i���-�-���'�����!w�9՘����.�yøU+�H~tG-�
���;��*h?#��OM�ӱ���>K�̄�z�\Dɟi슂$��ޘ\�Y��׎(��6=YK�SEs�𠅳��y��y�O�O�����\�*�B������V2�[7�y^��gh^��5��O�NS���N��0��\nY�����Fy#^���-���O��x#:�,@~�/ХP�Oc!,�2(��<M\3�`۱?c��!��m����v`�!l_DY�cd�e�6la��{��tvJ?��=)-�L�����v⳻���ܭ�Ѿ2 �yv��!0��u'�ks��g�XRd��UDn�sV[&�9 ]s��s�6�[{g��v�n�KG.t����-���a���r�r,qk��"Gt�!#+�pu��%,$����u�OHeF�6�\�:��(R�� ��E�D�����)ˈ���|����<��c{F̏|�g��δ��\���)���i�[m��y$ �C�5La�ڞ$m�N�w��*t	����!��p����Th�V\NO�J+SN�����0�wP��;��Y�ކ���R����¬�^������~�HIeeJH2W���e������~����E��iN�1�<��?�k<�ik7*�ҭ,_�[��-ih�[ۮ��df#�3p�2�#�W�O���3��ZX��K�D''�2J�9�OS�U7�W�� �#��?A �lF��N�q1�����jпt��9�o���& =qg_�i>�C|n�*��)tn�;�Հa#j�Z,>i��y��D+ڸ����C��$'������E�*$��S���|�G�G�F��%�fCf���)׵*g�I��R{Ü�*6��{Ք��T�FD�0F
��ؔ����f����U>�jK�]� Oi�V���ϓ���O"��DE5�Ő#�ѹ��d�xV�*��Ng��"�Ž=�Ȋ�4�i@���9	}w�/L'?K��2���M��_�U�y
�_���ط���>�o=5Q�0�Il��`��F9��J�ȖW��j��=��T�q� �f�)M�ˠi3��|�h��f���ȿ�
���`��.�}�B�p'+J��P�PTpv�'pj:����Y���Ljp}��ǞWy�?�4�f3��C$�}rtq��t�u~��pʕ&x���4QS��V��q��y��0� m1�9��ۚ�������~�x���j�l�#$�}�������*��/�-�W�<��q,Xf������z�3�\&�Ɖ_Q˯ M�2}]P+�'��.bp��.�R�D�1vg
�G}���g�lf��U[�UU�!`Y��Dl�a���tBZ\�k1j�F�������-z�b	o�^C7�n�����Ԕy7�V�f���?�D6 ��d�z�$��z��s�$�0�S1W�OB�=ʓ�g�
��BT֐�de�!���7A�u�Ly؍X�e�6ڈ����W���`߈�E�{r�N��z�������irl+8\��n~�f� F�2ӻ����7f�U&AD�����_�S��G�{˩ց�lF���9JO2&'3��̂rހBIک� 0�nG�oȾ#�ە�8�*Y��E���@��� ֯�3�����P�\!�#�#?b��SM��]�F��v~�Ӿ��!���@y������j��'�W����ŎF���3C�JO�7u�8"���4��݂f�]��:P�YU���������E�2ed/�L� c� R�����&yZ��	��NiU��ʴ*I#�[+��}-5  �J�j�A8��u6庎�6�V����Da�l5U\�����s�tpK$�4;�*�gD��h�㗯文x�[�(���vZ>��ع4bb<xy��[��2A�^[0d�.�׭f�����ý�]�E"K�'�,��l��{fp�\��2��S��l���d�Eԉ0�9�ʥ@e��/��[��Ä�⊭%��28��SĴ� �d;s�Bv~�̘�瀸�C:��22}�9��t�A����B2�ɍ�*���-ƙ˺7�x�V�F���lNE��a���9��в	�-����ۿ���jI=2���j�
�Ĵ��7!i�u̘#��o�f[�A��+�L�{Ίm-K~E:'4�T��������q�8��h��m;U�?>���� ;��?�_������'��v�1����&������\�t��<
�p�3pWFr�� ���y�|����;�.��^����X�W����kh��NHj��`�F=��.���������|�np�A����^f`�tf����+T 4�#[���<?X0Q�J���L��d�܅ϲk��'�K���s��Y��Z���c�zE�]�������S�oo�jJ��1�36Qu)�݌�����WB��� �2	�O�ڴ��y�CkI�f�۹�T:DG�I�]&�̟��f���򹱂̥��?@%���s�>�U����1���R��7� �/F�߉zYVm;b0Ц�w��u!�>Bt=��T*�l��(1����[?"��|��Ŝ���x�4Mr�����{���&�wg
��h�(׷�|/����fB{P�Fm�4gB	�E����A�#v�tq���٠4s�((S��2��Q_,���C�'�޷E�P��U�����1`���#{���j�
K���M??��0��b�v�]ޣ�FT��Z�a]3�Jn%Du��ӣf��ۚROp�q�5s��%X
��_,x��v�����*_�[C���ZJ�;8�M�= �����&���d�ө�"R�|�hu��C5����I� s��/ip�5 E�V*z �G=��|��V��\�;iӏ�A�u����2�͚�GsKp�=�=����
K���ݸ#���X(c�ܳU���9�L�dI��Ž��h��%C��st���N�cݎ��N����\X�d	��H�e�A���?�T��3�Am�5�u^��ޯ��^���+���<�d6ogi�2�+gZ`����c#^�BM��u����['���62��� G�+5-��y1�ZI�����J�}��fY��w��=S��a8?�n0���<FEsR=bąϞ�l���i.��A�%��o���������L��������tR�C�`+M�s&���H�~����X���ٍ@k��o�~�qc�t{��?)��U���� N�8�E�
�	�Rn8�!y�n�p ��::�g��Ґn&�1�Y�!�lz`����	�a���k�����݂�� I 4�'��ә&:c,`i��o�X���� 9�Y�WG~�����.\\�w�,�f����";�Gb�'�������FJQ�;X�yQ;&ZB�$��ף2�Cgh~S���*�`�L���<!�`+*hM�V"��|�k�������؏��e>��U�/��ڕ0m�`�["|��AӪַ�=�^�:R���2�r�����P7V>{鴶S!��;�R{ں�,J�U��!���>s�hn�>��=�	�2�e��b7p��,m%/�ǳ.%�%�I�l��Ұ�o��)���9c1��f9�V�b��@�@��jpC��9
_�	�MNy����;]ø&/i ����[&����DMߦ/.w��~-e�EDX�Js"N�-���kM���� �N`$΅V#�4�'ye�ė-�Z?��B����"j�P����/ŋ�e��%�5*�rX����=�i�ި��^@���u�ż��jl���&[ O�Y�w\2����M��N�#�ӛՔ%��$�Ŷz�|�b��+G���Vb.��RrQ+-�T����ݖǙ[Q�q�>�I�~gz5ڐh�-f�эڽB1m
�=��-�!��SA�I�d�rd��W墭Z��3�)������C���3�?y�!����6���x"����(q���e]"���o��5�biqu:�x�9Hs䘧���L�Qł���K��R��h�=Q�c���Ώff�hOh]�C�,�o�|�=�J=���Oʘ��q�E܊���Zy������eWi��e/Q>w;$�Χ����LX�B�LL�ѐڣǕ�Od+�rÑ�_SUw�R��<����A&��O����Q�S��2����;�.���6-Œ|Ȳ����'y������3$g~�%Ni��>�Q����?+)��2Ig�;���!�>칹��Z����EG���H�Y��RI�^�EP@���A���WT��Y���le�"I�	3�����0�*\�/�C�`el�,8꤫lO^7�"#Ey�5��p�g�Hŋ���;-�\��4#�\�&�YY'���'��j��ڡ�R3[Xk��=HeZ��3��X�0C�R�5ˍV�v8�e�`���I1�q�@-�D���=�������(qm��/j�Ƌ��Shz`����o�WY�R�����>��	R�>#]>�^8�0e&'������@-�!dp���݃��nH�j�� ��W�僺#^���ɱ|y�=�Tn���W��O�����=n���OG{$C�tE��g�^���$����R��hZZ
ȮtG��Ї���L�d4�P���r�?���*�}����1d�%�¹��C�Jl7�����j&��V�V��!�� �#&׿[��
���mE}&g���{�޷Q&���^\0�m=D:���Ҙ��旊W2�]�M��4R>ξi_;ox�X�xc�jw-��xQ�1��0S����</��x����G����0��~#��W<�]�X��i]Ca���/Q܆����Ja�kݾ�c��瞍Bt���
�l�ֈk��'R�	���)������3똒#�C	�|>��l3���#h��BҒ8��%���M���Ɍg��x<�q���؈��q
�����Y%��e!՜��k7}��;���8���x�r�X�}�"{�g�|$�I��!�WY\�b&(�Ɛz�ϭۡn'���]�K�2���k��@��=��ͥ�ρ/"ӎ�R?���N�� _^��2����p�����+	���!b��ސ�A$��}���Z���U�">���m$��5��W�{��!"I>1}y�� ��g(�������<T�'5�; �i
���	y�N5���MĎBi��� �����@�u�z���^�.�?)"Ҥ�J�Ӓ���}齠��4��|ܣ�{�!ka�le��*
x���(�y;ZW��S��Nj�t�5�@��əPRe��63bD$��?
-4���~�t�lDZ�e��6�>�途bȏ=����gr)�͌�u�%|�쪻 �XIV��1I��a>����\h����V¦{NlY���{؀��Q(�^M��RF�:��u}�����1�iMF���pw;x���}��
����M�!N��㨏���eY�_P�������!x�Lf�]�t�ǉ4��
��$����ޡ�K��r>�(�{���o�`���x�x�v��K���Ԩ-Alq`�� ��U��h����3��Wo�sgs�k�[��3|�]�dݥ���X⌒�2'�H@�]���zη�e�&�\:��x�)�(j�;�?��@>g���iZ?�N]��<�g�����G�W͗������h\��l���qUe�"U�9%
`���)��'<AITg5YXӫ<�)�b`�O(th]��h��3����G��h�U��w�åg^v�m�\�˱�<+��T��MW���k/j��5J^�asy�p*>��X����Z���׏{Q�)c��l��m��l���i�� �#�s�t���<��f��/��l�p
�?9��uG�pf�)&czޣ�E���^�2M���_�+��<�� +�%m=��IA��*'ad9F��h��wi�z'���"�����d����Z��m��R����r�.K�����7�UU�ޕʛ���LFǄpR�b2�!��Ӏ�K�cE��R�� �`W[6���-p����a/�W�����L#߿��-�,�#�W�^��N�BU<!�FEm���	�>V���/ӽ����P`�J/��%N�o��CZ�U��H~��a�<�N���ǜ�����L
��yp�b� }�>�P�H�$�?f۸�܎�t�q�"��5������J:����ٱ.޺�a�s��!/0�24}2�˜t�?���~PL_C(~��� v�}lwyt1N :����!$��c+��7����]ɩ�os�'�$�6P��nxop�Nh.�$}C��4��>��9?s���!��B�x��RM���U�T���?`I��ߴR�ak:�R��w��u)J��*|R��g'|ߴ�M�q��j ,�X�?��I���[%� ��,	l�Ӓl��:���r0RG�C�Z��T�q�s�x�!j��s��̢/��E�۔�.Ѣ
��.�B���P��!v$�叞p����3�^`�`�ۨN���J6�W��}�(���?�KɐAv����#�n^ �қ�5���$�	gĽ-z4�vܡ�dH2���5,�@�G8��xH>#i`y�E���DbY�$��=� �F�,�<^I������qn&����B����`ňd!���(A�*&�������4�}�5<��貾@-�b�qZ�)[ݤ�.P]�cf��vn>G�4�O�����v,�=������1<D��1�y�G`���������1پ*L�	�]�������5(���0��w��S�RE�$V-
#᜔�~5ye)�CV9˝w��q�{�f�Qu�#T>'���d�X��auƠ�����Ţu���g�N�p�����f�o~H��#��Υ��&�O���ܾ)*����V��%J(�v��o'��g9�x���i|@?����DL[���r�y�lD9���ĄIR�>�����?$�b�|��H4�t0�|��ej��".��S�.!g(I���ޓ�L#s�U�N��� ��S@<^��Z�tYA�q��W-|R#�(�״�4ԼZ��Ki�|�D<���nkG�|=�J|��	�����6̰U4]��Q9���O�|&�&��d�VF��ˑ���f��=�:oS�p~�TW&M~p����ӃM/�0({�R�h���@I�$�7� v�bB��l��`~�  ��{6ʳ�m��9im��{�ӗV_oYN����&s(�M˲c�0�l��˒������N/wL�R/��
�g0����
��d���A���ll�^�s�W��3W�c|�W��{����i���M�
�K(�&,��J�r]�{:��~�I#��$����k��obqaߧv82���Y��{��>�%
���;�����IM/�p��pj�y��#��!r�W 	��� �(@�U�W�Lq1o6���vH����H9�,Ok
�A>��.�4F�# \���c�s��$,r`b�,�z��V�;9*��6��D�@b�����T���0nX1�)]��Hœ��W�F��}�dd�V�:��>���*	*�94l��f�`kS�!{i*͵[ۿ@�ԡ��Z�߸;�.���.���H�s;�V�O�°���$u��	�Ca5��s7XsC�h���B�KH���|̓�6��t�f�Q�
$���H����NH%Ini�v���� �.7�id!R�(
~5K���k�'d\L��g�$�:��-(�~�F���W��갧9T|��J�.������ڙ��W:o��?� ��?K�'�i$��=�,P`T�����>�Ј>1�0����_q�o���l:�����i~�h�kO�삭b4�I���}��{x�b��CL�����l��Z��M5v?����`� ��m��v��&-���o�/V�2@Y'���E�Ͽ0��HO8f���γf�;B\<,�d�Xp �����g�?�m��� C/���z�Ǩ-V $y��ӌ��X���Iw�7E/7z���'�/M�����W6 ��/Wۖ�	�<�*fPu���7`B�+���>7�3Q��VX���1���K�?���֓�H����VD$`i�NM�x�zOܼVF? �-"��˺��j)��S��ݾz�i�w��ԟ�;����[j6\�Rxo<*h)<�4�D��U2'cMD���l�����9�������R��3��Y��
�h3�ss��� 5mq�/Hb⟔p����*l��ṗ�s�hOֳ7��U���u�t��<�(U'��<d���Hs��S��e��ԕOK�4�ND�����
���_l)`6Vs�m�v��-��[V��a����{Txk&�	̘A ֳ�����T���wd�}�M��͂���k"-9y��M���*�c��m���]� ��lɏ��BՆ��3�,�k֒����c�	�i�E���s���`!������&���(�#�.~�����b�y~�˜��md}h�j��/�����5=�2�q��o�� ���p?<��t��)7i�Xc�p@�S|3��EժK��@-#���W�+�i�f�w��yY����~�X���k)v\T�Bd��2��o�ˡ{���%s��{�#��]$40��	��q�|=��7+��;�<���v���/ (�)[L��;�A���Z4�\�MӾ:]+�;�N̈O/��YJ��]�v�W��:�4��"�w�,���"mj�D�|?�ȩ�L�L�w�Z���g�2�Q���=Q&�_B��.хNY���a�|
��1�1��S�~7�ax`(�f���]Wtw�f�ԓ�����{�Ϝ�H�}�'?h� �ZT��S��@է�(��.� b�o��x=�H��`�7���}R!���S׮�u5�V�Ȅv�\_��	o�G!���}M�LP61�Ԓ��y��^f��ﺟ�`�[���6�I�F��i�+�_M�yy'�DL���4��W�u� h)��V�QR鶧&J\����7��(�1�e 
�d��0�`�+���F9o�V!���0".@E}�9�=K��*����P���I�v!CdfRv�����Y���<�L�cUR�{���
��0u��W�����x����x8�e3�Q5b8v���mw��N�M�s�h
S"�l�|Q+fR�'++����O������xgg��2Re�ǚ�zpg���`�}���ً��������=O9\�E�^�l������u�o<Q�T���5��`"#J.Gg�Q�}���f1a���<���;O�)�I��\#ǝ]�1��K	U�81^�tG�[m�T�`p�O�:��
;�W���yRh3�Ȗ�A���N0�I.���.3� ����_U�cpf�;��v�-6�~ș��c�����䍟��y�	�TjܖBg�R�si���ə^C�b��N*1���f �L
C�������{������/Ҋu}�%^��1��*Ue��ڣ���t�sw��h^���¼7��N��Ԙr����(���V��*����qW`GG,��o~m(�`�@��J�ުF����Qʴ61<H�w<]����X�,F��T� ��R_rM��q�:`����:;��6i�@�ǀ{��9v'���m�MFR;��q��莉>t��<�ă��7���ă�r�x[U�i���W��=��q9��lmMo�ju���4B�`�l~�)�D�T�|{)�hΞ�n�-�ڷR��pMI��v��I�`��\�o��O1��de7�)X��|�M��M;30��.0]�`�*p��p�VB8@��<����=���b��E�������ɜ�{t�HL1��v��![�<Aq�U���j�Kq�{7+HOr]r�����E��K�����r z�3��x �d|�]����Q��?a�w�fk��t�;����+��tEw�"�<<��,esG������Ρ+}t�T���9US�x^*`�n�=�cL�U�B=����V��B7P�/MQV����#T�% 5��ⷿu��kav0M&�6�L��L]������O�y�j�1���� ���V2�Y���h��8��B��j(w�\��G /_D���Q#��_S�U-�ު�m��MҸ�QI�xݧ�9BTec�� 2��no��EK�g��T��ߔ��}M��u,)�0y��cסns���@��\�6��E�K��뒭�#S�Z���u��x�L�5-������m�Я-���� EܙQ�S�O��"PXQG���!]�ϓ~3��(��9�]���8�G�`��)ް��lJ�tK�ߛ*��3��+�"�z��jp*��"���Sxf�a8�������z:3�K#�ld��dwI�o4��#�Ԓ͜�b/�D�b�HI��ԝU��N[��.�[�?Ωd�GMOS�?)z+:���A��ۣC`�;��Y~Eǂ�%g` H�uQA��^(�1�0Ѓ��w�YH�8��z�3�~*����F���Y8ݑYr��%>R���9�5��g�O���J�"�{𖡡�|�D�B��-X��#	C[�Z�����{���.���Q^�"��b/8�è�
�2S̵�u��!ķP�2�E h�����h��1�jʘ���7����n(����Ύ�|��3�`�N)�eP�u�����Ƞ a��̋�iq����&���-}T� !-X��l!�[q���@�Ѕ��_b\��?A�8'9i]�#M3��pts�c��F0�z'��u�$����V\�ˌ�^[U`뇿�^�p�N��F�=�I�_���\���e��E�?�>�7Z�%4����ˊO?����q��	��Q�hq�+���D���k`J��l��Y�����eU+f���G���_���^��;��6���s�K�����I��_v��_��%������ ��x|xUj]�g#�]~��`�E��ˆ���BU�l���ak��	CN�0��ek���"�^be�Z�c\,�*�3��N�I�����_��-����w�e�7��c8���y�d���W2�p�Lo����Q���s�B[Wv���,��2� n�1�q�� �r��o�B"5�����;\m�AL�\�D|덴��IE� �kz���Г�}eo8E���Z\l�\{\��^�P�X)��>�za �����\ܓ����b���W��C�q����f��� k�h-Р1���u�z]�.��V������)�E�.y�����ur=K�׌�G��gW|*)d|�zZe�Al%�cQ��qv;����h�k����җ5W����|-}���z�.�G������ڛ��t��q=}X
��$�U�W�FP�V�@��:aj�v\M.�p֦�TQ�:
���kP��E[��o0��e� qŷpq���^�C���-�9<|p�^5�4��n����ڐ�o���J����X֊�� @��`�M����{J��R^Tn?C]�N�#`�k�fx�Vت��4m �|}�1�뛫 �M�.W�\�s�Qӫ�@���vP4��%�Y��8*7v��u
��"+J��kt�ū�^߃�;�]�_�~!�SS�w`�24F���SE�����I%�j�m���X1/��9F�詙"%r����H�le��v8͝��[��+<`!�	�{�p=�0�Q�J�e��,NA�=�R�/	��f���UO���/x����o���ӑ�-tL��1�C�4�QĴG�]���>4K_�Ow��*ɉ��ܹ��+Yˣ�ibz�M��Bޛ�gI�M�@���G>����q="�5g���e�L����U���F2� �>�F�^��8��9
^G�!*F��+�>�@�ƭ�F�T���>F����9n�����9�I�.���Ϧi��S	���p"�-�X���_�
�C��\]�ݶ!��P�S'�^��s�n�T�n^~%��-�M�(u3��Yj��iL�I�PO�*����xH1rmߢ���dX���L��o��٭Ҹ[VJ�3y�)��=Y�%�|(6��n����b�3N��;!�vQ�F m�>�1�ƸPV�u�K!�oD���C�u.�e��Ɵ�<<%����E�K&�H�6蕽W��P�Td"�����Z��\hRn;{���ǭ��8/��h��Z�}~�z9a�7�a}��2v��>�5JJN�V+�!�.3�7<�"{ ^�}�߂�ֺs��rVnJH|�Q��D|=2�v��#�TC엊��.��LH��l�؏%�d�L������ǣK��a����x9$]����f���j��)Rj�8C�ynj�6�h)̃�\2��Nnu~P���8�yO�,I�x��2�DrW�Y§8fAo`w�2�kJUV�%���tBy}�����űz��D-&(�׼w�2=�A��/�Ė�����e���r`űA�ᘮYr| �%�i(|�����"Mhf�e]_	�u,]����M#]�.��D^ �n`l$]�oњ��eߨ6�_8��ĉ�0�E1.<7
�[�8��
���[�^��8{D���B��$���5�9��b"���R�7S`����ִ�4�_��$aب����í�4�Iw;0�R��@J���v+έ,x)�~�"P���2h�@��|��izN}>�Z�5x�Z�I�QC�Q��.��%Ѭg���U� %[�X�Hԇ�I/�`F�D�-)�ǂ3D�/�\�O®v�`���zP_���~@IQ�`ab�o7���s����̖��k�H+X����gMI/zZb���e���J�u�Ûq!����sD;���7�C{f�T��=?Y7U������{����0q���?����8�����b�(�/X���AI!��aɩ#]�*��.���ɠ�s��#(*&C�xJY�6�!_DR\Q�F��9����! T��eU5$TN��H�񵈙�`�h��7��#깎|1�S��oN��F� ��6�|�c0�=q�(��C��Β�4��<i]��4Q,q4 ����z#=�7z\�s����0#>b�lM .�I�ŗ�k>��Ψ�1�<�CWP���K�e6l����S|�%�p�~�t��{X�daq�J���^�.G��MGx�i&��"y��Ycz����={b��ջ�/�U��zv;��xWsŷ �\�:`�|�6�ex�ʭz�ITj�U2�-�V��KZ@��i��4�E�ꑠ�M���F�-'8 ����j��f������Ĩ����1	� םG�/w����^��x�SmU�@�&�e�:�e��O�g��J�j{��D-�ص��z�zs�i�Uw�T�Z.�P0Ip^�qeÜOZ|Z_���!|�$�'����s��q喧�D��h��-���$pu��u8h\�g��f����i�ƭ�������!��x�U3DL�T���������9ߵ��j�o2�y�n�+N���M~M�*nܕ����0�Ϋ8�,�2�n֬�Ʋd[�^��:P7hh�d��RhwߠZ��5;9�4$��~�wnV(m���c
��o�����B�v:�<|�X��3�����dt]hR[�����ʉ��2�oҍ*�=�'V���[ab�^����?D�һ�!c��!��ݻ;8�
��]���9�?Z]Z���=��ZYZ��W�[��ڭ�"j�-�͈�F�J'ڙ)����p��'}�V�C"��+R�U�4�%	��{��A ��8=�h��Y]�aW����Mu�^���)�C�X���t�� hoA0&���v�gj���t�uX(�`��p#��OyS�a�*5Nљ��=2z<?|�U����&��:�k����ӑ;t�����������i���?���d`G�2����	���8�#��Q5���A����݄�D�m�8�n��-񭀅�ZZB#H����+{��������PFHg��:��x�T�Y3��~䟫��(��"8l0�%,�5K
f��Ӗk�`Y�L?D�#���b�PeT�����c%~��@m6�|��1�|2q^pl'�&�=ǎ&�q���+��a��~�>��g��eI8W<�JLgȬN�!�̑@ha��d�4Ax��ք���n�ɾ�r�iV�)J���1m�t��9�p@��݉�ϲq%�m0�.��A��ӣI���A��Y��3��"���e����.�����8Z�Y�wN�m�@Q���(���M��FM�)���\ﾙ��Gu%#2����91ov�������I�6��&���t}j�d��y~�S1���y��B\�&�FC
�c�q��ko������>��N�o�mټ�O��Կ��vd��vH�߫T�9`I�]l����?���H�E;`��k�9o�<#�$n�Y�E�4׫S��ٻz�c������*.�u�nl@�Z���ih���APL�\!��mnf29�:��a wy�+z��f��AsO~ʡDPy��qm�0}�xP���<?L�8��jy�����X�}���1k_��s^w�-8�9~���~fKq)��|���+e19#wC���-���X��ab#���:W��$�B�|� ����T�\�k�?����
�a�/f�#;^�W���3�;�ٜ��㿛�0�]w��EH�nS'xeqNKj��uk�j�M�b��}�=N�:ѿy�h=��A��R�<��%+qU>��rwe{�<Er�j���ЮIz��:�*��ǽ�����Ԙy�)��C�O����0{j��EQ^xuߔ��/�l��� �LF�{�z��a^P1�^+̎�|�|q51�J.�$�b�=w������VƇ�R>� S`M���L����
W�UM�4�`MO3uA����a�$kA=U8m�����V��]�?�|��|�W�⪚��is�IF_��������sF�lf*_�����c��N�p�8.���yJE4���_��F�-<.7��һ�S�8��Tr��E�Ǯ�ǄHADt������1u1�����"�]������<����a$LѤ��S���iaN���jI)��\HW %{��eH��p�}N}�q�<o�6��ɧ2
�I���C5��|y�D׸!�C���D�o������ �M��E��Vit�0�>��3sϦo���f]�����M[�ۋ���-ƕ�"a��N�甐M��H�V���0�x�=64EIN:����p��ht �]`SDRPH�5��w);/��1κ>��l�D��ANJ*m\���3�ά,w�Ê��U�(�e�Y\}�.Ww�%�,(b~�2��n3��P�u����T~�]��5�w��ɮ��u,�Ia�Kf�O*Y7�m�� q.p�
��f�ه�_��j�@�r���(��Qh@=ћ���Cs�����2p�Nk���b�<^�St�>ͭX�O��%B �}tg/N��ϝ��QL���JŚ:�~!��M�){����R���W0�w-��<�0�ǰ�<��Ԝ����}MhS�U�߮^�<[�M;���z�(�md;�j�h��N���L��^��t�`��d�������P]>%h����ܱ�q�n��X� ���w���L��FwC�ip,� ��$����AX��f�W� r>7�4�� E�$Qu��ㅧfǮ�w+�!���G��)��h���C�顭U��߮Èe8��|8?�ء��+'��Њ�#�k��T��茛�7�z+~�U�i(2ۓc�v��1d��}_�{^F7��&G!�L�J<��;`Qg2j�k0������E���m%.nm<A���!%U$,��G�Z�Ǎa�uڰ�#*�̋�*^��F���u/�Sv�$v9���S�U׹�(F!+�������DO��[.2��"�oh�n�2o.�[q�t���/�+#7��M�g�c��{'"e+�8ï ��T�����߃~����$9)^=�&��lT6�'o[]��"\�Ұ��_�NB�'֥� �@?>ͣ��,��ü'o��[1��D��T��pI$�p��[�`��*M3��S��.	ǡyTu~ ���������/ϴ	
��ͱ���i
H\�>�Ӡ���J��؂�v�;i��Ԃ�B�>��51��8@�{��ȵw��d&ö)}���6]�n.�Mi%�8�f�y|t�c)�[U'�jl���}���&Fj�	��b~��bu���.�T��G)^X>R�����O��V�C��k�z��7i ����13K&��rT��T�}{�,��~�ޫC]���CoK�c0)��ΖD�#���{��aR2��Fn�=�hl=�[��2Xq�8��V��"�dؓ�Ŵk����U�Pj���9��b�p:!����T#߸��ԍfa1�zP������D���F,�����k���2�#�� ܂�����&��P	Xa"Ә��Dk?%2��]V͊Tݬ�s�4�3G���JR ��l���(��Z�c⚉ 9�����9��y���|x�핝]���Ь���"	$ܿU��1E��o�'�N��W(๼�TS]x���Vh��ɏĉ>�iMG��ÿ���w!��s,�~J�W�*�ջ�=�����OZ���W��#�������;�m�����dS����w��7��}���9SY}r��}�c����$P�E��"b���i��֏���񅡆�֠�0d'lz]n�[A�(\*��6E^���ڴW?�'����`3m2 ����1���r}�q�-"	\G�#�y�#���4M��Ws��R��[�/�Z$�
�j^�y��E�e����SƝ(��%F���X%8�p�ו;c�ٝ;��s��3�+.gOO!�j���A�G�?M��?kP.t�����ݭL�4/K.�Aw��:}��"�x���=����6ՓD��Yd�΋z#[��+�Q1��T���b"R �6F�w������5�{X[�]����Rw�B�^�mn��e��h�X��D�a�́�v��>�%���=77��3���Z�gT�����\�wah��f�Ok�ͽ�o��}Z��n��/h���f<(r�)O���.� d�u6u��:voR�����dTQ�u�.���2Y��o,؀�x.2؞�x��
�D85�璻���/���,���E�Wѭs��	QN��,b� ���Y���\/��\����C	e��]���@��0o%��HB'~��Ϧ;�$�P�����e����>�������H�_��8O��Pb�~���[�����9����R<�uۦ�����^���:Ϧ��u�k'�;K	��o3 Tl����s ��!,���!���(x��,'v/��aRY7�aBhJK�d����1�&Y	����j�L=�i������C�ŅsIu+�@���0�r:)X8<���v�%p�* bA��0T0�ӀZ��MN�뤬��9�h�J����U���ۆ���e���
�:	 n��ȝE�8����ȩ�<1T@e�ddU�|n��g- �8c+O�i�暃����"�}��Rg}��l�Urz�4N��p�6�;\�=��eX��2zO�[K���!��kv��>3���9r�v"��g[F��Bl�L���SF�����b���8��\W4j2[2��I�Ѳ�N
-:6��l�H��X)7����;���c{� ��AA[c?4���Z�����7�hI�+>���ŵ���AK�8D6װ��6YR`c��zf�v���|��^��c�� �]3w[�D�5  7��R����ڛk���ε�Yi�lc���Ͼ�R+�퍻�y�]y�J2+!�g�S��.m��7������|O��wh!�<��o�����'J#�b�X�U\���Et�4�q=�T9��q���;�2�ee n�]��|l�@���=Fvι� ΢о�4i��{� A�
�zv�M���O��d80�W�D��ä��fЎ�H~�^ 鹅N�zЮ;DS��c�]���ܣ����I��%���&)�	(�Q��i� ���<�Ld��)�&_��N�!�m�$���=������;������m �lC�A-{fL�����ѵ,~���>�G�Ǜ�J��`�mt߭�Fā����� F�zd�jm[U����d8L�6CuJX_�	��)�gSm+]a� Z�����l^�C�?T"U&�:��l�L�݂���V%0��T�l�m�k���c8|XFy���a�"L�VΎ���I�������3��j��}��j���+�`TB���3~/]4q��k�8�Ek���B �0;/��M	�-C�]+aE���
��]�n��B�`��N:]���%��+=��ã��g��i����TYoQ��o0ڲx$]��KV��&j��m��\$D�ÄA�����5Q\�!6,;����=������(���M�Q�m_x��Pa�O ��}����x�ʊO՘�U�ܯB��ɀ*���j���=t��Ӎ�4L�_Y}k5�V� |�M����%� �y��/��RɋW �*ڢb�:}�ض���0)��q��-�T����ڎ(�^�O������$k>����ڭ��8QS|w� d)�e�ͧH�턄 �:�H�X4&0�F���5�B?�!o9�:��"4�0<z@�q'��tu�U��C^tYx��X�sJ2����_#������ �V�j�<)��A)$b��]�@�N����,wJKa��W���&U�4�xZ�k��D�ed�D��
B}�5j����]ס��Sq��.��b7ۃs����Cz^y�%_����i�EW�Y��ɲ%�b�k�׳��\T�̮�����s��=d���Z�%�����S0��r�#f����h����Ր-�6ErP+�H��ű`��x��e�l�06��Ka�r|�Zz�r�ï�l4�q��-�K�Qz0�O D��I	�*��]���='bj����q0<��Æ���<�f����5��������J�tǐ�c���T5�M�,�Ť�RkRCQ�s.�}�d�W¢����'������ja��x�"jQ9�rL&E,�H�	_�]tO����׸l3�cE{��c]s��%���ҫ�(B��L�8i��vk�OC���9�*�
�����7�	�"(2б�.���8?k[|�Q��z
fIu0�3�ḧko
Əe&8gs't�0H}1ۘ��h��}���@|!f��;Z�)������P^.��P*�172'�;��bYNGa�q_�:O��X��K���U�3ˆ~�^���a x���Iiˁ�Q-{��ڙ�1�59ʱ��m߽I���bu�2Z*<���?�m��D�if5���Ð'GB�ź$le��R���1I�0S3��}���rA��(�� }��J\x��$�$lw.y����- }	7.��9-�ѶH���^=��5��R�FX����M M���,�oU��MHm�q���^��ի/s����;WiKĭ�K�e��~w�5�wU�V_5��pH�!_*P� V���K���|����r�\ƊL����v�B��V%J�d��
���S�f��e��"�b!K��������]2��v=����Ic����"�s2G;� ��/��@I�T�ɷ{�sM+^����T�L�^��7DQU���AI�$�`�p����9�)%3U��I���)J�w��M�nu�S��Fو�	��k�5S�	9� ��`&��f9.;�Ff�����S�ЖN�]�;3������~��ګ��,��-\K|	�7��]���F����TH+
f*�Fr�q�����ilB�~f��(k}k��`�^���;�PUD\s2�nW���*�b�7�(у]b-�1ã'N@+�9Y҅ ."�p�+��X���`L}ݾ	�'MxV%�������P\?9�]�d�0a��kA�PDlv䁰M�܄����}j��u��O��<�|�WAE-�Ȇ)tL�qߤe;��K�C˸E�5���h���ۙ���0_)eab��Z���@����5���Ǐ��j>��3� �Vׇ.51�&���i�uDy3�3Z.#���U�Φ�/�U��t�#F��.��������M�;���;��Ma���Ɉwʓk9��n���Q-�nЖߓ.^���S�얆��w��c�B�ܑ�z����v��^�e�}�jĞ��]),���5B��[:�bo��B�KB�y�<#$p��eҪ�,8Vr�����+��A�4u�,����6JH3���6.���$T�%�kQ��>����lu��Ѵy��f�mM&��;ԁ���k��<)<��6�dvvSr�W����Kv��8}ya�a(IC[�V]�,�����r�E�=���m����q#=��Z��:�7-���;�R�$89jvY�R�`�|���hA��mg��S%���͈EݨAY�=�'�~���*�-�d�6�?\��͖*���B?�]��q%+>�|���_�j����s7���AS{XL��ʫ�w�v�<J��ꢉ;��%,�F''��.ڵ5#�RSE�k-p.�yJ�*(A�!��y,z�*��p����ˠf��,�lx��>ξ�K���s�(L�j���M�������;�֡CR�V(��m�:\N�\�{�v������R޲�vz�ts���/����y�.[3���ucv>���2��2/��s�aV�څ�,"�g ��x��@#�8�7��a ���	��lP2�Ȩw֏�b�n���Q�R��8r�$	w\�|<_:6�Ќ��Lx���)(�%ND�����4�I�A���T�\���<D,�{O�����P��|�cU�=�(߄@-��0�����ג�&x���{�8$�ۧ��M�u媧|��R-�]��e@�}�㧃 iU|!i����L��SNg�-I�4������Wƽۤ&X�a���N��f���N���/d�:��㗈��P��s6�u1fk��ә���<d������)���ĺ��ݙ��p�C ��&	�*R���Ȏ�f��%���3�V{ ��Nq��e4u��9���`� ��Ύ�QÂ{�Kbl���K["�Y��o�+$���Ba�<=Z�VŅ�)����.g�j��>Z?ѭ�fU=n���*Tc�ZS�cR���6���*�ߪ<,D���8���9|؎m���}�֏u�ȫ��}@��A&/�(��h_)Fg��߃���d�Wi����9+�M{UA�9k���á������Dba��Z	fB%�y�O��}i�l�l�=FѤ��&iΉ�R$��u�5�H0N������|*4� �w���=0ì�&���Y�����qc����^�Þ|�%U�t���3�6�g���a� *���l��!R�Q,�H�+T�F2���|Z�oG
$oI���!�l,���_�����w�?pĪ3֬��9�~	�y=cM!,�v��"9԰V_sl�ǥ&"���2�?#�OR�2�ͳ�ퟱ>�\�����i���N�;��K�'٦�7���l��~�Q=���1~
����1p+�W�#�w��/:������f��8�eRyL���W�v�<�)2�i��U��Q��^��5Є��Lxr���q�%*��z۩�!p꿌N��՚���$8X������XcP�87V:��ަ�s#<�9<dn��>���% �ǌ6޻-^�����z��%(/��,�����Lt�QIY�R�������<u2��?��Đ�Ǎ�3ʓzPKX
�Y��}�X�1pf˹M�L�����*0�4�+'jW��Vƨ�k�"4`qI���	?c-��]@Pd]��w���e��/�,�&�%t��j�ϕ"U�Է;V!��������`�0⤻�5����b���Y,���\�(�Q����1X�l~�w�AD�Wk���x~���	2����F!�PXi��`G��'̨� �]�7�v�ڄj�90zS���H�ّ��gL�9�@��ҺWҏ�ǆ0rٗ�T��Q���Vb�o�}��җs���N-Z����]��N�.�ؐ�~^�{�i���̬+.�m�C��C�_�����A0ǐD��|���c�}����t��A��}U�Z.:�5�6�����0T�hN{�,��vk�#��w�q��D�T]�c�#�نM�(��:�}nCSO���<9�g�t��9��*�E6o%�Lm�ɜ��c��I`2�x3L� ��
��g=| "�ƛ�.�r�����air`�V`N�!�>�`�%ޢ�e�w=���U}�uibG�"Hڔu:��@p� �9|x���	� �hYuw�]��7��E���"�������D+��2���Q�<�
�xzưw�(���0Pݛ�����!�?9�WYn��t�οG#T��*���\WD�?>��������z����0���g��,hL��K��ho������?�\��t�3zG~����^+Ǒ��r��/�Z�L�V�GBN&v\<��d��!s���^�*i�J������Cr��8���z�q}�2?��F��t�Am	NR{s��f�ԅN���g�U�Q%��>ki�E�樹��j:��f�X��RLtf���MnlU�33�Uz�l�&۶[�0c�R�3��!�.ȶ希cӡW4+�RTY�pz�(��E�m�|{�۳J<�P����:�2��ꮸP�+���m�j�i����9����-��POHf9�_z0+�}o�yR07��������J�-��e���������+��w�j��SL��� v\�p��n*��2�� o�x�JDf�F�IF~�#��3�mL���h:�^ �,�y-ř슫S�O�B�FiF�`[���C�ҳ�� �J��La����]l%H�~�
H�1?t��t v
h4����[�01�uKh�iނk�� ���e��*>/!L�W%?7-���&�v}�i,w�����M鹇>d=���%���Y��s��..�?��W��l�90��+�@���z��};F;�+R��W��
�<�N�|r�0���bcxpZ�gձw,u��[ɋ��7j2P�_9�-<��X�)J�K}��s�q��E�����g�_,7�kYDWN׭�A�R"ψ�������\ɸ�{Cq%m5w����T�)���
���ܛ3AA�J�aҭ��-��VT�KIHv$~B�����o�5�IJi����$'�?�bFl,>������c�'U�@�9B�)�r)�9s�$~�ή2]�(*����+=6�
�7M�4<�<W��vV�WUN["7�1�]�n��	�i�LF���v��	�������z�WL�������Ѧ�1��뀥tӀ����.B��y�q3tcބ}$$2g�\"�jq赘n����R����� �m���X��C���Xq��tK�����Fb�����O�q�5U��<��<}��^�uq��
K��1Q��k���~+=-�B��r�,7Os�=�U�Ճ"��5�TD��jR��!|�U5kXc��/.��\\��q�ĒK<�b�B��Dm8�n��3\�M/��o��L+<��렏�����h&�Vj�M�SNA΍���G�ht��>��X`�PlG,�r�ʄ���e�h�*�\��tc�K_ka7�ɟa`���t��^�,2���^�����㰧?ƣs�o�Nr;���#�Q�,��Y~A䮻�H����L�v��Ɯs\��>�r��Kg]jS��x�d�ԕ�����]�Ndð��WtW������gJB�t�'Y@k�P{�i�D��r��IK�d8��g��W���I	�g�u�h�� N�άf��x�Ӿ�8yE�ڤ��C7���91��ϸ7���Y����%1�g�:5F '�$Z�,�_�U�(~~�;�EIp[��c����=h5������v�q���̳���1��N�LoM�Q�d�(
qSv�0
����K��)�G�3��B���[{qэ��� ܾ��^���.�=`�4nn�XiY�-��(��"N���Ρ��%�& (	b%ؙ�6��%��;��9��kQ��:\vژ5��ڢ
=̅g�W~�~��\�o2�E�+|���'Y�B}�-*#a�;~�����z3]�Ġ��Ͻ��J�^���H,�^���T��ga��d�j�|�2�����u�f߶�O߅���2�y�m�x��ԫe��[BB�m�9�#=�؎���>���r��M�Y�`��/�����-R��l�b�iC'_��M��Ks�>����-�BA�8�Z:��������j�Ҽ�>x3��W>vy�;q!)�E�sp�1��`�_K���� ˁ�3{[����H��&F�;�5�Sݖ�r
(x�՚-%q_M�vv2�'��F�HxX7�C��@E���k�J�*�8�W ���c�Y��׈�����[�q�PX�d-K6@u��$u_��燆���Ig�W���j'��!������6=x�;�USsU	��]��A�"�#e�"݈4�H�E)�[��%��M�ٺ�tc�jfp=)�!�B�4�O[�)� ����M!Q�X~��TyC=�_�?��'p�+$x��em/� ��\&;�7l�:��*\a;�\v��X��`k���̝(��!s�>�Nf��x�٥~�� +�����}��3�wm2�m�����qN��O����\����7P���e�ֹ,Ol.�BiAƙ+R����&"10��T��q	a�lW����"���պ:M˜�O���Yg�AB�ٌ<G��2�Xqm:� ��i�w�Wu;{���6��E&�[�D�sy6�"��T������1UqӁ��rx���DB7A�@��k��-���g� jM�jpH%D�t��!h�;'���h��F<�^�~�����/�[�5�'%W�d�ċ�̞�x�a�PoL��W2	������
%nS��E?Β�{J�ը��sv�R�r_�@�\N@�����
�4m%Y5w��u~,*g�i�<�'$�^���p����މ�}@{���/z�F��5��#1}���\��?E�NB<�:��q���ˑ ު?_w���S������H�
u9��YC���E�����v��:�]Ed��<����V�'�wY����^z;$��ІU߅�ir�q�1q��2H*F�,���w@���LL��6��uڌV&���!���lN�����@_�Ϊ�%��F��փ%��]^St��}lM��뷋2�!��BM��)P����˻����bV�:�P3��zs��֛yRz�V_�1N����q��(�)�UD!����4��}C����Of�4��PO�%��V����ޕ�qKA�Ӗ!9�75���(�%2+��~K+�
��fpO�yz����Q�T�3��|�[��;.�X]��3-Sm���Y����(HbS��M^�mJ�]�����{f"����]qcP�r�Y"~NC~���Ht_�{"��j�{Zⵉ��]��	UO�;���	�d��.\]E_�*��|�KT���U����4�_�Z�%���O�0p��"���\	��P��-��|4�-�y��}:S?;�H����[.�kj-�,3O#��#��`O�����E�:�䖸a�|�QyEf��p�J&������_�u���f�1�k��j��#)Z�OPo�la�0��g
�`�(��Z�mX�~��k�"�,���ժ����Ȳ8�S͑�i'Fq�]��k�#���mB�:|o�iU��:�S�_s/��\�ӷ<p�·a`��l�� ��[�0&�Q"2�0��?��������%A5�A�s�r�E�{�ƊYvGR�F��(�0o��&7�U��H���[�{k�b�����Q�����*���'�^�9����FJm�o)�� ��W#��������ԑ=��h��v���3��%mKi�EM��-�ѠߛЁ�h�6Q���<g.���y����񢸻f��D#��R��xڟ�zKy�N/"�7�o�R}�D�c�y�6:�'�$,���������r����(]�Ϟ�64�HD��M�g�9{��I�!�]�Xy]�]��e�F���=��u�Y��T��.�Q�>�0Ln��%	�Sd�I����0(�ߢZP���c��NKo{	��=+��ӕ#ы�;�h,��#JGp�f���������'��vs{W��O�N�Q��O��BR����wlG�d ��S)��J{ͱ.mR�Rݎa�'��?��2�x���i�jH�� �Q��zzF�||�J������]+A���#>��v�#_/!���:5�ж��?��>����T�1�S-��ذ@⺸���ś���%G�߸����$|4�`B�����,r`�k��������#-ǎؐ�b�7$���Ȭ9�u͢qZr�+�RFQ�� Q���7����Kl���
~���K���l�>XP��`�zXv�j$���ۏ�c't$�*���k̲q�f4�D��R�c����X:a4�p�F|�e����le0��C��J�Ö�#d�Ա+c8]�����bqN�6m'�v1��G@xFO����G��:,	`fAZ��y�}aBK���F�r�W��	#_Z�1�1(93�u�i�Q"aߠ�WHu%��m{�W�ꄑ�����:v�*�1]��/8�����r��`r����"4�����wu�7F�c���Y��H�x׆G����Ù �ː|ŰA׋x��{�+�[1j�3�`s�(%&�����m�(��2GB�M�����:�7�KOd"$�MFo�]O6(���j��S��FlVRH�`W�^A);�Or��$�;ۊ����! �Hii������L?K[{�n^�6vg��y6�'��r�R@!Р�l)�o�g���4�9��7No�,�D������j��'���tǳt���L���ww�C��jw�1!���E�}X����4@��r{�3��#;L10��4P���H�W-0?���<.�u�憷�O��!�F��~==���3�}��\�h>��e��o��Ict.����s�hL!O{�5�E/�"�ٟ7��_M�V�<T�u,^�u}���
=�� a�:}N��5f ˨��	M�&�Rh�81�f�ed���RPt�P@ܯ��OZ����	��K1��[:��|xi�#SE�����Xo珢�IC'S+xt p�'m�);�I��e.`��( �╺j~�Wܞ$�w����"n��Y�hZ7�{�׼������{���BS���K�B��i�ui� 6�B���P�){<�Ҭ�7ߤD���cj]�"w��E�=�Wq���NX�Ǽ�-�?qVn���VНb��E�ln���������k�$Nhj�eQ(s�lx�~�;����pp�����Q��Զ��ȕr�O��Q��E��ae�h'��ã�:Z<L�}�%Hr��ΔN��8Y��4�ѱ��,[�6�v���	@ �Sv��Ѓ[�|��U�N�@}R@�^��� �*�91���-����'Qm�]���<tG�F|l[&>��;��ɀlZK��8֎m� Oy��C`�d�����8�.��4Y�%�8t�o�\i��au\Z��h�CՏ����]o�p��E�^�>�d:\�=(T=[��CSYVI?%�d�]Z�RxМx�ґ��V���q���ph_��#�Ɵ�	jq:�H@p�w�c?<������e�"�}E�լ'�ǵ���~޸z� ���GVN|��s��K4'�3W�P7�j���p�G�x�[0��:�.	�S^� �˷�/A�P���Ȕ"�x�����tH&|�x!�D��f�iï��F��l���@����;��*]������Ŋ۶i2��r����"Y1Ӎ�ծ(h�������~���#x�3�J�c�Ӑ�=|�$\Ս�~�S�ZWcnR�&^�h�-V�+ŠP����E?i�#���-�6�u̯ƒ?��yHWa�7A4�0E"�wd�L�\�/�'�~�k��6�eM}yT^��5���A*6��y�
r��PQ/d�-u��qL�/A4l$!��g����n��a�&\a`�I��QN��T��e̾��~D�K*�����͆sUr"�IJ<<j���፾�>�.�{��aTa[��i
���F�`���v6�>M����O��1�dv���p0�~����'[5��Zʭ��b� :�~kbb�^�Ϝ���0f�0�D��5!>����y�J6j���G�rl�
�85����?��o;����'м�=? No��3B�{�-]#��4�B��7��q��'n��(G�(���#�/���x�wQczy<Jϱ�8���5w�M��ش���G&k�,� Du������c"a׏���������A.�3��r�(�VB �=��7��n��±IIa�fʣӡ�m�Lr)Q�|�a"�p�y%��y��|�=��<��$]._����/���n�����[����}�Q�����t]^Z3G,u�Բ����U���;��[�HP�ן6ԅE|e,�Iԇ�����\]��ƀ���$�L�$.�v�UY�+�m�ƫ�+f���q��(��pna��p�/HQe^n���)��Wd��c�"q�gg���+I~c:i����	���5��<��r�,��1Ӊ5�]G�̮�ȵ����`���y���p�_�0l3XJo.�Xd��W�Q�1��N�M�FLy�(�W��.����XzG�̩ڄ5U	��1��R��;���{ۖߡ�(�����M�	��q赅�k0.��+Ǿ�?h��V厺G��Y巬���$&h.eTTJ�Ƭa<��f^�
jҹ�:^���6���Ԙ�J v���m���o-�F�%�	�T{�Z��}��o�aD���@��e�\�W_��4R�9��FH�����@�>݋+���F��4ڐ'��OB�dݕ�餳Ab��\!y�%:��$� Oxm/"�����C��7�/Jv�����^��7��e�_�ک5SG\�N�����z/Yۘen<8$����>3�a���qML�܌v��2�yL�+��̝$��Yԡ��!��b�9*�!N�)˽6��Pg�� (e�X~��F��=�����S���Q��U����鉮5xa��Z/���wee{�E�[ñ�D�P��m#?`���}Q�L`V�xN����<�j�C*�:Li!�5�^V���%lQ��Q}q#��.��"��[
��բ�'ds���5{s�<�BP[[L�L�չfJm��޵�R�jw��xg�=�x��c�QS�C/^�6O6��Xl���ARr�s�UZß�õ��l��Ϳ��-�}��K{�P|օ�}8N��s0j6��$�X u"�JR�MR���M`�x�(����$`܊@��,�G��@�hd��ɧ%�>/��2�M���È���KW飴�)$z�X:y�H˴q���pVU'���-�1�7��cBzV�r�#:x1�f�,�gxw� �Ȩ�,tlkm��"��zr�Y*�?-�48�W{V�d������X�&�N�:��4�Bb�=��p�wn�K�{���̽Sv��թ�Xs1�Q���GKh�t�,�+�|��t�����q�#ɾ��`{&P�P͛�Ɋ4�WV|?�"�0�\�10��0�Q����f-�ܵ�_����Hc�ϔk��=�^k�,�����U��F�	��n�f�Yļ�q�L��?�x�>'xU"�#M�f��q<�)x���� HpY�2G�	oA��7�&�2�f�:0���l{����K�v	ʺ�3�6�!��se�t5�,O��F-�l�S�R��C{X���)iI�E�o��@R.�-=�]I<T��3IyZ�����R�Ș�k��Ɣ�WT���eA�Hm]@�0-r�%��ރ^:,!�P��:��7G�0�br����ҝ����� ��j{fZ;D���-��6��&�ߗ��t���|���=���!�h�CG�q�ѡKz�d�p�ߴZ �8��T�x�Dq�kr�.n�*p�f`݄Z,1��UO��z��`���x�`�����]j���D�`��A��"���xi6��eV��Ӄ���;�͎�0��L��o/l��/`<����8@�1:�[�d\l�b?W����CU��q��F��nI(t�+y����̷�3W���2�ʮ�[C�~ T�^Q��*�.x���v!O��x�bObqZd^\�F<g�==�['���{ҙc6�(��	��.��������J��4��G����/�M�`_77pWd��<�l��Z�h��ݞ��8~�� �{��M��D��;B�A6�p�/�x#s6�}^�
MF��e�����͂����k�H�d�ЏZb[|����U������!1�}�ŭ����N�J��:���tf�y��Ӌ��"�� ���D��p|Ђ�E��rQ����o�͏7�5@Xۀ��9q X��č +T�moUVR �.��W5y�'d�",�?�`y��4�d4c�5t�W���K�@��f�u��O����Cx2D��u���TC��$o.���������n��! �f	���e֠Z}���=Z�E���|V\�5�QN3h3�5'y��U�f]��|��r��,K�G`Y̚�l�V�E��Kw�7��N�?虵�i��LZIϥ����$7�g�}�P�N�Ҥjb�}n�/V�E�R��F�\�v��a�@��W�'����*I�h&����
�(�Z�	MRr�o��[�����=�C�fl)nM̩4���9�/J��M�dp߿�l����U��B�RU�3�"�(�o�w����s�3���-'���R5�G�PW��L�Ѷ)���ʍs(����N1g����/��<O�N�z�]����"�%��u�J�z._�r�wؽ&�4Nu�C���![�����/�sL�o�u�q�m`X5���O���m�ߍ��Q��iJ&�Fu��s���M��2-]9S����=1�� �15c�sܑ��.�� ��6���o.�X}�e������\Ix������U8����l,�=��<*!�N�xh�[�Q�Z�I����n���Q$� KyJW�k:t�&��(��\n��f�z�i}	t��gu�Y�M�o���s��u?G�MO�y�����T����o��q<���PPM6U��7�s�qǛw�<_���X��O���)�����]�70��d��p����;�=�IN�%����Xl�L�K��O��*��d'YjO��[��J^s�밺���ͯ:Y��PN�����167{nǮq� �h��2�#j6�I����)�>����V.6��}^ܳs��]�����͕B�o��ǁ�+�B�y�-yu�l.o,ny� [������!ec��k���j�.fn#� �wT�؞�IA��B�g�e�0^n�+[���n�	`o!��.5O�K\��ۉ[�u�yM���d�jf C�z�^</p�#
B�:��4- �h&gu�-�����b�^k� Ⱥ�4G����d�L����bR�f��wF��J�Bx~z�����8Ջ��7`�޲�eN�E� �%a7~3��-��߮[��zM��T�A�!��M(xhĿ �G.kw�����dG�Ma �mM?m�J�<^j�fL]؃�����ec�*�v���k����(��.�(��(=�g�aH����	{fs�C14DX_���6 ��+R��/���Ƞr0?�Fݹ�h>���}��C�;��Jz��=XC#&�'z�H{�c��i��f�yP$~\���u��R8��/��{��hψw�p�Y�M�#?���]�ߍ�Y�-|u�b��ʎ���C��Ztm�a޷����>,Koi��iX���H|rE����3�Ui��5��2�����w��ߙ���4z�7<nv�9UP]$�B<�,��K�|�L������*f����.#�2�*��!jV3d�R-�o�P�Yt��(h�v��d�&����$��s����?;.���Ct���+��
����{'�բ����ծ@�N|j��
P-$r�[���-Ixzl
%Q3J���a�=mz���Ysd�Xy`a��%�y��X��{�U;%�TDu�cD2�@(�\7_�h��*�ƒ�h��6�f(��!�()���:�x ��g���Ӝgdcw�>���4�- e����,��C������~߃;.�3f)}�X{���ty���m���5u��5����wF���h��%��ʈ���E���.�4���=1Z܂���^r�&&�A�]Zf'0DԥIY.�x������h�Q�5��C�"��� !#ګ�Ÿ���~`S��6�y�b�O�f��,O��r��Lz�־<���7���.��jA�ԕ�aNVo�I��&��n-"��}ؽ^�Y�dy��ү5�O��e�˞^M�ҟQ�l(:�ю�)y�)n䡰T���A��B���'\���dA�
16�!�����s1���`RV ۑ��^@�J!�>:/ �y�g�����l h sD������b����a�!��`)[�G��q��Ǜ�[���� �EN�DBOP�����<���'dJ#>7�)��0%�Ox,s�d�V�	��	߶��YzQX5D�v1F�Vf<]7!��f������/�� i����I�I�Wjpw�|)����x�WN���W������j�粐z�bc%B��H�����C]8!��U�p�|1@����ϧI�|��(b�}�I�ܭ��3��04��v���3�I5|_���Nh*�0$������0M"�C�1�3����tx�QB�6����y�aP�;@�W�;� �{��F�|99.h�6����6\����d|�8����pR���F���Bw;#�^��SK҂A����Ԓ���{m]��ϗ��Gߤ��P�{�ٻ>�luT����	���;�Ï��L=��M�w�w��0�p�+7K$=��Z���:�VԸ	c�|��vN��]���;��|G�=SV"	��������&Z.�6O��.D�~;Oڵ������Tr��4���x���y��2�ȶq�=-"V���(� ��D�ӣ	��`�ܔ�K��'I���ҳ���B�_�G6Y<��ݏ�a��M�{R3:�ˬąB˷̪�fD�	$�<����)N*�ft�+�6��˛�+���	��v���\kl��&���M�['��^�� X�U*6����p�6TE�Ӣ[�`k"Ts~���Jp�h�ex
����`ż�8�Mh�C�_ՈGut��Kgm��bIC.��s�B���^�^��k�g%gcb~)ρ2N��:h��)귬���d�Q䞑[SXF*������Fu�C�]1ی`��:6��NX7�tI4_i�dܸ�
�����l��	�x[xk/���3�la�Dx�n���O;B�����1��*�qo�����/��W�l�,Zoy>�9����dVW�����w[�!&0�+�q�L�ऽDF�jx1K���m��q�$��2ԛL��n0P'3��|������#7i���c"X4����巓�L��چ�s�T�f��Q�@褻s�OL;��$
�J�y?��lr���Z��˗�T����"��H��ur��j)�h��5~�?�e��nD4k�;]:q��G%⯋f���Xa��s���2}]WJr1|(F�8
e�~5y���&��0{�d�%�T����M\mR#�ߕÕP�Ѧ�.����;��R��$j�Jm�����;G�Z��@�� �=��q�Ѩ^�VWI����H%{e��a�e3Ĳ`���ܠ�耲����*�$O�Q��I��.i]^w�(�W�
���ƌ�4G�K��B�Ǩ�/��jC�!0Hh1Kq
���.ېX������O��RY�`����w5ύ�A`9�<y�zQ��n�(��	����t�*�P�TX5�$;��$T�U*�2��iG*��Z��+FBoϯ.$� ����#}r98c�O��g�m�}oӳ���9�C�˝�E�DiQU-:�n�?�O��0�Z����9c�g�n��jK���c�h�����z��`y�?U����ѵ�b ��β>\�nP
���J!
8����7�� _�s�E\���b�~�W�ͺ7���5�(�@�+���%��|\��c�a�-3��ĥk����â���'��H�b��&,gh���l^���ig_H�6��)u�R��;��^���f��@��Y����/tj���7�u�csӔ��L��	�F]�T���H�}�]��"S�W�6D�)Qe�?[5���8;}�Eɑb����Ь'�����O#w�to�vm֒��u�3B8S
ܲR���o���Tx��F���_כ�Ӌ�� *}�	r��k��P�J �rG��k
"D�6;�?!����,� cUP�����IA_z`�z%��Hg�_ڤ��hg�)�u�������4���f���W�!���C��ث�9�Ş������(/���v7�zp\x��2R�5M�b�_zDQ����ͬ����^�U�I���%׺V֕cG�}wF��|idHI�W���r!N�K�Q���Қ��.o:�9��dkN�׋x�y�ţ�/쇹Z�R�r���xV��*�T��)n��/�ŋ�s m��Ǵ�V3ň��hi��;W0@sJ���ux��^��F*�Z�mC�m-|�A�)��"����ڞ�y�����1y�KyK�%�V>Q���uG7y�9�}���,Y�Ӊ�Z���[?D��t�1��=w����8i�_Di� b�Q$^&~����h�[�sQ�mN�\/�Q����]�Y)�/�e�S`��Z���Z�td�tw�N�C�-��>�+x}`e�iǳ{�+;�a�|'ֳ�;�NJ���������'T�^0[R��,(��G4���3�v%��|� �4ZچS^JB�Y��.���B][�}�i�)7�c���}M�e$�������C����C5_M��J�k�A�V�d:O���� >�Aȹ��2�R*兆��f-��O��"�F��e�::�}.�h�aD5�63%;�q�ls��� 0,P��Jy��*��(E�*�`��7&���mҪ������X���_*G��;���waе���?R��$kx�,h�C@%$*�[V�]���6�w��5��������˹P�wR-�l�c�}�t�iN/}���說�'���aգ�Nr�}�v����©2^��8�C��s��Ba��3�g%�k	NWj෗O~�x��I=����d�Ɍ�j��J�E:<ۼ
]�
�;���^�O�,E��;A�����OZ����%~��="j)Ӂs+��Y�E��ܸ��#�|�%��U�'ڃ\�w����b��E��ݮ�<�v��s	k��a!k��oO�$`Ȝ-����)�tհ1���J��ծ�*[LVQ/����l�钇�}��`��
݋A��d�d�h�Մ�c��r=��o���y� ���|9��@�������b�j[�H̞�a�m����b�T���P�>P7�6o�Ǣ�u�k�������h�٫_l`g��u�Y�&������%\k+d�U�����zH{f�n�,�_ ���*�6�^������LY���q�ma|1M��L�`�^�7�f�L+2��@�lH$4so[��q@f���СĘ�UՋ`��l����J Hx��Rp����A�)}b
�k[�����l�7��O3�+��0�H���?�EeE����4�L՟l��:��	�e*�`<�W���rE!\1y-�y��ԯ���
�gP�����^��T�b�8��	I�Lj`B�A%*?�QtIʚ;��h�0��<f�~�̡�+��Dә�G���Ž�FBFߏ�k�wf�� �>���|�O��E7��=�2�k[(�D��_ÌL��&!�;jJt�{�1�~v��=U��y,��aW�E��^����6�s��C��dZ�?`k�y�u�.X�)��#1;��)V�V���󗈄��P�i�%�%��ΞT����~Zդ���dʏ���d�q����=�M0���Ἷ��^��7��:TiG<����zn��,�r�X[x&�S�a�}�Z&�i��P�˵��^~V9aʜ����4��$���x�F��9x�Ē�+NpVd�	���i����ܖ�V1J�meN���:÷ؘ��#���`U�9�/���1�D�����0�J9��N�����%St YV��pX�6�Gld3���PtHy���dFy�.���x.F
�.�|.jr�
�d�Nau4�� td[)$�^PęS�Lu:V�p�D�͊\�5�8��$�K����(�;���v$�l�ׄp/��z��>�F&�vu��Wh���K���MM���A�6�ú�)Zs���ŝ�t�����+��G"�YzWU'���6�:2�z)�wЀN ǈZV&Y� ǧ�p7-����Bob#։߶'� Y�K���Z&���_\sy����N�h�����ǅ�XX�/خ��$1(�"�;��>��$d�e���N�>D��9$2ճ�9���'o3ꕲ"p�k�ȚNn��w���v����bc��N�E@Ђ��hwZVy��[/	�y�����&��0oIy0���Je�1��@�	/�0���{=u����f|k��]��ǒk����?MG���2�@2�� iA�	£��謪���gɛ�G��L�H�l�a��40�v���V%�g�1GeN�fu����G���WS��*����ߏ�b\����\6��3��dHR|�f��sދ���g�����cR�^��J)Ӑ8hN"E���n�d��=)���A���mjJ��۷f񵝁�0�;0nM -ɾ_*�,i�LAWU���wyQ��2�����Y�8u�� s㯚��d��{�`����T�ݏ7�C���R#��?"[��<��L���f�!GbH�م���]
���+W4����0rJ4�7v�w~���K�u�q"uC7.
���)�6!0ZP?O�\�3M�9`�j�]����bZ�w#c��$$1�8��P*��,h��v��MV�D� Sr'2R�W
�^�WZ��ž�C�I���vƳ
�.G�����^�u�5m����f=��̹�1����2ҡ�ϊ�X��A��ŝ��{�a��.�X&F�6�C1JooU���Ǐm�d�ǎ ���O����b�>k���+w����ֹ:�Ȱ���<M$h=~�삽�i �Y"�5�&N�qL��ƈ�6�d��~Ԋ�1�	R��cq�8P |�MT�ws����ʄ�Q5�)?d��G/�G�Q�*}���o5�r���l���9�cw@�kX�B��D�]�g�H4>�}���[8��C�y�flq�݂�	蜚�����3�3'M�^���%ؼ��;Q�?��P=lo�fn1143�_�yg�f?����YO�Bn�9��la!u^�W�q�L��\WbX����<�	8r�r����F�=c�����&��5&��g�{t�je6%��n��˿�*!yQB��S�4[������4�[{kq��8����XTP�š�e�� ��5~	d�VVX�����%a}�K�]2/?P�������z�-�i������;s���L �R��~ۊC]���G�Y��)��(i�8mW��1.J(Q��������T��R�6
XV��1v�jS,�����h�n]'1�����&��1��7�1��kICV�uL|*+�5u\K�K�y)UWl ity'������UF� ����>/f�x���5Ӗ�y�I���[t������8�9*�y�=������mp8Ig&���*E���o~���T�����rH^��%�Za�Z�c%l(n��3�o�]�]J�l)�yQ������L�H������Ŷ�ɂ�������:��@�-:AA��vF�ͭ3�����@��_0l�_`n��p�qΒ��=��k�lʶ�}�M�\+�NsdG��R����W�j�������9��R�	6�?m9�`툟������@�k&Ȉ����0r=�N��8\��mE-�"e쪃A�{�q�30��C�����jhy5Q�i�G�ݢ��d�@t>2h �xr���Bm5cU(d��s��;<[dj�D�f:6܏'�>�x�J�4���>I�Y��"E�Pq@�_�[{Z�y̛���g��[v����q�D�Э��;���/>�W�BA��3����q��U�$�� ��U����Nt^x�6ue7���T�ɺ�8�(*Ke����i��+�DI��G<�p{�Fx>W��؝����F_o�o�PR�� >3Gz%���9�TTH�vH���
k/�3픡�wz_��b1��TbG_O���sE�vb��?ih���!4�9+��?k�D��� �qZ��vĦVU�� W�����gk7�81�_"D䕗La�~�Psa��,^��􌉕���VnXr;����:���Q�Ϸ��Gy�/���vF��n�d?�H���9�$w�6��?���d����z�GC<)&C�9�K��'c�؂!��ꌙ����������^��+����SV�
�%�=\�y�`k9�ƫ���Ch��2��bLj�#�a1�sm�ٗ	�;�d�O�$����"��(�2x!��~�@x�)�<�X�������M
��Fd��:g�^�\RM�hKԷ}/�]���*a���eD�zP��&v���y� ��M�Q���9� v7��U�.�#��+Sn��VS��W��&,�j����ѕ7_���r���xD*�.�s�F���Z���)�X@;����Aoa�_�t��7�V�A7ٽ��E�%��������W�9��3�$��/,~U��q_/䘍�ͣK3SEp��\T���Y��9v�f���fp�������e$z��8^�h��a[�T�`a�s��r&8��tu[PN>ʳL�����h
�*I3B���>�@B��q���u��t��?�g�L�����S��I�m��^�3���R�k~��8|��xk"7#��S����,j��|k%/�?�ϙ�7�!�4$��O4�U���t*H��?�0���h:�}��̫牍�\��6����.(v:S���j���:����I�ي��n׃x%/�m�_�kC-l����t�/��쏎f��dC$,�X�d�_K���3u<{���s�	�*������ ��E�Ae��T��1��(mO��Y H��َ�)����4�_��L�xz�ʔ��o� ��I��O�7��6e��

�ȡʈF���͊>p��Wrny:��Ӄΰ������X�a�mF�O���I������q��c.D)�S���|ܪ~���"�<�#5�5��j#������$Gd��}�8n0��ǙL��/ԵtMVf�R�	�%�D�a�;���?����%JXhؑ��<b�����ݶ���$��;ټ�C#-^�
�Ix���T��L��C�ZѺ�w�ҁ
�5�&��85�l�H��Z�$Ҍ[�J�G.m5,����W|f�(k��y����医L�� �FF��_2s��I5y=i�A���H�O���O�ab�\���
�ê�:H����ѵ/+��/�E�w�/_� eޘxI�Ʃ�v��L8���>s�E�`%��0%������ΎG��E3W3 H,��<2P���/d;�|�P��K9H��>t����QhO�K,���tE�{�}H��2&�������o���y��V�0��V��5��}=N��aŉNh���*S/���+_6vE�kc���q�u�B@?x���I�MI�daQX�)�H�D�zT�'�������)�>:o�������~�,j��#��s�Qҫu=XF+m#�Rh~�����_C�L�ٸ���ޒG�vw"JՅ��El��������
�=� ��M���0�7�	�XJ�a7P�nN�Ŵ��K�UtɁYd���s(��T�_F�q_�9i�x��������2E���xy�Zѓy۲��.�Qٹp4�S���Q�������\
F3cD[uW�cp����NT���r�_6�;ġ.p΋r�+߬<[�5��̠�c�{��9hN4h����8�ݛ#�IS"��g�S��H2�ǩ�ƜX�{KW�o��.�Mdh#��^��A�tlO�`�;���%�Æ�ݛj=r*T8S �i-���B�mc_?��kXm�D��jx���q~���y�A&I��#\CpZ$�0�5p�#v^�8Gr�]$�]x�UJ(^�C�i��_~�O�Ĝ�wA���`;����<��wbuϾ��P�y�I�-JWW9�������z������V
����x}��"�z�7G��*`��K��f�w�˫�p��v7��nI#�%���o�ا��38a�5X���TV�ZY���!�j��x���zS�!*9��ߘ��4=}?ʓ�U#�t���~1ۙ�U�<��-��\7�`R�%�/U�d�dbZ��'�ci�T�DM�{o
'�]��e��ِ���:�>���-�/EO�	�[-0�j��/�#�)�������}E��U1�T�7��c��_�6�p�F'>�&�5��%&���x���z���_������[��L�P-���~ n��=��9^\34>L�zHNu_R�[2�q1����Cm/�s�[���$�ۊ���`&�Q0�ɡC��&x�B��e쀔�S�H�3���~�VLh��߫��F`�i5�/�/��`V4��\��@�����R�������=���uj���ߦWS
{(�[S$3@��?�W�Ix����f�r!����d��
M+Gn���l���%1Y���,sC���	�d�-�>c�'�I���3G@�~��*�"N��V9������w�LG�B�j�<���� ^�HE�{K��?Ů�dKd�^�mT��S�qM��2P|�b����l�-������x�|���r�ed���LX�/�����i��ܝ�v�o����"��Pܿ]۵��Ñ��}�i+��+u���r����7.�S9Iv����@F�Bv�vd�x�ټ��Z��B�Ej��7�G�YY,(��8�:u��ҧ����w�L��t�P�n��I�v8���H�,�� %2��l�A��gӫ�*%2DL�z�Z����Ot($~��b��G׳;��ߎŉk5�m�7�?���3+�~�3��H���E������e�Q �҉�lX7׋��'_�$�۳�� ���V3ffS��o7mT�N�e��*�L���R�lm����m>��ٙ,~��검Y����MHl��,dI�Vq�8}C�p>vd��Z��\Q�!�����^��>��x�#"�z�Q�h�X�@�P䃄+	%�ۇ֓}�e#[s�٩!�=���Y=���ĐY������g�!Q������~������(00���(���XtW`q/��Dkk�)b����Z��v8}�Ӆ ��.A��l-x����������.W`�/���\�.����*mj�٠F���}�:�ఱ�޼�b@��zF�M?v�:&����\�h�	L)��
N��2#mj�Jt���a�*�/)A��TZr�˪ؠ�K:l�qC-��7���6��w~�~�jWZ	$�4��#0����ڤ�B�B��$-�i �����3�*'6���<�P\?�8�4���1��Dj
-r���'.�M�⇠8�(�$,�IF�3���\APCX�hYg��!�8�����r33�"��aF�'�`V.��/oś���]���I�c��ūnw�ff����Lu��Yy�Jɞ�Z�����v��#��_�ԬK�k*�l��Wm�;Ҍ����/�������o!-��	 ��Ù����|�!�Q�>��Z���a�V!���2�|�DwH��|TK��o�Yqќ,K2�zk���m_�a�{��n:�)&�E�#�#r�[o? ]�����%��7�[T��o�Ƣ�^Y1A���i��]�Ze"�y��>�H�MЛ�Ğ����}}�� ���P#Y(NMm��}x����JT����/ԋ4�n<ͅ�e�Tr�+@��%��b�?��������W��V�wn����|�g���P��a*E
2 ;�`C�ϨFB$�U���H	�z���Vp�v)ɹjE3�-jZOa���
��a� ,PC�wUO����
0>�O"�PV�n�V�un�"�^G��upiD�#�q���2G���{t�jDD��(���)�g��U/��͊J���"��ss��Iy�H$Н}�|�K��Qy��.o�ŭe>uJ4N��J�W,�����#1o��b:���V�7
�ӑ���0e���	!��tU����M�d"}Yd��C�G���+M��kUHBP��KGnW���YB5P��v���@x�>�|Vb&(�;���"�T�A*��	d!�%Hy	�ܝ:j���n멩� ���K�Eb�\��"�F��6%��C26{�! [���ӀZ�DϬ�L��@�J�mƬ1�r�n��]N1A�����`x���q���«(Z�wk/MHpWY�8 �]1�Qy��<SI��)� aCtb�<7V��k �@a�՞Z��7��h��7.��|c�!Q�>o���1�y����l0e�.3�ٹH��6�?W��~�� ���b�9S��<+&d �΀���,2x�%��u�Qw��<�_��n�Q��#��o!\v��1��;Fm��#w�'&������i��N��L���p���LH?��Ky����uMLi��/j8��ǲy���p�~:ˡ���N�i�Ǯ�E�im�w��$ `x.Zac4|v�[=��j{}����.icYFJ��!�s)�5�1Ъ�� x��^�X#ӫ���ņ�A����^�a&fk^���U~�U��%��J�Օ���<�"�%Rm#ѧ��s�]D�oW &pM�;���ko�C���8�m��GO)g�y�,-Y	7��7���;�^��}J6/�������ޠ�� ���f��i�Ѐj�ed5� y%<��جL�z�ljUY"�E���L���Yo����Կ�w�;��m���k��Fn�"8��9:B(��B��C�FÄ���A�K�U1�O�z����$5�rfe۴[�`���B�΅c[�WV��5�B���s}�a����Tqu���7�)
�r}<��R�G[�������kr�q������$�W(�rh��)�i�X�e���{*��:����E��[�g�����mup�SB-�)GQ�_O;ۯ��t���(4�>��y9�t�L�]���)00�j��g�ȵU	� �}5����X����w�M}#�Ë�N"8��&���ߜ�4�D��J��B�#�Q��g�Lt���K��+r��N����
2�vń�]�H��v[T*�)�L�`�RiK{���E?�6GI�_����;�j��|l��ٲ�@�vRR�����n�5+�eZC�H���xSr3-(	������̄a��f�6�����-�$r���Ԯ|ƙc[���_v+�~[��=�k�m�W�V ?���?*��sq�!�*��1�k7�C G&�'��NB:jY�{t��*T��J�F��U(xCU��Zt��ߛ�㜐r�H0�Fv��
�։����)����c�5�ۯH,�(��u/u��E��ӛ��%°:��PA�F��e%�N����L��P�wU�fZ�?�(�u��1�7��,<���͛���E��'��[�`��b	�8_�&��V?_��e"q{�|��d�d��d��"C�܌�N�,oˋԑ����`��1�6
�8��Q��k�5��H�Gۙ�<�����M׻�\�YG{̏d����F8Rc�$lj��~��/E�K���� KʷY�/n�F���a�#��;�E�EG�uߌW<�,qĽ{[rZ�?irP���T�;���F%VDE)��0��ۍ���o
e����j1^�
ǅ�k�X�b{����4N8�!W�g�N3�00�8�tr��h�\�M��AF�w��},�*pe���w� u��M.޸J����Iss�����Jv�O�@�xq��<X<�J�x�8��:�R�R��uxLfꝌT0"�)�Yr�^&E[^�M�q��Z�گbEr�?Ê/��R��J ��V�078���>�|aR���r��!�6���)����J���^I���#D�,��AxDQA!I���9<������AR�ª	]p��������9憝@��NM��-H�/ �����\v� `�����g��O����(�T6	K��b�p־�70uπ
���� �����٦B�})�K���0;,Z_d�v��4)�A��g@l*F����8~P�GN����(�$wYDA��~M��Г>�x�3dȂ�o�3؀C$(���	��W��R�}�V�:��O� �9f��'�kj��?ؽ�!"j��	��S8�����i�-2�G���0�������v$j%z�|�pc(uӛ�C���eIo:��N@r3�,$"�K�}ゐ�Wx'��K����/�g��ˡ8m�%���o��o	�/ ��]�&n��pL�C`��M�/���y��D� h(�&���͎��]-.�<l�%�5����sZؔ���
�n��H�~kC�1�Ӳ���J�D�6������9#�-l �U��v�jK�{7���rU���8�1��6�v�Q�M��}y~w��R�S��v�j�+��TAl��=�[d�q��X�GPn�9�co<���}��H�� 9H-k�����y?���isT��D�<P^��að��)�W:�a�w�
s^V�sO!���$b�J�su�����PJ˫��4ڟ[q�	S���Oe[��\r)f'�[��]N�S,R�A�����n���D�~��O���G�1���=.� �ᗖ��+���ȑ_Q�R3Ch���K��X[�;���W�բ4#����=u�9��ZK�dݤ��Wo�_����7�)����P?�~��4MV�j�a�I�P�MO�����?"(vdw=��r:��ca���,j2�Ƣ��֥89pƭ�3��ނ�f��ls?�P����YqO��>�e
���ͻ,��b���P%��7���:�9~�j�=T޾&�k?�＋��UG�F+�d:
��5���G�w����Ty����T��W:^��ĩ�*_�ۮ~Z�<bJ�]X�F �@7t^7o��y�a�n��f$��m�
A$x��'��)Pg�ǀ\��=M�
ۉ�Ik �o��y��GZ2���R'�	(�]D�Y��и���:l�s����8�~cY���r,<�]�T�����:�r�W/�0�:Ed\%��'9KݸI���4� �;RE� �s*��~��Fm�?����\��"W pxSUwN�����Bvټ�v�j�w�P�]�_n�md���H����v���+����g��$[F�	�]����f�������R�6�(��x����˫�Cz�Tm7�γU�fp8F����1�mFH3�E�̢�w/3����@��'�K1v5}�"g���#퇯\n�T#��ک�T[�8�F��\ov��+WU����P)�$�U]Ғ����/
iu�f�&~+���>��a�?�"���+��5֏,պ�:�V�E�-�1|KIFߪN0�Q�p8Oki�E�~C��n���Ƥ,F����a�?_��&k��I��	o��,����3�w�Q�(\�Ɩ�'��Km�3��|>�B�[��UTJy��J^p�$}\�l��B<WmM�@ੑ�H�2�ko��= �O6�����r�W�3*t�/}�H�@4	�v�*T�s�(���2�*;3r!XӚ�1�i:g�2�"J�����ޯ�w��Hp/�|�b'Y2'��ӓ�C�W�+?k\�]�W��/�=��?�.��:݊ŸӑDG9Q���(�"C�hK0�rk7�
�>0��2��X/aZ�>�����ۛ���a�žKi���Ǻ���������Y%UdY}�T`��(kf��Ϡ�}��4��b��C?�6d֩���d�?�OW�Lt�ߞZY����ȸ�.}u��n�?>�X�LƙS����YY6]9}�zB��?~e�T�� �s�K:����B�����qr�`["l�ME���d�3��6��KG�o���=X��!N�ֺU>���JMZ���V�RU��!QZ��>}�V@�;MԚ����N�5���0�s]��l�L��)a��j�lظ�U��Q6*����6�r�G7���V\�c�i�`�sѺH^�34��C0_����u�@`�Rr�V4W�v��@ĸ���-py�GF��%J����Ç�ݼ�5� ����F�p�Y��5�{��(1�=�v��\�L�G�N<#����Ie�1��b`��C��&�n���fS�}l�gڐyT �4��xb0,]'I�ru�.��wF��{s�	�������V�R��$��]�BރjAP��\��:y�}~����SCUVO�م�1˧��m{v���eQM�{��t�0_���-�^aS�e1֤2��0�C{h�_D/U�5��Zq(�UR��=/*�3���+"�\��ݫG$6u�hx���pV�a�����Xqz+�t�X�O���|��S�f���O�=KK�Q�.��p@=�%1m�`6��c�S&ܑ#�/8�O�j� ~�4�@�3�f��)	^@1���Jb����2�[CO��4��  IU�1S�d����Q�̍
�˼�S�g�D#c����*^c�qO��{�c�Y�$���	�H�`d6=&()_��A�p^���:OJ|ݑk�n�}�i�3��ʱI֬���b���^w:�X��(=� ��́�=�q6�ؔі����~,_�v��5�z��;s^�Z@�z�C�&FJ?��	T^��8���"��\��A��c���29�6,� ه���CLSH�j���[��30��̃'��*�J��u�x�T7<y�M�Ǯa��h2<8�d�U�����z
'Nk��y�zh�3���ϊ��$F�_�+Qv+�T���A��X� ����%��$��`?���W\��J���?�JM۞&�W�I�_=�s��@�z���blF��i0�=�{g��N�w]���(��m>`����s|5�Y��\\�M��E���J�r.�M�h{�r�&@�����	Q{���Z)�ře�$�޷e(v����-�	�z�L����nl��ߴ���/�Ұ����K��b����h�Xa�<ߠbzl	Yï�ڴ�f�:����s�P�n��~�SHs���_!z�8i�\&�VQ�6Y��0�G��{��r~f�\�.R?�Gʱ���&�g��`O�G�਍/�zO#E#�ve]Q�Q>�'
%�~AB�~�	}.�~�.�����Vt"���j���J�B<e|z1��tIz��S�F�g4R��+/QhrhOA������x!�)�b�����!$����\��u"`���^ q�D�*eo>�"̹r|�9������H�#w2tnr�[�C�i�Gȟ��+~�5)�j�9+����Xk@���ߘ���AS�!�SF܂�������#�V�K�����og{[���7-t���gi��i��b�l�Z�k�Q��c�w�H�X�'�_�(�dŀ8���+�@�i�K���k�9;�P�s�J
̣x�F���-^�)a�����-���@����
�X�R#
���-J�?�9k��QCI.��� �g��P)��I���"��m���^gT~�D#�èC�Цw�S�"=;��K1*$ˏ�C(^(�G1��J1��p}/�R���FP]�Е}�Ur#>�}u� u�F�5(涖�	�Iİ�A�tB�	㺬v������N�N��Ų 5�8�8��B� Ȫ�k�C��$0���u�( �9x'��Ƹ�:p�|�:~�'Q��mU�˳ �����8�'�Apy�r�r����m�����l�E��Iw�]�G�E�"[��ͭ�~@�b7�D���S�j�#�a"���6����B�	ű�#��X��u�1 �n/ 9[ګ9�X|��ʢ����[� ���-��ζ�Æ�'\�������p�����ߥ"�|	7a��e<�Xg9g�(�����&�_�����%�e1���k�o ��Ѳ��W�~���T�p2��0�7�w���U�`�I�|� �9�Ѱ�FR����Ȇq�>@���y���:�ݺ�A��[$�HA�ai�0M��k����ES�>\�������0"���1�U����\"Ϸ���X���7���T�1?7�� v9�����H!��H:	����챚ۦj�������)�bȮ��17}�?�W�O<z��]> ��Zu���z���o!z�S��:u� ��������p���~�5�h���i��f'G�\���+�Pԋ��p"��c��p�A����3\=iْ �TC���w�UFy�-�x�|�{�-�y�DW]���3ҽ$��}�z���DT�����w�>�bN�RR�~��Ma��)�~[�����FEm�/���2�K�kv�OTk�����׫�X��ct���+�c��v�DfS�^���P$������a��8M���/��s��$m%H�د�w��)�af�4��W�Hb�U�4��%lyP�
w�,��<ĳ���s���9%�S�Ϧ��L���<ۮ�$r+�T7�6�}d�q?%�����e���LZ��������Ahְn+�,�b!{��z}N�2�9�X�A=Ҕo�<|Q�V5V%�sU#�Í=�U� ���}�u��M��c�"1G6��I�䱬�CF}�s@Y`$�7H�?_�Bi��j�oB�
�Ar�+���T��}}d0kns���;n�(ri�X~x4��O�*f�|�V��RU� �S����;sz4�cG��D�.[ �L3w1�G^�']�Շ��3��+��T�^��Lb�|�1�E#D�X���uIpR��_���!5��2"K!k�3UPd�ϴ�ݽ>������K8�p�:ʰ�q�(��=Z��2�Q��K|��� SiR�4����Jc�L<�iK�y�]�Y��C�ۛ�/	��Ky�J��M@۶n#�}:rrG�L������ְ�Dvڡ�7��[��F�cK&r�z�)�F��r�
��1�ɵ;�#m�"G���v_�sҘ�q۞S�䍨����sQy�Z(b�wKk�ήN�&��ly�U^m���q1�nĬ�y,�B�T5�
��k��h�ѵ��}ݯI�]	jf��O�y��RY�_�w�k���w�`�%>��̯�)�@��)�ʦ��Q�e,��γ:=��#�>��A5m�ᑒ!��;���p�!
�D�Wu�f"�
�+S�mgBp�e���I%&؊&�u+�^S���F�A�  �=�X�$̲����g���˲�ʪ�9�#�8?�i�7!�0k^�4��������U��_�����'n(�3�G�C?�����_���>D�=�v[ރy��ͽ����]5��-���KK�N;6��#䀩p�F�M0>�l��x�]�ب}=��ȑ-��^�1�.�uG����&��qBPn��G�5&D>~�D�nZ��E�%3�����\��zD���f!� �z���O%�q�貜��X?ϰ x[z��TSzl=��zg�_���;�N¯�׫�`DRaZ���Ä�tk��Ug���bD�#��*�.7_��$˖�����(�?5U�=&�)��T�����'9̇ ��l�]��0�������;�Y�=��*�Ep�~hv���oOf��o�"�j|�X��e{��L����:��C����72���?�����"��̎ӱ��[� K�c�3f,`�9��>Db�E��Y���z�kI	�Ԝ��?�?��ux1ô�k��v�h1�?¦e){�wu�]��S�q]j:ۉ�� ������3��ϮZC
���ʚ�rk.�/SRsQ���f�&�S�8UJ���g+Ìk���Ǫ︞�`%���)�$�
�+<dj%�Hδn��6��;�(�F같��1��H���4��8�L�<>�]��E���E�4�vy���!��oY�ې?�OFQY8�Ơ!�M���A?��!j(�x�XBYS>�.p;���_�K ��G�B��e˔�H�,m�9VѽJ�}�k �J���L:�2��΅ 0,y�COp���= }rڸ/�$�>��b�'��lʘ<���(o���_�~��.�ޖ�}�<�茘�_!�(R\uޥ__W�U�h�l�����^)���]�O�h�=W4�U9{�����u�\�ÃP�f|ܯi�"��!�G3������ա���N.�q���9��v��m��E�A�l@TZؘHvl��.<*E����,�4t��Rٗ� \�%~��&��Y��&��H��8�*dJ��5Qgy�1<�5�h
@*� �8+����u�ba���(_�|�DzKUʗ�g[�PW5�*q;�v��*3����w�b�c��1Qqc{��`[�$1�VO@��{�ӹ �+�2���H�$��{тE�Ԕ,yd���i�p���A!?4+35_/-r��9�~Q/�6M'�,�����$;`�=( �~pB���7b��ł|�x'�E׽���Lܣ���3�iV��i��K�bvx|�k�^A.�z�z��W��
Tz���Z��L�9Mȣ7T
���R�#����:olW*��;���V�:i)X{'�u%T���4��e�%���#�Py���7N��4�����^�sk�ޣ�i��1�2������i�ھ�5���3�8�)jb��V�y�݈ly/�ӛU+T�u_9#��M����5���G��i'��� �p�<��Wӻi�J�<��>UC�)�Nd��|+��ϯ���`ajb��PZ�}����{(W���zK�d���Ыz?�&��N=���<�)�������ʆ>��X�6�u��8����c#���ۥH|�H�9������u���c/k�\{�5���V�%8t��D��b3�2H�����*���(ԁ4�i���%���y/��(�Q�'8#��ւ2j����=d��A&)6o���6�tJ:@�];o��}X��������ψ����a���y,�9���"�(�%\Ä��-H�`���jQa�l�@�u:�����]�-������Ñ����͍����ّN��Nh�S-f,)+^Q)3~� �Â|�[����W��1)���j�>���y!ԛ�vD��L��yD�T6���o�b�VoҺ?*�4�׶"�!�?�(R�Q�#֝�lx�LM���>������@�	F	�u�.c�#�����G����ӈ�S�s�(`�� E��EUId�j�k����H7K�n&��b-gB���u�6Z�|Q�Z����U��DsӲ8S�R\,OA��Q����b��w?��ɠg`�B�o�S�\�Ղ����'(��)�K�tI���BZ���<chZ�������h��i���v�@0�,dO7(O�(�1t����"��)_��G��My�]Y��)�i�uڔ���(8�]���24g7n� Jdir�_���x�{����B�2������z�)��l�?�D�s��oC�0X��R�L���T�Qшh�����X�H^걤��o�­��ۣ��jL{�`���ƞXyU��+R���,6G�����}"]����WU��\n;�`ß�Gב8�#�Y��:u��m@�}�	4�fer#��+��.���MX\��&�6�8���O!��z���������3�|
|j	�|&7�a+�``�0�;i�WL�[�pl� 0��Ņ=�����?�~8�cONW���>4.S�����Dc=��5�9ο*�ˆY4�Ǖ����ލ�G��	߱T��_w?*7�R)C��?zWT0�V�4TY�%�#徶Pq���v�I�n8�-G�M��V/q3��Z��N2&��
h��-I@�;�D��~2��qO��e?�+	��OG�8���m�I°.>8�5�!B�����gZǠ�������R.0@(��3{��w@2s�:��&W�֑K������o��wc_`Nأ��A�r��� �ϵ�^�p=�H�wSƘk<-uk��^c�f*?!�mdw�W[�'����
�����z�B��?aը�v����z��Q[�u���@�X��9r�M/����B��[4�tn�|yg`P��X��Gzڌ
�L��S�d�����U��b�+�^��~fx�>HVr��,Qu��M�/�)7̤N'�)RV�|�܅�ŧH꜡(lZ��NՌ�]�������r���m\g�B��r���9Z���"��|Xo���s�3c�� J2�ڣA�LQ�N�l�E�@
��ٯ�zᎬ��^����XBܮ�a�L�W��}��_-�Ɠ �e����i�i��Aab��S�\��ÑS���_�Tk�Sp�lC��6>	%r���
���E���V�Ip闎lv=��W�K?�6#B5�Xp҉d�����@��=�1\��~^�WCS����e+k�N\t�3@Eŋ���t��\WS=p����X��Pi��~���V��d
ѰT��;�8�]�j��3�
�wxG>�C�O`hhR�<�	E�+��~������&�9F�?�1�6�55��WX�tc�X84���5�"��2fz���Z��A�IN�>W��q�yuo�lC$�tl�nMQ���*=��i0��_��
Z��/�f{iO�(\�Ng)k[A�.��͹8�|p\���Diw�\��Sy�DS�PN�
P[Ɠh�I�'7�+G�.�����0�G��]!?�I���[�%����L(LE(&��k��O�븑.�~:�i8�(���1??Z�"FWW�ݛ� ���p��f$Ԛ�-���N'!�f��1�\��	�q��/��]&3+d`��	4��jK��ф��(���av0d�l�����kS��TPw��)���T�����f��Ml�*���6��E٠����5��u�e��TI������y��Y��΄(i�2�#8��$� v����Qҋ#���J"�q�Y�1<g9����0�?���~�`E�1n@���z6��B4F[N�ݣ�u�NG	�ޥj'p���'0F�f��f.��C��:T�O�&��<gJ�;�j-����CN�mga�rj���$�c�3sߓ6�b=j���~�,��o7~ǿ͂��#m����@?�L��5S���0J��M ��`?e��qHcE�m��"�H�h�Ɗ���u�݌�(W�]q����wvqrku1Y,�0��c2���NS:,1�~}ޅ�&\nA�0��{��egt"�11�����lMBuw�zv	����['{�4�%f�=�����?���a1*t^U��x�+0uQf!O'jk�T�*ղ��*]����2󱕿�r��2z�>��GLFF������@����ҥ��Ɯ"_�6o�7y��Yڙ6=[��t3T.�9t�q#�f�ў����3���ѣ�qa����_o�H��'���o�����D����A��0�cF/e�R&��$�i��y9\%u5�I�����J�w-�B���z܄�/u��#������g�=+ٮ�b�J�4�\X���x�|\��z�h�t8�d�����ʥ�u+�����Tǖ�m����x�ј�|�QЦ��K4�A�I�*;`V�v�w;����z�!@�M�@�v�����Ϊ���%�'ާ�űVS�!�1_G�J�F뜭��ZǺx��J��?����ز?�7�x�ۍn�"�Π�9�p�6�s��O:�I��؄]�*s��q�V"G�Q]R���޴'c�g����4{;;�t��
@Rn	L�n&@l=�?A-��zVk%^L����T?�(�ˡ�-�wx���	,U�*�>�Mjw8�s��7�(`�Q>�g��f��]@�r������/��$ٛp\(�ې����O��o�hqor����k;2����T�����|)��6�[���B��]#AM٨[�/���w�t��ɶ��Z�My�Fz�}�<�CN6��>�r�)��Qz�� ~�I�P���S46��D���Yޝ�J㝇�BS��b�_��1���بs�3�{�`4���Qab<�P�t$mVJG�����;�R?�`��i��@R$�@�A���>p���;<��)܁3�k<�"iC3v�}�ΩA���7�n
���9�@�Yӡ.h6�-h��Z��o����y��k	��N��پ((R!�oh�2eX� ɘN��<:�xfq��N�$�ׄX���%�7�a�C���d5GHwJ5�z�ccVG�\�9���\�u7�z$@:G�wd��%0}��=~Lu��=�rZ}�D�j���K�Rr��s���,����?���P���˧�$�yk�������bf���4�r-���տ��j߆+��d�[��)��&�XӦ=G^��J�3M�PCC1��9#m����TY�j��������;�ml"2��q�
��C/��&��i���S5:�Lx�����kTLR��"�x�)�U$�;A7]Pϥ��5�z��%�g�weC����y*E0R$��ef�,㼋�5XU��)>r9�A%�ho��8n��_�I\��j�o�$ �
y)e�zW{��,��,�E�X,��|~�t|�
�����6D���}&�Ќy�,��X���㸨�0�q�H<�Z��H����˓��c���)Ϳ�A˫����R�2J��V��-kY��9c� ��w6<��8�:���$�7�I�ٟ1�����Ia�	N�J���,8�d}��6�`�m�W�+���?ĥZTI
�x�k�u]Q���4�0p���D|*;�f�T ⌂���Jt.���$�d�e��Q�"�:z/b
ʸ�������Vr��p�4��D]�\̑��fAhL�8w��Ȧ跂��nmT~�w��Vd%6J{���՝�|$B����h�B?*Z ��e��'Mw�E���wئ�>���.�A�Co���i{��r[|���6��o?.`��Q�UG,F�ŧ��A�M����X]r^-�����ɬ�RX�r����c�����e�cv�G&Q���9�_�~T���6��aT�5h3���1���'�{���k��#����\C�a���q�[\��W{yd?a������O���� ��P��ˠ�x��ĸ:��"d�	�}�����ޗ���Q!���Ɓ?��B/�$�^;�F�t7���ZQ���:.%�͕#��G���m ��`�kv�B���Bq�h�z��pZ�X=xG�4:�����6QӺ�E�RN��-��P��*z�2oFU&��;&�	�jT ��g� kT�+ �p���Q"p	�p���}��fn\7��}�ɚDŌ˷^���BRh�,��కW�Z�D���w�?Q����}�]=K�d����������.��Cj�����iy����y(U�]2]H�^�o�h"���F��JE���zO&�GN�$)��������A�Xj,$\�:�p�dU�ĢJ$ �:M���ԡ�u�iVz7�]J\��c>z.cBUӓvz�z��tj|�p���%� `�H��Hps^����n�/��q�먓z����#����l)��ş�b�����=�x��g�z�_3��8���D�h��.%F1�W�w��ޝA�!_�_�HR0,{��.�k7^��?�r`_�gK�p���,�T�ҊhwsL��;%��u����\�bح��R���}b.��}ZoVR��;���Z�}7��_ۦ��S{�e�%�)�P]:�����7D*l�W��v�j�L��T�8�(0x�� z���C�5X$��^��[������/�Q7t���N�0�-� Y'Z�r�v�"v����q�J����~�`g����e�=V�e[ֲў�t�h@�����������DIO�SEV1���?���#��!�GL>4Fdl��,�8�"����uJQ��H?���;Sh h���Ve�D#�vm|{�V}aī�B��{�u1�_��m�����h�Tj��vV��J%�"8�޳���Vvb���6�� �("Ǚ=���߃�S�U�Vg���30p�%�J2�������
1]=>5e4��Яq�o��*݊8�hjH�"v�)V���C��>�0z���M1Q�c8e���#8� Dm�?�|�ĕ����p �P���|�����$�.2�il�"����g\�*hԪ�x�t�c��m{�u#�,��z=@��D������.�F��mƉ���Y�0I�V-,Wh�)�3�Ϻ�{�1�{(�%�M�lA�rEŤ}AFj�"*j Z�QK5��ה7r2�W�U�`����0V�D�{�G˕z���?w�&R����_��N�u�*���|]a�Wx��4H�%t��@Pto-Fr3��?�tH��uH���c�:�=`�c�0���T����U�
��9�?�++�u-}FXL����]�5� �3^�(N�RH��P��X� Zx�S�^C����6���5H^�byܛ.E�^s�a|nF���imX�):����&���k��3��9�S
�.���cF�X�nm0ӄ���c��w&��� v<G��~��{."�C]�Ĉ�DPo��z�����n� >��{�㻷�h���m���=B85R_+���Ϧ��T;��=�M.���R�vw��(X��/i��2�kID ������.y6�J�ֳ��Na�g��s���pq�f+����	?O��+�&{f������̮ZQ
��X�5T�54��|o}Aͮ��ȵ^*K��_"�����x(r�I};WVG���Y\M���d&)	�p0L֓K]�~��� gi~�;沄yF���R����k֫�Cӷ:e�o�o��\���*|�R�~5M,t��/ a �uLi2�����o �#N �s����q�Z�>,�K�f�^�[�WD�d�*Aadf���P+�6%��S��G��T*��g�r�g�&���C�f1���2C���u髭/X�\�&����"n�葉�%�Y���$m��8W�>�$�dj��<��~<��%��۲.�H������xH���;9O'���>�N�I?�Uqm�qy*Z��/�Q�k���^_:�,�J���ڄ�,]�.��0�/(���&����My���O��� j󔠴���)��D�FV梨�z�JCz]3�^cxKK��&��Т�g��b(0��mH�F^R�#��kk���}sv�����h��Y�B,R����X_�V�'���­�&y/�A ��h�^�p0�|Q[�/��΄@M�l�8='��{��Yb���-�p"+ �뷨{l�J��}ے���}��+�"��E��b��c�K���N�}�&iU����$�&� OToJ��7�ј?g�Ҿ�ݺ�l���Vr_��o�^�F�c����n3yv�������׿�U��o?��3�ā�j���Q��J�5�S����L
�����r��s2b9�����|E���]��N�{|*}��t��jDTdp��������>qI/�O���ʇEҞm���C`�rR��wl���ѷ��p
0+�4��ͨ8(QE�eF�k�wqq
��ӑj~Z�t�>��d-SO�-�䨪8�^o�=j�.2�owBE�+{/Q"��'.��b�h-�_��~�����>��x��ꌻ��L���e|��A�S�3;��@�]�L��J��H����]��?��H<���RwOx�V�}E�A�N��;�\T.?I#B�xRvNg?����8^G�Q
U�JH�=�l`� �I�NM��-f�����[;M��R�Q6�K;\�Qv<��[xo��Mk��vX��_X'�^�r�&ǾyY��%Ů�2�X����xgk������+�XU<�`޹�M�Lh���K�)��l�� ٰ�\��tka��|������uʏ�/U����?����7��D��/i�K���9�!��|��K��1r>❅S�S����	�CJ�U.#\�	�,7*0+�e�r&	��og��[1B/�\%��`�y{�JiE�S!d�U(Kp��d�آ4��n4QHt
x�2��ٷk�C�M�^����Y�l�d7�	l��t<R�\6 Ln|��$�f�o�����R�� l���AOY�M |-�Ü��o�''�F���bP�������FnO���~`�-�U��!�;��'��ypf6p"��K]@� �_~S�b��s�� �|[�0��3[�yB" �h`In=n��sL=t���`����ɘ�>�a�\+}G3"#M�`��j�n0�.o!yH�ělK�$��ɡ��]��<��eKA�
�n"�H7������33s�����ڂ�K�[ʂÛ��87@���d����!�)�IM2Sn#4^����3�x�+㥽�˘�þG�����B�Q�uF%������F�,F~�ޯ
ĂköT�B�CM��Ԇ�I�[������*�b-�l�kN0�;��l�����
�HkQp�� �F�n��@�q�Z��c���� ������z�`�p��P�Tc�ž�y�ĽQ�9Q��%�vp�!�hK*�ܨ�i��t@��Q����o���Lk����l��k�/����(��V@q<@Hh�N�\WPLV)wD�7��pP$��y��|��r�%�^- h��V����>�8��}X�;��σ�L��`S�΅2D�@�:Oߐq��;���Z�����/�8�\�ecⲞ�Yo^����Z�cN��t�m*�Bd�ɘZw�ygU��Q&9���.⢐�t/�䜁�4tv�+Ӣx1���?���qZ���k�� ��zϯȐ�?2�=!ձI[�k+g�UZ0�㩖�� R>��o�X~R��O'�+����D:S�qo��{��e�-�f�D�t�%��ݱ�n��$HU5%�&�� �Fv��$6���R2jz�����	�?5���x����u|@/S�����Ooi����ρ��L�*)a�����#�r��A�c;g^LDF�m=�٨�"�:b�9����U��"L �U��#����
4����#'JC�V[F�V��_k��e%!�?�����0��:1g���@���M���cSPwT�YH)���;�������qu���<�6�mԢ:Xm����9��_p,|���!����$��LZ�7�*��RQoή�*�w')T#�����CdI�maxdʢ���D��wHdb�0�y�fB�9�OF�������[e�������N~�\�'i�f�7)��|��N�c�K�� 0@�������[2�)^=i��ӧ�u�u,����c]z�L���&�I��']Tx�xp��O� ���y�Agշ�%O�,�����(J�d��y����J�[�h��a/�[l+�1�J2��s�[Kn���5{#.{�u�_W��s�xR�����g��Z�	~V�[Q�z�Q���["�X;f�8|�D��*�=����1�9F�5!�B�q��|6'v��3x�V��<�VQ&��Iz�/5�G�v�gW\�,����|T3���U�D"��P�gc���S��Ts��J��!��4W>'5)�D\ǖ���x�`Pz�2�զ�m�k�mSXM�F=s���z7�u"r�a��f5�~wȩ:MQ�v�\Y�vyRnH�C�BB��%����<E8z�ʆ)t�[��v� f����v-" ʱ2�[$��F�)��FDz�.�,=�k"[:�`�X�GH��1N`���À%�X4n�:S+�N��&6�4\�4�!;�{#G�G��5!	���T����'#x ��?מ�C*��v�(`JB~����m��L�P�Z�j�/�����[W{��A��/$�9���lg�}!?�5v��*�lB�P.��ɏBVF�)"t�T=hޠ�J�TOc<�V(����O��j�+ŷ� t�P�V���"z!�]1'1�Vݠ��ng=W:6�;�j8Ld9���]U4W�7�.NQ�s�R.Z��D3�~%W�x�t�L$����;!i[�����lr�
T�9��b����qӒ�ޞP+�9�P�ƣ��m�����[R��O��W��J1�~�3��38Dɗ�bԯ�2�7H�}��\e�cy"� 2�L��ؿ��m�������� ԙP_�>Y��+l�jۙ���u^~��/�PI��H�,^İ�PVl�|P�?Pb�C�`��W�/}\��')`0^�2L�X�)��"Yk�q���:`��: `�H���E���Ad�|y�7K�GPY8��2�|�pNb �um�D��@�mRo�t��""�V� �oW?| m��V�҉m��r�e!�g[S����'
 �����gd�Xd7lnՐ���c�żJ��@���lU� 
�i'/6ٛ��}��uQph�o��ڿU���w�݋��m��D�7���ؚo��Zu�N2�u���^+e�L�����{:�����`Ќ�D(+|?k$^��C_��˛���Wsbm��ȡ
��7w$�_�*����E�*/s c���h��N~�Z��!yj������_P;y>9B`p���l�Ӣ��%�S7�m�#�|l����RA����~y��#.$���T=V���A���� 
��Ⳣ���t��rP�0���3��ĉq���-Zj$��K:�d���`L�}��t|���:ΐ��e��A�%	��ѧv����{��P�ǜT���5�G��������1���L3r~#���������\��2�����-=Ȩ^<�&)m7*��Ѡ�%��L^��o�N��h��tѠN�I��ds\�Op�
�9�����?��CV��Q��k�ӫ��1o��k�W�.<m�B�a�R����xlOY���2+%-:�����u�٨�������h��K���	B1���o��Q`g=�r�L/�8�)n`��v_�F�˛3��w,@,��9��lˤ�N��"iv�Ŷ�\?iM��Y|ީ��섆v��\��PD~�����o�dM1'��W!�N]���p�T���;0�����9-�e�e]�9/��?���E�� m��<����c�o晋�����돉p(b� xŚ1�|�B}^�g����3}:����	��,�Va����a�"i:���K���kt(�kS��0���0��8{~�M�H�K�"�kcOr�+ަy�����aT��z��D�����)ob�m��Z��9}�7�~G���y�h�J`�����>���|�|K�ꎎ'�N^4!�f�t�N�+�O.V7��gj��s�'waY�Ͳ�� 4�	�w���t��c2&T�/�俔��Tc�Z�d��S�lX=�����#�i�y�����*�SݬŒ��5��l�c�Ä13_�lԿ~�-��Ap�2�t�ᓅ�HNa�mY�y��k�Q���E�@ԐN���1�~�.V������ہD���6f�e��e�2�]��ӑ��[G�`�E33�ۊd6�b���k�#�l�վ��&���.�|�L����WeN���.�׌��
Ax�Vi��角_?4'���q6|�F ��M�`�"�M�������@��&W|���T����7�8z�������@��\M	!�����𧓞+��Ld�� ��u�3�kz��g�U�(��,�(h�ID�QЃ��lta�J�HU:~��ɰ)�L� �#6?\��Z
��\��K�o� ;H��G&HE�U/�iݛ�kw!c�*>��rS�^t�!�V��&{�f���:�	�,�V������B"�hm��CW�K$��@���C�Vz�H�N �L�tW��r�r� �������:����$37�Ƒ��/q�:���=u��n�Z��n��ծL����!�L`�s��3��{L��p������_�<P1x"�_��g#������(���&
��7Z��o�cҧx僄x�����j���4Ƨ&���?��` T��^��֮��"~����q�9��"2��<d]��G�o�c(�:m�Ҏ��jT�}�d�{+xPϳ����G�Xx��38U�<i-㊲k�a��2�j���g�����'7k�P 2J��#��u�S�'������ގnR��JG�-n�b7d��X�	�v|�]2{z�����hA������U�pΦ�����I��� ���:����%�)�Dt+���k���?HW	��p$yx��KB"n�����|lô5͒�bɄ�u�P�LCI�:���u�`y)I�7��۸�܄Х��9�k�^��s�R��p|	1���4�\	N[Tᒩ�i)�x��׏��U�"AU	��Š�w*X��]�e	V�]7���f���~��|1�z�/�Y���*\8b����B�����FTP�lƇ��%r�RK�����Ri��-m�τ���Xt�u%�n����I�1-bƀo#4���:A�����N��W��I��O0����C�5���E1mv��ҵ��*/}:�o�$���:��ӏ�y�~����UV	B1T%逼*���A�X&�8s<,7Qu�������Y��7�צS��i����V
V񷳸<��ru���%��J!�~���0��,���o�]+�;X�c���9><ǂʮw���!����r�w?O����n5�\L=q�I�31�����L�*�s���za�T��4¶�d��%��, 䔎M�e\00s
��o�V��街���s���^*�=͢G��&��x�d�Z,�.W���ТȻ���t�E2�5�L1����g�|���j��K��S���?r<�B���+���$|��`�W��J�f��P���������x��wo��9��x�Ŝ.�ԎA�c���Tp����،�O�Y��Y�#�o�z�u/�򣥜�7x��9��NawW&�2 4�Ylf�1���3��t1\T�X�b7-�نq����uU���G��p֞ +[���;.�m��\\	*������b{X��~A�9)S�})�ᡧ�O������+ ��gxG���D~l�/�I~�ȵ���¾uI�]_�q�Q'Ν䀎5d�������*wV�ۊ�L�9�����R���ןҖ��O����h�<�=I;a�b�˟y~s��N��9�dg�>�S�,i�э�*��^�Q( @�V���N�[8�l�E�`�K"����k���	
K5���G�s�� ��6��Sjn� ('��rȲ�b�o�Z�Km����»�CEi��~3��{bX��>�ǹ%X(]�#�R���#���S��S�6��;�f�n����>QM ���<_���^�����Z��OE��8��Ͱ%�v1¸ΐcOQ�
�V�
�ɉ^�W�ߜ��ß����qL�?"tk� ؘ��!��5Bu��.3؁�����,���ߌLw>���GX��ׁZ�9��mwn�C�h�b�'K#%���J����rc��:��WZaO-fn��t;��^�Μ�ip+}f0^4Ӌ�)�w���V�du:��˔��$��O`G�۴�Ab�����wN�ZW1��?����㰌7�1>����i��}rx�`/�&�Q�H����5�_\T6����0-���Mмʚ��7�z*@��!搌)tih����~��ё- Y%x������
�1�d]9�N���ꗃv>�_�8U)�$�b.�kO�����J[�>�A(��tU*�=r�.�����jt�;����B����Bi�ܽ��O<FoUu�*?�-����!3XUq�n���3�\{��u�g=f"�b��X#�'^|��>D� �,NNa<6����2�V�P���;q�y�(%�2����G�y�<q���{$�{2�a͊�\em��ѱ���-&Hǭ*��Xc8�a�A��!b��N"�$���!�Zg�[L9�8���f2{u
�B�ђ�}6���7����0쥼��*�oh�0D"앑1ҍ�ߝ3����R?'���$�M��l'�����;G��x���b^h�܇���P�����/~�;,c�R�lmf�:�̏g��IL>���ڹIY-�@�6�/դ�1���Sd�UD���^m��lz$�����I�I�L�O���_A'@�K}��(2UX�F�&� ��#qo�w���m�:���g8ߎ��*V6'��>��A]�����3`N���55��Z�p-��%����	��mI�#�p�T\��Xz�N�M LY��f�V�l�v�
��P+��՞3bh��ә�<�&I``1�9�ʲ��"	�*5���^�еߌ��s�GW�P�y�6a��ǎ���v�!�-�����}�贈n�{F❓\�9�#��̈́)$�þ��a�S:1^�ܫ���}���`��()V�4��}���;ܢ$6=���U���o +�o]C��S������2�>���0J�m6]��0O�}HD�R�g�|�u����Z�'*�c�A:�=V�"ޙ�9z��(Jr�i��d���8��R�`KK�a�_�	�Q�>Q���Q�^��fDult}��4���I Wa��8f�������*Ģ6��3&f�G��
~I���0*��7J�ʕE#�C������ם	�'�]k�옝����
r�j�lK>~�j�U���@}5��q��H<���4h�0_P�EJ,�	��A*��݌�'��ᲕhD��N��vr8��S������h{��<|������Ķ|�T�
��ю�Xξ��jݏ�f?���QV�,��[E�v�LNN5YF��wu�A��|�ZY����`b�f=��B��/jzA�g	�x ~a8��Z��])A��L���<Y�ZS�Q�N�g��� #P}w��&�06Fj���1�0Frl�a�W�G����B߰FeDR�l���q���S
zD�̠�v8v��|܂y �^O�C�L ��mr�����$�ʟ<���2�/
(
N.Dd�!3Y���Z��K@3���Ȍ�n�;T������?=��|�+��)'��S�p(~kDAZu1� V��L�]�nU�u������5�O���W�4�6�Qm$�VS��W;@�K+Mǜۀ ��_j�� -d��(��k�!CyO���E��V�3��3 ��s�hҝ�f�<��$ls������+��W>�mdE�9ޖJf��^����"2 ��6��d�}����V�4�q/ڕ�_��x�������s�1;�u�2�+��#5���'K7�צ1w-�Σs�gw�p�t�\�e���c1@-�� de.d�s�u{�K=~��o�C��|��+oP����Q���HȮ5�zuϦ�+n�lda�.��^T���μETpz�y���>�(���n�ɶe�d _��{�P�)�"���nY	�ȇHM�����!RUL_-�*�9�0r��Kwv�V������N��)Vv0c�7����vN�	���ȿ2?��D���8|���Hx�#{�@էaW�o��p>�qL��i���sԺs���4b�(�çW�iA�.9����b�[���kʵy<޵T�V6�R5sa�|�j��#hj����d�d��!Σ���<�Ku�[���6�(�(�gS�_�9)�,�k�T ��o8�I��e��a��"M|��k��K�,]�G��8\�z7�.zKo�ϊ�[����|�F�]-'�Ϩh�v�ʾF&��QZ15iζ6����gn�ڪ��䱅�M6}l��2ʃ3��3�#�+
�����c; ��c��Ɛ����^D�3K*�׵ҋ���?�I�6T���]�7A_��>� _�a������3�=�&!2�s��c���Ϭ:�ի���:'��xy��C��\Ѣg���Jmy����ӗ��
��`w�tCd-D���]�����g�؍��������j��}�]�5O�)��	�[�k�a�U���}��2 ����X�+u�����+Iv-0��=vT�Y7��%�C{>�KLp4�t-o@c�!�7_�>L������a�
��Iܠ1IZ����L�wyڝ���.17\фH�W�[��S^���3��F��U�?��4v^B��Be��Ǐ�Z�ᤡ{k4�o����H	�X��c�G�R�i|.�)j�G��Y����_��<�����ݟ�t������V0��(�&:2�O~q��sR�j'wp�q�A:�
�
,�U��#�;l�"����=5��`g�Wg�MM&��$���]�Ug��� �h�p��!��t�x���Z�M�@�-��eP�f2��Uk;�'�b�kZIH>�#��?r[?y�6�M��9mr:��H�'�&�*E?�^���9�mM(왪��6Q��?�~WY�	�|�qU)��,�m�9i*p��#~�c#y�%��O�#k�q��\����lF�_�	+v������y�$�}�=��>���U�Wy����E�.��w�b��t���q�Kw��,\ѿ�
 �Y�����C��m�t�U�&��}"ܘ@Yd��]k��x�S�3U�c�v¾��QtC
�Y-�|�Pჲ����K/8��:y�˪�$�	��(VD͙���`J���j�,�"���
�e�Ȇ�=�hM�[aL��"דѵ���i���m�6��L��K-��;�H��_şN�}az��;�;�]	�d��%�ۉ��Y�F�U��;I���{�+]1�m�<$�ܗ����b��=�J{��;N%���D��lзI��o8X>����3d�v�_�t�F���Kp(�Pگ�=F'���4�_�g��|�3��1۝Aۤ�$_^�\�+b6�G+|2j(�m�A�jH�:N�>y�,(��?�ymI6ZCл�a�X�{7O=㊞�;��	�+Ɏ\�]=�d{�	��?.�U׺��|#�ֶd}/�D�8T�� ��\ײ3;:�����x�-/������9bɣ-3��2�,����*g����?��h�u���<�D��������b�-��w����U�-Ƭ���K(�� |��Yf�t�vس�G
O��H2�H�
c��߈�6�)�f��6���x�:��j��)��s6�?�ZOg�}b� �(�~�>m�a,����\��L]��������)p��<`�~�a�+N�ɮ�3 ��l}�c�?&���W�B�`��|Wm\ؕ��[�p%9?��挏%s� @/�X�G����u���G�q����:`������M�%z�ť�;&�_���%�0s�ѧ�/��T�K�ޖ뿖fr�iUHJ�!;tEE���E6	���'O8���	���vW����
Vh?$�^;�B(�A�"	2��I�)�&��������|�?u%O[İe�&"F�'���Ѵ�HP���T�7�
1��Fޏ%_���̟�Q����r�s��9 �����DɐR�N�{�<��ػdW/��#�#ץMeJBl��$J�J��T�Ќ��w):�p	�Ί$���' �X��)/�@[]�o�
�����o�����Í��t��U��a"�9�ev`u&�!w��%wx���[�G��U�Ιb��҈�6��q������U�1�>�_���#��3x�\ӱ��gUHM
0�=�M��\Nw�J�*4jČ:xc՘�g,F�T4�|/S���abVs��� ���.m��sePn�=��J�
����_�B����&��DK�ux1�a:t���@�v��t�_1xa.�jM�{�5�<L#�.EMu\�8)>�����ɏ��xս�5����<��U���ꝸ.�YYo�����Ķ9��ұ�'{Ƽw���>�A�0�����%ؘ#��S���(."������;�q�|�Ժ�n-,%����
�3��7�,�?b����@R�3�p�[����[�����$��"z!_���c���5�ܹ9��1 "��6]��1�����s
�g�"����jw-2�����{�Q~�־J�%�-t����:iW�|o���
<SN��lV���r�h�������U�O�M��)�C*}2+�k5i�f���@4N��_1��σ�\�f��O���>ka8&t��ɠ����Q��hIN����c �������Kpks����[G� ��,bOr�R�GjR �)Mp�G쀑Bo�E⡬F�����L�~z�����b�X����I�U@D�t�I0}�A�LE�������D-�[Xy	��#��5'�ɢ�%ד�~*�׽<<ȗ]��HSP\��r�b�4Sz�2��2Д�i�Ɔ?��6@���\��s�c5��;C?S_�?��tL�$��*(�QR�#�H�~���iN��XB5Q������Fϳ@V2�- �6�r٘jWV#��=G��O�{&����PR��������߆L��]ݢa��Z��~�re��k%��Vo��7� ��nyB�)�*��T̼��\�Y��s�vˣg}|O=.PT�&=8s0�j� ���;E5��<�Q� �O>T��Rs�W!����U��}y���{ZB�KUa��p��<�`IQ��z�n�wZ]������Biݸu�S*i�6d��\�,�sL,��a��� �`�ψr�-7>`�cL�ApX�wm��y�)��8����I�D����c�@)h��㖿KPc׻.�n�"?g����Y6!�5�yA1[֩�S;n7t�¬�}X�rx�^��VU$󹜛�KKd�ڼ��։.]4w�?ᣅ\dEEθk=j�4-CLb��Zb,��86sh7S�5�|��ҸM(��Ƒ��˖�Nu�2-���J�H���ϊ��o���b���0F�"[���������mG�*�1��9�SO�$�pHOj7��w�0R�6�@,)�4�V�#����%R'�"j�%%{����&N�$v&�v�d�2[�v!k�|���AT�v���1�uo�P��Y3���r4p��1���P�3��@�{�h�����Γf|o���TH���{2w� X�]��l4���ecf�P�U���&����C��E�6�6/K�_)[<l:�(�t�oN��b`9��ͯ� ��!�zC�X���T����VKN�ܬ��קv�CԱ�����/�nq}���V1��Ǭԙ0L/��)KT��ym{�o[c���|Z[씝J��O�Md_�߮��D��
Q����L:�LV��	�ghoT���YV��F(P���A��5���� gq�?:��bǯ�ҙ�U	n��<�����qC�\�j8I�V��%���b�-��S|zL��@C15�'�|�� ��!&�z=�Ñu@P�(�U��� =�eG��$�o~�Q<RS�BmL��}U����$��\Gm�mu-_��Ksބ����#Ș��8�g3���:�dO�"�f��-9�(���\���b���v&��&�E�ߝ�m�~'+�T��ζC� �{6��>�$�7�����3I�:{N��:WOF�����w�J˧G?sfTm�Js���P<#�f�e��8�!�\#<��t����M��[`\suAF�_�yE� �n�˴(T�օn���8b�f�>B.`���Í���Eh<Y'uT�;b���K�����e���4��5ʉ� 9 q�׎���Ӵ���؈/�4B��l�����T~��辇���O|d�TA��H�u+�O+
VT��}Ʒ�Os��k��<;�e�֤� L]��#�})Dj������E,(�¥���$1�L~���7��e��sÎE�7��IťpɌ��ʕ�o�́*��-%:a�O�����A���[�����=��O��.�%�m��K%�HO���	�gm�.�tL���A�]�wL�e)C�N���[#�*������?+\<2u�՚��H!4�a�y�S��8]�����z[������D���kC���U> ���i|�zny�?An�+��_e(ޠ��Zc3ޚ��O�~7'!i�ޞ���i��d��ϢJ��I���t�8^��b�@��)�m^{-M� +��*�g����+��Y�\�!z��S���ص�v�s�%�į//5�s��iid ���.�WE�`�"_Ұw�4�8`gj���@_t�'����:.��B%3�7��O�]�t��
�v�l��Ĺ����)iM'��$��K�be}SYǾ������lLV*OL^��V{�=�*'�#�{�̜�m(��q�	 ��°�iv�J�v���ŉ_V�E��CWl��������wb���HʐhA���3W[>�~I_��x�n�%ݠ;����蘁�I�8����"�W�6g��ނ�N\@ƃ����{��C�ц߿�y�pa|y4G�iU$X}& F�}���)�K���X0�q~�Ze����.�n�7�����'��j6�}���>3]�7�yص�2RDiO�"�\Grd8�+$h�[݂��x�(%������r�z��4�=�1�7!*��.�JR�G%t����6��Ab�3��[������-?�\��z�*�u��K��/0;�a��n7�Ʊ�P"�3�T���/��uXrE�T��c;�T5-I�]':SqO;���Ā�!>�$���D���^g(5��ǯ}���i,���|� �c���0�^T{��I��!0���_����iM?\�� �{��<$ɟx����뉌��Y~$�?�]�P�F��u��]�4��J��ҩ&�y��}��pS�T,�Sa']�U�1��	7�����S��@b�H�7��뎥Ъ���<5G���4��?�_:��KqO���,��������09��VV�+$�)c�A>�J�rA6٪�e��%Wm��`D������ �Ng�e�l^�5ՁYه�)z�e��y�/�~pc�1�"�Q�+t%: c������s��9�t޲Ŏ�S+Y�͜�D�������5�����Y�d�ϥ��I��V����x2&�ř��G���Gz�D#� �Sy]!�&��=7O�-��>��Bd�>e�e�Ț;��x�l�q��1�{=�["5��	 ڐ��!O�L)5`�) pö=���W���a�-�1o|�Whe/%H���Q���[��]F�ƥi��_ gh*�:�t�
 q �K�iB�����������PJ(�}�LQ�>3��*����bG�Z"� ��:�Z�"L_��5��u���.Y��б@���*uvٸ�߻������ ��@_�кEO[�ޗ�c�Bm.���@G}����s��>�	uu�P� Ҋ��d��,�>�1.��`�g�C�O]d�yG�n��������y��lo%s��r����-ђ�pz�1�[�G��;41��1J��ۨ�sD��ԣrq�cT9Tl�!8�8�7�HA���	�i��w�st�20c2��] �,��+d7���s����4h�wpO�����9�e�9�q:p�!+�Y�'$۫.�O�<L�É�>���BD�V�eqU���������g���(#a��v8���c�Q��ZKěL?��&�~�b��q��x!�'޶�4�G�)p~NOwc�kQf��=p��9�M��K��4^��bN�?s�zz��t��*��~Xi��4�j(��2[��v��%'�ܸ�u	�7���K��%���e��;Ԥ5��A}c�Pg���I��ZN�G�>��S�M=0�#rLZ�&h��o��U��_�zy�0c~o�:����m�d�5n�󆹓'�DӆT�)���`ךS,��[�u��8�T cvK�K^"z�4�_	���79�%���tGFv��bq�y���T�ТC�QQc���!���gt�q���q��]�(C�~�����ru�4:cM��Pb���b�壘U�AU��*M��v�R_~N����<cMe�ɀs7$��[t�і�q�����V bk8>{3Q�Ǒ���t8�9ԝ���Q���1�	��l'�XW��W5��a�_��Y��_� '�e���f)~,��"�7��-#��FΦI��aN�E��]	��h���z�Ғ�p��<�bqd���3%2�����A�!�3Eo����
���鼁��Tj�3θUc�k�p{Z+����a���h�?$k��i�<}� �YB��髅���ߜNA���m������`��l�1L~��Wٓ��P3���-��q�h:�o�v���,��ar�W2�kfd���֠��T�)�Bݮ�x����`g�����	���E��2���Cۭ�nr���\0!Ml��JYG�:�6����.[3U��N]�'	��˝����м1����8L��p3Ċ��1Ej+��;��U�ʓ{�7d���m��9�@�K����V^���� �em��Ž,��g�\C�4����AIG"���?�xd`_�z�����ÀU.�����Lc�?T�J����K n�혗�[��
��������	�6Ӱ�J|&��\�(J]�P�+g��*:c������9wm_���x��
 C��Joq��pK��R��s5���}kVT}Q�������z���R�ӂ�����Т�4!�o�ӅΏ|�9;]q�MN�&
����z}}���[a�����|�~V�Ϊm��]�j��s*�#+9�\ټ������^^�"� ��x���RXsVve�u���%�j��ǳ�J��ct��9���R�f9��P`�D�SU׈0�g����2<XIO��M,�kEc���U�&������0�[�#�׶眬�#��Ͷ5�WU�FA��S�"-�"ެ||���$��pE6�HΚW���[�������:(W3i�RƩ�0��R��������������(՝��d��+[%e�����-�����R�`'��	����+����:VP�_��*AG R��X#�r;���?)
!$����GL�<�0U����W���|.��-�Z��D�bۛ��+<��c,�\X
!�T��w�C�?�
�#�]k}�*q�����e���,[���;Y�;��
�ĳi�ckж���2s�;�d�?���S���oVsj��i��u�~�jL�M�?`�=�!q0��k�:�	��#�����,�B4�x�*~al_�#�B���>��@��|��,��+oڹ�\�Ꮼ�xi�hV��"}OS������3P���9/j%~����%g�Pzn�U�D�y���4��Tu�汼�Q-[�]�j�9�=����Q̴Zg��sh��(n��{4���dI
d5xt��QX��0Y�z�4Oy
!�B�d�Ȱ������2�+�z��jñ]�%s���<3iV��g�SH�������}P���r�sh��� *��)�!{��x�+���詶2�S���PjCb,O�Q����uL��_�²�F)!��_TlFK.��#��k���	��5D��r�3@4�,�+Ҳ|��-���Ѹ/ҁ��w�P'�2�,�����F2)]ͳ���-!c���;��ݔ��a]=�鏼��S�~�AƺR�uϧ�n��SNbl��3��������A�A\}qB�#�6�f��"s����K���� ��˹J��)Q��BT���B2#�|�B�-Vx�Ra�����)P
����XSM��^.�'����J]���j��u�8�����YZR�r(�"U�ŪR����;��a�Ǭ�^^�C��z|d��g1���� �KY[oi=p֜4�'�Θ5� �,@��	���r�P�FW`U^S�����~S��J*^�B�q�.$�0{�T�T��o���WK�;>���m	��'�=�FO'��a��3{�82��JqYJC[����3�4�R#z�|����tk���	�ۙT3��Ŕ�9��3�_"q���"q ���hl�E˄Bq��������x=�G��fK^��s�r�.G��_����\r��&]�8_��'e��>����jo]��Ͷ���z�B2ͳU����"��D��hD�;���n��`��j�|�r�6��n���4.8��mf٠[S��J����b�W:���vO�[I�:��Y�#��/�L�g����~�
��TW[;wS�"����\���fV⸎��!g��� 2��MB�� o����"�=$[qW�p$J)�ԅT���ն[I��x15���v+Z7��Q��f4��c�_�NiFi����l\�o����У%d|�\�s&��'�ت�K�c�;�@A'D���;%������%�F������:���̍~