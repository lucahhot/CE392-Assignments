// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
nDWy4YuUt62eRLLcQlMteKHT2k9xN5dUyIocHe+xsMZUR76Qr1QyvlRGWPMuBdz2
/7uIvWHCk4KqPsPljD/Ucbwb8oJlcGvFOInU9OQJXc7M8kHT0+Bx5UABmEckXkbr
ML2Y7CrhgB5tKeexSpFZ6STdGielqybScNmS7USu8YY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 31072 )
`pragma protect data_block
UV28/HGaZxs8EqzfAZSeZuEEENI86q9IhWfIAyFge3bF1/8QLfIrzKQ/TPR2T1lI
xUxWf8D6eyZZ3it2IJyXzyQoCtECD/M0NZhW/TmlHUoaAKgoCzREAtyTQF/gEPzG
J7FwEb7zBahNvXWls7bc4Lku+jqSw8Pdiq7Hx86/AvLz/UJqv9s8FjyURrzk52Yx
uqhRERO0n5KI7mdqlVjquJU+iHWvYSaV1qoFkWzs5vVw7blfxMWtC9HekA9XPs0X
pjuNCvE0CCYAAgDtu5r9rN7Ac0x+FzvHf+T+VDx6Sos5ta7YKtC4YCWHcTzejwKn
L00zYBUDGsCNXCwFPvoVxam3MOAP6IYtNGfcBrOEzTUghuWQ1+RuGKxpAnYN3fKK
muO3aiSVjYEVoj/unB3VWLSAy3qX7utUUGKcRrDeUIFQqCihzjfWthrR7/UsXGBS
q1Ba9yg5N6ZFMMwquLczhGH6VUI+TftPz2SAtlnPVuLDb9FoPCN0JB9WF7DnucQ9
hA0ZukOUdKWyAgsyKg3Rjfdrl3YzRSlvawiXYHtYakk+omktTts1LNm98zc+uUEz
yqUJJ38ZcFnLVTRxaMt8+/cuvwHLvUvWPMCMnUG494P71d2naZwml7i2Ko+6CNv1
bAHMbkG1Qpv0ujX3+xbzqsK1uRgrQRJAK5u+m/HHHb5Q4jV/q7MGB1Ipmv/TVNgt
Z8GoJFFMU5Q73DIdsy66c0YIwC1pkP6RWOvWbPv9ppfIGLjqJzEGxQsv7x4IU5Cp
gznjWDTvNnljy4EJjq8MnGLgd1+lmlPSqSPnGh5XHGwPKO22aTfGwb1yB1xRxJod
jroZ6DuIi+wubv86L0saG2G6w7HiJfeDGS+5/7tlEMlGG9FDQWzBOkI/+qi30uzw
ktQy6DIS/g5cZQGi0PJZC7iaCjJqdKmIs39szweCh0eixIXWM0JhFqKyo5p/sf9V
fILGKaeWQTvE34bNpgglBhG4iQoefNKEHpEHCKcCZq9tHX5jWCQrnNg4WxA2/mRM
NDkH/xBfRxdXmlgo4A9A3vZsTlWKo5fjuDdW1XKTdJvskB1RQ+hUOZGoB/qxSNOE
/KWVuUNvy3EnayXwgZn/+elc3riQHBB5DBjC7OWWscZcsbxLfjaqdFxbQS2Q1M58
WFzCDWW+ne+CNRcGAKy0QvFR8rSvF5ivc6zTzKS8sRJgpJX+tdmVtx5vUryCVcJM
mNJP/xhdXrxu+Og7CDkoWdlEf+NvYzx3S1ncykd+3hMzg+azwoCn1Lht5BYMwQf+
RHXbF92Rx/YAOE/bQizzSZUfowWPuAqAgeQTXXTFtdRnmJ/2FihNR//mB2LmtyTM
zffJwfxL81xhDMvAlafKCMMGg12iYgKqJb7z9AaOFvbRb96joske4pwJQCRwcRXp
ai9e11FO2VLhhKWvM9bhihXG+cfwh/AGP07uI5XDwseJ4nAu1c61zno3xKPjj1TH
EB0Yxdy0sXdiWyEe629DJSqmOId+VS2pSuRVi33PWwaHK9DIYh8ebFhFQM/qnGF7
+JWnKPLCsDgnUeWRBNez8PFNyG2jY0BINe6uu7efLYUS6AYW6D4GijLUXtASSKfC
RN5PAr5yktJdo+1iyICLommI5Lsv0QFxD5iWu5FiRXVJrMFv047HR85KzxSprGHI
Pw7pLWNMOuNwd6nl3oi6YjeB29NaBel42/qVy61FGmkK63PNSSjQttUNP344pFe3
40QkI908Ho6VZ5hDrmkIDXOPd+MohwgrXEEW2QuU5EHZZeEO05JlSvRyr5yQciZd
deCGSVe+Z14uBPfoL2BRoe3+qWzy9cAGczpNIudG6gYU9BhtroNTns+EWz8FqqiW
I53sbT/lezmci1AvVPWNH7eRv6nd2V+BBMJwRxzeE7p9xQx//A1GLPxSILf3oTLP
DaqCLAT2Npgd8eKX4vRbwORJgcm4zcZtZ4w2m9gQDPOoQqev6+uiRBJHDAxWGgG1
qvcYQxU+DxUdNMag2f1lij273fhrkK0PUti3FZGblnH780HsjBwOKvfuOAcoLgue
V9uW/ayrz9S3dZVaPFegGUb0Tf38ML677viR5l+4cit8M5tlzODio/dJ2la8sDOq
EqHkmOlYjke9/VS532NI5Rs6xN9muLK7R9Vcru0dN5UVvYw2VFDtqexNydvxlBvE
kUV169xHXmSIkT8+lLzWH6nm4E8Jvd6zVRT+c6pkQmHRghIjeTv+/e1cvNQnPmIn
G5XUuuJI6LPONidc7A8p3fMSCuYtfqqqoMykwPfQqdf85GQUj44rKNzzdD18Gfxw
8c4yhqNZgnXeN8emM+JOm5vDJYAVAhl4ALLcnek5VkdD4AXAYXcx3sElbbVO6czM
HCTDdPeNlU20RHCdxFC+i/F1fU5kL2iQjw5yMHJZG8pEDo0pogOFC6a1lEJUj8j1
Kn4qOARjZ2o5yh826fFgw07LPw+WLsbxt1BFrAWhyMNxt24A+3Qi4XfIkTzG3Ivo
kin+4tqpEOHjaXYalVYclPPOzZXYf1vp+HI+CJ1MZxmWTpr3b3AUz6QmWnpeI45h
T3E3DUr3ze5RfL979XuNsSh2g0Wn1QNrt8bbhcZbosDZL3SptbK0l76KQyZweByS
e/QTWqOgIcnOpv3/TT5jZiSaUxBWiL1uvMCAxTRH9tfke0fGfKJRNYnuuiAaw74n
yy8BRUCJx6O+bAzTqwURyL2E+nx1NWaE9b+6lAVnQmDtwEDnmesmEzdBhypf2zVC
jGzvGmW4ErUfJ8fx+Xtd1rvSxtZfsu1sa5rSO+lixP0falJXTe70tVB7Sm8JNU52
yvLtlzFeExYTjVOvSLsaRA4jQBxGtaoJcGGJD/QxL3EtCYw5l77TaHw2llbN+rr7
OjaTQI4DoHaM/EmSjtOaQ2jgKcbmIqcqCkGuFFKLxMKNDgx1H+n1sqrjokciXgam
rdei+vq/oGBC8k+HOO7zTJ0oG0tH0KrvmOhX13uMCnMV9NV6nqqs4fO9g4l0rgoC
aJXwZAj7Cn+PcHNCtQbPvdAvo4BtqhzsT1J0IxwspyBVzrzki2fQEz5jDhprqzCN
S2mQrVO903OUaSWtxy8SUJ6AEesRK2VJjVwy8kbUa6SIs75SxXpd9GGnrzqwOsXl
PFSeE/Qws+UJCKRnleY/JwriMm/6EmAtQ8mvvE3XIMmB09blS5QEWcKhOjmKt2wj
/lDwNPzcN3ysPVuJ8/xImiuHs/5TK6PgT+JRrk/TwcIJWa+e+9nNn5Zl/CF4AKhq
HifasTEGavse1bo3UMnK9Zy9ceVuKemubtTJrxMte7jGU6FZfbWj2TbwhTe+TtUM
wDEM8TeBYM6Y83S4ywwlRhb1S5gXHq5ZwLDvq+xd+1ERjP0Hiwqpm0J2Bbj929fd
BY050Uf/LU0p5IYe8SKmIVGVGMi6K7LQZn9iFCAbNPwFg6lDm8ZandNDYOvbA7R2
Gza/VrP/7zTuM2NP+6XKcLDTo7vqoAhzhfO8i0qvc3795yNY9ChG4/T/NJS4PFCl
J8khb6nRX+HacA9TBcp/6VcnPFRP0ff2B6PvX8NTVUuRTYn/QOepieXPTDl0DO3H
/xEJratGL+FzcwyElUh1HFYqmU2CneX4Z9zJyj2TJh/V1oRdzgtlvhMxAoAymNU9
LfFK7NBMiHy8iVrKvuw88JiunkWE8iu5pOuX/XTn8CjNyOMu2uERMJwdrkDrxEEd
4qpzT1HgdLYr0JdJJHJtvX+BHH094n6FSYl/14zHJpGmvhU1FZizVl49mKVWU9Hm
diwVn3NbfFDSVGsqSfkFNVsYs+4FQVeWpBlmTxK6PMDjDo/foDy9fZKPf3TAU4O4
lXxBJxU6RAHx4EbycKw9ilWoKzj7YG/wkc4vN/0oeu309YE2IA15X1Sadhl6ar33
yBU4IWQ5K9o0BZJKnKT9j4GqrMvDaAzYCPSn6abE5tvUhIRyXmgI0usMKGcppZhx
jne7VhpH8Dc2OA+kwocPJ85i7OFv7Zban5EUDQsAtuCDCWnv6O6vCJKRVb+xGg5i
WdvftAIpSnprW9Qc+49Xq3mPQztKWTi6qzQUZ+9xaFwpumFYq72GZLVxgMr0E7mg
YmFUTRZ+EyenPV4HPNCZN54T/jXpnPRLtEfqdPB6uIMYQGt8xanw34hl7ZJbINOJ
UL4utnR0nhOs5TgTz1Ene26mk85Mn7vT76OPk2nTrRmL3ADLxDKxtavkUv8RD2+S
7xBGEcDhqwSQOBNOu/Ax/BH8Yw6O3z0oy43ESMkas6Bh1VDuOtLvgFgF2LHUvkrt
io7SHaaQzbEHnZu2KCA3xT77Irb0o7hqcGTrpVs+CxxCZFX8uhuYqEpwH+zhukYc
C1C4tf3RBT44I3cl9b8VNNvpjNxMVWMTGab4f7IYtC5w27bOGm/caZVgHv+2Qt44
EPXcLcWAq5NVurEQxiuw4Gg+Cb4iWyF2PSwx3HKQn/m2HGO6seZm/vv+VYEXiQZv
yMn2JkiWaCicex8I+ZHFi3qnnEKpn0+717P4KW8b0TileoRDtMhs+WmFShQ0k79c
CE9Z2I/UC4MtMCUTPDLiYFXY04L4/AZB9aTjtHvdqgFawMiCmWKb0udGOJofhH3Q
T5bbFgS/mrWLNemZstIcUuK4GZguPI+5fmJAIpOI1NczQDNtksijr+wEJgCSHCsS
A6LyVduSCvEi3zQiDFoIqKIZojS08W32Y2iyg9ySh1Y37g/a3XNOF/26r72PSIKy
tKO9e5oS+LBCdXGW7Cj1vCePDc8ssP3NznOasElPJYi4ORdEXbuU97rtakUTt7mx
8q35IAqCOon7F2TPnkgsq6EAPxzbugrFkGip7dAAyfwlLTnpf/FVy8s9J4yeV7S1
4TPmeENTQ/NpFDSyvL0i9YY1pG9FUHz5CVOFYYTCrUWPDceub7O3mLyygfZjXBkS
eb9XVE3CiCYDC3ySH1t6dgUP0izwUk5p9sgEMB8ii+e5n7OcT7XROhReWfBLMsfh
YevbvhGmnJlUQqFZnL4/u/Wz2sZMg4xZIgOgJ3QUq4vV3/Ft/qbB+plwwzUoJXn3
TVNCeJvGD4izJCLXljBUXACnk5+SOolODfnTHOgfLYrXlcKafx+OyfFiV19iynJW
E4AR02EBXnX9LwaWgurMJ5VlRoq/tS1L5dMElmv/7oGKJp7U/bHCF3pOi4/HbDts
yPcyJj7FuPbUmDCxPTHBuj6MquCsxaQFY6XyYyejw62JYmtD0Ga0N4aCWeof4d7i
FDNyYdiwE3+s8YA+v/Yd+mHS462JJLNZ46JXkoo9IE5jl9bl4ouQIlT16sj9qR7T
5IBSpEGXYSWaKgUz2rwkJDRhrxVisey1APy2K4Uzrm7Nvnxxb1btAIF2wRxOt0Ep
NiMg4fX1VRFThi7i5J0jojKqdFJljHNa12I2e16iHsge2Zzikq9kYZ1eTkAxshMs
tMFe0L7rPVTXfGn0xl6q8ezbtjoS2eLnjlk6pRtZWyyY4x6SK9jN5GkBz1xoAxSi
y+FeeypWu5p7araAhj97V4nGPKNmQAWm1xZfaI68sYM4l72byiy9lE5yBl+RlLJD
1IB7ACB5StV9smkoBjB+wR/lnfyvxYIm/mFUPUaBwniKBJQ5Q9krTY6KZAs+jeVv
uU30mwvMc5pQJOfKu+bwenm66Pv47iyT/Me4PktqKbEmswnqRWnyDbi76LPfklvL
ZHjhzMdmpz9TffdYxrXNYF+ZXMLwYD7V63enXsILBnEAq94GweGn7R2+8TROXws9
UwIVYvfRdvCIly+RefbSKHBsQmO8W1rmo1VUmLTeK6/BB7d/63EtIXpAoLotx69P
aAXTjKc/yiQVN0v0BC3rnhoJBZdcChhG6OMhl2RF6MgyLnLs9k77O9vnke/yDXWT
hsTWiqd/Vjj5E3Xeb0beOPVEBPP/hWiwo7mfKk3v/yAmmqTNCf9fv+lYa4gXYlP+
pMaIqte8QZgxSqJ6PedtlGZBNHZ00LPobVOQ/+gcNJpH8ihKD1i2mak0fR2M9Mbw
FmyspehcR6xVUJJ0DgqF4Vxg/iVR0PKvGGECECleiGZzW6roikjfd4jU81p4w9Wh
ODW392zsszwyR0u6YcC1kA34F/fe3olyTDf4oag62a52nRnuSElOc6UDwB/AGw5e
JNhOgJEyWmqS0Kt/i9XwflF6hfiSAz6+x98tqjYVcxO8277HkmC719Ylc+oubpFw
sSy0SbJS8eeSPnEToQOEwB598waQLJ6hi66S/WviqddfJGZhtnCi7bebDjvoThJf
yJyD0pg05E9ZidJAaPXO60O1y3hsn67JxcQi+lm2/V768HIV8r+T2M96uRNsnY69
IeC+5Lp4tupStsYLRWZ1VR0KHUSrh/P5m59XnaEqos0PvM6YvZ1Dsuj3hSiWsLfL
Lshn2FYk78Lgd2GxKudEf6Q8q/9wkpsiX1zFDkOFpV9qqakzghqecnjwcYK6Xmnz
cBojShpJb1rn46pYEYmzU3KYqAfcfFLKtLOp2lPBebxg2L1AYs/sHaRyHlZPcsDG
ftSV2AW1j7H+6rcfYrrbIJwodoEn4hnzCwDTl5VbEFL5e7J79UaDuwM1RqPtEBWG
S3/IFe1QkatHhs8aYWiwacT1zaH8miLkVQ3TnKczgrxbl12/vxg6di4HBUxrrsEi
JKd5z2idPveWr+8zDvb1od56oLjgyqGjNfHgUdPM9Bylw6D12xlZ/Jkl5cHc/KOq
omvFMLymBUge62D48t+HeDd2U6G4hsUaKOkVmhDpH0+YPaInye0tLrfhydcvWOgz
+z33b68tN4BtHj+ASkLPwKnOA1V/Hl9rzZ0ixaWQyDmzBFTeD7NF0UTDQvOD5GUW
nf8DzV6me/uGEnXszruv4oVzBfSA1Tp2Wp1tWDFkSaZEGKssxkVqdN6hqwUcvKcg
eDmnBhnj9N/2TAbppcRSjFCvHmolQzZ5U7D1rWAYCwK2tec3YILLEvi8XRUBq36A
7R7haZPVQh/MHyh/Vd3lPDvu+CmU+3T5cMYdAElI29WdH8O4cjsHkEEjjrpiB5DL
sv4V2Eq82IfQfbg2N70LpUcP2uMDL+ovpbOaVKREoaZ2PacZO9fnhGLBDTtUDI5E
kAG34qEY5VNjUQmdSnXyJutxxUBgpDXcfBC0TKHdaCWHGnkbEdCi0y8ph/oNTJiX
oHBposnNJSM3mxqn6hF0JLlCwEF/wbdgXOifPpoyOE+Ow/LeNZJEOpyBnDoI7UmR
td0ziA5dc9aX1jqxeSFUmesy/nzVAaCY4BP69BBBOKwzbLiHWEto+HxusC8wzsnj
SigGpge33YhS/p3ehUI8Lzga4k8L1jWSBjAY3yOOGA0w5LmDNoa5uvYUqV2mTz6O
I0yCOiO5lGyzLXCyRjzW6pPe8dccsc84GGbSw9dJLjVKwKkXpYC9SXeQjIjR3ybp
3bkJOJI1ih+aNH3s/B/23LgOo2rXPkmxbipfz7kpzfny1okJK5F1RAJV8PB9qS8e
dpFOSFmvr6byCWps1umVBX+JI1g1F0AamzpF8vDYQLai9AIfVPmB5V7cDVcTXuJj
SJ/SSeTjw1kRUQPMJbyAKttxv6TKxhPdpW8Jfq51sHRtnOC8mDo44ySkVEBiFGLT
ghazd+vv0PMpg55b2w/+QPg+CIwPmtTcnbkSHx3WIh4dDgDmNYfh7tLVT7LM1eoF
eRv6J9QC+ML2h4yE3EcoQAJklyv3W/UZxns5ZE7OqgP3aZYLEvy5S8kGC23xJx3i
7+d0WcRPPdTub7ZGaXVLZX0gLeGm4iwEvY6xFpYOrJrlAqsW3AdwSRzeRPPj/azC
tdUqMzi7weyYvT5vN3zXLK+GPspcsyj1tyCFJIYBSF4PajFh+BowA9tDXIYxUu8N
Bc9cb1tLpUbqfJ2flidPr/0z+amRS9Lm7uc9y2qKYR36PEQaR6o5f1lXTTCcKe5v
5HobzbbPQpJodhNnd1+C8/Lt3LlCQr5fi6T7AykNMjWsBVhJr5nFp/P8QV99KNtK
v/TpEgDp6Ict9m+8RzGdn5dRogydCCEJZD8ELaYCStuqidNfgZl5mdBMocftGq2r
khXmi2GltLlSL6Mvwg8+VAULTEUHuUzhC6SVvgXFfrPGyXYoceA4M+YOkT5nC5WK
GvfmvezqmItbowI/qaaePNULOwlKOinqWmqUCQG+hNLF/jbMQZEGMYOIoonDIw4I
Z0XFWqNYCpTAn7L86d1y1DW8mqZ1Pgz9eA+W8hEYZ6ACkRE8RyBipzmmquTg7dZu
kTE70fffLmAk/R9potAr0oixMxU6T2/1MkacXmRQpSEo5DQf6RkIuKtoCjBubd8h
6vJnuWJWHUTucKAlNnVikI3mOmquRwiO2WFBW7soU6j/ocF9ck7ZPoIGDIUmWCbK
R/NcQwQsS8wchpASyyOPuxOpVQI5P00ZulKUxdr5LQY1KxIvX9yfNsDuDJmEKf19
q9V73TiVSqkzdi+3XJCyEpkXmqfzpDyXQcEKnMl5QSU3GXJOQRQRfOip2GC036SW
6XcOmbVykjYlPfwWGEtJ1raymKUIvudEMIZoIbXyirWpE0y4uPl11u5A/w4Nwl3T
0f1YVpYr/8dtSTuzldX2KTuG6DHEzzPeFUu15IPryTAkUEX4DoyXcgvuNhnx04cg
ZahVh0JPzkKzlsnlQ13SJ1F1ZAcw9xA9w65HMUMvXtbkxLIhU9VVa6fy+rTzobWG
7ZWKaFCm0E+5khX3u0MM85WaIQpytIe21JFTpgLxgG7FbxlDj3lZYZFQZQadMz/I
PWjDhVaYapL4i2iSZzsvl9Pxt1Ixskg3L/0yy85eyZBp/Yalu6UKcLZA0gB4c3ae
sqgXY6JQk9nAtV6QxUInJORS+m3vrn1lCPDFkDS03QWFjtJoQUSPMfHRN+EaYn0f
atIjBWN3Z0mY7PFTi7jjNTc3+BsHuFJdVn1OJwpCWak59LpcVtge1YMkUt+Cm0ZK
X7MhptgMtxRVeMimOUxUTZSgW4VvqQFQuCJ1/tP69nnP93g0ZMXOG/rSPkP47DYa
sHWpCwY78vw6W7nG1nL00jCFnHsFizbJxNPgTfQieuCf4qj5zvgK2llDekilwGL+
9F25vz1mezcBjAI2q05fWr2LrU+97Rh6HjKTpfyJespZ3you24NiPAy2CjtT9OT4
2METOzWdD7RM/gsYxHQY1G/FsbUBs0WSKeS2qQN0/wPpK/WKHH6KA4t394bQhkYZ
2j2/4jADkGAj1NcKrps1rMbF8zdYjWKlNKPSc7QhFYsWRTSssdY2HuAq6yug7xt6
DascL3bH/IzlOH9sBBmif1Cb7h+BHoIxPkXWH3CWVOut7hkg0RFXLmSSiN0mWS0X
ZDENj3yO+AV/vN30qUOhr7X2y3Bof0+Wcp00kLFNJo4TrhQF8sDx034ygJ/tpryn
KHboipe6gYjogNHOPpxJZkKhLPyO1lOjXy+yf6Z9wvoafplA0GV9dzvfomq4JetC
2BxaX3OjzNQZVQS8Pk0BA4Ib5hFwfsL8++CnMK+wCMLyqB+joPoDO9v491tQoEsv
ti1WCkYvat0vT9yrJoV1oeydKr/zZ8mBpfpQl64jROFroqKlIvCKJJhkjU8UX4v4
JGLP1ndmBxTteocGXIdKJUvzEp7sMFhJWegK+/nxxJXJQnczmKVEkPUyUDwQ5pFh
439DDTQ2laHEg0US4Xt8WjFBozPfRDMrEHMxs7aD7x9P+7qiQuUhrSM4udv8MYlm
x8sU8tFyITL3Brvyr0V1IdjruiX5Ns557Cboc5EU+9m36eZg/GB0HUxSwntBCk7c
uqzgY+cgfF+XzVu0MsVML2rAPBAO3FGQJSHaf4e8lUuFihWNKdE0PB2cahAXF6C+
IrpQ0rTjUcOiZxwEonFWXT9kywVgbmHmyyPz01Qk+T6NiDf0dAwLcUcGKkMxWEXP
wmkI5STKv4/jdLIj/6rAZly45uB7ooX+7SpIjsTLp/guE5mMqQ0RnfzDH3++6UvB
g2/8rrk2C3EQ6XD2pj1bRZBdJUZAcIwyjR/CEMwN3i5MRyNp3H09k2qp8XV6jAzs
surfcar5J7jZQfOZvNr6BDzVZuloAE0x0ZyLPSJa+dSSfUKI+T4pCGHB/wlKN2a9
FsbdfCYk/A1nw8nUIPyFkoSSntcphnhjIMoDUdzOUEvzWnu+wuA4b4xBEhUvH8Rn
aU5056RBhDkFSNnu0Hv927ZvnCP7YEboX5JeTnOK36pQrtw9MpqpE8JDc2S+XY3y
ZTf9kzKLZtTa0NJTTTNfoCF8M2AF6xFUZXbWcnQniY52/HpxOKIH5xIEcuvAOEZR
zyjsp5VDMzEUDKR15i4sZ4KUYn8iXvVfJ4JJD5FSuv/EuO378D6uU4JIY0LI3Vjm
xzPoEGCnG8l42iWn5OcOwE5cK521wkUHquKP8Ikoi0TeK5BlKoYDZQwHOxW8WMP+
deFxQ6mn99WqMEAzcL/oR4IOxy3g1AzgpPcP7uTZwVicLB7kz1w5P91B9TR/FzFt
J23pj4QH2GMhTlUf6sANVHcwj61HT+iNbu+WQqDNfYuid93L7T9UAE1qFjJ30mtg
eE+bTyWWTkmooGOzMC+mCDJU0soipfMG0/4LnQT+Rry/dCRFFxqWQ/Iigr+qq9+D
0g0CO35zTV/RKg+TwVwuCbjx2ZuDK+P4OmPU/c6lekySvymteoxfyrjI1y8ubdfd
Bpt5NtmbiAG43K+cuzDQHgp8YKBAEwZcqw8XL3DTATkAcS2I30SjuQqf0WGV6jOU
BFDM3dCO6LujkK918uC7BisrGVR1kI0tPQQyBecoSX98hAMECn77OSz7/B7gEWUx
psFicSy7IA4vq74+CaRW7S/J5bRGUpWpnTy2WMQHKxaj9lbhviPfze8FszL5oFl6
DkApyJcRCzQ99NByC2NJrQ/1uIEro2CHEyha7D7gg3FbCIzd73jOASuuP/sjYf7U
Ypw1ldYiVXMZaMCC14KKQgSsDgmXZCnA2NGFsaRLJrbjHTtGsC9+PYDHdlFT+CCn
d9KAuJKJVaOOZFBbkutSY1tRZ4HhBMLDhPyXyydtKzRDe759qKZQQW4DcIuIICpZ
oVf7P+JkjFV35jwz1f36D3bx7Cg5s8jwiIGjbK7o5/ycxkkJ7id99sA5hA9YVwAV
g4VXxQRMl6ZnR17fZOgSL4AuZvZewk1s37QJAitZ2P8y5WQ+EF7PDyPNiLyOC5bs
vrV0htqIZeYliBEudcDdOL8+awtOMDgNaR8wRJqq+Wgq6t0ki1HhsIhR/CHRb6Ou
P39+Qx0CB9XJdPztxUeLrOj2qPxXbWo8Kv7miPrm1uab8YlQUm4Btyd5+Kuqz/Ah
N2zh8U5rueJk/idcRIgCFMTW46LNSND4fbYMbulUU5H+bGs3B1+/W7QITumAFYYU
b+J8sVGS77eXBLYffOh+BVqwmff8jmjTejk65TC3A2b9GUkUH/SKLFKSd4rgJdxn
bg3UjqhrZHnINoY8PBjL+D4HTUbbBUVQNnuR3Iq9Buv19ac6c52SW/A+8Vsyxc+e
vWm3EULEKCPmaltsdG5tRhPmqegUehvRA61Yb9mDevuTpZ9a6oy6IvvKV5Y5LBQP
vh3YkpkFjqsDjL/13giXREYhu/Is3pRMfPA99jCVL/4nfvsIir49VBkXmkdHPyJI
d1zkNqPXEJQlDM93BHwUDJu+UbaY817WsHWFSeBL1tT4EflLDVx/k0EDEzBhORns
xVtElYKkLnFENWyOhcxJzCIpimA/gbjMktSvYTAPRnVNQ4F0MPphRF3pCDBOz/1T
9dcC87tC881i9rPC8kuNaTLRFZi5uZmQGBEZRnxkZE6eLjVoiUM8SuU6dOGyJVLV
Nq6KC1k6p8caQKgyWkwZiBDJouSF4WITu6pN0IDDoGfKVwBEMmDGJkR14iLL9SRs
qv91+3zOgXBd2T6ziADSkvKpKR0rMVnoywq0TPyiTN0FhrwTbluaw61t6PTqzwO0
7d+P4UhPI6W+K2CgnjxkoR7pNVUYB1EUMlzr4bsW+ka6TFNpn9ZgPVPQVgHUe5Os
LjCM9GD3uLT3jY5NIMFvkr36rsF2DMM1y7Y4SYAHxT+GEaLhAbiGCohTTnN1Quh/
pXuOccRV4uX/BJScScFhVoCZfGdLqiKtyGRpynah69p4iGJlNGQlLosKy6ga3zfo
iLkt67ACFD/IWuVi71VQUHjs8vkYX/+sLaq3E2qN/dhqv5/8INA/gY876M0VL1Bi
L4H5v1ADdjX9IaeNs9TuLXra5msnGX9qCkVxx+SW60IRu1GNryKT1D2p8Y72Rhv6
O59P4qgDFmRIbsa5GN1xgyaF36XHzpam+CLmOnpDXeMiDwLt3+QuoxabM+ERQ+gi
nkxJejJFPrTiGDYiuDP77iHd9/5sSqaywfRw0G9hFWfYW3Rjv0jSvkOE3+ssnon7
DpRGdBDoYP5coXWXYg0YGQ7tjd8K7CLWOFoiRu1PYyT8FzhOQx7wPuFzzfD8ExfJ
n14GDFXglJik8RZX9nXeoHvvSIL7aYCDE9f1BYkmFCB1gaejduYpUopLGWhuAx/X
RcMhsxnLQsOZKW/7Qjr7jvKFEtPArVceZm0LFNNH6wmJ/XsnOh+c2rWnMGEriN4y
zwkmOYsECLnUlgYWQpuCqBZKXkGbieexMGM/yXvS2i3yCUdoa17fGXoOMXAjiKzL
S2oyv5bJiGIFjQnKPV1QSIOVE81+bbQ3rNurws3em0WvNfFobyrCfcBOp2TIDWIl
h/2/zdanWDCM70WoIPdtPQQAO0oTuV1VW7CUfdrsqygMsfGMXYi723f49tl9+L8k
+QIFwUBBCB0xBveTtRA4yTo6TSMamSupCvSfG2BuhLwnV64P5tbUFomIe5jiRgLX
FkQycs/wAkbfwuAn5+qldjD6U022vxtXwVsxCZCow8wSo34LNyL/Df9okbmc2IVg
RNn9vL4cC7GpRJjr0bYL1vHb70NhzNkqmyPwioZ+JThXRPsWTavsFKI0B2ycscsS
TKVDmSPUiE83xnOLbKOsPsVXpdnOjqsRwrdMeSEAAiTRPmRE5rPlAgyiqRdGRusc
aEcbPEH7TQQ7hpgROmySqXmhK2VjBBIMzQUAAdk1b7fT0AHIvwP2wFq0jI3vK8pR
+/qJLUBkhUbOFbNFQNrbIg5K7G427EkmlCM+aD3AFP5KutslVY2p7MvVPJXqHHPt
CGvc5qS494zIjcdHuQ/1VUGKWqrNnVSPWmurr8boyryvKgYCc6T7cXuGQ0SW3g6C
GR1MLMpcS2ej/YxvprzC6ONaGg0QDvQUprKUunZsE3R0Z3eMScpsto9yF/Wxuqx7
s5W+8XrmP8dV/J+d/PIlZYGalso6WJcH5YwINfFBEDbS2KvCLH2i2M8hIrTLUv94
BeYrL/lpOTz3/J7VN0xe4tmbzZhhSJZEjIbWPTKqbnZ6munspT5XGm3do9gzfuk/
UiyjQaOhiGSQLUZ9gG2/SgMIf/s4VpHlpp8dNDZ9WKlGQIn+dGdt5HLelWZheGDn
coCe4RrUAsCaZIHnZ69idxE33lQwntWP4P5FP3724ziwnWV+dtyaWMvc3YHGQ/aN
g1Zn+pTovLDrc70vria7+/1lbwdZizr5IwEpsKRFrQ0jY2Oy2/nmpdteDGA42ObU
VTkOisiDtPPtokMYLIoGHIcg8XB1N6Xo/6/odVvD3jT5quLS/Wwi6r/JH7hKRQwg
bo5YsAJru7wwug+NZrNjC5h/5382ThJQH+TmpMI/WvZ1WwasTgyLOHVjABkUO65r
WNsl07tkL7dqwQGpN18LOZRfpAYjehtz4ew0SYvL/kVTZetgdAh3/A4dnEBRWDX6
J0Hc0NWlVg22Jvt9U9+TO4czU9IkDEZ0FW4y9Pbt3ReqY7DmOFdIobJYyTW8+Y2Q
t1fi7IVL8oSq2WDjrox2PQb04oDz4K6+VXGs4Mvm5YfLHh0csLHtZn2KSzaqgLQb
QSmJ5ZxsRRFtkJjcxORR6QPCMif2139IsJbP8n+eRJO7ssK5QIQ2QmHrP2f1YHAE
E7/Nfd1Poyy0AGaVgXTzffCgtS+2nzGLWThoJAx1PILepqTIno627JlTGFnN43t5
2Vs/WMe54yaIiTfBKeZPlSFJhniyXIkek4eP4d/FQ3c5waiznWceSLYQQH0pjiLb
80IjEnMEap7LLKNiHP/O4kWhOAY5OpwWuomgqD/MpFicAx612hodiB+UtReuAldW
rcgmKJqfRDbsZG6xhCqb3bmQJUgEsd+LzltdLbW1tqDQlrD/Ol7AxxwrWrf9trPV
gumvxKthIHHE8bPeznoYDciWAl7i9f8uGy7HONDYNgnhZnpYtDiS9AiHjhK0UUNz
L1NocDV/RT94cSYvNZVUPXunyR2Om+g4mvBDbqTd1wrGa3dUAj660YvqBoz6d8KC
0I5zq23aE/3SE1OS3s1umWoxk1Ly4GYVa4YoCzjATZK30gtsgGpZlnOrseees1du
AXeBPPz1+mD+OQzzFiY2iY9A8gbsKZEyAMhNVEEusrdb4+1Dx7ZOkyf3lWErdypw
W7IxFXjsbrc46SnACcudZZxjG2R9IA4CEdZcBdfwox8IV2K7hq4emVZp5mHoB7EZ
V5ej5i7p7KVemHbrlbFelBbeSDZcLB9pwKLLmMLX/E5BA/xbccYotmJBFKn4L6Ed
Ngb/dYZoOve+Yn7NaM6Zl3NLs+Se4qFRH/tEMfZQ7I+YiGiTmvUJ6+ZbfGcsqIuz
Ig0PYrX7biNdB9EuLxEmcqMf71if1PQDK2ASp9fFSp072p4e4CSRTgEGFkF2NNpI
wPAXY/nVQpODQozi1SBl854NLSJwEnngv7eLbPS/nSFec67FMMxPPw77Kxn0CZ6U
4fu7GhrroBfqyLnIhzHtNxt4Hzj4djIzHDQNVoO0hjQDvno97UBv+nk6JwwVR0rz
nMzB4u/sIrOcsGsjgM9tRrZf0zwuXBPpJ8Y+D2pJrge3bD6ZcqHh2mjTtOYBo7hf
hvqohdqLrNCMC1nfX77yQkor8A/nwFd4arWDurvr7RIWjEXyxYc6QFEoGT0kLsuT
3kvhkoV8S3MD5uwppNxkKJD9dMsLZGpfHIxmUmA+dnWy9eMHPzQZbNt3OrwHodjk
dnB1YqusgE9Wj9qpQQ/MW/xQqP6kUkqy/tcSt1Jzf2F4mUCETC+ZMXd2evBKKmhF
qRpw10P09KuqYyHfhABut39hSuqhWAV4M7RbwVmVUFIQ2FnyAQlr5Fv2uKIawZMj
QU+ZmYLiwXYaVsZht0wu5rIrU4RQS9XRmJZOiZAA4+0NBkYdmTvQQ7EPK7ImPnFy
ycDZ5k5bMOQjt/V0aIUfjAQ0HggGV1esxCKJs8yxdTYc2+5aG56GdNU20RpFs0u2
aCy3zhFVuF3AU7tSawQFE9SgsSBTaIl/uJLolvQLpin1SN6mnGLN8fIOfBLcjlpc
zTx0nVDAUh5rZpSNx/PnOCSFQsZuKopFCAehZUlcfkrMB8O/GwcLZdf6vVWJl1e8
+XT0IcpXVxLdjVOfqcJs1/ZDbgpjQKn56UTHi3rrmNCbJhhsMm1tUfir9GbFJ1CO
F0rP0QHw7Z5X60TyvLRZCJgIYF1DDRUl3y3plTEq1Hj71zNkSQrW2LvtHKjfyaJn
9xzKoX598bfJYEVFvuMm7m3gjOi8u8+IV7XU5mcbaRhTNqFk7vfvHsZCDxZYV0vE
YgYcp5pZkBTVXcIsHi81+fybQDxu1h/Hpy1nNzFnNt0LkSpSGPNZexXjNvNGi8Rk
VWPqPrFIt7k6QP9x4giGPgBPmy0QZFYpus+I8mQyk1pgm7sgmX03D9QDISw/Gffw
wgzXpDtsP6Ef7Gm/E/qv7hxQmn9pLsJNTwO7KQZ1k2XbOhWuE0dAihauesSh61Ez
o/OSc1LUB6a924SIXQ/Dm/XX1YN0d4/UZ4MlZUxsMCLaw5nDeadqUxIr+nN3plq/
3MQjnKgGIwr/zh0Jr1XDkFsbDEMH/v2Pv3mfMEJOnlvrnr/6GqGP/lXTgprxx8i5
R2QJ4lof2F2ksxlgkQcPfkUHU0BvkIIQ/pWrVWgox/b61Z5H1GZGbfgx2t8egCKd
rUhNvclcjGaR4L5VXTbmz2jq4ii4dsZBVf3js7sRJU42HdhguCTbnNK8VKCUstPJ
Op6zPBkSaHpMystbLDq82p4u7/ObHMU2fg4DK5TuYM1dkns+l4bI26gFjxhwLJ5M
ww1QCry9ejXtMHUu4FXtEiMoJLyuZ10KkhODSZk5dzD0zAGZItBRTtYEG12JAsTO
Hjr/nLN6v3fuIDs4P7lqg7qUB5iThFqbfUdCuXoMUO4z53y+rMmarxiUXN3FGyF8
zeVZsEuruITAUZ8BCfdXuT/mWxbEPkoEKTdjG3eXWQk2VXs6dYY9JiscrmYB1REq
BEzw5wyEV+8pStS0za3aUMh2TAg9ZiPuSNa/stwsoPGrHJQZ5+0qAw3snhjUHU6c
tpM5ADmkTKOthdYQlIh+mwnvFceJ3t4QSe3T1qqI60sq1UUjAYFhmmADFEIBMH7b
QTavjUSswpgdMFnhdcCuBTZWQKCHeaYqUoQipRqoVS+gUE0KSuIg/O/95y0ufgXo
8LJEDnozkM2gZoGK8J+yntoIy6d/2jwUZj+BAu/HaJaOhOS7ZESm/i7Dz82ElFHr
kvOlDkWXZF0gnqpWkBsNfL7cvNv/39PMzn+5hzLd31ur1NxVqbZ3BuHHdpgDXJRN
tDTNsd+3K7/0sFXW3cfrMu8s1rbW7g1hvTSjRxtyTdCrUmbvElANJq1bynVKsRiM
tLRHEyGEBhLxUdJCRQCehdFJKEvDPZOgEkPxOsy9Ar1Y0jARw3ZMPHRzK+ByR40y
MrqrEjwHD/XJyf1oOfKdf1B8aGb63XlBQejeEi2heib8Pt33f5Uxaz6ZMNzUcwzg
ik36qVNXiUGyCsjsN7nQQlQZuXcK8nt1+6ToCXtwC393UFaHWmCXRk5cHBQRxNPw
iZkqRzUzmJEW/96kv2jGoCNRf9vw8jjgshfl/ZMpSLKwuG/nv8FqUOcQoPujFi2j
kfJuWGxE2SZ38EpXlnlTvQfQKI9kPPWpTrU1nCsQKGZY/NsHnJXNTkVcGOiYWIfc
vvBKZusp4idjgqA7tm+6jRhQPSgQwtLDvhxDZ03aii+NSi2VrqwbRWkF/MZBKJWB
UwZ69EOWiOFj1yFI4tfFKhL1hQZ/G3AdkVSjwK3wcmHhp3dVDYt18AaNgwSA79ab
cJF6vUd21YvpP5TDaJsubKpHAXx2/mI3aazBHIhVmUUNz4YiWGbuCXFXYZhENU2f
Prb6LJB131tNNx8hOFbqhasBWEAjK6QXl/zwcQq8EvnbauH/yLbmRwbLDTA/oKgw
/Pzew2q3kXZkScOyDkZLxnQ5/vXDaio8SpEdOdv8zwQsASEmFEkd4FmbWQRFL5/f
eqauPT3OevRMlKuSN11fUVkaxP2XtgqhItCYJ6WFWGzdNl4hmC5xWO4sArsrgnvH
H5cIfjNOtEJ3Aq7P1QaV6UrgnaJEW1rwA6+/AUq3dxwoI79J2R7ia6XdbRcyf6Gw
QVgupuCidI1fT8yZuMutpSVcPrrrE5vjJWjEYgTandHXMjkfvt7OYXOKDYcrUrh6
XNii5HsAs49inzupDLaErBthQmTRvk7HfAAAIgtV/vEKLLO1YRG6uN3jABlFmhUE
IdnRq4O+PRtVfT8ZrI1NbNpkKxxTQtHE/WrR++T/zlDQ5xbkgZBkAmIKRQY9YRDW
Li7e9JT6j3hpJwjan/ytY4DPVTYAF7/U6l9NdK9CLAdfeREhX7L0jorPzVODFxUM
dt+Ur6aePk3C9BRAlIOG1BlYRMRZd89WXVMboivSs47HhhSmdWSy/ekpbwGoRleH
wdWFGHLE2MtwSOLAoP8sB0Kkz6rVbXZQRq/89kduTGlb4ZivFzHhv/D8YnMor8jp
EonWgk4/07fpFM3mx6nkqMdZNEYYOkdSGBx/XN3/+yq4gnhwhZqV1FJjTjQRzZsg
R0aPbJxxsvSe3wyAss/S8ipfPRjHkoeooBez9rjwHR62yjG4tjVM/jU3AXiXqWrP
zSugRJ8ZKa37galshW27GkHKpW5ZMQeRJV08NkjXGFWseMSeH/3mz0pMGaYweCvF
IYxXZQehlLFofNTKaZ1IgQWW5htknBZ0wTyCvu6bPTwk7YMf23/EShcqlJvz0UKA
G+DoEcaa7Xdm8zgH+ARUntwEwUATREUhr/4MsmvIDQdIbzBNqCu7JC12zm9aoGx6
Vy5plyWujPfFp5InPB3obI4romw4cL+9qJfikP4sf6ero5hqBQVbLl320Jr/r05L
fRHzmQtlwTd6+ELbdOhRCS1+aZwyXgI0n6AZMed7SrbnBSE21NV5MOBeWEuPWgRV
dxsmkULUIp7gu1zLN6smQccAmVireP44+6Gg+Hgow2S4Ea2ZzcNC7q8SyQnxxAar
WEJndScNeejASuEx4YSMATf7SZgv4HdAMIKugWSp5HLTviDm2ivJSrU4Hf+uFZ/h
u+2QVRxFHMx5LkqaDwC/fhK5sqjr47pM3AEsP2GzscSLX9bcONbt+hItY4kPzl2V
6GaGA5ywhY/LnmFHyZL0jd08K0CdqOlotTAlacPKHN6ZHBDt6t2+CkM4kyBzA+8f
2WDjRYyVXZHo/KLaQmHsiYiY3D9y5WrQxIDVOlAk4y2Sx4KdiZknYw4TnFcBdEzB
BI08aCJwNjQKquP0Fh8+9OMrMk9sRlMzGhuhhxN2f9FqM5Mqy/uIFeQsSLx333Xk
PUAKtH/xYzEL38pv/RYcuvU1sxne1kGJsMgJvnbrJIr2y1RuYMV3MSMwi6egybbG
JFdtw+cMXLLBleJdDn+WQmQ9KEV6mvGCpVwbDyzXrVBnDKdL73jU6EHWssPsldbN
6J9Sb6mVBn/YqsMPaFaGNvDTFxEst+zXDtqm7EIV0z63/TgTHb0bghFsJXPGRhOC
8ZfxLKSm1UjgD1QunAuhar/R41wXPtUS9zPz6vnVMlkw2DU+bwYRqMh/P/zr6sOz
lhdWVeo+E+FAIY/8AUFPmpkePqLgXOlMZwyRCm58RiFYIPF06Zpx59zJl2FBsSEq
EzHWh9ooKX0+6BDLe44EqKBhVnpcJf3BDmpL3OaFQqx4bvyaZsC7HUUNu8gl+IsA
q53E87QgdJJllntX4GVQvDyYjk/JSuU+K58EutE33iWsljKrHF/skawBRZY2aFg0
3fH6fgL+aF19Fq7j+Pl8cTYjzqKD5NGqvmvHqBrGdUVUIrUw+hupyGdnB2XfoyVx
wWYdjTW+Zeo2LcJ3yrUzJ0z5YrRH1UppEryiAEZH/Qxfd3yjKdUFsJ9cgajK0FGQ
LlwAbxXYadsr2NcYUGi8niJvswmxAQ8vrwmT7igCy1fiQTCUa5dyh1nsfljTTn3x
AM+HFMdScYL89vRNyS9fyLxXLA6X/2mbNG8UFA6taU9kSzGBLLdDjzHiAFHpcMsh
NZ3cdU7vVYJQOI6bcMQ89Bs/vzM9/ueaV/OF+nzABaWjnH4d0rqKTSxMklV0o/XF
qfvpf/tsL5QJKNg/DiEDtxkO/kzMljMV18/CzWjvqbNo0rDqPKLYGPRs7X1iqblu
NndHa77z9yMsBHgdDYlcU9//PNGXraDvx2KATk+XRtvcAcH7KmknfguUaVSG7IQ3
3rhs4+6Ui1xDwSTWnjaCP4y/QkdxTKFo5phJltmIZqiY5nyCreQfeqy0ZHUn/rYt
+qLNkOZznc7XzjbNy+tg0Ll0r5lcJt7umI5uHASszvkqELt/oUQbUdkIrE9EADOR
Y2vfv1VCmhI+TieodBBuo+dqhy7kNfqfc9cFyrnQPxtDcSD5sXr8F69fpv6uWEs2
c6C0UmcQxou28Syo8Axu1hw9mFE0BircUnXRxE63eean/KvXOwbLaDEAVKD9oECw
rz5moa2bYD393ZYAEAcxDqH9aZJPluDYEk6mIXtFmF88j+14au4boubauP0Ndj75
UI86JmgIxZmUipKf/obbaSv1msjNWgsjep3KN5ob0lLZBqdihE5JGSm7Bw5sxC2n
nXl5W577xQOSj74UZWJ13F+jdwQp7iTLB0jqMEGDVMUqHXlnt/PPLePVzEz1tpWh
liL1uCvdsMhQiEnh4q9B7JIm32/YltSP+HR0xWqmRAa3eyzBQxTWdG/PEEJmhN4B
Wa4H5S9JZyXnCt2lmfJcAf6T5kJmx6/f/a6KM0n442w5cbBUTHdG5X0676xnmlCM
brZf202T0uqP4+CbqzjR2AObaj09kJPvsdEr2T7Wwl6jEHbh7WpRQ5nACPLVD8gB
6gwgcAJ4BO8aAKusKemUQzXv2RmQwFlfMdt99JHxbxiKIK/NqDbGIKFmGRZpq2aU
dJNB9sBWIxRYnCv4KNZgyZ6eePA0UeGtoO8lxS+REyEeyCyG5993IR5F4kUbBZbc
sM/GlPpRlWWaZuiHheIe2/fUSlhh7/E6l5qj63xEGWvZ69oJ2G6dVSgzgo8uGrs9
54uK2C7gCF/YHkS+ZjifuMz0YfTGQ3Tw/gl5TI8b7CxWMImIqvLSHcFjyrnDpEDa
VnewhtJrJAL10Gep8RAC2ZBjfIMq9bT9cEHYk4g6e4bLAe6VfSJGGBXtBe+R6OG2
vjbRoN7vhzpjgADzZCf4QMzRoRfCwi2k/Kn/CJUK3qa7BKrYvxqoAAjuFwl4/qOc
v8mQAmmdcQz5Gn5Xmq5AwbZ+77WGM3q8fBVAQqGB1dwMUzc4E/ymxGDYjSJzEsHv
qifmVTVqt97KxExQmbebSe8/R4tw1xLRXTnovo/DjB4eZOIzJJPQ0OzAdoq7ey0M
qls4pDkpUlA2hQ77FVoEjBS+Gx9I2dxeo6GHJvIpKY/tgZQbKfoHsgK28VjKNvuR
JWHsy8RmB4MgzUQv6pTM3zIW8U7WPG8M6+Y9xvJI3n+6LvwOnGhJ9FDeJPEN4XY3
9sEtqEpiKMLCiGRVmrmz3OowNuIeMssj/J0ZffM+VKSZWk06hM75wiCKDgSC0MUT
4lBCGod5C21EGAjDel0YBPTikDDynaiQtxCKTCsU4R+SJCmmBQKEViU8fLHnQ5E2
FEN557o+RaKpaDCnqIgGa4EImbHd36tmSy1KfiEHjF7IS1qGZPlbPwMxPIz+gq6n
viBvnRQ3aBnzWPuF0T2jYP3aH8mDKdn6pb2nJFNlDke2bHW+c5um8G+wjntOdS0D
EJq1z0k2c9oE/fvEKgOlDlQ/a7Q9ClENVC9mt6V/+yryMoJYxGgNf0HbL0OMZDI5
Hvei8SVTj5i5gLcxxdvQF/4Pmop6BURPbHHYj899GuSgiJSFOuPjljU+q97ranSD
j/ezoVyZSflX4e0+qxxbQhg1WVziebsbbsdRoRHGmYBew4oUrrUpOUiJGdCSZ6rz
u/SqwkgRdlO4UcbBDmWdNSCpvVkEFzwpP7qZJIlCq4PTCHgGHeStZz4fU/m5gsRg
byz6MoWiTWjHXXuZscrGg4toj1o+cvVBskBkaPdzdvDLnYw+OVj2GliHsaOGG/8M
MxfwJdEv51JPdyWvoHMw7blLFKCvI1SkZ/LEQOIzPN5t/E5Y9QBz0vaE4t5iBRjE
KwJFi9ercdCcU4l5l9x+cLwpOJY947dQ/LFsvzCUbhqbak1ZebQxCC5eIAex4mkJ
KF7TorVLNFSXceHqefJr5KV6gpvYahWujJLoHiYGQ6QfjjSi7IYPtRFwXgCQ+mqJ
gkGHZ+X17PzeTO/yNQtF04Y8XuxtglHVmg5Ah4wkjzg3KXiU+/TYKgCpiYeeREAp
sLkCcx5ULtf56coMonDJcb7nMfjVA58wVQMUD5e5f6d6oNECQoAMQbZOYWqO8imj
e91R4p4BUpAukpeo94WLAVbHtP25RxhTiJzhQe76Z1J39iW4ktT645KN766Se8jZ
mNKETK32bH8gbTE62I3yIotlgnC9FLs4KjfveQWds3jlM/zz1pOxcLWgOD8r6nzT
28aiBuzVyivKJcLaG3TUgzzl3wnYk987rQNZFn5YUY2aty2QSJ7YLwWwOkge6txI
5TdU0WJm0z7gneXyTez3fvRFZ/HkW5pKpVybfT7BjMa/RtPI76QA5bOqLRT7V0jl
rUW69qNanSzudMnCRKQHmXIAlDDBUmSY+HONDYlXxIy5N1ChReauQaVGqytlOSIc
GTnDppmndza1IQictdFUReW8pqaGUIBnLVlIQauYPe+NQLfE+0U4IapGbGNDhbrz
Wxj3tB8mTtFyExO9fmDE8Sp06KHLq34s59diompYNBymrhNES5dz5YQ5GwP176u3
6GFO5cLtTBxe6Hh8M2XOxcGVY+zbe6lpA4kiC8hDpX0PsiD8fWQLRGIFfEMkUAHD
OgiSoUtoDvj+Aptn/dOk35gkWigI9c3clpiabc8URarr8MwyXO54EzWr2Eogt5oD
Yj9SEN5WFA3NXoYWzGSU4gyVGjjedr7uEGhoqCCuMOWHcCuws6CHltt+V0jAOvA3
3OU/ACBHLLm1sZ4Z3qVpTnT/SGOt9au5RzSO56Nf9b2wwpyLXDjyObLXXtlJue3P
x5yu4N1BeZdG6LyMatEFUw/424qLE5kTwcQwY0RkCMFP3L2soY0ZmF7ehLC+2IOX
BDdS/DL1wU0Uozb664alwVH8b5sBiAQ1vyntwvks5C8USZxku8cUmwKWLrTlO9ya
ZII6AqQWEu8+B6AvP9++zab3yT5LNs7ET+0q2f5jOxO4ae8EZzdDlo0bqcY/2y04
AlSmhVA/cn/c96FQG8KJzKWoTaplJBVlO7MjgJrgwOQAbdstS/NRnu22B8zrRDMo
dirlqHOBkYFUIFph82pWGNq2onn69Mn60qN7vUcNQ/yb5I4xm5DJmgZXGtfIg5GG
PPvPEe+onmnLoap5/EdfHzn8qfpEfKWeb+/dhWB74OEoMmSTIve8RYKP1Xi7b1Mr
pHClNZQZV5N+xqF6TXq0LP32L6inAPiPJXCuMA0FeRKcKU49rdkYTpVvtoS6gMl3
hPMgaSaiRn8slig2P3gB3J7fokAh/8xi9XQtTA3UhsOw1UYIQ+8QkSILe95/pk0C
FSc1Uzxcz+EiTgOGimigKhOqtDv4L3vYFJFQgRE+eQxi/C+3N/4G7wqfdCjT1Ygh
/efgvN5e10VXO2EotmHvb++59fGy4z4wj5ccxyRU35+K7Ut7S10P7VJloZzwwqqs
rOZEO+qzVg8Dry0kqZlU8K9c2XbOgAWpADaOngZ38ugovg+2tLPUtTx/hok6faXW
SWUr86u9KDWCO3GEIkcHcExYimO6okW/Q5tSXZJziOGxJdssy3zt7ufUKR8VUJk6
6CVniwAVtXiYk0fbFhZ6NHMHLj5RE/HQn2G3RWRMD+FIcDtj/EtwUZzR4LmGG23o
6XuSuMvccC9ycyeFiwoBWaIQnwYrJbKEyZluOLdUzuvqf6ZJUnMFUujHlEUSBZTj
pzxTCKA98CIZ3xHwU+COBVftJwK8vP/DdqcJegricLkjRhSFePtErpwr94FLg8no
z5QS/R6YtHNFR2FpSrz7mGEl9Npde99NtjYveSLamcEGlw3fUnzotM5mH3T4vbD+
h/ZSfwAzR1c8g8K3m1Vh62WaDmBZV5GaofvAfik0aSIuWZjQ2+KQWD7cJePqLS8e
B6olGRBjCIKxQMiyaTzyFF1tvv8dm0fd0gvaKhM2mztRAQq/eb+T7RlIDsTQfelB
as4wrs6+0+pPnOYZes4Ds+rgodj8aNjWQ/wGPLfjzUzaIoOhgCbQxR3ewVM9ylsz
e/ReOJJaGem5K+uXiis6iP11mQ5WSVJcvAGIPvVKymiygcGQDJiLG/2K3+YeHa9P
X2HFeEo/Rterd1NKUnET1J82vGqC09HUfO7HVmOuLxGsCERVNIeVZIuvmXoxVDdV
RSDLZtPCgGl/p/b7BOEgyQisTkptEhV2QC8zBDmY1gJzW7dhKvLzR3giVyq42BXo
/PFhkRvbOIsZTtk4l9VhU//bUOnWveo/0VZ/DUQJuCegM7Poe5AIyZHgVzNdBNUX
osd5Y5844AcGcTHh53/3DQdvFRn6hXY8uRD4nYPoUeUHcC+HdQi3/7NCdKGNXaKl
GLT/7V/Cwr36moXu4A2Hqjl5lFIFWR5T3p8v82lydO0maXK9jeTHgfAH7dmnhTnP
m8T7cVkPHzMOHHEQubmm/51XUJ7Q9Va2t/Md4l8ZTWV2XPfgfELyQyhzygcpg3Ex
qbj2dei/8TB5EENsGk5b/Xlj8oirzVLZN21e4Sk2Hjz2zMcFU/lcT7rrt6QFRUWI
NLtFpiUdzFXCOJ3nR4U4kbuECMHg/edNMu9r60xUwNWQacWj5d2r+2D4H2WMEg5P
mSKHoUoKfwn4OsN24BRV7jZ1KhQN0+6S7Lp1658DaHuoKK9odBoYmmu7acRuQs5g
+ISpF74+3jxfkarJ7o8GWyN3CQ8UZFRH13j1N1mRBl3ejWLXoBvV7BAhHbb3ufwA
ObIN3caRzTAOCawqAfbOL23jmVtjld4o2LXbc1AcWf3e7AsS/qanYgldM9P6Ew2Y
7gQ1SUZd56v7jtK9vF5/Ul27sUwlNhKAoTh3IolC4HzAJZY38gBFqAi9icoA8Yvf
y+IU/MwxIKmRUhyTkkniMMZ5kcB5ld4dAhwF8jFYZxj2vqm7Ftd/wHZkpyMOYQSM
jconw4jy+x4QjK2tsonNAoihzLYcpmT/qcrslSeEF+D5y5tAnx6jGJrOnZnOZ5B8
UDzC0+AGPpGCt0ZsBAsaIwi6nBMRF6wtrzauYVKiasDoMmvDMrfcUK2rwPLasbq1
f4tbxAYINVpjxIUM96lWzMPTZuabzZSYdnkuKju2sqZaSLsNTZD/5Czv8KHSEie9
nYJ+pdzQ9GSPDdtK/8k/3LI2ttPrbHu0CsWfOHkqPuEb/GMy/8ZBoGAfDn3AdUCU
xD4QZPIR5NPP6Q69IF0ol6nHbtP9ypGgZWg7hUpJE0iOrkh1ziMnfL9HaX+5PWZm
UMcwl8r1XbeXg/IoysLZaAG+1sXR+o/2EhveiBqtKy5bhAMgjEUfohEC/gdYYkmb
hbTlLccN7XZaKmQejFSbgDy5KIwrbTfFiHgl0pUHQdLhm/K28nujre5mfwCbgTXA
FSxA1F7A6y9jYSeyCj5D1VTkNQzAFTADqB8tZAg7qEG0nQr1T3r/xcvGvPmNEdqO
qtWNlN8SckI4rtKyblFxtZgWVD9jojwZGQ/zo5HzlqgFMYtazsNpRNePolf+e0xD
RDbjnSaf+HO5HnsBOzMtYNYh6WJ8m3VCEq1x7wRUqNkuQ7opIh3/7KyrpqUAoLE7
XBGJXGBVOjusfungxiJMO0hZyadZhsvMbRNZUDVFci8jREpOVC0qkTRa89SwFrHG
6eftzOP1Zrw0nNVipgmT3Zyprsg5Uxs7l9S3dU/0mm115L0Peaf9UsEaLJDfrXci
jZc9pl5PPLNO6kvKPAkUnDXZeGetIQxFw0MoWaSY9+K1sPkdxwvkyRAC1ZXNrYKS
ZdDcyxjajgMvcvx1RTIzol45UfrTD/ZzRAOiR1bUFiWEHiEOX+a4m/QActedVy3R
GGQuvIepvhSaRyulFszkOzy6Pt/8acSnQAE2PydIhZ6ZPgfi6pPMS8YKg4khrMj4
zWjAoCkZHL1mEAi3qIa5GAtrw8cQJU4O/IozdTxn+54FPJtYilAXWDuP+v8RJeQF
dQ1s6ZfSAazbHmeKN1pgm1b0wv6+H6syQncmayQ0WA7tDLN3pHtlqkEynCSscfQ6
IAnrUMciGw/WKSVETJMsCtFkh1qeGahhVFtR1bPGnv4hNpysd/B9FHeCydGhsPZF
fnN3anEkudtkZpit3/PlSP6hG+D+dVfCpINhNh6atY/3PY7wA2+EGgXogUYGSgVY
xxFEMSIyrc1woAAZu1Sz7RUsw9pMpdm1dcYJs0FDCNpQQXaCaxMxwqr+kMQOrCGM
61TmgOTzkkbzqfnyZwwf7PDkIrOM+JHP2FU3PM1eUoGDWuSe6+HhhLL6PK2gcRdr
9uCepYuz9ymNsoAivrsOi2yUF801CabM94zuuRvZi1LMq+xzDrSKcmhR29Ng7LhZ
KIhDGnD4N8+uSkin4RvP3h0hyqXBZ2CmgZQF/8ldtNKOOPQ4qxexla94VQhqs4xt
sDQziW9Ri50en3sJatI1fbK/8gfxTrYG8agXrrB3ZJhNwqQLTbam2Sbxlm9mdIrC
7DayJYvX+wB9+YDt6C//US4h7vTyBnPotiyKLb/QMbuIVaFYhLiQuKlGMhOJKDNG
/EmNGBbTgUw+iwb7gFgbCtSrnyTzv5tLtA11xWD8dBi6MjxyzSqtrWDXpKlOEatG
1MaC/f4mT/NycClzuaTWpnYSnyJggIQLSHibvcgwv4bmTUqPlPxoBKseSv8LNscN
BwStfXjSU55WHBzuk/MG+FlNrkRozG51LXXRhWmWSFfuZEqzVRRSaUMDn1R/vBE7
dBNWVBuGCTu7NUTOyzXCTN/4kcig8uyPw48NrqL2ITZvuw1MfVM2ga62zhdNB+nj
ZY/myE+W54HqxeV783eStCeFUv+jfnfhTX2IQrWKDyZMG5jEkHKBuwsW0jqAGUw5
d7fDJfx2kwq/W0vNp1LH7hgqZVralBzpbccks40OuZ4REXGbsqmjCCJyGHtFXO9a
x5xsFWvoIPmwmHL1C4gK82rGL8MxGx56rYkyMJC4Tsx4cfwjK/8S8qrgnNUzgd9A
4uzaqlQi4jkeysruMAFOALFlpf91Ah4VItU+1/ZjWBCM56YeJu1FNawt3wSkfu+K
zHWr5wRdeTnWzLQaWHocKy9BSO3JNS4GlJoE/zomFT7aCjzyhsmN6kP+BbHs4WPW
JzV6eeJBkhSRVJSnFJYdyHgudaFmJuWAzhydkTobssk10sZC1qKlyIADPpygSe7u
A/ziCe4AfRdtCAG9EBBrENfI/FhXG3SKvTDkZPfQAcroF9AVahY6fw+qypGRVBvX
sBxcb8/jrWMVKjeR792GP1aqrcg9eodIWfi8jkNyCQFJL5K9IiYX142A3fnYuKOY
LQwrTwa3kkPaI4k9joQ4ePh+tNalyJUTkz5Pu4zsDehwzGpW93U8Xhi9Q1phqdb/
coQXk+jCPRCfRge2RuFOarq48+pVYdtJijhebg8b/aWgHu2LX8Q6WzccYm1jcuYq
T7goR0KnQSTRoWbQVowk3rVAep8KCjFv4/pZiTRgeFBYp1a13THIKQPYlytDPB/F
H8K+S+z3vfMmpevxGGaPk96J5J/nJ6YJ/9GBbHDOvntylC2tof8FRqqElOpt3B8f
8TNMwhpCkQ5cUg6uQjaxdyTXcEfgPBh3w4NU9EAgZ/LBBW4+F9LF9jxhUY8JKyUF
zRv8QETtpNNOI5IsMGUe7FODgv+RV76rKlOrKdkRMvhCA1sMb1a+JE2Jo3kuhizq
uTzUttxwa5neADcUYxlkEMbiT5gKPuuXVBRxKaLyog7KNQ2ii1JSbWnhkuWhE2/W
d8lvjuBIvaLKKqOZ6Zl6eyAxv8oVU31A/M5DebsXlNkXVRj7ufojNWk4UelDApvn
iQeGm38cpHIwzkpEPu4uh2GfyBcIcEeI2ejrRm1LqdbI7LdKk75zqFKBONCMAnju
682usjE40/OFD1fmWxhaYUeSjwonZhk/4SHSEkup04pHVsRAcdj/L1AM77lEz7rf
pqIQgMNGFYM32Hs/eZclV4pkRh7q7Zz1hmA5K0YzHp0JaGCRpo4Zw4lzGntsS3At
3igCDjyFguqzY5Svtizv8HgbuELvyblrQtf4g7CMtqt6+whNsYVlFne6Q8g+Qbm4
gOMZS44RYiqwfQ6YOyaprRjUAJZRgoJa898gx4+xNjQmXadE8yUQNj2nRB1i6dKr
p9JHS9jKuOOjl5dmSJVXtxxAjomWLTRiA/it1zWu0KcVlGgVRaiwYr488C23/5t9
SiELv7lR86B27E4S205yK4ZQewjTx2TPm4BHU6AXdYpB7pCsc8P8KMn0JO7RSF4v
/HSHMGbDttrRJKoeuYvmoMI5nZCqfiYJ7hNdxszAgYrA/cfpe9ImvhMi4ov1hq4l
FcNGYTxPzu+v+h5FNiALU+JvSNDIRB9Us0d+yzjgqPQ7yDsZnxCGxLVCzf6cJCQS
VDM0CdqEUX7kM5ATE1jIBKugwR7klXJDGX+Mi6ZZS8v711FQM8b9ZCqX6VOHP/fG
5KDJnmqXmmwi1gGfvWdJpOkBR1sYcEOBa/tb17O1CPl9V8wZJib6TEzNIj4mJPpN
DIajt2DsjVu3mSaKsL5JfD8reYG5YU+bcgdHdswjT6BTs2v9hBqWWhHk9IuiV3GS
0BTQXzv1iCL6n3B/VbZ/CemHSN+JGmfOxt9LnhRDTETtnpCFXhnU/jeAuNnSmNEa
URuCzUuiiO7mXHfs02C9hAivpAoEuPd7Yj4XXzALK/hBpYW7dyHB3sQqc+nBYH06
tPqdotqGaLmzbswJ3RWWVXGoFyDcrsaPVHqY974VuJaCK9+0X3npg4CEwFXTrYgi
3oBLiu8+OENpqWdJqcSQhJ6Zi8sTKuZEjm3DVeU4ljzHr49fjGFJONBRUrXTmYS9
cvCvqq4vnlACrvMekNpNTxdcdcmP8xx8V2J797FzZUNkHICJIXRMM9t/l1GcwNd7
U9yztInPBqwrHMmS68d9qrEnOsQeCoBrlXZxw15FCw5MnrWPz6XFbgt9WCvAdyCK
l4Fk6DM3W0pA0Yoru5q8hRtl8kXNV8x7qiSFQ1CZm3fodx8fm9bnxz6OySYhzFou
M4Y97s7g848IhDjWLh9/re7FpN+8RTCsn1Q4+vacjd2wnMH4i/eBZfl5LSQz63qW
Ut1a/0Rm5//BYi+FRINxCYwva5dWvyfEsAQ5/5/AEZZ+jFZLW5Uzdahtxk96zWJQ
R9VImcl3b5xO/9DZHtSfv5ZA0EaALbO6Zk9EiGSZ8gsCIHKBtM5AWi+wNROfIOqq
9upfTmbEjFGfTgrXJdM4cI4eBwGwzNF2JrHmI0UBeRLClOwRa0Vgv258vUzPVtKf
PjtNiSSVdyAKh/8QXoyzzPo9ECIybdlo7KjYhUCCLddZWbJDk0JqgWpy2G+XEXFk
E8RdXsz77u4OBPr9w/amElvUFbkfYL7ZndakcX/RtyT1FJb36jo4ZsT9JfQKXe5g
xYor7G2a0WVmZUIJhFQ6z9pNxttX3j44yWWgHg8ol12YCMHI7qQf/QEu0i5/BBv1
rJsvGSGjLgtNkV8XKPJLDX3IbsfTz1E+LJaJyFjO5f6i0NCLnPmnm5VJ3sF6wb9p
z075Xn3oOzy5SfBN4J/u8iT3M5yap+eYP13RyPUhApUiyGBn8Wl9zFveHruCxk6w
HLbyRkC+4blLaWJCnh7ylqY9vKEGggSj65+nZm4sC++/w78xZ1SXs2wPsUjgm95M
QsBpNqCQot3uZDsw7O8zB/jSg0yy3nWE1aQK20jTJxpeStoPLJAXteKrTCdsFeHy
MHWWP5lIgI2yG4f/h+6MmZ+hOr5CHTN408xeae8edTOOjVQwCXzRy/K2nSznD+Fi
NddXlnbcNM4pHk/vBQLw4KFOF0bnA0oZSRYFKsRUYOoL3j4/JljNGNs08h/rs/sl
Y52pGdx+eO+0EUvg0AEoU4PpF47DTV77E9dl04hZeVqK9XaT+TSAvt4veJeGRwHW
YjXIFPbz9EAtZ9avViNEkoG+H68vD/CGwE5SprI5QJIYTIMLQTeiWlxsK7hY2XaE
x/PqwjA9jGQKqWY7QLYlG3fMSPmyRsd1wm8PR1tv9V1Nm3OYiV2c4EN7ptuwO1MY
msb1EXDWOjtPLWNIlt9C5XPcoo6j+HQ0EkVznKwc5ai0iUMYx6mK6tLuMW8qUFc/
E5oNNc2sWiZhAmToc+LdAom4NQXpl1cxBrO0x51ENqv5U94YzBNZuM1nH/dNpke4
Bl2pd1ES7e8OAHbsNVqhLI/nhArU5yGIUg2Xp15nMzv8dv+9dVdYVj2GB2Xmq/yz
WhEYJUEsoT0oqK8GIoHCZ/uj81idSHsjVCBclbzgEmQ5LrQgI8XYcqGlRf7OFG2w
+tlqvRahk4VZ1haXFdKpGelIfK2PDg+yxpmKRk7h6WHRCnXlOpB5/m49ytOqvwbt
eAEC0J6y0iRtmJATvqwUkRegZrYfw8wqtUbVJ1St7Grx2EwBkknahAlCvnkm2Tdz
yU6SEgasofw04DAS01h97Xvqm+w6dFKymlDjn3XRP5zHEABpHyhqVB+toCQ0nS/z
F9ZesoxgQqQ6slG04yOorY7GjUFzYPXMrnWdkUXaf2F4ypw3RNUuAsUna5ZJuEzp
wDubLdeoE8mN5gdHKn4v0kZfI79n2B2Sv2FPwxOc6peHR3uIbazlo4hrIhUvLzP8
NFamC+hfN/Xb84fh0lx2Po3jOqwfTR/kDaWsoU/QtGI5iPKLCVP7KSEgb/VLOaGk
oQ1Z/F43KSPG7LgD11sP9kVO0QEXwOqJJuXDCn3S+FCE5DX6xa9Lcf2pGMx4GaLY
ABxxiV+sMs7Qm5OeyRBzmJnVYSsMRcKaytMsKXWWlOyZ809cJdPHC8nqvcBlWwlf
d8rXSq/uBRQO9ZIsasHe9p7COC8fO20TjaONpPnaLRT7qMFZH1z3QhhALClCVPFY
HWwvcMLz7Lhp5+EZfw/IyLFIfP0n14yHpUPo4Hm2J8R/QiFoBzgWOn4HaPrJJbIa
JXfIwIA+FLzPDyNJElXRxf/b7VfwWvpTcggtjg5c/HMT1Z+tZNDZWoSq1hPE5EWU
l+KuyupLhCeNyp8LOAFIdtJrKcUUlrB4pbep0ZRTBM7KmRsx07PsggVzoVFI8LCP
w/HKJb5XpG+yODhpqapYzAhPMPHVsYGImlf8USQ8453AmGr5M2YTlNkY8xzoAn8Q
xVvTEakKrop5cKAgqXAtqKvynk2xcAoUfutFSEABMq7udEdV9/4yCOhKG0HBrdad
qtSv+nWBKbdR0mj0ha3hIWDqWIhSy/yH5DGCV5BzR9k/a3PBMjPnCIm62fjPPwmM
xEbDIfRaUqahN+34hqia46t//SRCfUFupWn4kMUuJ+Vv+PDM7BebCckT2FgQ7zUi
SP7H4z5cU2SrNHbjCLXIaSlGpjEkXAGmw3iV0bnAmsBan/cBfm4xJqhZ9Mj6XUaF
zEEIsb5u8y5hphCKJaOZ1xQyrCDMcxGPYTJJ7uyZ5sEoAQYcr5D6GyeX7kIhdyoz
Ctc2E5cTiPPsKUeAjIqpvagwb71/EglduiWPQOhFamJb5TfyHHroH3jxr90JppI3
fjm0iWmMhNF211qr+2WuBTDqyqP2QhgpcNmJ0V/4eS0FrFN5G1gplJEQzoiq74IE
cs4AcvK54UJkhW1x97IJTgvvMt/fo0S3k7kGHgJAvh4e8dt+66tzOKTs1DngSxIU
DSYZvxGP/uBHF0UhD3iytMg2oKe1nTb7+edbNalwSS0h3n4F+Zbl+9qjvHZXav+5
UX8LfLHnTA3GYe+h2wnlfePWIzMt4OPlcIlWiD2uJRDz8mrnhRZxXx7rtxBlLLvB
buZvXZlFrXDRmh8Ljx7mqwDW+AsxOAStg6ag5YkxJP3PTJsxedexeB9mrYlrA0Yy
6PwxP+nWO77AaspxtfrjwNWX6G+WjjcvkPy9wZCZTebLHtiNPzAkaYVUWAXvHwNG
Q2OrrTIurgyoZeKOBZpr8yhWpv9muypGb1mYAathWjfFUr+2fLRG+q2cqaWcOIxu
UeI6YmzT943VIJvjxh6PEAf/hcaeXU+wfLWcdxjhknRJRJITf5iv6eQOd7cx5ggC
1nwukdDQBoOY3wDw1PneGgUJB+U3DfAEloq4tvk2C4Cb0mCraNjVFiiPHJMkPTvL
OyxTDQrKEKD/aBWtSqVSQGV/Ii12sTdQ1bAZbo4fgqbaCBFngoSCuVlpzB3GBH9p
UAioDKAoykSY33bUa3bq9MsnWFE0higf/MsrGs1NeVA+M61PVTM05tDK5f6cGdh1
obfAqzT8rFXUtJ4Lqt7qaNDD+d2xF/+IK8CAtGV0kduf3O7IYHthPHCKFo0jy9km
Hr3h3DS5xVt+vicZtYM6Vqd1qyC0e0fx6iLQl6+9nqVk0Bb0d/cQQy/MzuXHBaJ5
z2g2mKIh/yJY+OqEsinQ0tzHv5Ly22vgym8GoKg3UQhuHZj3bp4iiuFAWA6E8wl/
0qfUD97QddeTI6OAv0m65xZ9LwZ3IAck9F0oEe8uBNfTwNCR63GE1AXf0jLMel5t
NSmRkGyRednaCfNgw7J4d+5ElwSibviTgO/2kMVgWWft/xNTX7268bAC2PTkYbGL
z5YAEdFrgH3+65c5qYbUHqJNk0kuhSRotSOufh1MTfxa62HLSRRhogJ5qmV+kPQf
fZ0F5pqGDGIKHMRZbJWMSE0P/c8AlnlJmgVTpl9XoTaeuxpDivxQisqbODvB72WA
WxIwNFsNShQ2mM4EVVE2yMNfqUFUlYbpNXMwlYlE4I+XGPEtn4UYPTKdMJsEy89T
aaZbC2gW/jYKPkBeMmMMd0dsqmq31RfN+jQgy3UaDSWTjfpbchodfgp0LizCGgfs
eQs8jIWgzzMd3af1INZvqIfqlv/gN3EcLLR1ZEYgAKUUvVtyXA5GUl3FfndYSJJV
ERGK/8cW9OAGfamiYjs4vLvVDzTMkt4QS52x75Wqsu/sinR+1CSP570kys+j415O
/+bGXkpSbuPkA3JomPLJuqviJoVosqdoACQtfrhYrTHYTgeURYkPNvV6fzACn5zw
QPBl8ApIHQWwZKph3cbJA0Z3zSnTSG3q8f3xDMzT/+HQoacfNUanjNCGDQ2WQSZQ
/U0AfginklwWUNoxXPvfLL5w1lMFuAw7DkaY4wzBQqFZHswkzbY/JrK6ktQMe9hO
cLmxbcMUq5/m1AcWpsCl+9gLkXtUV7xEXEu6mK0hOpyf+SynatVISPqJIWJMQIyV
sxGFqry8JoxN4odzkg3xOIZAiluNDR3lWGqxtewYJO8rWHhao4scoSqdG2oOVpDJ
XtuDm9EuEhUZNe4Bc8ghdJZ4OpbzAJxwK2MBVlQdVwyOdf4R7Qy0DZbUvnK5e5Fx
4GeEpJ1vwbBL3xF2ip6hwMj6LkXQM/YGvRTqRnls8aq6XaXt9OnsmV9W/IURjOE+
elXkrOR7rqEpCWzxugd0PdwcW7SXexZWYCljIXKvhyWPAj/WJdwXkKhn54IBdZh+
alA/rCQhbSVUA45+fs20VRzzHbGWBOkULgx4fveY14bnUiEmqaGg82ev09HEXcQP
5v8+mzZZXjGcnj6d0MqIJvgr/6aw8jsFlnzyopNzRfWx4kZDD6azYbtFIsPFvUoC
oFn/33JZ6sI7lgpWSgZgNwozTIK/I2AsU7Rn0ZM5HYIZDDYTcqZ8uaqCLgh3XCkJ
fcjIcIY5H8ENAT52OFr0TC3j7F6uBybcDddASdet90B2pejBJRs2ZBdkglFDrHhC
MvyWZJbogKBZodzSQshIffRbqXZXUlPGlVH0HF2xhAsSAHJNGUQPmjXeLj4yxEk1
oEoKty0txBHqaFgB0bZNWJ816104QQ3Cdu0kvf98qI1LoPeJaB0NAH5Z3Dl1A9dp
JV15N97M0HFjIaHMKeqP7NCPDmug6rIzNI+YH0xd2pH8gsHS3keKYSXVELsQCdgJ
4fE5+F6Cu3CUFlY0cI0DKF3Sh5Dv10a38vEQgpqj1wt2loOAgRaRoDsTxJMgcGsG
SlpuFcxadOUp0Ar6dHI7CwYnIrzb8Cq8SR/yPfoXEJxNBa4EWJQ+7SBysbRdvN8C
BtYUF82o9UOktyxEIUHxEjh0qHxXToOeZLxRFdIlT904akre6hDn13hP+9+3Lsp1
TuPYW8p9NNEDMzELtTYcQNi34LUe4cvcsXMh0tzHfRyQAVJc8OPiza+bsw+8SHi8
VUhLfa871/pIpu2GKIG/3C6gsiEop5x9tVhu7q+IptMtA9wuGy7ZKMopASnRO9iP
I/kxHfXJEdDClesQKmGlFdCwbqO6nbquSR5aEG/oGE/e+r4X/zorlR4D4aUQQXu6
ig7qIY+pKfaRe/g+5rQAniLhEod+Po2pHzL6LO2IXyoshI2x9puVdGzi/9KSeZsr
9WdMrxcEGYs0/8iNiriY1mnB7NN8P9HPAFzAlhchM3PH/fHpQjbfosZQ/2g41OMZ
LWnb3z5JATewdkX7NONvsw9cLvQ7ldzsTF52DedaXnWABO00HeOOPOBg59W8IBvZ
g+nBvkAlFLeFQ4CdpX7NZuTeA5Hml4+XQEA1InWD0RVb7pWU2oy1q+H5PkgkX6lZ
tBWP4YzamHARsDJrcEbjTXCbAKKs61pBqOTnmpMG3LR6HV/s6ZjEMbpTYm+Zjtz/
qqjvxphzD8GUPeFoV/k37KJa/WdR0MtSpTOoBvzMTnDDyHJ64PjyEwiwLuGs+3nc
sBHnm1ta443mqhdb0MlMZQ1NM+LosSB8xw5kixEH7nEal0jLbup/Hg0563UbW8mP
rZTNVPFcwiDchmzc6VKtRhqGDB4A0vu2hHeVHWwQ1/eARgUZO7Q/+jK9qjwe6rB7
mOTtMYNZ3SCZaGNUEuVuXM714wJt1AwzBhsEjauDb7MkGXx6kj5z3on5PhaARSTb
pX6YW0YLC34qPy49ArLkQfa7JNBuDp5vVroiL6mEdbD7cqbPWHwXmA9OdUG1bpHJ
wgObgdKDQqKziThkYl+XE3DhJUrHJ08Bv72Pv3Rdh4YY8u7UGy0pj5jRZfpvExEg
A98LhU65iDyoVykdCHzX1L+kKwj5QcOz3DK+atbXj5WpVz2zIu5/04ZJSUq0YcPi
dTN3r35Lt+cNV1X0TYt5IWMkgENexYSSDqs6GPUztza92xgx06BQ+kjR07tpronr
l5Yel0SqRJfUmtlhGzQNAWYSbxS38BD2XCPT0Tmsuzil1bjavDWd+QYkQivkBn4i
frhCEQdiRwUyRQEUaz2jkm8HMKie86++x4UW1a7vd5Ck+RQYuzlfxHuJ1aPIJirV
LIJd81k3niZcjj0Clrs9Hdvh9+thuuz2s/+hyFGlcCdB6QIFvPXardl9Maxfw2vS
2JwHgdZroTzJhPkQsdd8Rr+c9oOJ/7ovEp6BXJpOy0ZS1tkfrB2O3JYHwCkxt6FK
TY4/6c0fSNPYwAqj054nT4Xy94+QGSqcQ7pdvL6EgHZkvpDyLB2mH53rAFQhlJ8W
nKfX4l2VAvkX87ICF1VYzMOFZVOzVsdnKR/WAhzGrdEXtkYqqy2NGcEu/pJU5+7G
4oqCA4lEWq/EYVgtJk6p03N3r0YSB/w7G8Rx0hNXioMNS+HczVRRIQNrEPFwK0LY
bD0Le1DaG2VkXj68BcMUcZd0pWPO9LXhmZaH1Onmq3g6uSEN7j1N8QVbZRkDJ7LQ
wGYFw2gMPxdQdHp+hD+cHTpl8ce6IjzC9/cYDWLDr+SSle76luIbwYqF9l0CeJlt
OYCl4aermrBAMeYjw2OKN+K9WtUn871L3MVs+DhHp6C4TlvjHFcbsJN2GyjCRQ3I
ej7jLTLtiL2jTak+2KOhvMI0Dxmixnd9ZF5xBGkQpHxapv6NmnZsg0hrqnFh27ef
h+lkzNYAyAN9N9LH0bDBHBrwVeMPe/RqNBwuW3/KJ3+hyLikY9aHoarzjcHk0XAi
KyRcxJXQfUPCsKf54NtxnJEJo+wif9/GSe5DPdwpEvC0Au+V8POqFpb5iSV2rzw4
NgktooW+AOdJStxePFWWrYHV7WyUJ5x38brw0z/UKgsczFdrUFrxJTveA1WKtGHV
vDODyz6wzr2ibSOOCMk3ipWiTSbwUkvJZug4UG+3Cyl1Iqqc7TBiST2cgojm1nSw
0+GPE4otn8a6JXpOfAPgoS9WSPYVcPGGbmMF1IIaS8CidnFZbAxnGfGvr/iPtx9O
YxTa1QWBR0p6bHIMIQ3CpENduZYc8q8UIFkRv87pywfe4a46O4QU0cKR5NcA+pgj
/Ebt3RS7FjsCP01C83PZlSw/sR0eMjC4KQB8B9JwPywJVTdE+jJtV4ahdpPRv3bM
339Ijam9B/iuE4OTqL6CHCo5WbrXkCGBjCKZZdZPpw8WSMyyzVVmh05sgEORGh0j
S91nE209EnE3dT2K1ELk8z9CKjyGFCSSHVKDhVALGXG3+XTpwPhbVw3eJB+fdYVx
idOAbE6Pa3VR5+utxQ7gYwK74K475bQpk4kIr+NlYly2OXIDK8/Q4ENH/9gvlIpN
QWtvIQPWgsmxeOQMSWNJ0xfYrORzAIcz5D7NguOmBIPN3j8ae+vxaELCoqf3sqVE
w5ArJvPG4s0B4HDpC/SorPSgNEBs+pbix61IaFeEdzIUYqXCRYHl4pqa/WbSLgAX
5yQNkaPT3ALWPfDp4fxukVXG4Kgvo8H66GRRA0uOTrwbAktWQUwSkDY3FWl9YQ0j
suo+rEckE+K3++64OkTz3vItoKRWafa44IAzaBETdqTEqKnqDX8J0zP1VNqjPDm4
arEPsfHZMUmqHKswynIrdtaiHOmezKHiKVFotb4AH1QRq+G/DGMHnS/T4XyqE0tI
oaZY4KK26swhTsFyJcFtSD2J1lGQ0JPj7UwbWoS3BAoaVUW8wah1C1Ja9Ozj0tYT
Bs6ItktTPujzWD85Ktr5EF6NCIEEqM6i+kNY1GmSe+c70MW9ds8KB9bGPohxwge5
27MQ5InEdfqWTfU3mS0XJiNJZL93YoDN24edsCoAOdYyPl1VwHNul8dNkaBavciX
RshvtWvS3D7yFqlxqjeXoKFwJSzoL/XOujoZOoXBXfwuZLkWfifqPUUW/KTCLfj1
1vJ9rYlyaYMb2PonZK6KLODXmcSC70YZ7viXqw1uvt1M6RnDag5GtqHaVVsRz3dB
Fkp2XxH9sdKTDVarkTKaKnl/DJCEKV1jVeo5s3TQG/COfC+E60qozeZYVJ+yda2P
SUME6omaO+X+iwQu3R5TouRn38oH9hHgvABAD2WbiKj4/yjX9/NTULuSir2V30WP
/03AFPTNowOUoN+ioWUkZf0Q6s/4s/ECLwN7ziJp87d/N6AFTkjiDDIjofCLVmX0
1OlfMiaz33C5r0mS5DFZauclk7vtqXOjXrLuNZ1qTPkbFcaxf33hUMOJQWPArSYk
hHmV0YzW3s74OpyK3ZPVpNL4M+tB49aoujrfNBiz9EJLBZcYw5DiMeGRt6sNwdbW
2trgNlbcpH/L43bSFpjr9dfp5xyHV33JSbgKq+6hvlPbTY2oejIrjsV/eP0X00+Z
nOkhFQUVsILWUlvNyfNozu4u4AtgxdckzUBdAIhDFxhW/aMF1e0lPg5X5j8PUee4
yJp86qxknoen23xgMBON5iyfUj1CyGcllDrJQGn/n5ABpuZvf6KtoDXxp9pemabP
PuLK/h5J3zwBwZ8Q1PwhuK6Af9mmeJq+XXu5bAEKXXJsgUKN7mU4eQINiOE+3k6z
jZiyjvZyPGGu0B/g2xsDTdEPzzsM0SPOXtFjzSWEtV5YAaTnzprHLoUBc1UzkbCy
3TO84BjarKx3qUULcLviHgUYyJ4KV91Oo2jRU6lg2aOpPclQNW6FItqIoXD9WTWl
KfBeuRhmFMG7LPh9VWeEqGvR/A9/KEpF8sotEaGakxJ3d6DwJOjeFra5949xTG0U
7nkUCkeZYWk6Mcpu/p8Y1Aa3BZSAYZL0FMkPN7sShW4aCWeLKwSy3dz4JmuCZYX1
VTt7qm86Cvng0s2A7o7GKfb05NutB8woPL5k/dLFUsveSa5hICrBiiLYMiYB5zmD
ZmjUIgf1Zg/QxC1aZLkuIE6Qbl2VC/Ly6D48JPfPwe5ZiccG4jY8/OOvnxw7G2BB
BJ8WpjeqVCXeMtc192vOfj5Rjbf3HHbfIZez/B/2Pp377eCFRM/Q4AaywkyzMzLT
k3EZV7dik7JuWr+SvtMibOHo5GzS9/Q4VkBI7Ox/8Hbv8gdrgLnONimeSgcJdhw/
tcmG4Klz8iVccYhZnfUgbVVD0UyKI50oXxake5+bpSEHC1nl+6AvUkG5M3JQEHpO
F2Cp2FEx1jS2Ka9t3bh3fRGq7b7g092/XBvG/thJADmKFSxXqEgWgdRN82pBxyLx
CKSTZ6SGalsuzS3ZbIC0ane6aMcx5KH+lxXNWlP3RUOLFzyqFS0DXH/4qslXBhW/
xVwdtRzbU316IqvaC8DZJ6tTIHa4uVUe78x/TkrfCMOMXuoMTit7UOWEzsme2Q1W
pHMZobJFB6VFkcnf8gqWiEoWjYUWHESiSkOiFMkOfPsytSHniEtpd3LaQlWdvs4G
+3OeYG+fM87UvHMGWxSFt/B9QpZ2MnTEY3zTfD13uBbecJ+XHQEMQuknim1PJoOs
PzpWVBmVqQJY772v+Pp1l+dtwRNYmiLDeWxfVNyIrlHXpqeByXUX1WZ8qTL6Dl9k
cT5XZ2C2xhGcdg53m9JgvL6zNlbh+VVNpTW5ZcTiXc9EtxKlCRwrGQa+zmYffTP0
Tqp8Zoimlv18htKa5cfllKUU4OX3X5Mf/WwhfsJMH+noQMEJtQEQ5TxT5/6EhkW+
082POPDqmaOwIVsWEhHKghf/kimjFCbamJVQjOehjxGtct8Hy/t8PY5mmN/o3JTl
WXRDNABcJqsKnsFn453ZLoH7PvWcfqwbl17k8ZIC0HnR7A+Sljh/omvl2XYD8dYV
McR+HtEC7XlO07mcYGr3N2m3rPO8yul0c95Z211MB0iF/9sYunnQhBQ8+8Z4GZ1B
KEeGiyQa2uMJGHJzFbOrI0ohjJHqwrdmJ8UVt50iS2YdY8REWkzwP3cg1F7PobQk
HT3zeWcgKBh9IV8K+XydCpxs7UtTVdcR7uManpqUcLJUjTS/DRVwEw1z3uV5ntrY
XQywgoxW8GTfbXglZlSArc+bAPfvtuy5t5O/+xL/SYktLxNFOnHhKn5VapoI02tJ
rh0n+TgcdCXX3b6gmFUAod9qQ5R/0HQSDasQn2UjcwSZktjJUsW5yZx25/Idaoie
XP0aRUX45BnT8K5C2yT5zHRGat/IuY8Rgz+4fA3iSg84m+yDDoYa/LBeBM8eGNAe
Cd7+gmcaxV9bcjdpzyslmwuhhIuRwk4ZUFJY0wdBCdX7K0I9ssVjeijlRZPq0/RY
3uP4IlP+klhCC/JwiPYfY3ncZabwPSYb6MvJr8BkKbvTlaYReN+ycWoibE5PPys7
SkGSzbGn9LnxxoqgzLp8XJwLbxC1fhEDcN4MIO4t1gsel+eeyTfm91xd306rwyKM
8UU5WMogP2AXHITTyRJRuV2mHSMDxf/gR1Pw6E5FNnDyufdbh4Sf5hOimQ0Tp/Fj
ITU/SqAbOncx8rlbk4VeXOO1mknUuxJWumu9Xjd3KIPDAXs8TznM1nGAW0ndDVDu
tG/x09WuKSkmZNXEp8j1b7sRdYDkjZRd0330cOMuNjTcBoUyl5yk0LUvMyz7Cn/e
VhYwDj0LhWA7qFK8QIQlfPckbORpQvpiaCpXSGXAuEtyvB0w3rzUhnEmT9J3C6AL
EIGwgRrXBcICZmasYWZvUYUSmr/W07ERfhp388faUMZovpKFqzKWrp+hrILONfON
YyYUj4Q5JVC4Io8w2NlZ9Rc/EljyA7tFY5qV0xJxnpAJvqgC0ZXFwAfSL4li1qp7
4U7pKI3ywdttoXnw6ym7fsOeqVUAjurruCH0Txop+kTFSLLjGT//rETTfW6G/3RT
CxTZb8XJn18ghR8uTaZ5PJRh44luQ2VTn/6cgRcs3U6lh3T+uw8UTTWlDXN10wmY
TgIPM4zXwaOVfttpE3/EzlvmpfYrnOFG7YXBNhzeflG57ZfUAAjkDDS0CeaTU4OA
krXTqj4Bqn5qAXFC271BQ9rX5hIvFQMFYi5cQ7ag6UHSSHIe71BJRE3tXfkQEYkx
T9EHTvpAKODBnma/NcZChzhWkPSt9BFkZQw2QAWnQp0vW/WzvJMYvXS2m4UvoMYs
4vek97Q1lpUdGcQsWflv0k/GCifhlOJjTlz4sHudbHHjQFES0B9Oc6hbT66ig1vN
cT2/VSwwtYwZ1C4Pnvsd0GZ5/5UoAsNXTkRwlSPF++pelF900FXxtynn1TXG/WgD
uLQSCltT6pC3++HT5k73kLgvUWqD2sNVoWZ7IbabNkpAzcN6vTjaevt2466cwx6v
UQ1BZYCrlDvDYqZ77hSxRizgCFhjoM/k5IsiLMzzT8gN4QEFJogxHuI/KzC9UXzV
S//9KRn9261VmBUxrk+pk3iWUf9I1AflgyX6MF3x998vvIGyclZ+jFcN89tg6AY6
BQr52y59MAzf6TDVTgrDeB7DndL2Rrxol4RIQ8CgPnQ9biHupcayXyGOdVuqBqzj
Xp4MZQ/183XZk71OlEQBnR1MrawQoi6G+KrxYxBTvSuIypVLEWaL0NQUsMdtL2bU
NzQBmcGS6osRZ5DDdpvjynIrSnfSLcR6IxPF7luB3yZsiGvNAAEQQaCtRQrogIm4
W1niH1hxQ/55iA1q4MmAv9qvBkSj97Dz1uJtaD4dhu32IAg9ecVHFMAEpdkM7Yoh
eFVB7bXsC/yWLoXLT/HDV4LLOmJCweE6+OAC2upKH3TUKGqLHpOU3FCV3ghNsOMs
sYEUTqUKQohxVP1qebGLnevFE1S/fn64V/gmQGRf3W0Iu7OjFafyfxmXML6VFpId
qXG1qRWQoGWMWiigr+bHCcgmF7//z5WGRV4Du8FeWTdOR5kJMem8iOlj5g5jh8Im
Hq/peLaP0/jgHu/zqc3Od75tFuDHzSLeSWE+gfAPc8PN+2g0qjpywhfh5eX3tBFD
C9YujNXbWCQV6U4kYRu7MwxeqWmPZIk2KIyLcfCDbtoocS0U12/xlMh8OLefZUR/
31Ekqvw5H/oV+b1QSBrYM01Nbx9cpR0h0v4r20fV7ZnInV/WK20ldoT03fPA1iOl
bu5OOyj0ABimvQ85fox8gnLhqM7C2aIGTxBOS5z9nIoFxt8sjxR7s9KASrpw+xB7
7z2BLvgsCuWITTYTJ4+PwBOv0sZxwbKuwkEGIZxn/WRHIxZMx6zpizUF0g+K+0Ht
0Wq/Ej6VjonYrhXmTH8j4YZGZvg4Pc+tpP6IuKwUMH3plLElQ/gCBgmH66h/KGRI
S69ecEuBXVLXxmw9hWMZq1qJOQc4Q3m7rQEFVmT/5pgcGt0d190cuM0Sh9KIFM0d
JR/kCALyc9dotPoqsbpjtiQb+bCmyprd8a8oKdiTtpCWiXVggQTgUZDLhLnlg2zN
OrCQJSUbsgNRCZFrhQ0wnib6ZJAWOBfEMcfdlWf2iTFIvQkUTonPoNvOm8+BOJuQ
qV7/15/3zXbvXlvtFoRy2YRDgV0kOFHYONxXHv4oMGlAlnM6NvFj5xLadITY2pMc
Fm+6L3KWgDQo6Trly6YrFYeDbCxH82oL12Cn99qGOQ6JklPuMnMfbxByrGU9kAPC
8kQb5uVxHQ6jGo6p5eF+orihaoic/TDWNnsTh0ZBH473OAkIKexJXFdQzuDXq2RS
04iL+n/bBWEZLNj+MXyd9g==

`pragma protect end_protected
