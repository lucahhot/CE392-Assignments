// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qKilkVq3wqd5KcOo00WutOQzwvsg/p511krv3mOe4JUt5sHTGaHVDhXsLm20tjrXPpAQbwyhWX/i
Aim2xFA5ol6tm4bvD8NnUsFgLkpt+bCDa2blWEg8AmS0Ld0e7yilKWqmD4nszc3dlS3yhYXgDq6H
duVskA1raFT3CCseVv2N68EPwHwihgWdnBy5CFqLdhmc9jd+DmcInooc6qc4rWZj6FK5OnAyvOPk
V79nKeAfS/f0QOmOE7rvxGfPfqz/HB5NScvWGuVPosJvqsEvbfFZxJL5Lz+mOzbcljrcLXdr04a+
WrkbsrLKSu0pveJVjFyJfup970TgiPo3VvbUzw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 121504)
1Fjaq+npQAMBpGof2QURazkdkxJcn3YSF0jDbYj48nPCZmkAijej5HWchxGv/wdJuPA2y1T6aGif
gyneuo6HbqTCbe97/j2OQgi+ZkvYvDqvnEwzHpp2yHWZypqW1s9+I23wyp2Txt7cfa1NOMGCSlRv
szB901ocXS3Mg3kwwQrkDVlyF/xwX4FMWEK8YaJk6SnzaPRL7JqbHAkpC4s/wT4FoerPi2rQuWEj
1eDBgePj/p52qaNLburnDQqhUv4kf/DON/mrnC5ji/qDpPRVeAYbRJy4JAiRCA8mJjGiHfQhw1Mv
XGjJwATnGq2LgHBJlKqZTj3rSDWeWJMbUoJjVQVK3F7zvoT/dsDrW6a9BdX8NgILCEy6/vifKteR
/mEdxKXFgLtKIzG8KHgBa38JIa61ucfGfeFX77vDgeGxj7ffqrQzk/9Tcv9cB73Z00yWXqWJ0Zy9
mD524UrndZjef/RYSmRKbFms8w7RWVelOvp+fUuHyp+XaNd/wqKrcySJEcqcvfi2KbJUIHuIA4t6
yEpNZw7+AtL7n98wuyv184TeOX/bzeAEuQfC4zB4hQcdNxPvK2ilL8A9iUf8tqYTocvHZqvoRLIu
oQnWHkXgCE2uHNBVdJayRG8+fnlx1dSwfUvpn6FOpYo92m/51ChaA68h5pvhi/SC4qaHzHwmzcLd
iBy8TXmktmmGYCqIT84FsabV4lhMKXwJrcy2AbnvVTzdMuOuyo17D2WuNZOFtqGhp+BKfrGdlIXy
ooPJ4fHYZchkH3XGWFx8I7l3+PqSz12PZC88m/7dw3SfAgUu42H4paZ7gelp9kl9aDEanTOI6v7F
Az282inw77Pd9BbMXlFX/Ej95hcGzt1G/c1Xizr+htqWuVjmhjCj79JzePZ1K9j4ZqHOtdeQ2+fc
OyuYVS9mk+IOLOk1hDL/yP/IkuHCtIX7FlWJguPHNOXiOrUTXL0zIFKa1j3EOLiH+v3pSM0tvh/q
OxCo1maix9I5DRm5QfujwN1oO95nTkaICPwCyie158RkVI3BZ8O6w+cZbEbHnC3zGNwx6rzMhj92
8hyn+SsXitkVlFeKQtH7IIFw32pfE5cxnFDZW7kiIgGwj9oJ7oUcqvZ+68ZXJZofjXqDB4JH5Phx
SFy7ys14mxQupGex0ui2oN7oHHU2pEKoP9qoYDp8MAWRNllTw53O65pbWBqRMjr3CYBqlKktMMVr
hp9y/1HxGN0N4ZZ7RTOUYJDovl4NtIyjvc7uqp0QYPustr3QaOF/NpXkBscfy2hBAOD8fkWHuE5G
uHZUQX8WLPe07sjk1nb3eZYUnvnfmobHnY0YSdPl71zBhSB8f5YUT/QniP2Ws/b8JjUv4crgTHLU
6xMGeZTHMECZcru+9mBvWeTQFedJ1pRMVS+wJf554TK6d0C8zSWaSEy2UtSJjx/YFw43iO73DMgy
bw2tXOu4KolPQ8+4LuounhNcLhxT33CEKMfxIcOiFVv0gRgzVCdB5O1YC/meIykRxt4CzGuC5W2i
20tGhc8hEvkbta+AnnbBzElWHAgB3LtU3q4OpS9RQ5IKZv88Tc/7Ai9fGycbqAhrPIUneBNx9PB1
R8DIhheCc0uKWxM52KlVkIvy4jUjlzmrROhT8wx4CTZasnaTREOylyS0f+EzWBiMfNafnOJO2yLJ
AdMSnJ3QFKvBplh9l6Rv7mimsM24ahLLAwGWWISbR3/cK8+6Tdf4y+IqrqHTE8ptOP4jM8pznoUS
T/ep7gnv6Q1jUuwLhVUktZMuPgqhttgoxK+3wbJbUIyuZVAoTlJwV7aIvbR1vRHAaaW9BGOn70ub
5RMVE/FXszBhWMJoSHvbQtwf/tTppV20hGwGaFhPecUoaLP8pixE121rar+wwlDUukrDn7sLSN/y
U0OFxJghiOnRAKS0zl363qDW1lf7ZXCB+tH7RXRXphzZaDJNvq2OWHbXfLzH68BZz+EXGVrJA1yF
rDajnK33pGhUuY9Y7uH9EfU85S9YyObMVBZJlVGA0SJd6LvlSDQdFMsJ6yhMPImge/+oTG91tXHb
C1DsGa4AoAdInswGh20ncvCUqAvNRqFBrRvj3RM8jVeAizXvdv05PHR7qO5ti3dhq5GpDWccwUsu
aGiOKgxoc5cMXIvqPK7OISK3jBkJPRteHdArvJxOkbPO7UpzVDEAjFJHrwhBYLTgMfKNqUtRLc/J
mQ1PEy6SwsW3v18jUin8AShLXOxGVePsjbQuSIQZmRJmcTujQQpgYl4zYN09IM+rgfrScq2i4Ukb
Cce3lxQ53dZ9MJ7z2tkYLBJNGPo3IpALPrt34FLss5h6mmG+TUkYFvc0xyzLwzlc4JFde5tuFIdM
HubYVouz5hHnKoE/PLS87YuS6delbwK5RfpkTZcsNTWWHFhWFUfQ3dEM+vqNQC/RI03pJHMUYQvN
47YaPodAIA/wbKRMvRglWUdsebiw3Skij39t4gScHwYoBKZ03LhUBaaGdO8XPbej4El8OGBVy5gX
Stra6IKfiMBBF7fM/VWa7wCdH94+SNqvgyKAcuqcqbPu7tAXNiQdCykbZ6TKaw8a8l72vXCbUIl5
nsEgOHIdPTdm9ZcWrYnmCC63q3PEGncCkmHRf5Jyq5YrpZ8JshL9wIKNe510DSPtGAtdQkUfBl4f
n/BtdWpIs5oHKF8YzERljl58aa2U0h1raFTy/g5a0fLln71ksKpxDVPQoRxhxD7mBxLCWRPeK0Qa
TMzInvDcuB8JzxzDwxFIDdY94PrcF17+ymLSAuKN7kOP/R38rQX6uGsQadUNIZUpPOpxvreApAVb
wLuYRcIPa/k4C5mOO+VONEh/xS7HUouqA/uGoBT6UiUKXm5RPMDKwbgUHpactYzespHhwiHwpv3w
PiIqhuWJeXbSQR5IgxSBH1ALUPjFDPWN2KHaDlXTMj9TC3bIUp0WWMZWdseJWfAz3O14IDMRrrbD
0oB+950iz1k4IhdkBIWqjAikxHQbh8m289Ldh8OmcIQMtT15x95MorjlnWZ+qhCYWEHnvQd6aHlo
bS92a1F61l9gL/lM11PSB2T5zKsz9z1F5LxQbayfJX+I2uL6+BhSgOakuU3jBVd5AcSttEHuPiGt
Xie8A7wEOwSzLVqV5JlykBT4r0ceie3JkHQg+/T2zijpONxc8PXatfb2vdjBwq1ZEa3ue5OQEsc6
F1k8KNccGrkYNs3oHl+NuUlLKjZPuCci7ki8voMZ0DgvHwoijW+bD/WtBrkjOlP0cE4kwRGuuwav
8I7pQ1PYlnwx7l3RfTvgEilyIsiM7xRGyr4+SkL9e1neCCsPKB6hfgQBM2HPcVe+0ZYxML6Ils1b
JgD0paOj5uaOD3ZsbMgsJW0X28Yhf7zdb38ZTzfMzKR+zWPC+Ci4FM5mwZSdye2G1smKHcruQWVb
BwodRxmvzSNrIOtkEvZZde/ppLk5tC7pJycZ2vNxhZWSEqa/IhKonh4Ksr9UwTuufayqNuhoQA7G
u6f7iwokglQqzQ0Pze/r8v3281d0Xo0KFIzGMuERALPes9ffkFWrNpauM9IDBrQLf4ZRqWu9jEkV
9kT83zpdB14FSwTfKbi3XsVB2+9w92PCztnKUCelQgLSQL6DRPPDqbolOnY1/rzMz/lada6pgH17
E9GChgG53Q0J6fGttUBIfp8wAZLDTk0WNemiSOVDhkVN4qqD+crHiitPC00KcJuzIS8Cr98zcIXt
CIX3uR7HiIoNub80rFOsPr31V2Lu6KWGEgiMm1ewwE58mI81yS5c9ynGyMtSZJol2suA6bDdajYZ
+8ilutG2gfUd75xeHoIvSnwUGz2e74STNUEV2pJSH5hSgvRiXED7v9egC/1bSTE6Prey0obUB1tW
fnsvXUeGG2BNbqHxunDPsr0plBD+UAlg7caoyXTFcv43jTS5meN7kij2+3rbaTDS6jNapeHbiWq7
xAtZv/dzSnriIqMhMqvGPqBWb14NEz3wAed+in1a3jaNHbsCHO0ybqYcSutK3+bRZOozKGACDID6
mzXP5pObcyFnCE1uWMW175Z/Uv0HpAhY6mw7xS/iFK8hlKOstAC8eekITxZuDOSeTjQZolFh2j2z
1XvAUxfuirIZl3BjU2Tp3T0gnSL3+RYf6cj8XuxggWxHNXz3glSCGejKsHLeG8nWxhq1GRrLb0rF
8iRdO/GH3knfJhc76QtJQCKnsS4LYxny0dOemrHF2rLs/jlBlhlrpIuXQ1OR1bKFASgjzX2MPA7J
YZ9Sq2v9cufmRMF/bYOQ/ZPunjFyPHcz4d6HcoXh2ESveWqNwmdw2uyghefDbHtDGhQ8meL6+JrC
fCohTVIwboyVJPI/RdV5k37RSYmqICphvaNkGBdAaKDB16EXLcSmjR85d9Cx1FLv3oCS/mGCquPH
XmlD1Rnq8qUYsnHyoyuPHvkg34y5K1WwaSnRCWL2K0ZGbxlGhcRLqX8x2LSrNkcHt/vlsHXbOMw7
zwfG2DRxgHGD8A1z92vyU1ZoJF6JUVKt6FDqL5coczCQzu8CAmujlPiGdcihr8DYdZVCjshd01R/
IWI+4i1nR0c3jKf1Yo4f03HhbjidVAJQeN7JuqjHSRJt+iBZ64/wNpK52d6BR7+kFOCJhwB2zh1d
dgP9gx3dVj4w42zwfr6mnUJla5hujdc+bf8EJV5canP0Z4PVeW1+74RB9HmOe0MLEcw/4gQAwWjN
mv1FmDGFwIOecpSoq0W4dvB8B+pUI2rw/NYdRkqCT28qrLeQdp4fWOvqcYOdPL6k175Q2xyjEpW9
d5SkYFSrQv5/Pw9Da3PITY4m2WMnP95cwEjpbOPaywu0VaDN56DDjZ4J9kbp8D/Wb+tj0ZKi0G0F
2VP9LM+RUHasDpplouEgsKwTeEgpC1v5H40gRxPSqtHH0HpFvdQmB5ZY0GSN+bSozr0Uo01q5UF9
fEYC8tmsuuPLb+Zn8LpzJqbVg24vZdQDf7AMVnyNfq0427F0YRxixyySKHSaGGewxgbPkLNkVMns
vZt9HFELglwr/WXCiIrts+FgjfhEM30+70c4eaV3V7gUKG98O0vYFO8W3bZ0boOnpisVIr+s6Zkb
z8qIDD8ztZJOVxDmRMok6XmNI2SsE8wYktNjQpU534GC7Z2NhMNutzDWn6AT9tIsNzy+edw+A3Ku
6E+HobWu5jxE7hwYQSpU4RdpbzX6tGqJ3hETrbnHCzjtAUgkw9igeB8qx8rVb1qcSt4NxK3JSmz1
H+2Kt29xg+6D86gd2LhjXDdOvRKQwQ5sGKNZj6CMZlnY17Kfr0/X3547qtynJiwV5r199BGo6K2V
7F594Hg8OCSZHicNYrHr9VSHH5Wf4WtgI7RUGko1Yh2unTGEBDC9tl4lHr2RjwrmgVe0BXMZJTTj
1Ut8NgJu79FlfIcuuryyl3OmGFesA3kiiH1KkRzSK+oN3XIEIMSA5aXnz3tUeBJPaim/4a6+7RyS
/+wxNc6yynvDkekntIQysLw+d6Z9lHSEQbUrrwFrVkOzXrDN1h5DUOrNJVgRsHSDLSlyVuNqrOc5
FAkzeglBzR2y52G/XdFp0g1KHP07cbHYZxX/x0+TVMPO5jH5Sn2j5gY6kXXAmHQZmtmHmKNrJtGy
VJNxHDC/hnVPVNIYNkW0fBoQLLoM98cNSyDbDQ/9/YC2p61rLYb0ERylasFT2RjTgm8XEbo38avy
lwnOLFqJy1Nd2bk/jXOZTV8QOFmiNq5NB0xWBchrbd0UWzsaU4UqDaS95BMIkPZKUtUrJ0p+1GUx
6HeS+0vCbSTitwNn5D98yRUxCpZK2tAVBDS6CzdYB2u+UjubenSLv7piHTsc13ZJEdRWPmrWN7li
qf9u+1pG6BQ+89VAM79d/45UnWZZqh7+4KLRz65JVKmsbnOqoREBrT7o9U5Sr7zcaWzUjcT/4CUu
CitTBcji05lu7ScXqr+XaiMmNg5/iDxeP+eFHRfjeHSVklGq6hOLgQdC+4Y2AMecCj1CLHOCZB/0
JQ0nufG/gDWyJYUavEXeJWvlk1wBpzHKfKi2S+CAFpwcC883Xx3MYK/MzbomP001mJZ9g8bXs8aE
q8NW/3A0Jz1HpEheTVCtDkJmA6l8FnLq/Ix+4OauYl/SGZmsPMQlNl7moD9cqZ1o7k8bVbZPBCeO
VpoSXjUiFWz2clLDKSmc0LimcJ23ias6cDE4RkzVCbqpH6PX75ahRPxy9arHhbgeDTIYx0ilXxnv
4YxZMafSnmpwWUCABFkkQB6j9nJw/z/LbUxNfQH5Z94Xx8apPgq4jV2zrPEx07UlZvJXbMjHE2eY
uFIdiBSxl+lCbdiA0vQKpHqWf/kmT/mshWA7FqWxYBKW2KWmabmJ/hv0UpxB+6BLGb7JR8pIwbyH
l6FOhxtC1pZ99eo4wycTU/6XWesfXWkvHVW4oksSTT7Z+82peoDUBGwsteGXeOuUnkPtEm+dwyyS
YEa5BP5nK3SzQcuVTS5y3oZPDShufhl6DlkKB7g5EVSq/Fe+OfO+a4v4PgL8jeOIiVELbPcWc1am
1SIEDhLIBZmlXZW6c7epsYlNEdTddgYsRInviaTPJe3+gLQjN+JTcVyw+Vf3EJAM82+I1eSVdCH0
gu2by6ZpGZ5MRRs/DwSEXuCeF0AC58FniXBcZ9UeY6SHWPOGNaYEDGKfxSPhxaQjN8NsCGcWTXGt
DwOLY8+bZas3eCaORyDXrvUSuP6FtI+zk5YB4O7d1qEOQ5jyeIxuv0m9NpBc2aWH5D7f7gRV6/4w
A6UE7009xv+O8w+iPd5iiBsmgoJSCB4gEhNN790SYV2xwK7G/Pq2wEzm+OBT98ONcjLRbHdvzTd3
G0RL2dhrVM7yAfkHNqXqZWRx6k6CaSY5HGsqaz0if6m+YTwkaCAmnZmeGsNmYUBwycItRXOiQA+M
BSR6b8x61Ov3dibliuZKahrI438ETt02eUpJ+B79IRkEeVhp33GAqYs1P0HgbX9WZOhf/h1zLWYC
KGe/Z7Hnr2GeIol0Nlf/3bwaU8Z/zAipm1+mpB2wix6y+59rtVKSihxgT9DJNxuifNzRdOMxIy7X
xXP4zL129u81QyoYldU1cQna83JioqRCndfg/GT7xSEIKK23tW8Zcfh5opoUlVe7L6XfKwxh7uPR
ZyWMUgW+DJ/uwfq2bklMYZT+MtvU3qPtEnfS5ff9o+v2QFjYRZqNzWzdFya/ugdd9QdKlIBRPLTm
nX6Fh4v2DSS5K2FCdIKty4GuevmT84ugQ7llRSLgyQl3QZDMTPnjAjHe1eYq0Hq8bbZWIUIGh5Es
hziWaihDuu+2YrwFf6hWHoDzmAQ/tN01D2cOrqqxYri+7x7RAsqfJKHCu9xz07QE5RJ2yaFNz/12
JbLm8zxeDIM6ocIDRiVRS7BD6yd4iUfFTdHUASB9Sf03IqDzrttJNvysQzr2Ts+RdLdOc0zjCnw2
jmwA/suZAFSnPqbUoNIWFmIUMe1qBfIZlTixpYysS/hCGd8vdlTqKTVcNbp3yx2iR4NSQnEYw69t
fL21RCiV+9dfGc1n+abp8Wgf6M2L7EXUsWYnOZoWSYbeAKC4FZNIlIoECw5eAOprfAZXba7n0LGE
6P6FOsrDqPO0IwidxezvmyF+SSpn3lbzDIGZFFAuydTgM8nrYGYhIyzhuRC4B+ZTRDUc6CA7QkZG
iJljaJyugOYKSBpSOdvTXGqAWtBLU3SSkLqp/FJco1pcnjH1uE8SbYRfLGcRTvVLu7uwEda/XyEn
0aU8MYKR+MjDJ67P+PcuMoz8oXN1xdNmQ1xfDOq0VGsDL/wawTgt7790AiNsslbKu09FOz501+gP
MuW5SqGWyT+orlK1RAr06ZrFyUFn0sn6ZmhkSL0WrsM+gk/ZelkOBuiIJt4bxII/zWH2FF9p0dGo
GQ1j4Qb/xRkYhaGXrKQ8IYxwQCcl+FPpmhm36LD4xfPS0DW9WourCDUo5eswRSO73b0nanmrmqJa
ZJ90RbhrIbEnMWLyZ1vS06baiPQi6SdrZeB9wwwd2Sg2nD8ItL5AvgKBDb9zmnreJUvliAd8cVJX
rR4PCl50J0y32hwm5+ULgaNQQGhGVfKPfY2OVwXkITqpQRdkmm/nz1WBJOt9cA6z69LD95Uxzt7S
SxGQI7rqr6X2rQSnXRNKquPyEXLjVKzmRsRnFe33X3Ag9rcPWKvQ90HvYnCTuy7DM3CWZL89SBdL
XgyAp2aJTFyKDon0NzeO4ACMGa5NDYerHE9wkaTz543Qa3istYIsmbbs3eiATFGixTP2oDZL60WF
589F4LoXHzMlrTulxPlESZDjSG8+1liquSm7cFWa4LFEAOMvFvMDC6KZ7hx5j1emtMcyOmyyVTAe
56zkYkRO9e7wCjLiFDbTimkcJnexhZJi5TIV0HTiR850k8sIaZ/MJPrzHH2R06PpxCbEPs4Pxy01
uiSKF4W/xlIbFWCNX+hEHmHF+scvyXQRJ1mvmS2OnRnha01Z3APRQzSXl5JPBRcMtPfxIVaEXqaK
D8u9hAhO8wwdEythgjT43pK++q7EKpDU6WDyGyUki2VR+jBfIYhg7m6nGZ/DwlpO9OnRRVMNWeZE
8ModNXV77G6+aXq2BJPQxe2PDB9NucBhLKR2mLqiHxYAFteVORHLmgY0v2YwuMHzN09dSJhcv6A8
Y4LToyvGv8m4QRlRwY52BmYV2vKdbwGQta0beFr7q0g7Yg15R5qrFnCWeSYHx8a+1LaAp3bs6Pvo
Gh7OPDHWANzt0xW2vZcfHgb5oEJqjartPTOHcn9khHLpFTuiOAbujWc/5PLR/g8aJJBm938oe5NH
XF0lYyWC3V6SF8qqoJyozEiocu7/cwfw9FWzFrAfhjc9N4xsh6u58Xhe5iTGGexXVp7Uvpo4MrOp
rMIjIAhOCQo6vVbVqfFn/5dewWoLzigY1j2kXNUVISEgcu9D/Q/ccSDByghpWa1eSIfJ3ChEN2lp
/mORx+U7LU7vMmFm18Xg1gv97qRih063ZWzE0+vaS0eEZq7bvnH6Md8WmilmITBrKtfbPzjC6Rf0
06AhLFZ64Ie+grSgWP/6B4Wpvsv6/ilETpN/W6muzjmJcgWwdDDnFGSX4Equd3TiFY8K8IZu3rXi
b1u5/jQzLd0yY0hrP7jQgClR55WUhnQgAw14smAaX2H9Z552wcshlqA21QkFDe6Y0gffNgOIKJqO
1TnjcbkWIF8jx6wyLUgvKH+dgP6AmTxE0LCu9W1f8jEeY4f281Y0tYT9f9egVRKDk3S+Y2A42mIj
jLUG+IMHS0f8QtdOhdEcvkyycOh3aUumdepBDlMKrBfU3HKzmzz7NiVK1UbVWosydN3/mRfV12aL
JaMqxsqEhG0A0Drl0JYoHyUmSnYiouDsJlQvIjBFgL9OK+cXlqAL/kTLMrlR4Zt9JWZmj02vfQCb
0lZm536FCPgCL7X1A3R9TUckLRRcI+JKZ0jnzvDpPS0llhd+SclCCNxQXG8QmwviiTK+mSatLu0B
csvlLBj0u5dt50EnoVgKzNVQWzzcYWxsFF+DXrSd/3ISQ7M0z7+2MwuOuG1EN0Em9SPU6GucmaOL
gQSm6EpCZzIMOSxT1hvsOJdoesg9Abx+Bhq/Y6SYrUqhYiF/9Lkf1WZHp1I+uOG/+FazmFGOHmSz
d7t1UejC46zz9/CKXBqZOGj27hVTb/MuVt1Y7sdvEdAew0Aoy87Z+goPcUD3QV+CeBGwhK/2i6Nh
LzvQxqKMjRIfzmhyHbIH1hvkeFEjVN2cCcrAiKOiWIbiJn1g5XVQZgtzkYFME/JrVVdGShj2Lqmj
L/XpWD/nK7zhZTfarm3f98GMKKG90WysGwUyKSBOqCcsqzJT5vCumuznXq7iwnbFYw6nQZAPOn91
PNr6taNwaOZMoAbui3OhDaiRs7opX0YZFylvfUIlBwIwXSHrm5jBcFTUYSBnrJTIEOa3cBXpv56P
RhcCV9veRE0k/iCVaItQN/vaDflfRCKPv5bfhPF2JoJhMlQtrNGRxA7W3BnhrnipRnGqw+14vdeL
HCdoLlcsmXD60NnB/ocZ/tHAb+XPHfVcXotMg3n8P0NN0Xi1TZkex/kCpbL/7nONkSMRHD5xJbJ4
E73n61bB8LL/0PGN1vcp98SEkefrOmf849wQVxhCf4w2pn3UTiIrZ+W9aOERF0znx6Sr24jFawDw
m/0hkECVDDNoPzJpG+7pc1ifpVf+bc/jYsUKfvaHikSYi2y6KIaTHQiQ8EKidPr/UtTquSwPJsms
xgRm82/CO8o4kEXP9XeB8sQSgkRRrPdi0a8WFumS6D3uDpTj0sO/3mHlfwkQzloka7/QYyoNFpaa
Rm6rzCR7+qORrP5iu6YDUvi0TYLlqKiT5WB5ieZ0e22pgMF7ZpXKu5K0G5tRjUCW9TadMr6dHVwW
KnG3JF0Jpg/fwzN8nHsP3JMpL2snoRgeH6frBc7iYG2gSmcZ8K+NYsO6RxCO/mCiUz89XAxy4/2q
knBGwWrDOXG3EXV2Zx9ouKnAODW4aXJBZv/1V2MN+3l35DWpJ0TQO32C0Uvs+xWmMmCyXFQi6WVz
eOc6UkOJ+j3sM1RepMRquBmodtuaUMOa+8lQLEeMLm+XWOlPYI4qmgbcPBdFJMc1YVFrQ+Ydv7eW
OHy0yOrkvaeG2EjbOTDwoKdTrAtRMwqpq7iZq7rtNfrrsPTi18ZM1/gz7o24Jo/61Of3as+Zzjy0
jWmaM1VytKgFL8d60ITOrpbD0gzi14EsSLpd2jMmfPkrN8be4WG2NTX36hJfY1kfNED5Dzr7Qzuy
qV3klSyvDHrdARp1XkdfjMs9rebXNwiN1qjlLXliFmC962ESKauRJZtq9f1OG4Haa2dELlCHzicA
NUiytz/U2U9gOtaDBznf7KBfmyVjukAD/u7a61y8O0P6eKmbQtW9Y35v+0gPyO45Q++6dFOMxyW6
kpZNMIJqpypmQfX7hYgOlMlos5mMrgkGCpY+xd9J19b7PWqsGyxsG4MO1bNHydkQKc0ep9jFobZz
OJE8XxM1vN+wDVB7FeR2UOv8+T2H6AbgbTb/362G9RHqGawkjrrUdCIPvAN48Iou8yHET82Pls8Z
0gZUtGQthqPHkWRF1Ssc3+C2xS+U48QSyHJsK+8Ovrh+CFcmY++7qnVjchHo4SnSCSmnXU/ihDzA
WolSsnOiEt6U3XV3wCZXocWyMiEK1kDVRif5TglWTgPetPYSgQfPwPtxsvq5XvnP41g4Nky4nFMf
Dy5/NIvDN+jo+F/uDFh67cRNrix71Tp2+wOjLKlFFhN5d+2NktLvr5gdpdTv12nHggEFOcnvB2so
nmExK5rQvkfm09rj6weOfG8R2k0SxG5WlKpMK8yOQ80DneW9bQmtKAOEXwv+M1hGwHnxSQIlNdAX
b6/jD3UD3u816+oN2ZS2gM0rcT0X52qP46SK+z2jpIp6zuRYPA1sTyWP/pFVfLy6bnxTHG7KgrF1
tGqC8GmS/yyxOUWl4gl5B/ah5sLUHsvKQbNasSm6PyVXxF05oTkvBcAluuNUySYyOteLUn2yEX6W
rNUzWkYtU/XajXXzg1cBO3n8EnTaY8HWwNOOhcAsVst5H1t5MzQbDqPuEMrDTvKEyFXX6wpdNeUe
slQZ58ak6VGpJn4l6eVW3qyDaZX0QUGKk2uaoLmobupwFTEnCkiCRi0xgDuP5GZX3+e2r0YFFzI2
kDmu8rPsZ5cOivJM/MN9WWpASDynp1fQ4R5nD/VJRRrIcTjSxeHJTLjaSE3OfwxD40J6ZnCxDOIn
4yw1nwZ/d1c75qb6P6Mv9kMEjEo54LL0FxOMrDaml4a4FuG4zyGkWxnxRXr0HHFV300gEOMaZ4qx
444qvLHfn75VeJeNq7kgP0W6JGuwfAFwPs7IQfSISy9wqPjC5vQHnOuLWSk3ilPt86vW61gDqCm4
W4e8e0WYhhA8bBFfQGQ2TK7aop0AMI+wqQGRLRAYTR3ub8Fa1h4GqlDmpGaAMo35wselGrKwaglA
4O+J1JClvc6w1Bj+/CMobSbDaHF8JeWWglIkFdf6AsN83Xv6QKKGudoQLb9lkxPz3AxmTRnXBYhm
DDBxqFbOvx7NscBMKsZ9clhGVHrmss+7UJVGIP0dSSPBL6kTQcg7ROu6B9SJXqBNHph9yfBX9E9A
EIyRzIUFJsfi5G0Kin1lXKDFSkjx5glbuct90gwfePXxactnMEv+2sesXGrJUdAhOWTupukwCtpm
CGn30a7yebPO2CHy6zqQIULxrSJzuLiWeFmmLy2Bq8l9Ai0NC6FzSUvQZFTIBj6uPuy0cLvskPok
6+606gPrGT9PFs75Hx84NVvGe9B4TGfYPzaKoO+ADgpGMTIFMKn+GXjeAgfGsox/ubnjqf1HxiFs
NZK50scqjFFck/M/SLBQFhYCpRCPtVdjGw/0mQ4bGpzNWTRdB8kPl/aKcAt/mp6G3+tSC1I+KYU6
YBPNc6IQvkb/T6aZjJGsON8Or3HuAz5wi8usE65bXgTKMv1WBC47zkVTdqRnKKjN7jukjgs0SyDD
MVZ3fIwjpeJcb5cvcvO03nkT5G8uu9dDbQ8P8TyK7tnaJzf3mJMK4CvPyRYrE8Y1dfMEv/EXTG2X
ZIsOi9IVmXRKoSXlcRp/ldzWCh+dx9ktg0sG0U5XBUdm5lRoEp/cAqqi5peGf0AOxbA3b40JTqLI
UcOaHYxMS1ohTN/jgm18sP9ygtR78Fm4lKZuSWSCPN4U0TVXso+3JyRidR5HB/6i8McLx5O+thwL
CHF0ExwC30m+bYb8Z5ERcmNOfbbOCZmPLmkIGJJTUtrE3Nu0ZztZ1BqFUJU1qb5rP31Xl+vf2Ck+
jGxbNo3FxH4ffaZlV0q1FZzF+gE78WFrWwVGaOwrsbUt/D4H47Q2Ps/59z4QQ5p9cLHh95fe8B9W
12z8rKqXK4WHrefSU4xHnH84SUbR1xJS8YHPHIgpVpAjjglnNE9usIAZ6A5N7RKS/Zjy7YTkNSPk
g0NW9cDV9M1sJK4WgDsxBlgVVt0LqGcF05iRS+W1dlqry3xut1qw/KQkDLQJDv+QvNNPtUPD8T4/
vXj27wTilwhDYrbl4iinSX1O10899k7b0ggZi1BcTqM+FKjAYVZRiiwFOeX9a1CWLVmRL1Q5cabf
XSIxdqtvpaTARPXZYHgwSzMpDqXGz7Iv+kjGON+z/eG0j5A+B1c7jAvPIDs1gIkBXrbeAzzAehYv
xJ7pzVyimlB6NFVI8/u5aBsg2q2LE1hlq5bCMzo+i0k0+G6a9l/Rrp8/YXU/LDdATuZ2KXtawLBZ
0HIMo0LVida7efFbSXCireNjYfcSOMDg+JRESbYcGWBP9SwLe3Qb0M2ObX9lNUcOkYQz5k7VQwoT
YH/wsjDXLoAbq3SubSlUcGCp4ELgUmdHZpr7YjCDQbShrA09XgspAG+/r/FbB3shcGIvl/46jiKQ
ZPN4vQkHKMU+uvCWgxCzcoXKKmBaOT0wdM5SWsYkuKCzTa99APpgkXGPmHANoRX2W3Sp7GH2Twi2
y8xj3OuZujDYBtZ7KIxujqWJYkjUttSWi4q/IaKt6uSh60ArFsvZ68B5URloQSnX2pQXVNrwyYGT
tBTYy6KItctcGYr09l8IvdJwBJvIdAf2sYgWtHZCSQSZ+VYEaRCmFKlXKQgEjAIbVLSDwBF/I3le
FDIAGb6/YHrNDxI72CEmXPwXbwVDjqa/YWf3qqgB7d5pplGJUqbUdwDux6chqhjUHKyqzwJ01sW7
cwPzDYrjAnWt8LWyQP5k26J9XawXDFL2lGwy/BAtqzFJO7/qN3khCxrtdNEjoiBDbKS6J49lUa/h
FoG8dZPcZE9FHkBC0niAiPam8zuivvGyCJjNFhumFTYn2NeQP0YUUiTq9Q/55dmHSBBZDnMPrHfi
J6EM857tMUtV04B2izFCS/aGA5Kn6cIzqNtu1UWw3A6Lq68BzgxYLsPOzluOAlTTwD+cyrJoY2ze
P4qBMVQAWLtoaX0jRWKdo8Q9LIbO/Wy88MqfGk4auftOzyfNjJGrzYHxV6BrIuVdhRwDvEX8eeEV
9Q0HRGx+WdbTgDqFC1Q60aob4UWgxP1AoczLslcrvSpGChU2tivoKjZ0Bjh7v14Qm+9wzKVI+Ffy
zS3xBGyVbXToAWRXPHufNQHbKNmkdY9Uax8WEj3umO92t5cYUTZxOjaGDSbN01q5F2qHK+/rezb3
uHIe3VDoaL8ZyVfKVEIYgZar5AeY9k6avOMJA33jVz7K9jYMVRR12yfqlfXXjmEKGdAN+xR6JQJe
K4xTk/ISSwAo2eJEvy+XQ88ULey+UVRoEkVk8RA/MgzQ6gRG5HlgTM5lmF8LTUBMcklVBQHF3lZz
jJ3QEhtsk8CjIoI76/kFsDPu3EtojrGD2q7siQG6XBoP7hX22CHWb3yFGWY66epWvkRUoWT3D+Re
T+hXJb4bs2MMyFOEGvFlj0W4Li6dRNcRdqzlI4GrLReIW+X3PsM48cT6uGz10x3OwlYUGN8yb47B
01Q7TLSysaMNkQ2f/HIg7QEJbej+WUWQBkTRnSDVg8GGCm2trIwoqAM2hP+54aweGdsGeAp6rVp+
YdDtJIkes0AZMVGmvIngFrlLpn1NNqFczAqg11KVTImp6E9G7RqhrZwJjMwGDYMVyCbNZCjG+eg+
9YXGcxI3+WECjPCvSSBUdepZumN72bOi+nhxu5wN3X4FakFpD0Rll/Cg8hQZsUBNw1a4ASIJW7JX
nbX8Skf+1VyCweNPj2XONafi1GDtTjt7P3H89EycURo4PY/ASm6mUrjAqFQeHiPS9aa133k7CGiz
z4HkJMdPqYxSCcezr4LKD9ZWz3rA+as4fTLkgLWmI/2dT0Db/3ofMvBP6ZCfr2ggzuo6lbmkzXfv
IyTTex7W8iUc23BN7+o3Um4lQsEyMo9C3hpMqu5NevKFnOqmSRN23pdCFa5pSpWTJTXT9hJ5Zkkr
K1GaVk4a/UGn5emCrBQqQrq4NiOxhtF9fPcxYDOM6LjppG4BKcrkhsDuOQtiMKWw/KVN97qWeram
nwzfG8FivA37lFRUEZnx/RmbsChgZNKUH2o3KxNfidMA7d1es/rVuj9r/bB1TW5qpYtb3VIVsKc0
eRPu6AePAewHm2gBu9OJsA0tw8j9Zkges5vs33D9tdimHiCEXAW9Y/ER2f6BdPmR/6KycyTG2ZOC
YXWLVIHJagOBwo6IiT2u6AjwT2nhp8u8gTHzbCm8iTC64QnaotKAc3D42+UsRX5lHuqXTbKnFvOP
dV4FBQBnUFZowKSaOcBIa5zTgIai3qUB2GTpPQJocOm0GhM51w5ZO2/I5AIDS3hqip7muxozA5mk
ph273e/oiKibkAswp+oDCGCufT7gH9mo2rtZNZAd7OK5zV542u5QA/4ceQmAYL5jJPgyKraNnHS/
wl1UlssMu0OOFFuOjfpYF0X4dG44K+jKnQubsdTA7Vaua5+HMFgIwBTEeReSxQmWsXxfquJIvLDr
FlxmkFqcGTulWYOiPKe2rSpBxB0aTKpvKSkPx8ScqNiBx67smzmtbFQNRLEMCnHW+CRrTNkGi2fD
TgaLwYGMH4groN8s7kkN7do/XE8aSbCZfB8pWYNuQPolhJdCp3izWmYiO74id16AHuiKT0AeH2tH
iCZeWntvcMiFSj1CT5j7M20QiKDW3HrwAXXhJATjmhye+kHQESczXWxn6mLHYUsNetNtBxSUh4XP
XeHZJewjtR53CCU7kHKoUpUQdwClDLRf2mLUpA0i1wpYeX4oTmA/cICCoYzhtCjZjPNN7odJzEOx
NWINnAOA7T1AjlnVd5R/8ptUCngLo08fMqsJtm/phgiTtoQTwALkAC34Bl2Fok16e+igB+ZmprF2
pnBoUixH3r6X0S5Sh9on/r1aGGCbemKHxmKqZM9Ftq1SY9BuyMHB+iraTTGQ7RwDRe1xtvKN68Y7
M/+z6iKeDmGeSWTeMEi2HvePlcJO0ntyvpIUyLz6mo/Mi+fE/gwo77zij7EmZhyU0WzCEL+8TTkF
191LWSA7JCvslM8Wx57GHn4/CaNFoqpSdkRxEOgeqDhTthrrB6QnePSbwW020PZ+zHM5NxRSE3/x
UD9iNn6MUvnGmPcFTvWQF0JPdH0yTpyTf5orx1Ck5RnPHzgZEaEWvtIrmUhaj2RTtztOjDBLuHWF
cXInuWaIddyVpv7eMsri2NB8N5H1t4i8CQyUI4M2ccNvbeoxCJ8w3E5QDMUB+6ObZlj2M42Iw+8C
BX0ZPSGH2CI6mSbiW6h4b/80ikHJNmvZqKCYzXbIgbttc1F7APmCLdx1aH40XLacHDVBwCYYaaJN
tgQoH3CvIYYHfe0pEesdDocRCAWhqT8Us9hkPYRD+pKf4vax9CftqGlb7RiSNznOUt/QyM1THNON
Mw3ajeu2UsNG8gUAIDFZLJXxaeNhJlivaOpka2fcO3QNecYkUP4Deyoxd1JOuwmyGhIpa7KyE2GY
QJ5JLYpz5neBzNZh6MdriqJK+jtH25DrM7vViB3GdKPRXyWgWO0Dtkv5jQIrzxn4rlqNaPuyYovM
ir+hZqov/VS1xI7rs5Dg5otHziUCN8gnXxdW1XRO/zQ3R/Pb3pdyjfTjViDGCL0bpxM/LEReLH0Y
3uFEaHYJ1EtKTBkYs2pga7XLnH1RlAR6tvQG5Zw2Qq0/4kjL5LVV+rWwePq7tLuG747X2f1m5/fN
UOtHfdYDKQDYkUaKzHlLk7DCRf3Q7P1iiVbEfckJLAwinqJBY3MxKQnrBAuDpsfB51M4gKV+xQP9
GYrJfOcC0FcilCiIIiB2U2JgErT7zOOojsufx28ESD+22xDVA5i7wTfpp4wsNx1AURftlpqTqIb0
8yJQbEtN43uQLcxPmo2Crk5CNzK0rOjJF9U27xqlSxBUSPykjGDcZX7LFaMu61dYFI8WgbN7tPeW
oy/xmnqCHDx5q+FMQn852aJC2lWX58HNXNsdDp0Ph+Ej3Zw1zN/xylQBT+ANX2kGjgTg/QduJeIL
fJes2k6Yx8fBS7ssMtMHGiYi8RunFnerzqtuhqC9+SYd9fw+VUbXw+N7PNCly35dacngpT8+fCPf
9G5nIw4Lut81UtEXah7W08uQxY8v7s56dfndut6ilqAdibvr17hPByuQa6S2phn4WQt4n/lLBOwo
Iu9X1IaY2H7DS0P6fwY4dpmSedgmf0dS9izK2hweqSdPKXJ1ZolR5CmEK+LqEGRFcblfbNn0xAjf
XpLsU1HgPGQcb8YMY65CYTlRifEzsi835XmgqOyYvYhOQtWP44SQWjfIRRnX62votK9u/G60kyaM
JZ/SyxYLczuTltv3gATgNSg1hR9Kx/fn9SaotHQb9uGPdpFGOMlJieDFjeVgaXLHHKJAhkGKeiDg
7c595MBZ2h8P9UsQayHKO5z1FFJz6kMEdwEUeGEFghHHU7Kf7F3dDZ4Wi8pg31trUQrNhU8Hm8uG
MAna04V96/4gX6q6TU/ualiIJBOeS+Rf2LqDScmLznAokpv8YtIE+4eSHXm0idoLqpcQOnOBustD
o9y1PD82QiWqoWpymBuBZoDNFQrettHKQpf44ygRTNhU1kh4SPOezENaq7M3JcqtIOfQwOdfFVKc
vdGRCL9YYre9d7MbWWxwKE/g06paPunWzqgGEcxtadLLx0hNM3+S+jBPqwo0Y37DNWYIgg4VX5PF
nfD/mvFoSs9PHGm0iHtHXK2fw7KV7m0mEhX87Obb79rnvy9o9Jh1N8jsPpekul/zyREYBqqCxwTd
Rx5tsNN4b/XRzmenKSiOV+H48F6Qxigh+TpsLKTRjmz9lZ2DUW3YKjY0ARKeVgK1wRHDzly4SLqW
8hdgUsrAZC3j4mJFK0FLUVm7zDzM0tsctW9Fff0RGL8JAXl1Lc26wzE9AzRr+x1VhyoEdXrRn+tX
Nf13uqtF+dQtHvXgJQ24auacasN4DawcQSejmM7Qbs/UMNDQ0d9w5Z9xMP6W97+sjUM6vs+0PHUO
ZZHCRb6vShQK6TxlxG64ti/5PKrppfQXV26t595pIWS9Id3WgCuPmOD6x84cLX8DJz9t0WFPUARg
b5BSMt32iYDQlPo0U04mWTlWW1lfDt5c1sm9FVT4A2Jhc2+8+O/pZzYBB2VHQbfXdQDv5fek7AR5
KSjfVatxdZyAwT6ylGItbElHCvtdtHWLtDzg1iEvBOPf08ztCfUP5XXGq4KOmRafLABOZefyLoAu
rmoYkvkRdtn9Dx9jZOGuvF3pRKV3Fidg0xLlyvCaM9olNULAHfmFHe96YSNZTmvcmZIKPJtB/DlQ
vywofNijTXuHDYB2k0ieWIc3WJ9ngssfPTrk2x1h50xtU3Y8E6FmL0a1ixhSIGvffPsrTokVmJmF
Irpkgpwfag0/PgYOBwNrxRpiCykLvf2UTyyQNgw7kW96n8ROAbB0bi7KbqzIDGhcxqodly+pXe4m
OBR5xHKYwnPWh/TGO7BfieV6Ht61CoLIAz+hwKHknjBEplvMXxlNj+KdtAxLgjUcOb3SYAd9R767
sj5YM46XsBIsJBETk4E0WDgraZNQsU13Fz13ZU4a0kBr21tOROoA23PBmzqyP+TdArmBKDCqrPkl
ewEsPuF4k84FnwvTe7HpSjU6amrudvlbsapnzLiCXiC9M+zLKiYy5EPXubHS4PAT4MO+U3fQdOhd
Un8L6ZtxbvZTnSHhjnr05A/dOMKJ4S+/IFS9LuC0QbN/Wf8NBjSa4bxdztTfDK8VHw/zasrX+eBa
2nfW4LfZRFXBsADG4iyaERVQyy4w7S58YFR6u2nU7uwpwoVg3A3PKfBSZqe+wv7M1jGbPPLPgDMM
dGVrXdJF9AT2tb2dJ9uaE+3rMc4nAyreijRiD08P/LKe35CJnJYgJaRxXh4LiDInu+GLIxgafzBn
4UJhMFkexDnpnQ2liQag+YbfyUFJAnpso9+CmlqC1Tx8g8P/7PeyqQVQdY9aanGz2jSO/zj28Mce
9GlrKKCNtHVCl1MdWk2w4UzW7Spma2us/e2B5Y88BqvTJ+czTFqNpHnPhVbHneaOQZuDA79SW4Ty
CcCH9qJkKqJmxbZBY2bvQAD7vzN0gAb7bImBI7kEiq5b5bf29qndd1m9yXqa2fw9vgMvqo27tX4S
lw82OUzQwsM6SAPRVJ9gliUAY6klb4nhCaPcUTe1pNAp2CgML42Hwgn/H1jqCkMX6RMGchG5YCKz
c1n66qcZA+If+xQZJGM5Kg2kn3BLsAahBS01oTVAPo48aibtVZVGOq4Wjj/iR6uN6mitkaxkfsjN
x5vtcQDYCFJ+BJeCiJf7f479UNAbrxlJiYOQZ0/8I0nS50axXzgmjCBScV1stPj4DShaxBeU1Wzx
0KxTLhyEQMT9bRV4CkBjfocf4UZTeJln6WRuv1lBQDJkWi4VqxEDidD8NIgSvXSKGr2HdBlaX6Ny
0n2fe4PiGW7GmsoSb9jFfeXNY000WnHjR8VaWr9FuZV8lo3Nl6AtMz9o+dVvDtNJC/8ZUDBpVdh+
EFR+qAmtRQmOChy10ob6D1YdOAc9h2NluPNhyLgI/rFzuOfBKUfw/HuB44ZMlPPMY5MHjSssXSPZ
lbCQC07DaG6ybAnI6nXwV6xQe5aAO7WgBpBSR8FZGhcq46sqMfuYpCSsL/H96KGJhEVAZbjhJqtT
Ge8P3hLhuJcvGH7w+ua/aCLpOAzwkbfnKOr/6FstcvAwomxt/6dGrNA0xw0c81/d+iprqXWZxO0O
OFtbf3JhjkTBJTMJnoLRhGYI9Y+rtlU9RClh/w3qIQaOC7kB4Vc6ZmK2ckyB7q+aD7vvMsI7FWvD
rIondqVkpdtZJAx5x9G6y94XUp6ZNnU1pzUp2b5FRm+Ve537x3bIcXi1Qmh5vszSwvejz9nsrW7B
1N+IIGwM77kcpLdXVLfWEYS1EADAU+qK3e2myVD//DgyxlhWnHrLQfe6N6wOg7EoQ/DMGSUrSejo
M2Vhtx2tkenE5Y+Yl3p//Q++JqvEOnfDLJW0o6jjfO8RQO2tpm/CKx1nDPIOF7bKPuv27FtfbtBY
NBDYCbS4JI0lacOeJ8TkztN/JQzKXJK+I957vVsNG9C95wbSeqvVE4rFzuJfSgcIMkZeLz66k1pX
8ci6UJLE0LiZZQF4IECoCyFFgf9D6R3ECs7NINpKtniOweWupH9fsLdh4jGld0KQmwN18LYnXQmU
2MUL3SHjVV5f91ppLX+1JMRHrmEyhwXXB7Ps5DucARMs6XntExtZWVCjHdMZDES0KwWzXxEvy3d5
VL4b7ymiPTidmJ2JF6sD4LWpUtI1dLnvFbb3qKRxDysA6OPTtloOxaWcIrjo9bKXCkZu5qtOP6J6
t39LJVDGp/fok8IFFK4vNJl9DXBGyjWxVq1d6VKT8sM78Le+8DyV8G5Fib3i2oawMUp20NzIMp+E
Xy/483/IbfZc/vIiOxwNUvGhR/Wqm9bI73xnwuo/cAGXOXS6voPCHcOU9Nnp2Lv2rBh+LQHtorcj
AkP9sS5XR6/mSlEkJyRWchWH8V0eZEgH7S2FxtA/mM8ztAwtFcoSNZFWp+poZZkdWXUeE+BhqqSh
bFaEYURVNVmfGQHlJXxsYJjdabKHRZQrdKAxo73GrgIwGVVkm0Om/WUkvgmgWdQV44cP/p9BgCyt
CH0MI4tlLDizgCXWP3edQHAA28pe6MEJ5KeyaWfldtm+RSksMHHdUVe52cs1d5dUa59NZpJFXWqD
zUiJpZ/BlkldmBV/TW8gkEbQ6+fO7HRJYrttaCux4NDJ1ukpelewadYy+GOHMH7gOCDik1mrA4uo
u2TGWIGg+p51dY2X3MJnezcPMkfntNAkZ0YQOYHhGBH0EYCFDoJJKs6KhJ8Tib3viY4rgDiSMD3t
rGqeyZ0TXsITU34Tw72AUKUpmhwyTywd4oiMtTpcnMVaiZoIJAvDcuUxP+7cyuY0JXuNGMmDODUg
s4wRdIRdp9CN7rqchfVcC35gttt4UJju72UFVUM/ntwtTBp5FUYtAwgcfpaDkuiwvmJcwHp32MYu
fNjr8fvUgTVMmGaTq/uK/Er/mN4Z1ufPtZOYIpYbwPLSjV8zg48YmOqgP9KOO1pvHid2OeQSs22K
fOoyY/dnhcBt2Qn4GBImcnscVIUZxS10D7/ccTr28Aki+UqxuuLoWMoXEtFDk4JSYDaRyN+f41hh
MjCIZ96VWogXPtrCr+b0aPu8aBhI665V4usqFkr5pc7PbWkkNO4u1mcOvVjgcIUr6xpbt73kyQFh
25WU6OPT632GLFZL6f9MYs6zy1TKDyKa3MnodF/iNjCHJUGFm2yPid2LEPa+ek5K0SqWq+Tk9qJ/
WsPxgN0YbWeL8kl/FSWGAP2KfSkYegNxdUrY7X+YNUfFONqKyOenPsODvZBD762RnudaeJB9BgBx
tm7PecchZ7+GVNUxYwp7CDi1/7mGmNKyMr477boBe9XWaj3GK4lIFMqn9M6KKeSr83LajnKVzH7n
iaN+3O1qqfWTDRVgRU4qTpziS1RZ1V3pdS/Y6Bi/CalcLEakiL+KMXx+6qIZaxWam0aEAwVoQHhi
JE5pzN9OQdTimx7H0ks7zh1pKiqW47CgT4EF6lb8++TOmY+rxkQUCJjCDv2Xog2WoijccF3qVups
6Jwwq8bn/AkA4GhNwHv8JDcsPuztu9DRDQnns+CEKjIsddFOh7r52la+9ASdPHt70sJuZnk1d+Tb
vyvJEgQyNg1NcdG83G3PpLpUVejdlHtmQxoAestV7K9PG7hsdue+1JwbzCz4vWhs2BJ1In5emoGF
GuaHKuilfeuIOy5nkqadkzTCWED2IyAFxFBKgWYYrSVoJr3uTGyXhPNW0Z6SObxxqU7QQloMdt12
b2XLkscMr5bj+h1JRoBIggkQZR/VJeaAP4wUdMT0ARI0jRgHpdON931es93/KOJHaU7GKBy6fRx9
7S+XoBkssHj4K7kPunuAhbzXO+3wVqL+u+XDU1vqHUvELlJeb0Uv8S+cwWd96WyOYDWGS/TLeayD
d9Ju4cxqz4KyWHoW0I/pMiDY7b475trGL+c/5WF5hvbg50lDlEQt0m+3tCeRa8r9e3GNgoKwok7d
x7U+PWoL+9500yIBnVb6j1MwAGBpwA3gpdLe7R8DTX7KGppe2TwVNL1Rkq7RCWqRQUaqAeQcKDWi
bf15fxWDyK3tYJyzmv9spFHttfKKhYBlvsWvKwg0Wg8aMNaL6D1maxayaQqj+o/rEzHw1E3jfYcM
42ZXv93ko7HU5TERIghHNybQ/SU25DtfL2YGs/IfkhRlJspHqaaYiROHjJICx7gJROS1G8wF2za8
xzBPyFL55gTvZstocTZ0dseW5Nu2hBQSPzfQUz8XmPqLuox3gFNRhyxTq7ArI1NuWGNP51pHZDAv
fWKTSsj8XDOPzGkc9q4mdCU18dRoadkJExj9A7MCTcxZcWnl3mYv76pP735Zvz9vyoapjiGpc7Vl
JQfLu7gaB8W4sxRwGHpug0KUA7pQ4DPGYo//ObLGh4jkX5ulm/iAHDCseU58GvFfbcNA4YNbZB3m
mXqfAIUuuAN3rW8VgkAguOZ7S676vjd3dcjX5+uOsOAccDrDfzc/bjFdg3lmLLwXM3uzRUXUrHZd
esrUDRaPpjyUEEH98rlvNQpY2uHsZvTCXn5gWlS5VGqtVdv2iO0jgzw0R/PIXlQH1hz+FnF4P18J
uKfPg6lbWDzO+bbOM5LsDiNIoHGaU9uW/FRjwbaIWRPnezFcMgftmpuai76OS57arXQkHsDcGZGW
cg5bqLonvPMU48RhHOfLrE57XZhG6LkM+ATx/aXNTPZZYBAZlExpEEd3h50PpUVbfSs96HNM4rD5
FOBnvZd3FxtsdGf51DFL1cUWtgZ7lnSXgVvRsIFCYx6Ud7Eho1K/XNVi18HlK3qaI4IAGR92Cmd2
V4ddbXWQfLzqKMp1swc1xeJSLw1XXQYxRhrcWwyNtkwqRCNTM+u9QHehMSeJaHB+kJcflcr33abw
BWOqOX/mfCGAG3C8kqLYPFvxm7rahwFrkdNMIHmRMzCrnh55JQ6pWDTV8HRt7lAuud35riAVpvYG
O+tXEbDWTkRHq85Mgtz+DKpzwQHUMaqZbsi8OG/PWoUFOMom/EPrVIQwdAM43V3zFQrbE8QNcQRR
Ca9vMlkG2PC1tKTv9qvn9Nbedixn9aC07fnoo8dh5go+YA8QuWub+gLuocvgqv5E9iZQLzu122pP
VHqCjC2Zk1AIjAeGTEBN1m47Iu1pfP8+7uOKB6zA+hPB1DZlfHyqQeXhO8+P6S1eCjCkb+WaSj7u
lvah+gK3etjJLDdrK45WVf1gEHwN3ppQnMt0V4+Li3nSZ/1TNi47FvJb5jsKm+N4GjFW+WWNlaN1
wQxp/PNne/M2XAhdB9tDGeS2MGTcjQcl0KNKZvvkegDBMJ2T91I5Zaw5cCGVxLC8vEieMsxFvZrX
2bu45nqY6e0PCniDYLGkbHAhgvnavDSZXpHT13LAqFMqAn18HTGIEB9+ryU1doDkIxYhgxZ4qRoU
TaCLOS/X02MxiO/TaXlMRRqlr8APwIC58NUcFhU9aZKZaDK3Hf+jbcGxoqbBQ762T+D/ATFoBvtl
AEH60HP0m5rGI+pgAS5NBgpi7Qux7Isubn1SalnpIPcq/IdjDTF1aTgLhFA1OjUEdXKMy8m4eoA3
ynXvW5f6sCv/NCxhjp8NaG+N3sf0f2YBEUw8NoMfbFKO6yVeTaR1B04ulS5R8/jhwfyo2J7Gp9pU
sN/e2bmldig5gBiPmKqclHxB607vHjidUA40cVXqXkzp1Un26MRb+daDtymXFIwa3pI1HGIms3CO
IMGEUbtO3ETeEYNGF0oFvjhYQ7wZFApRXpWA/78X13H1ZHrRBzchG4Rtuh5kq1p4I9lzP0ZOZpXh
xdNXU9/nc66p/qz74i/RopPj676hPhtDFMoIdT3liKywmo6ev0xjLoF6chzc5i+JyyU0BpGdWZzP
NIHTEsDFXHoBVm14zUWYLtOqsGedO3GY3Eo0YMPsBh0TOhExbOFdnL+eKiDz3a6+aXzP52WdoECC
sPADQJFod9vDop5x5DfhOzZlcN40P4KWNSC2APGPDiXFlTWYLWOtXX60fMtoc07Cz/f7KK643xAf
CL/4yWDIbeT+XsEnU/KCnKmDNIaspDA9k2jkMvuCZmtcMT+A0JP/p4nVgWOh+jP+0VvxIa2Evuh+
7kTwvVGP1bYKl1jEfH8H9Wib+yUmJeq/IwPT6l93gTaGteIhbu6WPHRUJpmlpiQ1+UmxknWprkkR
5m9SexUf57qoGO2ZqzgoLYOv+BDpNWhEtxlolpz8z4LlPJeHwZubgyus4QQ0buU+n4Or/kmSLboR
NKPzGqAsmnoZxnzG1POlpssOYuCBZwn5zYJ4nHJpwQl9lHjsozE6+ny1R7uEqM6B5qL4V4i+XG6D
4dCHBycNzUcA0hOyugyooOUT+Tq+NzwLOv9jSE5/gCc2+9rVuQl5bniBpCxMLaeT2OC3Tz+nYwJR
vmOa9zE5CuOcw3XYPndYkArZa3ncqysUi8GPLHgwpnUO6q+MKApoSrDbaNBHFdX3Jds77lJYlyHP
0Ane1rUzG8aX1SlqDdVLwdSBCbec0WSE3W5+o0YPafqsjbgMUqHVHURQvy195K1grA0N++ns3KhJ
KsKtsPB8d+4QnWxiXdFp+9Mn4Ggdnq5mnrtZ0ARTn2feYOQGanfvEuVQToK8bkhjjleTmTv7o1/x
ufihltxcfvvkKbm8LlRQdcRlY8dFAJy1o8LKKVFhZ/zVlCPyrvRPv3LAqJbZV0OHgUs+bXlYVTso
0/qNseBRb7HcKGFnmjs5kYtyxKvg7ctCfcHrJ5v8w74JbpXoMud9D0EZtt2BnEIqTbZ8bdtps22D
wd3oaepCsZ8aS3E37uF2uLy9AOB6O74NSHm6XH3sQ3aAuQjzopdN+FxyuWEqP/yd8w0FizzF7GDQ
bYc9shQtwAISKvezkQjCHmlBfJFxS8gNPrPYfGwxXItztKaAO7skucHXuLK7sKWsf2buA8EQ/cOe
EtD12Zps+wJ9I8mWQqbVw4iWV+8AbgmOmFsqQR+6SE2Ylzvtc+c/FaWBrSLP79rW+rq2JodGkpVQ
vd2aBRXYDl+k7mdSP4G1KlKXxJvD7qafzsoxrQeEZlgAIBLJmYOgkpG0VIKfv8MMC13P7f4rt/F8
Ylnv2NRB5TDYlO++WnbwA/gKKs45JCJLw1TEKTpv/DU72DvUoRwGN0MR2u3a4TPyJcCOgGTJmE5a
ffX9kHtgjlSijUTGO4iAzHsD0tjmnTLxK6pPER7n2K4ksshnTaWNiZurSZa0GLPeuLDs5FN+0TG4
gU27X+sDPclgZT0km0b8tBWSh+kiWUZfC1qdwyPIPpvBfVnxdT13DYdUqNeQ4kzC04qTWM0RJ+Hj
61NeQ0N1NyXaoXwI1kKAYaOhidG3SKTMVLhJHG0O+G1SIMWy8H47MQbr+PpADiVfk9XLzsw/38oQ
N58ag/lMuQKKhAcrNzHniddcnBcuyGSALkRXtH5DZ800JjMYje0x5IveqVK4yJGu6134TX5BoMPy
Yla+IwgE1alTlgJKF5h0T8zlI9v0iNklEpdxTdWnDAbRmpUoCTd2GHklmwPGqBE/XrvT4zVTCINL
ctft+44rDg8n7Oy41vfVomeIpMysAYL06Ti//INQVBn3kLssCY+4Gvdgj1oNw6vFmXpYaCcxmdg/
DCqXGuHM60uOEvOXPvE2c+jKdkOqRs/0QOuWoo0ptr6+6nOYV/T5dIByfDQQ5aEuHcsS9CHCwM71
qucDwsVvQfN5JI88uncGREJm0UwMTnmZpJRajILBrl/T6ZAmo3Pky0ArjAN/QVzWVnpPXTfT29tz
pbRrPABfGa836polc3ub06mKe5UVN3ZuGXj9p7I5ogqOOKQ9VQt19nBnFCoq8Uofkhi5Rmz5ejmp
NHkY2NK6+p9Jy2GUe3a2MQsg1KLZhW2XrZueam9KFzO0BA+g199x01rWvkqPGtJ4brW2icPD0RXg
UNCwUVysq32eNVhEszVilT4QLRYpJJarJPC2lEY0ezbDBcOaoJJvDOm8akvJ4cp3xEdnG2Yj5qIs
tNFdJyOG44+LEijlLn51QPeuG6oWdcULgaBLxyUrj8ro+kz7KXrC7MEOtmLtDXFR1/iB46xToJNP
JhrEdMpt+7mYgYsru3dwhGAn/b078b0LN2ln1x6W5hOaqeoTL/7h1BgBAHNYvJspi/XQtUqTEzas
5j9Dp8T7HdTTDlZHjWHYqsYss7ItWYjyGiTQTYw6cB0u+OwmqFbs4JoClo8haFn5JLRVq2rH/Ux2
3O244vdPmQcE7UDh5hRoeTxJ77Hep3m65mc3+wMZykEwYXYnuM+DnUU6zFhVEvyghag9aPX+cT4w
4HV0vFJJ0SVDkbfgjTUXI12xU4m5V75v1L02RTkBjzKuS6UJLY6rnWpwWVpM2IBJwX2w8BC8UIY+
RgmzLOsySe8xVNWE2DcrSQ5TL1SNooXsBjUW0lcWgy9InqeGqFFIcrYUnUOwlPTUNkfNFiLIq5+a
OnPq9uqtgxsO7NKh9as81+Rw8ui7ZucBNxqaRm9DsWYYy82jvv5hhQKApZZXWQ6y2wbISATivyon
jWaJe+GsqdJqFsSF2WGr3fowNj3GXav5yaYk0F+q1sRENJbyoS7VaFHRPNAVWuuMq8+fkc2qa/pL
3oRtKCS/mCSsdES3MChn+PqsJl2P7/fDWrklzKK0DyyBmoyep9VtjJW9ta3qGTzOmPxZYMfVnRXU
07GG44UKZdMRCt2X29+2gHHpzz6YXG/uMAILsH7esc26miiQsSoWYdsnWmP/GCkT0hfjnT2UAhBp
rM7+o+lYI9ogO+q/0nrdT254DQIqv6VEJaMRSFWFRBAMj5TtvaJKrgcnVZYgHOmondj1FFwqmE2Z
jqbxYvd+o4Pqd7Ectv4zcxAtZZsp/UgZ2+0ckjpzvDXL/edkG15ayNIc2k3juIjJk1BrPXsE/zJt
PKTa8T3wq3vlm8cvIhZD4+3wROf/FKmrYuR1i+3RMKAMygkListFxdLqNhKAAzXSCq9dYBunLMZ8
Oxv20lk/V34aAOekY3s6lCnPquhN4E3FCcmvaC+NZtX7nfmx1CT++8+gD5V2OQZymYauhIH4/XFD
otPRI27showtDhoYb1O6aFojjiEYa2q6p53+BGyHOVbdVyb8d2xAFzajTw8V3edRC4GV8OcFtY8q
XCNuTuUW35EjRxKxiRPNwKCgBAzgVGfELBBx9lMjDdwOPLKMIpoQ0kq1B1wiclrjmdjCING5FFoI
Ptr3x1/wr0iKZuaNUdnAiFeRc+Bso4cn6sXUPhafZdc26VC945upjMaqxEdHbYtwbEz8BsaglkbE
LX/GoB6viZbWp0l+7R8t3uzUX3QnVMQ9CE7KsbEqPQiOkixD9w6oMEb3MkO4Dr2Q3kew7NIRrSum
pdWT/pUoBDyNo6mjObihm0aSY84/tfT95BN6YyTPezYNV3p8xIS9GOXYNzfYeOxqDlohrojy5EYc
vEevX/XQsy9IUPghzWaRJqh9yTNuTJUcDzC4x+PcjPUalcl4zjxbHUdIRc+valgavkHWI9WCobmi
SiSYBtODyj7L0esmeyXXUvc7IrZrvKFwTK3gtI4i+9SHphuyGpofMudLXqsxdej8Ci2P1ZS9aEUc
8iFO4HxVMwt70vTU37Y6zrJtjGx8gvePK+yJ3JOm9FLcFy+tomhhbSySMXFHU7oBmqTAQBBYWwG8
F4QJkg7ghrgYEELvjX53OiNZskLzaIL+mBscSzSlqN4Wpmb63atMNEJ5OTAlR9nMALshh3zAbx08
VfhZDYOg/XFjcrfsAhpmzf55E5gFanEfECdSsb5sLrX3mMh4RpM/aBnc32Km7DoVO6t/fggP/Bn0
37C//T0tOQDojXmHj2835ix/Nr0ljMYymTdAkNhv4UsTrg44ths04MOTjKXib31+AMvShTSxZ44R
kT/LI7h7s7KFAB86CzvoJGQ5vah15BI2Y3LFbHZxcL43LWeI4HOxPToiCH1F4jGvUW48xRXRF+Di
cu3gc8XaaBQ/zK5uEFRcooCKNH0j/fS7oPhmWTiZnj8iI2mX4beqNDkcmJ2RVuu9/oFo6B3lUXLQ
yUadIg7wGpgMa9sGTsB5bXgPSFiGI9jROQUGPpe7jDD+mWDdW8IHUkg2ZsfLecZ8Tn0fLsG97vbf
TL2/I5Co7GRp0uS/ppb4eHUIlRFNqW1rgzMzsuTgxxwqXFzFnlEl7pw7RHPIuOnbqYIBFZplrbua
zd6nbeH4PxThHUQ01rYge5FGQWdxyCJDscyRnhblsRjgRODsjsllx5qi91PBQwE0D5gPNCcrM9cS
W2TYzPrith5C1GHZihJaPwKM02RykWl6RSpyt8kZ1lW4opORYfH7aoBbxbPWcl6RZmXJp4ciT6BF
DVmapg066u2mcVjfh6NruQL2wp7yBlV8IDHJUYWaeVBA4OpHKn6ytiRw26e+TqX1Zls+/8UsMxVE
qjt8bNGjjRz7AYpmzzDSRzb0JD/MokhIF+HuNuy2r2anuyIvGT5Qm4DxcgDAmFlomZ95A0s5/RSo
4IB6GxbTrx/vPFnrWh6EEvWO84hhsVTEUjgO+3/QxM2lVASdsm6ck188Zkqc/4G3gwNY7iytlrIM
V+SDKNsLGRj95tYfYKmfLeFBaPCWnAF2eAtBqREEJ+sLjSYjFVII2VoPyCOY88lNqSn3uAa0+9ma
FK8oKLoEzh/5414TYXiXqudHsaEmg0EVoiA+PCvgVibOpkCuf9CDIwtHLJkxax3QpmkrJUedkdbJ
Oo9ShUpKdJtPISSTMujxSyQxqFZx1zT9rInpxn132NjN56lSn3rwEwiz/sd4NpcVMMpn8epM+5ZY
IYZJnTMQCTxK0WCDRfpL7I/ynzqbkTeoSD1uU3iJykpWnrjNbW7aLjYDGR7086xrBDU0m+ofNiyZ
kp/BBUUpzKajn6RXz23DyO1iPsaMRZ/sKDFkC/hf4Ji3ak7D3YsAYTY72pkJIqAn3XtbUIKb3ing
N5w2D39rm8tLRvlFHGKq9xeRp8aS8IENGxoV2mphzpXmaruXEqY6Sjh2CTzHrF3g9k/lEmsMXyjU
7/kLlbjIg69hvUMAe+9wy2yrbfZ9ht2FjnV6SWfwmPIX41g0YZ8jJu+3sMZH6h483DeOyks1hjnC
l8Kf1mPEQ7Pwoo1i68OvRSa5cuR4c8vnmqhQ6OlUuz2zYvMMIscFx7f6yPoGgCULu+lCEucMwT5P
IV6lNaonus7HYsRDGdTVGfIIqZ1pvwPqSjzrejLIKmNRPqoevqb00MFGx8Lud0aR22QHjbBMXtIo
pAs/Vl/f6uL4HQrnn8FSxunM7BUziciVFeG5s7DItC4MsFpbrBXvei7K9niuZQh0+a42OiVDyKon
UsbavuZxIyml0uUYhj7VuvpiwCTBtxWmUvrqRdZmcHr9c0l5ytorVV+Js1U6NRPIelsLIBswfOV+
kdFlEjgZCnZ9Dp/uFlILOi+pxX1VjLtHgYy1/qpzXN4MI3kqQW7OdQ6TeJFBc/P0XFJhT3PwZ7uL
6njhRjP6oHZu0lXV0VfYNl3zrQx8MPc0Bk1QnWeSbSuH4APU4I6MkY+w7mF4LoJCXSZysECAmj1D
wTaIyB90GdJpwaGtKrdHRKQXZJefz/baK0nVKr8F8J1mdSWCXhzp7SvabwKVkokKZEuxJXEEdcm3
A4d34x2+h6vg6kemZmr8+2NoT5JxL//jJ8AUEN1Z9a2Va37nqACO7Z5qwbGYp5R8w3G7dVY6OfEJ
b800/aJUzT4/7YcbvZS4eZB8yw34k/oS/WjfAK8hMxDMIKiVaeRmjz0x4tz2Zx0b3d7X4g82rTcM
Kc4V/yqXk3lPo8sixRbz9x4OBSqqtddFDWgaFhb7vhGX3zs8IhsjUZZmVPRU3lQpjjfXoIC4UK8Z
bcENtzYCCT/S3ZdPDueDJZLiPdKSyaw4lssorBhplTuYFkOhrQRE5spI/Eoim2Nf123QOPPjleMH
r+vIm9lCr66u4pnnzuKEu3vSIRmliNWgVcqanEpFKc1qOajyBF5F4n6ldlqILb7HBo1oGMMlLGp1
ZTKqf893M6Ew+raDTi7t8grGjwPbOGDXRcig4VIp3fznK8AkGsr5TqFmUXN8mMQuaLgyjmMzJT1k
Ogt+SjLYeRl0k65xzz3co9ex5czf6PDCOjRLQQQuq6wFu28mOVRl7m4eO5ZoOnYFgFZIOyKlFwnS
lwz6zpeNEBeLbL137Pio0EcagybmJ5uhmCggN01tEr2V6krR2q59nXJeMo2o8x0wuIaqYQpbcSsl
2dZ6D0NO8QkV2yYpwfN27Cia+Je/w9pKnvPk6jc275oXjUuWDFtufJyG2WUZtyFrRJeoNUyUjFU1
RXrBgyu75u9NoM0yOymhv9s6drxtRy4F7yHe92MdrXdGCat1yKPOV+2XmdPSFzNPLndcV1PVqFZ+
xqT6r5kh7a8P3Aof0lGZK/JDf0+0BpdT14quU495ML/ZTMrfcmR+q2Ywt3yM8vOS9Mi/VWuT9x4E
rrvbxF8bBiQHSmRiYsAaiFrelVuzJgOSqGG8y4g6pnu9/qXX0epeSIFUmeqnc0Zp8vxAj7g2fsry
8bFHwkKTjg2GBtITUFmIM5YElgLHQ17PoYfzxOBFFjqoWxS99K+aWCyTTnkvXz1vHTMXf335AFWX
7OC5oG88OmYLVblfzvErTdthMorNn9YIDdUF6v3/1A/OKsxnS4mg91Q95L2awiy56hEm0fwgXcwK
F57Y1K8FpUV5cdcZ1S6SNApWlqPLDTAIFKFO11yqnWDaxrm5byPVyAmRYJA91mhCI45/VoyoLEcq
F0JsqQS6wbAns1OPNpT3HGUMC47JpxC/Ws+AtSX4MFoj8oZIUY3oeWvvAi8cgCk4EcFKrc4KTWYr
JYQIA1tdFS9Nq6OO6Wym0eA6gwAzSDN/legHxW6yeasWc0nVEz0985KjrZw87NR11gzg9TBMkaQi
gUCx3HwkJz9Lx50JK6WHcDlXFxTTK8ss2t2WlfWpRlxUTOQ3wtmmKMkZSKREfoKzV/S2JnnRxExH
L976dDgplqoQnTI4dOhqN7QK71gSsAGkBGTQmOOXHGs/of89wa2BkoAKbdo3QV8q/mMwpG7869LB
OPqhym0YDwd5PUMrkxzakpvr8wRIL9bmIUDThbWyDgoIz4jEWB5wQzdUZ467JCBqSyABvGJ92xph
wGcJ7qRr21CeTOoynAXoPXrIXP4p5ri+8kSsgoH2UMAI8jxJCKdE6wgP2IamQxDF1Vm8j9y0/1kv
Ts3lVwA8rMMJtcDFo6vwm6exC/RhSywHi4x3jf0ZMElFAuEodyA5i7K0QHYw1TIUFoWcPnRmD4lT
QkySciATOQ006eZ9gL3MDPAAvUckeKKht4q/By1dTcKJhp+4foiCXtMxazjkslRH8J6VDsw1iOON
rmOtGBbqJDmEprJ+YjPLKKB6EITuQXSpW+C464FvXAr3BAH+6jjwLTRCKb2L+Wfsqk/W93Pz42K8
a+bbIcmZK3jryQkk063iC6dJOTJ5tdQaswoRP0wK5RzvnkzJW7KnmPRr16QqngYrcXkgWVR/w6mx
BBEWmCZosx/djWWZbk09lvxOV5/HNjH6Gm6qqRLGH56f6lB6g9/qMis3AYcS6ou6zPFnhSLTz4Iz
WU7xeur0gECrK0/LZ6/TW03ihkjVxq4SYy78KUqtHUAtKxSPl8UPDeF2siDn1RmYtMQWeZR0YY0x
OSCLBclwNtqSeOWDgFWHpC5hu92P1Vj9nhdstB97oAklsAW/sxoJ2ukpCaj4JgxXcxMMWjeJLt+f
Kv+QqKQn13b0XmCIg7GF4Z0Iu0e9F7piZQTCgaf+p6ES1JnZ3n4SnjugSfX0kNMvkasRdEIMnRrB
P3neuBahcy/GYVgoxbkYodPad8t9BZby5BFezV3Y8UhKlnfLyXTHouxB88nCOOizAQsNnUAbKVMs
BdosYhH3pyd9B3NTNo0qvTW+qXGsZlNBoYJzYvnye2n0I6vqNIx1Nspnd23cA4D/3u8xdT2Dzvnp
XuQrvK49fvi8MfkD6xINfOSnS0kJMLhtW5YBJa9QJ5Fbnq7y5K8JWgoLI0gkmGaqISx2W+RKse8p
5XmuH1C9R4fJiKqZ7PxYHuvyCPZTW1uOdNUQQNDYQ5Fhx193QeJDEQj4m2fxiBkOjtoI8LbIZYDD
7CLGWsQtPGkCazJbDevLx1m3GaL3LDgONPsmNX+la23MEBamxgMtPOK4YqGk7KrxnPREqQpFUdPj
/SrJPbNMWxo+7kcmBIvg5YQ/96vZp/vg6Vo+dz+6av2W6cuofWozpmG36HpcMfWuR/KQiaJETOpr
7HLiXSFYB/gUCYdwks5jk7kV/V47OfumYDQaSM8xELP2NqP2kmstv7xd/+BXbEWpmk9ZCEXCAt6f
otp6/3+rlDc0/Ek3oVRO4si+27s85wwpA0VqdIKAwNq6XCjscNBpmn1As085YW801mteAu9nuflV
l71te+toE1ZBRhx9TL/Qxz0DEhE64iWIHqrI4Fn0N79ohUCcNaQUutNCOykgee8jS1cz96Q00nVl
P7G7Otg6Wq8RIRq6p4wa9XcV6rtZhdvM46SrTbF3DxocIvjmQof03Y0+M4INnbqr2TtuFp60ozc1
VpSAF2Vp7MoP/JW43pwzOC3WxSOvn+xX3KsiUK3sB5zYNF9tGCgvSkoYixbdNyLU2EcL4n6CPx77
PSDd9L6AwdmlsJzhy1Mqq+Vt00iXHQiMaBlBkwmjv6Uf4e+VDGuLWgTf7AljjxNikuh/l7HbF7hg
Enpzmax6jFfRoF/zzx2UR8cMm+qXG46UZZam4H4vzawuFe+ochqPyKeANJn34FpmewLVluJFVrEQ
ufHUxUcaFVXArgij4Dsdim3yO3zYbvSELc9yNGt2cbGFz18X93P6yG9Juk/RUhPvEzFncdvhjnG5
XeHNylezJsv+33o69WvkD9iCPEvpogvd75ehGEr7+Tj1x1EuTj62P3BpYGkRaU2KL7ub8qtGigDV
eyrr3fOlH0nCDqmkv+xYZfLAsUjmhIYN1Ndade+tGtG0eH7u6buf3vVCUKKvaNjjkJBW6ilnsAvY
iZq4QQQEkmDARBibjlNT47IzSXq20ZZkbbok0Qf7ce/6N5FXUQVN64cKi0fwGsQ0Ue04/t9QTyMZ
I416ILLnBGQA11dvmduP6AcgZjWElFLMVFzSJHcItiioQemI6T1DZHGNmSu5D6cGWEJ1fwmUdf6k
YLT41cJRas0ynli2y92J+ZOkKu4clRBmFsFTWzLU1pe+K/dBHbrE6uxTLsVej+bpP03D11namysm
ASR8QFGdroeg3NR0M0dGa38Pi+HVrVx8vq4OHlLubl8HAQMTZTVRcvSc9DcAijztdiOBf5Xw5Pxo
ai3vplP+w/DLvTa3dbf1n27OhR1ll+2uYWMfivWUHK/Zhhk3ILDkCYbaV6XOhKpHYQAQFJtELmgk
0zb/7nYwcJ13TGakKryI0CFXYfTPr0/KP83t5b8SmoFlJSks8JhakgAcqYk/ZuSa49ZGPNcvwgR8
JkWGqeLFHPQLcpEenQnQyGK/KgF7CMxT6tt2JQvzIZU5ArI3KyjEmKKo3HQn0M7gLvbo1MIFUAUc
rjxiSV+Xi3CqbBX3bA9aEmswe9BMRmGNk/9uVWw0Q7Yan/uxSqSIaUUk49dBk/GDfV/FUdxc1kul
4dEOIhzEM5ifo3sHrqYV6Lu8U04SSd1PDpJ1EbR5oAMQeMI2EatRmOz9hn6N2HUqDeg+Vb8tzNaz
Jafe7MzBYRiUO2YsKEbg/a7rmhjYweKr1OO9Gk3v5gRysMbywjlZdtyZjzhkO8Mn7ntIiRBV6SRY
9BRtV13HSOZ6d8TNP16Yv58TQ1VbJLVMwsPgvAsNslnJwRHDEGgRBB73jSbdFWgoDBygxt0e7JFk
gtM6wyRQgghMaKrqT5CzEB4GaNYbwodRTJ9eYGVyZ0E/131a/KU91Bj9AfRXXc7djTVzcf/sPBn9
RkYrHcziVF7W83WERgblWj/CRY1SE/gaez/1PLir8HOxpcva3DcRE93vzeQ0+/Q4qhqzPzTaFIWu
414z9LwjMkoI0sG/gy2GQgww5MraixSWTZwdTf1zsA6SwYtMQ9N0U41j0x/IEqQsRu4lAhxmUt5d
WZKJo7w/B9vpmCtY5AC1LNQ97dzGSYoRY84LRB333uB6nQ64jRrJIOp04vdvKUYOrc3fbbZoEObe
ZVsC1Th79NDUtUp0ETdRo6YSXSJw4m/9GLO205SEFu/AAaflwz17dxl0HnOKI0TuAGNJrkPs2+d7
EKP4X15slSIKMcBVJFY2Tj6f7LAGaAak2udrgiTgn/m8BTldecTvPNBx8GKhaItTdl28m4KGLhrX
KFlU+Vwy64344QVenoXpu6vmXbSNeCuALl5PhwWqAWB5GiSNSQyj5D0htQVU+7mXqhap5YV796sE
V6KHVUVDCg4jcRtYZBRT2lgnRDjNrLyFzihA0MVD1gScoSt+R3CLIbfzylwFwUiCRbGPzh5I2aZf
NtieteWvZOqKkHinq6Blr3SfE/3CV9RLiVLxJbWkZhdrIqifkAPKSnWe6hR1jLcI4aMwvNQ1wEJh
Z+5vT7Z7UUVoTc2KCcN98bKEQJE+jyHffvc//8gkdbvqM+l8C3hAQDLGXq7URfP3Vm6mTkfEp2GG
7jqMLuQxy82YMsfTXiO8vYrn6U4EipPgtszaBR3Q8Fa2YfwMz5rpOtMT5u3prwlkhJXgMhQ1wHJj
GVC2OsOuBQsFNQZ578cWYccBIxv1tL0g//EvhueyNn6crg6FImQQO2MdDUn5h3g4rb3RP+K2cZ7r
a2aXGH1JaK/dqVH5XtS2kNivX/+sXwW7gcOjvdteLw87NfQWSDTRyT7ZAI6tGNQ4zBXdQvLOoY9L
pg4K6RmQgQ5OXM3PQjJWqEyE5ZGOpHaWWPXmWX39Tr64WXS2SD39Swe41QuMGLhaQnG/gkzmT7zh
kyPswzN2bhYNrcwbpk1F+Xjg1wqyLJ0xIBFeg6LfItrKJhlKm/aQW7IOxwoa+qVQO7Edeg2q8pF3
KkKQv73YI1jBKB3Cwwv6tWufhvhwqE408BPYJd5tP6+O/a5eYfGZts/Pub4WQ4hghTJOE1q8lasF
vBWzNV7WRucekVJqdrT7z1CBYaVIatvvXdHIu4ToBm73DAOwzuThUe8q6HqJx1qr02tNi86+DYbh
vDO+5sQ/sRsgWqheFn/0ZwPHRr1C1/xEm+gQoOv1udUvyGoSRU1nyTSyg1AyU7xRWT/D+X4zv3tZ
EuRqedIVmD0TDtmC5ND7/wnO7eQbZ2BPEbXyZFDFnheCAy77gznpC/OMCjA5aY4B4+C31mzDLFs8
xF3WrcQvBsQlDX6dRvJbDLy2w3OExwR+toNc6L00zMh84mVpWHUatOVX3sE0mhGvXHiRbD0ci7wt
EBjqXVxmL3C6GLPjqN+Qb+PS70pTK6BL0yfhixC4UzgDyWbGlXEGqA2EqUNIvgjLSHK6rHekPiTf
s2vyVPalgBTtORf4MFdjfDdF/AGm+bj1qXbXCxzUL1IZZC0g6wfZVnuB0D6cmshdWFdULPGJfqQy
fA6vaiLOI1sby0qG6qIBKNSNsz1wUihJrifjr9jeiKQXYcpQvgrQk/+of38P5IH1SFGENwUW4lJE
ckLLaBUyistAArKM1GjueB6lJLX3Ph5PkDz+ti+J+UNXVvhDdPnE020r6R4yOGzItuS69RB39k5z
JslnSIqQETyvz4kjdADWP8GyhkjOUzu+VF/JhVAJDEJqikMFT+tFYP5rvqKilhzalMLh9ppC6ZCG
lrIk8yhqJdZjg4jsh9Bxsm0m+tLuNH0a191IaxDnnzCNjqrEHe1nd8tA7972RWwb2Alqs8cz3xYD
Ta+8u6HtpWik17aJULRG+dRGD4e5h7mnG2w3R48YFd+NPdfmd+13MGA4/oBRmC82Qw6whwbflZWG
QEhk71zkdg3GXB7z1VcpbONewlYh+lMm5pBuel1sdhcZ9ctT7C4JPXb7fM9vWPk6uiFmXpaLC5Rl
axK6piJlZ2bGdU7NhX/c1VWFYzS7lWs69gj+vS4wpj646Gm4dsKiZX8bUr5uCuU/kY4z6Dg/bxCd
YB2jZAw99zRq7ijtOQnzmOxx5plhqyLImyaLxCBJXF/Xk4PD3Xmsa/803Nt5D+mXngNNtXAN+IW3
mY6XasqRqotnHNc/jpaIz88AEAEnyEWTdYdybcJk/C866Zt/OgM6SIYriN1EH9jq37k6d6NYdgXH
XDKqlxGOC910XZ/rp8T3xiLTjewPwRd2tTe21TkuvF6S/rS51I+R1KEFLJ12EfJvpi7VIyypowki
qTd2cH7gDQ0b+Kdtm0QGV1GkqT/VUlC8X/0UVYFF4YDcD9F9qE2uDyQcSnnfWWw3070CuTPZRYwF
a4osCPAGxhWwaCuEGbHYKT0vwwIb7a2D8gNJpC5I/hwRfvamImQcEIYsX33s9kEHDiUcqPBRcIUZ
MjrPIBVbNyYG4KFSNj7XR9cDVCYgPwZZWtNSGyYerFeQeyKh7hZ4XODwjIK/lUDVOZ+AH2URNWFd
yqkyNb54jfzN3PD04TrjsGDhHOhKa+5ftmj4p67abqgIBCO6PnGOOoSfdOMk5FqBeiC2jbyxLMuh
qh6z6I1ULrITMIS+m+MkAS6PVdLt4FOSAtpEc8qC/bZhL3kO+47cfZivBVSBrtq9CPeK7s8uJAmA
GNx1nxPOJLC4itwDne6C32GxkiBUi9duL7ILfeRuCL5GzCVtRiP1HCgGXlX+lXEw3PKMhITnz6GX
sehErhEM8SIoKjFods3MX+ia3yDo/F8SBsTTC2Gplf+oVfPM7lKLTuZAfxuS8Oar+nbDao8RRqWh
SYDRd8Ak+yF939UleK5c8BhPLyM7XOjQ5/TvAx9NPlTXWW4k7CHIiZi9k40f7jQzfLLjqhL7ZbHf
do4ZtklwINUDRJt2dlyPUgyn5ieAvKqWv8r/7yXs27st/vtklc6sFUpv2f7iXUzJ0RdT27/Cfbot
CkMLdRM1Nc/4/lU8Je/ELT6ePNnfO/b+vHuZe/uCM0pYaPeO3y6moQOISihwwffkpDLIjDkHLKta
nxcVXT7V9aIrl4j9a6wJZzmfDumXC5ANCXjgYZUahmFwcL7d3amDdV7BZGvyx4X8ofCLvYrGc7lu
73VE+L8HpMp9z9Cv6nwInXyKXyWd1ffviql/uyjk8YExVmuEo+8BwCv7Fwt4QWWE1Pxs1qF961Ci
1tTHbC2+GVPd9448TthCuGMzt8VJZ11q1+UzjIQcqfyTbqWOnEFPWzIMRSVKdG/XxFVbFyZvBgVF
xzLv3ca1GM+FmtADbEuyTM0EbMp+Dxr3HvyVxlvDoTmowsfPIHsMLy27gqlNqEOM8VmI/pBTYrBs
FuTIBcLjI9Szx7rW4KOIlzDMO27TSBfEVo0bjLzjpM5OBU28Ea2DuKzNGwaBFDZ7Vkq4MK4EM5qn
DHdLwn9ez9eXoD5qKyiWsXiq3FeykdFwxEmXO5NmH7kLwZWNCW7JxZi3geT0Vf1cGS7UUoxsOLCi
ZuwzYFPAGeGD0MAC8r6q0sba4U4ZPame3bAh+ZZjNGeWHgcitDOtmnch/V7fiQ4CDsJEHV4ht7hc
saufnoUNBsbOgRZmGNQ2jPLcrT62lwnzDZi4KRrDD4JmicSEb5mIMhN9CzDl3Zuxs//DINb+4wQc
XzMHEjjSn3wPpR8WdITdYxW4+xLMSkV6F1irEXHea1fVn9MxTJYEo0+vgjNt1L24tOCABxsWHC+c
APefyd4dl/aZWHNLJZA6bWSQZed5CcitxPoSPY9RMrdtBDP6dFgy07kwz0PeT0Qpo/sXuQfz4kup
5xGRqCBKRP4/RpQJyIcAL9ZofY8YBErii2Gy3NjhsMT+BrUrU8FWIKvHz3YNlAWVasV9p3nwVmEf
stX2ORtdd15wfO/icI522iufXjPnzvkBHEjMVcHWmPtZ4dzUy7m+rsIWz8bFClOBHJT0zWwbgdts
gTkONLiOCSi+DeXY4wllFDvW949y1yeU3rcE/egZ4hDvX9peup8L3rxEv36WUc26gbgwCnzZ/pyp
3nxKITa4X2GgnSYuJoPIsRC5817vifrSO4nTM63hLSTv/whQ58X0lmD8LmRMPh37pi9ioAmzu+23
W4wVtMqr0UIGfyc7dHJVz9ZfsNFif7FZl5M3B5XI1QHnLrId+lgDtUpjb+fsadztbxy16Xy+dd7a
hNSNwMrOZwPNlkMFjGEcuGGIr6Jt3tNSFG3XF1CAg5HHxEJm2s9CxYhs8PXENsTgd0+pehEVOPcM
RwV6+RqxAvcuG6TOhzuPgHFAmXm/CMj2fzK8lrrFTNc1KxY3k/JZwOkI/qh/tqQBhD7+qG+utnbd
gs9XdFv5f5/Y/fqjuT8eE/MhIVrvmqhj740AU0bhGFZhH+zRxvdZwmkENqAaDKM0NIfuZhz0rL+t
GYMWHzLWbtS/LKX0t2XrKQYBBakrxpw0/f445DoqL9yZt1bml1+nwOqFjrQfZl6Hu/Gj8mw9zVi6
20LnUod3uGreuQ4ciY8/EOE845alEeVwT+Sag+AqhMGRgH114LFC4yTjfJy6GJv3G0uezbjRoZ4/
qRgevzUwYRmFfIwmRFnYfdVwgEdmy3nFBa0vYzj6ar18guiSupH7TIUjPT36jDxqvQGtFr5AVIry
auCi9wsaB56k2+u7DNA/Z7u6z6PaJtnJVghW1b6/i3QoUZFriE9FsYAZIcvNRvxrDVwxWSxapgqt
xAc1GQAQSWthqBliBo1jkJhden+M+tBqB7E6Utj49nE8R5x8uVguzmzR0t3h9e8ol8O5/CPVTj+F
js5Evlta0kyX6nceOGbmR0AHc/AXVfF/ZmYxPjh/8JXi4Wwpwgtiw5zAKaX6JieDrq6vu2ALHkQy
5Jdj/Fge2Zlg40Ct8SFLjXaDFmYGT/KYXigwrZW/sTWGh8JGHytTnF+nU2AzqxFgEmwwN2jdOWPw
WnHSptUOn26oJ+1Csv0KEbUyBrgdfNpefFw+9OV8T/pcl0TCcWZvbK6X8UJHYpHdCu9kAFikw9NK
GsMLkRD8RrI2VzPxWZxxneQ92rGIkVpQmVtdc5XokzH1+BUI2fuxEQuj8wHP1pZSCy5WzWu6g+yE
hxSVO+trDE4SaKfc7E82UMh4Ofv3kuww6Ue/rrzXyZ2rdre1qWJCNuaFLbYYyiJN3jHTE8zQBL+u
3VJsgFx6ygIdE6yM8rUMylrQnW6+XvQopGR7DgcYbZWqI+n5hxWlD+MU2WJ3zFJLkko6LQclM8E+
z2XRc8svQBvuPdw0OlVP/UUPJlIfDCXqPMACwcvE2dr92pcYjYka+xbNvbaj0s23NBZ3rc4p9olT
SqxXq9whQTqxhZk48S3HkJ4O4huQR9Kg7d+0EdtX6wdZQPnSFC1pkSRMNMP2jNTizKpEJUHzhnII
lDL4MY+IizXgm0aGSqguSNXhEY8Qn77i6OH2LypjFdN6LN6Y/jk+xl3Ngk3ahatS8ruaEibJyYJM
G0pipRHgNFX6f7k9DNI7aBnrhO5Y6FAxgNkTa/F1YFC1lZH8Tc6cOoG9Eo5Nbh/mJrNc79IHO39W
Tx19XmExYtCV4L1KAZVkD5iEXHHnQdc4Y+5tZhFVryKNQ+MwWiLC4bpEmbFuzAb0G75Xi+YXCbyh
5XdizQvdDwu/s8chMQGQtBIASvt0uggJYpPRu96XKtUMtd6sJ7CMrcguXnOT2FHTECU6KGW40nTB
qmDISiArHY1NQBD0HhoLvO5A0xYEarpY5/icf3CCz6Rta0JRLmzMad+RR1v9wN0u/jIzUdax/o/D
v4iICdtW0Gp260bOMk+57uB1GsMvOlE4AZnmdDfdqbvJYk/uFQUFyfJBm2XIktarY1H/Tkt2I+MO
JRBkWZOYn373CjXicPKv4nqzsVHyjBCGW4gx+zd2ogOjg+0iIymR6sIS+VVAwurL/Io8ilbSp15C
jE3q7ePtRu0rPTrx9xcfK4o/5fEUR3NGsxmhp+26DUttn/7YhaeHly1StWaIy9LMNutvFc4B7dxe
7rmNTDhwY3UDcR54Pj6h/chBgDjR8ujiPNYzI7okh26jGlpvywhS9mujyO/OFK3uzSegnMlgIoYt
ITMPhC5ExBQpyRNQl7PC5+cRshH50fGmnFHGMNVIfgM8Sh+AgGnYk+/C63VzUAaQughD31aSou9n
cpTUxxWMDOmYpQAd3SM8XW86MHyNsyyo+rXZ3OvjQGeMjClX0T9GEOazvoOgdRqcJKBy8NAkocjr
O32Ob/PBe3xMt8ydumG46tQzWYcrpdlylxnTWoCjJWdTIyrgFQ1VBg2P9HHmwXdO9SFeEwcQoQY/
4yhYkIofLs3uK7MWWgNt9DVVQOIwGBsBZZBwgJFR/qC/xTkHI7HTBIv7yq7Rx3V/avC9a5tjDByB
8ADvFOl1kHpzPNgegzKNlo4ZfcBH/eS+1zTBY/CmZxYM8KpnMqDjknaefOWIiYLFOByt1Prr/+9F
Ldm05tnCA6AIRlzGJPh9O+BgOKXX3rdRUQSnlo6aSPB/PjVJpNDuD6LE0TOvUhGNpKvZ3qH5oQCG
3MCEduWANgOvjScuS9whhW+NBw3aJB7x/mdf5DAi+PGOcOJvrcFoNg8SAM8gfFhiCq+1ODWIlojI
7WggdKgV9+1cN0uirYvTVxfB9JLQfUI6S14KuP35JNfLlmEIV/5MF60W2a3fPAFanx1OZgsO5PEc
XfeLHQd4mfSf77xdelFzX8sn/TWPCteIRst97pwA7RjxlOGGYdhDErNd5tanHQoezA9MtMvhcLAK
YO2IZmCAT7W6c5ckoh1TtUgjwvTD/99sLuiiDBR+eZFMbnMlsTTxyWI2/F5bgDeGHf+HKMgFEy7z
neAgjaG72187+hld+TwF/roj4yVSeE8PY2wmw/j6mpyAd8ZC1z4qKRxTNaNzaVuVa9VgLkMcQVfT
J4B++9WY0dofIP7cLce5pT7ajfR6nDQ0AgceFB6QRBYCZnL9K5orgq5Nj2aksSBccdAlKh7xSJhz
Re7nP3nuMz+qicOzvAwQCaGAahEUZ3DT9MLmKU2zc4CBC/+snGP3QeKAD5YXxsXIaoFaZGdTVbDM
Qft/Ok06gRgrPZqNpQ0+xkQayKzVtjliLGbkr4kYW+IipSxSXMECnQPG+L5rm2zVD4RtiOYHrN0g
7Zux2zaNnXtT4gdC98CWXSId9cd5boj4T94nOEs3vLylMn4Lwk3yFTf7u+FNbugm7rnW9tK9fFKt
d0pfMAikcP9Ol5FKmWD2mSsQIXdE351auUCL4B2ypk+B196YQYFQwArB7SqKvXl1p8y/3TAaqFXB
vSFCKUmS93u64vm1D4BN4TXiOAEQOcE1t8YQa2CvZCLyErORRtlJ1lChL0rlHuCjmaHph0A1aZ22
kiXcw7r8NIkEA2UFkdlj7AX61n0SP+4igQx5dAljH0Z7kDfNPu9JFwTN4KsCqQfcImbsWV8EyvQu
9OupKqDG/kT17SsUPxN+SF2yIu5Wc+Kbj7gEoJdE/hu3mo65TIDows+gY3erzKO7l5hlYaSAtIKJ
dS/yjOk4k2BUoQEyuR4mVoF+gvkfOlJ58eTRU0FS8Y6uQ8WIcJESAgjoPpcNhx+icLGwnlPI9xeS
fPKtRTC9CG8SEB/jXSRNC1Z5cHZoGXkAZaKKoEtHjSDMb5Ryj4wiqoN4PwuqLT67PsKMVrnXy8KG
QW/jaoaTlMPgillLuJuoE1UZaVjwCz7AAdrRQ69FxothFCJvoihmDUbeta4ssrr7+cA3DZAm23gM
l9ovRCOFcjUW2XcYH7foz2uLG4AFuRhLOQoHYSrykQqgfwjV6b6ebl5CuZsOXf2q9e3JXX1xDbpg
O+GboVvNP9+MptDzGHrOaQQ+Woba+EvewC3QImsb2z8AAlmUZLShcVz4UZ3GsfHTcdZ+/0TNjruS
lI+WGWe80R9Dpza4xDF3iDGIIkq+PdFPxTqZKuU3NfFLjyNOkG4av5x/nDqviQzKt18Tm7fb0mle
mk7ipGjElSorQZQet780GY6Cb9GH9sZ0tujJggHRn7J2b2UMEYRqQtb7wDqrOoXWuLqfc1rXfkuf
Pmy7JU+wEQEdS05O4rpoVEBZIkjzqq/dUOgU9WQIph9pbf834O9QX3TCv1iv1O0S7Pj699wJ8rY1
M4fJkVIhiuyU/7E9Nm9+4u0iK47Q7m58m4G9AGJI3faiGtjdv9b157q6/1FUVWBHeNLYPMLEbl3L
HasrqnjYOwYWf0cV52dSkh0LeFe5MbOvWSZoVCwo+etwoYWaetnaG+h3SUym1YWTpHzeH0wmxMw1
oimidh8Yds+xJRiHhNZqPEAe/yHZxQRhCqNaKZa9aJI0Zb+Lgmi8xkVFyiUlKixcWn+WxIBesOE2
5O6WmKDqSxvREtvnFCiT7b66rNRSMlghYw358dz2iHYthd5ecHkLqsbSOzCnlUEUjpgQTfjELxxN
h9kNorDqPY8fgq1jLgXZNWFwFc/6XjxDOZsN+Xl97nK7ObI8Ji/84tKcpi17K37oNiO6tsiRIu44
ry7xHzy5/lvb/TbQ25N7fMrYCDkT7uv2M5llPvaEvE1x8D6+/N85fATxBp1WJHF4+MManJp9XTTL
milhJXah9kt9r7mK764CDGNqnfGDrt7OBYSy4syUavkgQ7BqrIY/V1BXPTXioFEAH6eBgEPRwIiy
kZrg/TeBIDzM4z3oqOrOHSrRQWYuAJjswxWKJFD0J3mIk3thf69zaMowyMPyTsLSC5zV9/bmQHC1
Z8yKAecT9cf+ApwYABg5nErNsGaML86CycmQx1K8ojetZCBILCxpkH3u1FrMJtk9MrX1QnuWZaiU
ySwEgqRQ0e+DPaoLr4k/BBtz+atA99/LP7NV7kuzViPZarEm1xvIVhq3FeEB+DF8L7j63DoxoaJT
8qq4UZK2rdwo9MzQyzLYY5Bw89NOooUNtzrjtaMkBoY20Ohnu/iYwA8om8KYqfTbuHBHCUsVODgt
vtC4sk/7QDUi09HVdtvXtVze51cD3X/sD48jaWYxA9JXPXcILZf7R927MrBnKZvCakCn5mXFD80r
v05NCkyv2reb79+jJJuC8fhKjxyfQoc5gnN69A8Ga/pnYOFZA7Sigt6yxL1WKqMmCwKuso7/EnSw
KEGJP+lPRPFWzLAM1GnP9emlGJXzVxyIvpHEhWVU39QBd36W90zpT5Vi0MmWgmlfRkxTm854b2+X
l2KwpxMXJ9yvC/6eLoBKU6zIFegBUu/dqOMKKZMMu4TqQ1acopaZCmMGz/G6QCFzRiMCsBnfoHpI
Y421Dt6i9744i1cZOOs8bAhAwdsyB/8Rqo1N6nwzBU93fGH2KXoBx9y9H4HAq4rksOTL3Paz/n2X
KW5riQf3Db1XViS2JbCSDSgVwPrbEMpOJllMJjZ61XA2+PSG07Ihl0VyOLq2bqywu6wfZIEgIxEV
P0HXUfQNjqvlt4f+qYMyBcOcXhrjXgpYWYLxP2N/p9lgdGqKkLfJ5lGSnwhcC5KplyNWHLxW23Z9
4BFoPCkqLK6qbJ4KbKrb07uzdS5yzQKQbjI3bNWkzaWIyy0a5pmEabAKfpjrDrP4xh2cqbSYUbS3
XXPEN0AELteyOKMoeb2nyv/kLvxzfD93+3asIJV+JDvAfgWK9TkhkOj4kR+dFefWpyR1HsWU9AXN
reKrRyo13gl56mSGGaz4ozQ9S1qnfv1J543WgH+1D2SeVuQJ3NhyT9jAuWqM8KfI+0lkF1KkoWl3
vmL2Q/sscnVbHt47uLoyzF2Zhf901NbapJSMtZxQNrNW/XTJgK5XbqQs9AJd2FoMcHkhKB8jsMiJ
gNT26tY8mhMcPzIaroRf4wqJolB7j2nygHqHQTasRgSf/MlhLFdKTnAicA4vWoSDM5177v573VZL
J8zU+QgZMGLL28ZMTbPHBUd3I3mPOeKoQ1i4tPfqGlb0ILuYVGFWdxSsBQD9f5pKC35I92239I/k
XKHXsWUse/ffZoYJ8MJQPm8YQ+nhGzTMo/+RbrUUjgY8lmfHe/D8heH89dPdJLRHUQp3wFx9HcOE
izSIeP55IxxvQnFt7EQNIrW6H42IQ8kNZunBQdkxGU4ztLe9YQwCHmEQrSpFmNipka2o5yaBDkp2
qf6p04XS+ePjgifV4UT6Cgk1OmTLgP2wJpBWvajjJQ2RFTpbiPIHBNipJi5FjZr407cPYgcCqVCC
2+XP/fCiEG1jhGJ8b45ci2ZNR9yGYvlpBuTeUVTo8QVevt7uSwSMFK0OVZu3/tNhOhbNTItZWhMg
TfHCa3DwaZ5z7W9Hdry9DC9Ua+3nBSItClU4CRcS0iy4s/NHx20LbbtfL54ZTeALtdz5dYdvG9Oz
nkw7KiZnX2MxHMPwy4UEfhslyHEZ75KuX8e2QXoJi7TzVCGFp9sSLuVvioWzQ+Qy0tgJ0FSYmZG6
eSnxYwqnzGQGQm5r4nKB9wVs9ruTorb5BhRzu2pmH1eVJydlPl0HSetRR7RonRqvgIcdK4gK+T5X
gcwPhCrftw5RLgNZHc7Zutdk7ITRl2ytzU+xt2IdjYlolBig2d7pFsUVlb7ocasZs/B3vDwRZTHH
xaIB6poz76FNLKip0o3+7xKH0LsaIdJlTfPpck+wHFW4zuWhoWZsm9s9D+Mwz1sRYFYqMMxJjUsx
WYR+b2Z8wEiCq6HZDii4Fz37KgwbXU0tSMrvit1Z8yO2yLoY/qsu2lvmqzBmvGHiBIZMV2SyoVOI
PAwKsTUjZf5X2DrhhbecD8TYx8wRp4JjB7hIsu92HBA0tR5fL/iPHCXDNKOuOcSGNoytaRCNIwcT
EZmY1OgTc4KgzRHhkiMWmDWZtWWenHBT/6/KsHRJEP2nfri3TjvwnyvHBPZfe1WMBk2j0QC2iK6L
zvXakRRfq2MLDApE5zBq+C8j5YWTHEYkE40OjQxboaNBM1VeQ2N6/snIxyD3pl/0JraVPAJfiSyO
Qmks/t5N8E9loZspQQn3WxVp1PkaWltzCOdpemR1QyMm2shqtyEvubbk2GGPQDrw8Kc8u3+Fm4oK
Y50u5gB/CEc9mECutYgygTqRKs/66NHbPTYg3hPbmvjUDIxj+u93vOA5laWvXYoQ8+aeKwtIINWy
hze+Uf1+RK1v8hZCIt1ik26sF/4CYBUt/UPzoiFsv9VuQfZ7hYNh2sKGdd9A1exZySulHWPLHk1l
DPgc8b7rSBbH01sZORLMLHvnTeSDa5oNGFW9IsXgIhcu8h2IgEadMiU1ep6AvfQeakmBYaE32skQ
fXcgZxP5nlE4eAsuZDHgcseSW3WAh69BKMlNZYWtNOL+KIWDw9+3cAxb1vrfEdSr4+Mj5JitF6aS
xTn94ZUIvCMxopas/XPU46BoHv+1y62g8UlfGW+2aaxZU2cXNtUp4XLD1aeHla2vFW5Fc0DZm4zF
8IBpaJf8AD48FlwmQ2HUvuMkCWgk7qMOkp4IxgXVHQg7b/fzzc9m8f5Xum6HSycdIK+N3pdXoE9c
Tt0Q8VnX6CjkSA9Ka1sdQ/B430mY5vsfCQTbsZQ6wieaTh478o3ofZFS+UbTt5CD4oQRhKb4N1/+
5I0uo85iZdo4y8Y4TjYXbY86XU51uVZMshu04yT1GrIjzDTjvVUfZg4KfvLw5T9lKUROnSHm7KKJ
McelT8BOdypf0ez6g4spZzgbMXUxxW9JxF7DDBhVCmHSoSujeczo/ohw6/ddfBpl+rEYNsJpK/nh
KZpeKKU7k2VOOo9jculoIWIr/eE4Y6vaDDPzQDoCPshk5N5C2ho0MfvvfbDhNbLBIo05tbvVopHl
EyVmeUJm88k9/inct9hKqr9hGCpfwASb8ur2I7i7vQfpPnK5SlcHJ9KpzJks3KalEZjhk2iSCQLW
ZVQLa34mM2KLbaxYL6l+JCscnT9dHle1d+jTzAUpN1WUjIwUUg+3p1iWDmUO8IAOfQsCeQtTBMGk
PmtrflFLZCMJj9TKSEcOgZvf+zSM8UWOQqIUjwUM13/a0cBCtLm6vbzsssUYs9vRXdULlTmsr0TX
HY/LX9kxQ4hla9KN+jP3R10fNxm4CmkucTlLF/NI7HAL9ZYsZPAtGemeZ09X4TuTYHgNSPDXobGe
uHZ5JZuAnisYRWShLGpPJhEKcOhXOiKbE1bHHFps1eIgja8IIl/xKhSh9TyDOVzcWnWUDb7nHWfv
pbQw2v6kYR16OUeiEnHcrEeHafWJZ92YhWavvi+Qv388aFXdooa0I94gX2y8g6kJ7TfJhKHN9YFE
MIJGC6RRK9zyb61FQthyZQSGBVrJbPBpwACd+EN1e4H5FpEUpFsimDCw5BMBGJNhAHkIxgk7q/i6
JmqE8qEskWr1iEvWD/JzqtB2mv2uWUyi4TMV3ED8A2elcYaHqBQwPqvck+RAK0mBJqFTKfjzz7/c
jix2/KWs0uBAFTPEId9eebX05UMQflcyTE1fF88JfK/vnKEYIBUAQQy+UXBqbWszlGo6r4mi31lG
LaU9aVvo1+5mZy9J2nkEP1EPTsyRGXjQhQZxLDjAqXfiYSP07zuvH9Lv2opb5ornXpeTzbgf6hwh
Q0RsYxlJIwT+UJDSATVuJuFvZYvvEWu8kZvLLW7s2eLEbgYVJYBy6mdWeLf98V5AvSwm4lQgFm50
THZBge79RfMI4pHmMSJQI/NqaNRPGEdHm/PYcYwnpQ0fH6JqAw/jtHHezXqUipxb6vq7Tr1m+A6N
fmAtRZkiekqXmNnnX+M1IrNFYkqX8VpkHkId5Zeo6ak8+0KdGBRRmXsvHScmWT1hPoMuigwRJlve
mVyhy57Vk+s1Q9TmeO/cJJH0vUhLOwn/BW59n1d3Bbc00ZxeyRNYqlcdCDNA3ipRYl0bXMX5aY0P
2u6B0L+tmv8gBfQtodcqSp+9ebHvDlfsNcVlNzTPm2w+gm2dNgOJ3uH9mBUqSe/UJTSNK5YDrhQQ
o7QfGYriFvogDEMsr8c9nP33UWPugWGdcSF18Q2SMFA03vBwBC/Q3c60FiprtyceewAWWxHLA9iN
ORUilcuNEMMpM+FfZLxQcEPRj3rPjSfwes8kicJ4T5/752He0uKu2MZiAlNz+8NBrUuMMo6E6Fnx
aVJNexKWtUGVvI+IZW4LsVjXKW/D4TE8Qa3D4eY9i06b0HizpsSys3eoXtgp46vHGLT/sEjsf6FY
IZ/aURyrs0MOTlAiToK6NefzcovIm4fGzAF4lxYusuBENwUYyIeGXEhJwKD4v+HhwZiG+lZsTxZj
m9q6cuciHjZlX1Ell0A4Sh929kC7/phFjQKX7YXCv/TIr8n333edVGNGR2K0ruxEzrr9eO8y04qu
vZc6ulTmJhVNUbPYxuwHpd1p/t2utg3ZWQTlmnnICKhBIrcZkQJyVEwupTvpP3jQsbeDoOU/kgJA
JZU0LTVS2VIAbbXUcpH6WLHGy9F6xibItklefnRUQfbDIm6XO0RZwFtNZ1ECkM5Te3Dkn5E9/Z/G
OKBwKkVz5tFz0jHR3XeWpOcvdq1w2Y2TztlvPc/tSOqVshENEqrsZaNYDYitp+zeNAGSOOYL/EHs
u1fBRFcJgpSUf6IpFrFY96GE9vmw4Kuc1VfwY1ysDzuHcVV7MQtw4UQheQlIUZD3QhytVuveQnA8
M8+a8Z+eksPfstB75zxBUH25tRBiEKXT1frQ+bxqUtP3vEOsUGx8pFfmXx1T212tFSIU7S1Y4Xro
GNubQICyBp3OjadugLecctl9xkwKadbCcokmLrUWLjeUN48Q9Rc1h1zwsSPen6nRlDfq08hFlUoB
QfY0VnMpqgV04Sz1431vschvtCyHqCq8eU+ug6fU6fkhNV+qYU9EZFpMdewLrBqDm7EI+veWPoPH
Um7TxxBH9w8+z9vAzt4M2/VO60fnEtWHGIPjvXhnVMP1a6qgKm0ImEUZcYpX6oHp7MCWWWqn/Yat
vOYBB8D8Vithm2F4bgVEijfKKMGmpiz/3MKPGeGc3281wAEI2XXPTlJhnUU7QpcX4BjkpedaMOg/
jcdjbm6+M0bOzjv1jyVuSB0WNWjOiIAtmiAhzUjeQBAALl7zHts0pypRucUBP+Na720OLQs0gZNd
jA1k5FJptaF0vIfShSTMJjhPmnHIAeT6uYBL84jbeXBF1TGxPfvzsP+IZqjvQMqCPzEi2kJL9f7E
8Y3R9AKPsFhLIw82BD4zERN9G/Hh3l8ac0201zlD4MKk90FI2DOz6GP3vUgYK3cGXnUdc3PZWjWd
ta0/h/Bb76PoynnKYNkkrt4BnzsnqB40f3m5nRebsd8JwcVikTgU7mWFwkv4Ft1zseh/NR95V9SO
PNLtcKQipn+zEAPmpcVccr6jRHgnEYtSXwGda1c6DLHJE9ZUCSstThX1RWm/1ufaSSJ9W+eg/qua
Ylzw3LCfHuRnyU5ugCJyG9GXXR10jNiZQZJmZ3ieADnQqTcZISs8PUvCCP6cydDlIkjFi/rYXcNx
ujBkMuxgo/J0dZx8/lDS0ECziz0a3LiNAQXIKnMs3HNN+gUsvYWa253H/5BdNlqixtPKxtv27jg5
GFHOV25AAOrkqd8BmD+GSaAZdjocXRhsyzXpBlB0cVvZSdSAbkyiLEHJPkIBZNUZ6KjLJ1P7i3dJ
U3u59SJ9IyGb3rVVpETyxLsVCBOkrKpuQf1dU1heBadxeeuhLaFL/Bpqd8omlH9q1u7MKoH4bzoC
KIOrGKwGtds9CLHQT81Rs5gIL4mrJLbi8zH4TgPFfnFW8Zs0riWRhxcXq5QmGNGfgjv6BEHhR2Zj
G28gH035T/77DFM+LJdoqQq8wGBmNAZBzWrA0XOpqdiA82YJgI+eHPK5YjopOVcfFSs/qcH2vhIh
i5+iVBlEC7R8Ww8t+LthZ0fL3PORdTMpdnOg4uR/wP/honZvgAQQ4n6hP+5QiOXR4UpyB8g85iDm
r4Mjy4XVgTh67g+Mve2NxUAUWO0iaB0XL2VJG8CQFX7CoCPehBFYbA33VSuCkuQiIHyDFaCR0ThD
SOwdpwNU/33XOiwihgs+k/ED0Eawo4dnfBFmhR8yfHBIrst7qGKDry+bbYZqKkjeCSuGUInbEew1
6N3/h4yYLkkVMXvYs4090/H8Xf1Ktxtte05dxhKxaAySwzfze+lvL61COjU7rt/7a59SjuO3hXuR
mknrAluCr8B8BNPS4Nm6oo8/CQJbBx1EXaA1N3QKVzg7hUhb1kFNbDxVY52kFdthRjSG0u0rm9yE
ye8j1xhaYiObgtKJ4g9AAAX5s8dIy+mKmiW7FATbuzLTp4512lSMe8r1FNBx2VfHaqWVp6yIMPii
D2DaijaeL6HFRvOk/rSodI2zg452trdFQE6274hzsJG9fjMKTlptmTV/SCLiCcsvRfo6TBlqh+If
NRuT7uiXDh2FRXnZ48KHEsCNTOZ6K1m/57BQ1ThZ+oaOE2BvSfrbmoFL4hTJFAQUJMo+v5zOM+d+
btxSkc2yHf+HkGqHpn6l6su9nHdMiqQKsl7KwLZ31/jAGUL3EqStGYXEGHC3Fyap8tEfKOxyAXL3
ieHwoqIXLHuTZGnko11Xd76vfwIzTQACN6xkdgbZo3Qxw99aM11aWIEa+SJQGjhZO08+Jg+9aEt3
zqHGY0jqy8Rirct56Gtkf1x8o/LBCd+5F10cL9SLLzYRYlH/tpUNSqbud87YPjrRjEq/l0oZi1B3
R91h1kFWF2nV2sNShmebZeK8pn9s/bNVoQEjwb8E6v2VuZEZVjeltMD3W+DiIo7Mro6Dbb8cf8cv
L+IfOH30G/buFPwQ7v0ZuZwh1cTILrmyOKelVblh3Y8hA7dR7QTrExr1WwbX+J/JuhF3CBj8GmaG
cVyDoCZLh69k9pkU3TmH8phGC0jLL27cni+t9LhmKDOE2SY7GB0fvp5pL9q8It0+XD/crDohmGFx
6V/Aj1+uHoBGIHLZvvIVuuSH625nYm+JCkA1q+TZy/rM1mIsmm/3SvTWVvLQEfAMBG3aCVOpJw8w
T7HGK3fU6iNIeUMoS+3v4IsZbljougSaXVF5KUluionlvuaVa7zireiE9DSwnkABdyQ3izeVUpEe
0LX+xPeY06bGRNBrqtw+5+v0jdlFRDSkprgeMdMyPF0j6+TlbxLiAJUAQhKTpkyaQptGSRRrc68t
Kde8skJWMFe3KJ92ns7wu20rlXOZrQrfEhyKZ2pcqaQigX3ABs9iX4YQpvhEDhvsiMAtlgk7StEP
3DD8fiHZCgQLf3C/Df1SmDYHq4QLfKYKOX9OEL0Nuvtelw/6CHh+wnRse+hyHNJiAugIashGREV8
q+YOhbeuoXv/pSSusFDsfCgyZIj/kdzRQGH69L7VBlvyPS6YNvpRx4JESuMvPDlQk8pC1EH8vfMY
YCGZG8mrJbpuEnhX0VY03DA5j57ZnHzCTafRJEJE55bqe8i79LwXOAmWpmlCdPYWPw/oiQDQhkiJ
ieD6ZQ09P25Sc5GBZ+lYzmQUymnwkwn1NMLg9t3DcFacJsl5Unl99zAxWuznD3sUnsL/po+16eFD
oGni5xLcIOgw/yDkKUA0lVYSRrBNgu9doYtA0y4AJi5jQ3rvG5fniMBvz/BbGb5MqT89azWbu7T7
xAl40C1T29XGmnjotCSfGpoDSG6NrrTdeJR3ZTNha4oA3PKsKvJpdkPQU1LLqYw41a/V8OCe2Vm9
BjEcUi3Hd3k59Rf4ZYPvMzJRSobETFFsnEgpl8lEmczTNm657pXSiyiK3RVXSo1VWBhD4Ez4wejm
FpMy/5sWxwIGAxzR66cCHd5i/9el8ydME2YeKNbK0LOpdnYyvGIhoaxD5qYEF0zCb6UimRSO/cls
oPZIffz8BfvsqXvj4ShGWXxcxZIYI8+k2KdliSBBlrZyFy+fbfR6aECu6fLK1xBcliANiFfdSgMb
vZvQ1wcFfgCz0t7FU4YSYUzgD5zGQkDQlIoKyRr8z9Q8Uk8cLINypuFTW8VOIgUU6lrMZsXMJJKi
r9351DDa3Wu0bLRL476QT2/2XeuIuV1lYwIhpwXHe0fbwpz+3K/6pswWPhgULgRwTvO/YgF6K3Ey
8RjIie0Sfd2fhdUFLa/YUiz8/A4xxj80n6Ppmd9ob5CmjRoASsF3q0Dr+NM+xVAVaxRCah4DiTak
Ea9rzOdV7HnbQlkV65dyqC0naxjTSVd27ViTcE5HK0e72wR1XGMKxEypw/E81ElB77nxxkVSSe3f
npWBMQj4N6X0l6EHQYFsymZgsioPfat3QS6caTDZPnceFpmz+pTc9h6poEDr7dlfgr2aPbLYA4V+
N4DTkmgSnrdbjyVuKQHzkjJ5gy26T3e5p2eKql9a+UnJWmybQ1dsRYpJWczAhlpcDhxP1aN+gtSV
LPD/n6yGWRL8hiakAjaKmrq4mXA5cNgG9Koj/gEZdSJWv9H5Jp130FGg7pAW5zll86rI8OMVIYop
pLksFJRBqgGB9otycNMYaZM5QdiJVVH4aRJruLhoIUw7hIWyST1pgN1b6gY1sfaS+KsPEDJYDKuS
szGHgEQXsKqtkbkgVYS8aNfa85eEfTTqG+sIsdo3M4441+Isb8fIJ0KYmaXmnoM/HzvIoab01u2e
1wY1xxLgGhTKIrHR+fpRhkMYfO0BVmGZ8SC5VuTidjd/NhLJk24gLSpJnYR5RcilqBBmhJ7kJ0yS
DS95vsb4wn4Ug1B1G1C7OVwCB+IUKKm7RKA+imeyswd4Jkrq2ai43CJafSEXQ+i6zea1uJlFO0CD
Tcdzy5fFdgHGF9uvfOYmb4AGWm0r/12yDjlwCgXWWtsqMm++fiKKVZY4bGCWSGWsZIp3Y4jy4Oi3
Pumubo5GgSrdzJhei+celmkWQdIYIWeDIBAF6y9t4ng20chyWRnOPMZz8ImBpEX58qWiQEgmJFGC
g3ZDxK6M73RAGEiLgi2/BegwwzLtXlzk9axiFdokz4z093qS/g2vBqu7Jq9So1JF+2eSPzmRV2Fm
Krw4rv8BtHxJMpABH00SUsbwD09ZHdnGKjBMW8B8066DEzoVKU2NGX9rDwwMJwAl9trHVuJ/Ig1p
OZlOE0HV1st3AryAEBoLRZHYsAteqKpUqCC3+pSGRtx88VRo8VMLESmTUlxyFxwYySxxqi4KfLsF
Iv0/xMUM1qkcX5RmgxNfANDTOhWJ8nICxKMG68mcEcxAHICewlB4ct3huzjEivh6hkNzz6bp1u/p
jfsySF3630bbUc5YTrfy6jrNVWOcLI3VZYH3zlRl6Odh6KuSiPV33VRDF2L7EV5BewPV7ZoxR1aD
jZwtn3XGLR2UF0o0PLU91YVvvHA81ymRapAXhL/JthN1Z0F27xw+xshaz3teXmfrDpp6rvHB0YRR
so5g9x+jmEkGN2ccoS4kvMUcwSjIbIEc0TT+zBPMrRuFZ6UpJp1R25qKi/35s0u0smgFcNJI84Gs
anOJkP5iMyC6H+Y5rjMRPXnwmkjAFMgMN0s8XOedYZUnGBE638o/Ydbxo4ZDEHmYB4CK7vBnKvWa
IAbH5md9BPuSXUBNYQ9mO13oCjLpqCJVYQMzX45Sw178xhANkZunyDrDah4DihNohaf/StP3ukSx
84XBry8tnpfJ6ftxkRVfXkqajX6s4nH/tjIMeQAsZ9Nhd/1ULkXWejLj0HqbCTsgrj/uHKKPTd4X
CtzYlQihoCwjSW78qL/mz8vn7pGAjDBpL5ZW7knQIrLEPJud7qhaWRY0dQPtgK1+5xGK5DLg4dlt
4u/7uhFUXZfEAycNmW3RL5Mk+k7FctqB4kcYnBvc7aohJCd24lUzsDk9WSLVur305VI0C0Ehxi45
wWv5TXe4KP4iDa2rDHHlCMe4SoLfn+tVcffBrlTZg8pld8RsEuU5ckRCg5gSpkZQo3F2BKSgiExO
08JtvWB5xcCeNmdZjzhn0o2LAI2GWTgRVjRMQzpivw9daMTEOvixDi1+JWa1jUb+OY3+4N5s+3M7
zE5e0bLv2tLsZWtuDLUV/NlvAm3k71l3mA/2s+4hAD1Ro1tQQaIBUI3vqQt1FG9QarjpausRaefY
Vkb3WV+OiqS0OjNf3MAYIkNiTjuX0pbQhxIf+1uZnUXRj2bzyT/xebZp66uXMdLIU9FLHoKiO+0S
C0gvd5jt7HJbEAcNOz0f3pEFsRE7a3ijWZzrnMxe38ug75/lMyCqILDc5fazJC6izIXiyoP+7PCW
4b9bxP022wQbHS9SJlOMCGgmo3aio2Z5Mw84AF+EIRzioMHmOI7aTPYdtM2rbomfpDjpIbnFakQO
x4hRiqQuTnAiW/56olL/6zHwgwpgbscdrGqGIZ84Fs+1qUHXc7LbOnuRTlr39rREDw8nyzd24997
w1O2oglEiSKito8cBmGvywCqJxR7sNih6+bTeXQt4O8yBoGclx9BHSkYiHQ/yoFA2WKzEHwIkW+6
DPiywgEFHTL850FH/iviYI+o6uUizedfcUvMeraiW4dABOKkwtEh4eWM2my5JjPZz99/6ySVnefG
hEaspiS3gKhqYR/1aYHnyzwib2G3hxaZHLYN7LGLPaTjBpDSel6Vh7/BhIqEOANgWyVYYrUrdg+L
mr1GxI84evfUrJvAtM5oa8QB9pLCMvBCk5mzYlyKS5yhMK6ioXzWM7jpXYPW8uWeaEr5nGfVvGPk
59JyCt/N8V52lMjw6jhdy0XiAioVOloIb++9PqADS+9pqk8NHgAkIMAeWNgNlaYW0K2O+s+cEj2j
Bsi3CseWTNDvFVJ8s4KiJpWFQo3HCdaaAPecQQYzRUNQyZGcQf8ULZYTwoXquJZNFyu67bLYxsNc
v/4GwsJP9MH9nsRAjexvcrRALS9tC/rPfm4Kc7+Spnk4aMgH5dPjMceVp4Lw8skKOTepyfM2PQCX
syHtXsn2AWjjR6SwnvE4/sA/D20jIO0glGHhpUNPOUNL9iT7gjadtzAeap3iSUeP3seBxj4ZYf9a
nzRbayAWc/rT9TV/pIg37xqDquy9rTN8tX0CGpEOtr+cqyfNEZFtc/mNGZXV5EKaJVV4IkowfQTw
pNQa7XZtuSJpI6UkjN5V9OwnPIVwqJB52jF4Mqasnc8AbfXCZ0ACzG/bpzwr1UZoxL6rqYl7cROA
EeTiFI0GidOurFlg2+SHR22q9Vo2aLhWHAwDTHr74O10myCIQhe+vuS58diPqKXwfPWOBvmIQbx+
8eJhH8Mwi+ZAOPAMfcpIZcrY+apAWar8laynPemmsR/f45L6pLkxjuVSy1BBt3ni5WFbpCl7RO7H
qwZXPGZrYVMYjyMdojNm1IrZRaCKrNvD6uYxk0LPpHCW1pO46FcuD+hke/c36gXSp/t5opIXzQTZ
V/x2P/BaSuMhk8A6ZtnTO0pSm+XCssCaIAvw+UEAUf0e24UcnuFYJHlVYKwP7FY4/StSNJWfZiZ0
JOrRKk1MyiQULwZ1KCAkixqiIm5sscs9DCZoO9TO4hV72rX2rKBGb0zLmVs1rSSIE5tjYNNh5eEP
aoVQELR+eUZKYdlkjLE4kvgeoRH9mD0/zed9poXxTjg/H1/zJHuLZlbr87k19WLIAq2ZxST2Kn++
jq5y7OEezg3R8Fiv4Xrzx289lzX89im5ddBApxs67YkoAFbnp/zYGEOIpk6/BHgsNAuIPxiBEiOe
O2j0aIZWD3c+tmUydbuPAUFPqG2XQfD4I1dub/ItkgN8fnVA/IxX0xva7SUuFYXkO6Z0FPB9qDT8
WGbNN967XvNE42PPwKUkYBv1i6yTTERpwI34yRqnKgL6yLVK1pBX2MrcWcmQFrZZRuaiXXelF4ck
0tCb1f97UYKx3VFAE8XgPHAPnSJ9NuktCQwin8NPL844M6I1tZFxHL2JEjf6j5gorPBiWAxCtp14
CV0h1DU5+m3qp3H/3xmcn3uAl8nSJuUWjkdl66YnZJLyeQLwu6UP23aINUw4J6hf3uRsXm1TxnKL
U0qHcJ+GDs+ORenAfLLS5o1BWNc/2lzDdJdt3w0WkUBZzt7clFVGx9gu6oljigajqJMh+9t+BH+e
2xSEPFCNKLVhwOmey9ZSu0VHFn9FZJILSNA14/If+W9jIQ+pw2xFpaBx3eNSeqaW2syv/Zb5PDXc
d9VPvjOTKG4u8ITV3bhy4Fo3v/6kt6WLslOqW0FwTp+iPPTg1GyTss+50r7jRzNqzmqL1p0N+Rpc
hGhjzZMJ3XOowwPnvk4FrO/joxOHHLKcMOJi8ypI4esJxO0+pMKSeeN3w6v29CehupRVo4mImLBB
2LskAO6/8cBgnD2g1ptUUSl6khDkBvhshdGgeUbd0Ejog2+7IJmTalvMdQ28qV+u/1rJhhvp9QIT
ajCityVQl0f0QJ/BBZsFsQqh0UoMeFZwMiC4WFGJhTo6mFB3QYTpEmRa4oALwMMbyMCRHP5nnUXH
cpb/sZnsM8GQjJlyPk8VraVfBBUpOB30aQNhC32WQutJ22vRpHYgcJRExZQgpuzq0m17YvVxsXga
CUKJ7u0bMej9HYsGSP/CxL8vwpDv4ZKwRzroOWbY0z6VOMR7ieexBr4WUww5sHQoUw+5qoWUb5OZ
zKTyUHaDSjkdKt0g9MWSIvsxR6LJBb5UjBw7BtxKZPAIcNPZRopAQWU9WHH9BhJhh0GYVpHdtd0a
V2t35cq3+EY0kwqDsOt+Z9VDeyziK51fZH4z+Tb/ceBExCwELAawgipwihu4RC6RPQr7+GLW2uC2
npFru1WpcZHXGmi57xqEEs0sThE7zUtcxwodRuBaw9Eqff4x8KSOH0vYgXGtuQIb7tg/x2J7IRhB
xu/chwUvKNo7Ph2MT71gaD/5rliI8dv0jzf7j4BdlsGqzbXhWLvJ+Ydy4pnxWXoXHpcpsaX/Seiz
YU09G+7r0p0DPo+hqnRY58ADbzDlpJ5gcDI08mnlETFAOQoKccnOEwAb2Zmv5YYaCk+dciCPXyHC
AkDR5MjfX/oTkI5ZUgobWMxOy+TIZTKx7Emv21i5q0rnm08F/pXtq7zulzd/tymTfaHtKSFnW34T
VWOSHy5uWuH/rHmy5z8SXLM5IGmyG4MPiQFomYjijGXNsvPMWyXC/Oqeg8hExNCEeGKakjqGo59w
MucwvTH7Zp6OhRmDIZJeTqlUK5YE8GGiOwTy1EVGOEgbkQ0HNWwVMs2zOgFGmFythWWFgi9oMAXV
3DDCclsYXgIhMgjAJ0M3sOdFk7nQiy0/5DwsTSFQ3NGx1aT/wg891frUcbvqP85NDa51emIja2WF
mrswSYnKT5pv6/s6tUkEDc/3W7bv2AZ6gz6SzuYYmjw1wCp57YkIrfX8lHE2hsfEjmmjXYN5UBOR
DJgcNtPgoiWhAJRo/pEGDogcK2NvwlwDrHT0gvY4Dst835kEQ+j1J9kyCNMXNxeT03a5NBBvPwRY
aoTeQfMJeKDR6cUj7pFistalWQwn7NDSdj7Kqw7iNcG0m9db4Pejg3INqDHErIsLScJ8UG426l0n
Y2UZkNZtemkCSXqkOw4mrvrIzStlX5IYLNOIBpMpP6VvZFZFG1bpX1IUk8UEYLafcR+njPA4PliH
z4QmvC0S4wHSQnLfJ6qU5lScDhhvSocBn2R7/VTKF+0lTI8pA4WlpcqZ6soj+utyFBwRUu0gyrlW
/3wdoufkDQ1SjPY9NrPGhCTVncgyU7fMTZNQG4y8WHIJCIpnSDzXgnxVJ/qa1encrAdnt0ECBeYG
tTfTZrINl5MYs/VMdGL5GNyY7mT5qRcINP+Ly+NoJ/joPXojN/aE6inKW2iVwThDVyDEqcQU8kU9
fvKoZt+Dxg/OMksl102Pt05AyYrMrlE1s2Fvzc5xXYVwqnHBknVsV9jTdfIvMdJF89CpknFjbfQb
Hfu7vKBq92D9xhwd+bf4N2DZczmhcZR5BqDwrjU2anx0BbxFUXCCVpq1dnCIB2sBFrXnU5vvdWNF
fxNUcrRIujVlRwqFu60HkZkpTxg06hPX+UO1v6pQ4VWNT5MZhHuTgdvdrhTATtIL2HgK1VyaLLTi
/b1kamY8sw9LuAUDUJ3fae02xg0BDO+u66s/2psrQIga7fLzvKyIjBSUoSq8AjYOkz7O2VIDE31Y
LhiBPzlwOjgx+pQF3Q8sNb4OhAtm/fZNMY4Cw2XhGG7U61ir6p+6mEkDBdHsVYPwVN342zkIjBeG
NGmABFrWgtoJEFiK3/GvLigdH6ih3l4AL3sFJb9lgK7m5003XId2oE4w+FHDykQTjoGyI4SUr7fB
hVf2Ni4TF4d2MnVqbjv1HJoGl/fYLAo5A4MNXkmyPKQg5ObLzczV4W4YmqkQNV7nXdIWlkFBS5gi
S57Yr1AOeozPgcvTh5x+VqDp9hXWWvPjjqf8seutctUT+884M3oNpbvEBjPVb7dsmYwpq8ttm/Zn
SjgQvhwAc8ifsMCodWEOhYI3e7BDqRV/nvK3lgWjVbxVaNfPP7/Fqds8bgMTyLE9K/Lfssh8qPYA
ZisR4oKxCVT1g3381+nzHdjgqH94ZVAJCHXBtmxXI//NX87gNrl8B717qY0PW1bi/LVhj9qj/VrX
0dWmRHeBermtqLJF1cFtDMIq1cO6tMLdFHtMmsAgJaBJMWsBl8S9LF36aJUsr8BhrrQyoI0M+weo
ZltLAph6wDAW47mzQjMKnu4DoJDly+4uMdzL2V9pcANo+5jk/CdOUBvlIpfdq/MSqZhXPFTUHNT3
SWxIOqTNMTMmjvFGldcgoDbw9uyRLzUcY8yclbAx4UTsQP5KRYHqAshiQUWSiYT8roJcln5W1m9Z
/0MqPzE+Fs+X+v4V+9STaBJUsfksRW7ikzYoxpIuomcb9V+Pqv/1rh+dLe0ZZAdIQxnrvobCyOyM
7S3IzNJtTrADuGQnBDFg5tHDBlS8sE4j8obJDriZl+aer1UUu9TEejglY4SMYt0W03Xxobe3vrVn
qJzTpkrmx/Lw7UY35BHk8S5XK0zEee1AnRaEN/I4LbHVwu4fHKHzZMgNzazb/T6fdJIHLkt3yPhE
l53ToDN4p/IFEykqEQeJ5XxIyK9zgw9O1E/KutEtAVq1AAFEFGhVi0cjfbn1y/fk/AJgIXW9mqyi
UG5yqYzMXin/ehJgJl2gFyKSc35sdwjn47ipl93hQgujY6IGepzz4pslDStyt/qlM3iZxENLXIbr
gvA5ozwQA49CmgEBkZg+0oLqCF7FbhcCWtY5d/zgiRBt8C/ymjXBt19F/TIKcszLJkNXE4DGtM4O
R5WY20+eMU+DVTmZyWEUNnVhE871DtI38tcFw4XF4HaQal91GAJlgJCFyCkSRap0uTmC3EYKhTql
TnNBVkbPzYAToBBwQqq0J3Q4hs8XgDGSBJfOme+lP1avrMK6R7dzltgXlypijiaPmeYYM3ceD14t
O6WbLdMqvIcZ7r10p85ffURLiE0N9p1J0MTacJ+bT7BFzWaM+qXy8qwp4L92j9/d4BKRO1uFVjrr
VRx4Ux1/T6xc7aQK3jDWwvOTQse07ciAZLB46gUGYkYRm6u6zmFsXr5mjABe5aABd0j4lPE8B6Tz
b62TYitfE3gCQmZAJH3F6yLwqKcc+ggnHyHigzgj96ZTOP4U6w6fipfY6CfZFcVPvE6FM/vQAqSt
1+8NMlR1DGOzqG0C28A2R1VlqXJ4CDVxIc5AVtrpEOSUiWhQGkQKkJz9ktTc9jamcXIO/Q+TOYQ6
wcUV+T6c217J2iknP7s85NARI0atVMKKkpudOkWs3sLbmQEw6ERW4eKzOU0iwhQVbMVQEWByQ4wm
RqUnDZXa+QtyfegLh/UOQJGnNuPJ3CPz+ONmn+GedxFKrTy8hWqBBgTIfJWgMe4vkyCZW8SaJ8Gl
wG3A2+CU7RXunCf5Oa1DuULr1E4j7EylVZwREuA7HJWsqYT8kAmKILPhs4RVAqDEIDZS7lFu9vBN
leJrrY/OjzPv3i57aDPWZI/Ki3ZltRZ//Y12dAXRLc8SmItpL4Vug++CqV60ANcYQSZG3xEo1Jo1
SOH/TXgr2/O5QFZaelWbrx2/j96WvHGJiVf/f1HzivFv3KENLtpud7zaX7nPKW0dkf2O++NGojep
+TX8XAxLNfeaQV/cl5KV9+393lCqcIVYWou+RsH5TUpW1f0ynKokwadma7jjWuYnjcmOP7JCnqQ6
b6c3aN/CzEo64cSqZlu4vRjQoQNBdNVOmUexDDQQjqh9eaPthd0s9MZEsWBSAuGdJoeaLXoeJLdL
fHMDQLvWK0didqU8sU2sM9Gc0toP0vSaSt/Wp8cVgahbMFrefUtZTkmFtWGwQSBgAyjFx2Tok0i+
zzGtA75LUYI4lvyDJa7EOUymdMaCa1iTWpX2rDjsemYShc0cvQ9SuYz+Nd/dHnPVob83MrJaBYQE
WU1mJ+b+Tf2G3PWEgKiyaTDI9uCBANeCskGkpwr123udL7q+rknPLher4fBDZTqyY+krBLIntoJq
H/6EQtViaRkghqd4lJDCD8iZMVEXE7Fa598k+iv8/s5s9uyAtXMmaFP8PYlt3CEyoi0zqonmcgvF
b+f52pna4NykiAZR2i85e+BIJX5AzXibqN46SdP+VgmvLcAvhM/M+1MbYgRdICD345gOBiJKAjvo
1PlZoFMmttM4g5Kc2V57CxyWjbZD8FhPT1T2OpzrpvzXrVgxxMd2a9TE4aZCNWbk4dLWtOSYSRo2
zSXg+xKIFBEk0OhOnnUboFey5yPUaNRdZtRk5240b3v4DAqlgoTP5JsTPrNfuyyl3nbtVOh5bRMA
0kqlViD/Z7fPBszxxkCulLtOxiJ5MEv3hgIJHXQuK+bGqoNHhET5riH1IZ15kvFODukQBvsgl8en
QnkCwjTh7qfdBUjs0aWbjy4aSd30hcmFWIVZUE9dplKotyyS1TESa+xhx1w2BSg1ePMGhjr79n2u
YyjMYttKayjWUyIp6mTqKjW95hCmmFMnNweu5JwXUi1ADkRkhSinA7XvBYPwTqil33Sig/esNbG5
wnk8UFvFQtiOi2ZAsH78MSuJxqqx3IZ/0NnjfjAgMmYjm7KMsx9via4yI/dbpS8n2RaFpMjVwSSc
Za27iCkzKVX7KbUdQK9NMIL9SoPXqJCRZzyTZmMQAdU92iChsHOZin2eyLpspUsWhMQ/awWDiSgf
DC68+o5u3ZwlzFG2D2llV5OmSJMh8RcNv4uhvkgO7MzluiLbaug7Np1NDQmZUh5S5ok2hgGGb3Gn
8Ph1LgiKOcH8kVSNSNeMdeg7S7a6YdUgGsDAXwzDI7k8a1FdljOk9wu+MwrGEO/618YtNFTJeUNT
KTEvTTcTflgBtL/rchxJOWuBtNoJqLeOOKMVw7b8WKXPkVtMsaYpRBf8hG2aPRwGfMnErypSO3IW
EDjvQYSVYE0T7Mm38tVtT3aZZiV7H7Wo2hQVbKhko5VNhs5GWATrVr+wXK6+xgaaFdW0TA+ITRxo
YI5maiqDwUWEaqjTh110RstCP5T8mXPbpCHJlRU4i+RgkEnpQ/Xhzf7HeMEj1vI5Pr9z7disGmVo
XD9wAv4HjXNznNSX0hg6eGLKh1GIV+tnEu+5+s1sXhEKbyMzAGqH1QsQ/SQezHOSXCoqmhyH+7Wf
+EpcAty13BoaNx96deJqMbdrDb/R5lXvhOK/xFPX8lHCjoSUykzaic+fWZqG5wu36/WQuuw7m6qh
XLs0b/PIXSBSO0pv2S4mDuaVE5GCJFjN6jj7yUthc2vgNx+viItrHVWUwczZH6n0irdBgbZyITjv
X9E23UY0K2zu02wX4d3t8oQ8toX+pMa7ixG1o7BSe2ISM7/cjcMcQU/II4a8GeNcl5pkDBYpDMkc
CdPI5/CiayafIZ92xQ5Cd6+XKSoYUzAfDAEEI+P8rfKEx4dtDI9m0T5mB+AWj9MEWKwBbIaGTJv9
y3JMscXdCgAONPO2vYlTr0cdXjQgr6V2EbCUGkwA3paNg4EPVkLLOcJ/Tva3zjdzwFeZ7hQ8740/
rVP1NXWq+2VfH70axqiqgGg07HcKHefoQaywwt2avzscML+/85UaQErdluHEOSg80LKnccdwiGSv
BmjKiA7xUjD/Y8V5BoLYqg0hzAPWjxB/dnecQNMgrhY4DikJLVRCU1b8FAQ2iHM5wuMbSe8oJ3mA
Vde4F/2Z714rI3HI+9+PA8lBRD3vYqv/Jd7Nye+ZvQfA/ls+D3/j3N62zJRbuuqDpbvGOEUVJmi1
wmphNIZPMBP6tRJndH2ZfAg4EbC6fYfX3I7NmDhFBERhVaryNmczBT+Vdoxd8zu9WYjDzHcMnV3k
a3V42zqrIpqx5xbCzoBp5v0YGu316oZP0imHu+fnZHq9P1cp9mlCSZp0ZcQCkEKwrP0j8BVNjZCd
agME2mXIzOPfnsWM3qY5qK2DM0HLZUl5VCNHcVn8ICgIUauKvbO6dO88l3mpn0f9IDioy1zT4zVB
1yUTqRt7VG0qnGjhXyhXNgarEJTrb60CoCg34k4oweIUDcQSqOESsIUp/BFlloPZywTEIzQGgv9W
6py3s5Y+kVRn2pz0bPTqV3qx0nLoKWQttHCDnBP8yjiltc0WAphGLPVt9q/NR81qyhcoQzVGALV+
6WeEbL2Bq0Wacypec4lfhqICp2u+Lljc8ev7dB8fkNubLifl0s+BoNYxFR4oLbXpuSIzD64fN4F7
9JtcWZVVvH6SiXvtB+EX6uE/Q2w0FO6+KlNv2oF0X5GrRJnis4BRaYMUknOrILabk0nn49lCe3+j
LxZUvt2TzyUjFjlmegSE9/aZhKL81aaEAvU58ytXKutPGqtSNgrCpb5/KY1HxOJYP5iQJANsoeUj
cIHSClb1/ThuDqDgZEF9d3F6ukKDu7yGuqJvJivfL5NSDLAaf+m9ZtifkJ0SiUOy7o6wUtUnbXsO
/rziVT16KlMxQy56dkrjCn+zgLGR/TnLDaDwTfOigNQnX0Uu7kU3M8ZMXxUVG+dnJs8qfebel1Ny
l4Ip3qEkwKH5Twnh3xrLQVb1aByPUhfcvF1gGNvfrJN1y7DriLHr+mjBbHT89Z08AgjGhtDhEFyx
lHlB2dV0HJuSC/Ro05KcbrpQYu3adqh1zuP5b7i9eCqMcx+C00bFc0kgcawCQDOeyKbJyR4eZ7Om
coLxPFyCYVGrtKKXGIRl7ffIeu6y7R4HIpsc220Zs2ie2QL/1ckveE7M/842u188K8H1GoOSersX
wC5IPeVz0bTRgnoitVx2irOGjjFaPf42836mvvBXf7VlKcMvW4KLZcRxniXYUrkPJZMnr8NoUiHf
xHqHc+tSd3mhNWMQlCjnpIdVD+vn6jocuXMI7+t4maWs3VRc6nPHqt9gcgmXu5cWYwe/PW92tLkd
q6HbkYsfk2q3tB4OfRP6wrzG4xw183ZxCtGSHRfBNBB2CfL6yCir/nOsHEAwvWCx2yhH3duQFI3h
g/aBUmKuoEHlQctC9qsWEPxf4SEIbuEF+fX6dHne70DETnH3oNMoSAkkdSaT9lQ1DkXh+UK/BviJ
lGjf0BOiNas9SL25HQ1C3wGapue+5YXcCwyxB/k1EazN6lg0WzotBgqONEH3FXuHcu3NuajbVi7U
gZIwroe/a2Ycb9aj2ECq4SgPiB+yHmEJmsiGtV8zJaXbjKpks7RnYM9jwwI4qDX0fqLhJtzxd9/s
bOayMoFyiG6TpWZyrbkAHkN0LjeGqF9Xk5FeKs1orA2AWlvafvcjrZSA9m2dS76F1pyD6xPQMVxq
eXXCpp0wzUE+osgXwwsmKBlo6isS5+o+Qe9oVWOZ/WnA/eImHe5+x4+72BxJGZS1ya35+WJRGge+
LeYcFReeYk/DDw9MD6ksmv7I9K6hegdiBgfu3tYS3AYdkqheVVQNHumwfeZmgpLfSNN505hMhYDH
ZanXHd7vM9H05J6XFulZQmLCCl/IjLBkW6eZ6gG2vGExqldT51HqHbT2hzOq7GO5hCyA/tBy6A0P
ND8Vf+RIJfkstuIVAZPDWSlaFQHnnYFmvNtUbwLkPNXHzxx7fs+m4EK4yMdCHXk+oVGXQGQ2bHG7
0xN4aYD+akdej22opvx2noYcO2qwDIlolekbXWD3vnQA7joOOQnirxXYNFU7UCMu89P0XYoGChTp
90mgUolh8S7x+cRss7+kBPcYXgLnqqqy3wr7cjlUtDUgdgwdhlB9q+QSz8TCvZjtt7xPluS9cwT9
FturT1ldZ8Op996i3Z5mSEhUO9eXHOQZxoc54+wVhlqKLfAm2KnXfufj1sPgmC/lSLt5ZouDyKLz
G7PIQvCDdHz1ervUngWUqfaqcIKfSD5PmOxn4xRZcDmC5kGJpvsJ5mbsiKjgExpqDat/2FzlaXx3
e0Ea9E+ZzFV9zg8AKpbFO8LApPc4E8D45z4OVLlRD/KigkdWrlVKtLSrJb8ereKEsuJ5wzvId+pp
6PhjffMeXzUo8tyncKHTosa7RH92E77OEvRUyazCOqcls2tggwJ/L1g4Gv3FO2ULKHN8vZVXfIKd
9OB0Jk//UTdMCpi79trzoX+fk6qvYpRDMqrce5A8idvcx7pWDvgd+J+WcaqGjInD7aatSNYIpYvg
kUA4bJbqwu0WUq8DHyXBJcFsRgogLYrSNHr2y14wgwhQQuSx9WakFZiZ14tWY6VaZCiAdSIPQPH2
SpnX/nOzC23iF0UwXOafn1wqTe9x4gMtWK3i3AzAhX3CVCkhkztv4fe6M8fyCNmUKsVggviF6yme
5b0udQFNCMEmXArnizSwAa/zyTGyG52iQa5gyylQiIuoxMxZBnvrnAqjAYkl/DgevN8Fy0lq7EJB
D+duhUGFz1bk4OoUzsOkDNjPABvjRysvsryE1RT9bm65WjX1H68EkoHrsyA+HcgsgErnM2yKSXcN
f2TGZuWxwCIQbAYSXrUXDITQC/tHzMGEfRChut0yZPqeMKila4Qtwd1IMOYnKNbsOy3rLKT1fe7Q
DR5qOHCFV7dNJr932CfzN4V5GNFGo1gPCaJDA0RneX+JAVlLPjYyZ3x7WKL74oaq9wsfVaaqfSZF
XtIHDKNUu+O16aVIXlW1iNhSIWaOeaMkBkLGWq47AkoG5ObhebuAK5/QQdti+LWu0sn1B0sB71oN
mmKl0L5Dd+TxBFt7SJHvuVDfFRy7k1fqxOHvyi9HgwDO1DVIMKVwUsPztCtnzt+Y3mPbpxRDx1LI
ptKr4HFbbfwytL+RLqsUmdZGZI1mT8rfR+gGT71xyQQGub+DoU8BBKzZ/rMEJ0xW0ZnPk4TFQKkf
Ur41uQXp+1pMseL+9lPv2R/uJRB5F8Xd9JZZgFBhWxOluBkGuL7wUT7jp2/IKTX2v5oqo2e1A95A
6oYXiuO/aQWPAIVRrggkjbmPubnJGnpfMwp9V9ckHwPPF4FHqipwxs574vw0h76ekTQgzl/ntMOp
R1t3v2SzBlNhS9EEpYH5daNRaZbihAb9wfb/8q3pC1BUmF03277TBGS4FMSt933t55cCIXPQeTsb
y7fQIt38B4bKNZEcdOzH8B4g/GYr5C8o8DrLSeCHEtSD6kFE4YKLv21RWJtYE3vU7N0MX7lvkDZd
Y4bAH+9Ezj0SgFP2//wZffan5g/GQJQYFwEJ9/af6gdU1d35H7RCqg324PrsyZbVcB9MfBszyiWC
ts+cd8jDDfKDgSz4ouUbudA0NTAPaZVPqbzOyR6mNA57NOcPEnTjgrkO0qHeggnpHQq9bu/rao1u
Y8bwLFV2Z8Y/ZkQ6PdzFR328BPK/kcDHlcXVO9G4TIpLBj7CEBBr0FbjBGDi/Cw4OC7bKHrsdw0t
SW9d3mU8+ZR0ynAH2kZ0zY0xAgS2BfR9EyoRApdskS+3g2+0NoYk1RikkmToTdtklCqy0BkHCfRJ
xMtNH/iq3nFviiglgSBSjip8PVvDRysPlqIbREdTxvYV9SBRmsA0ICwujtT6TdpldscRKgqTVc7P
01WLGCSYvZr3QgWkYHppaftK37D/vKcFnryD/ukLOAcZhj39v9iHpV95lCKs4BCajnILEVTLtW/s
Xw++FnWpS6iQzsR84hz+NRFvUdj3DWndXv8l4L5+LoxLe19d9mq3APSzByB8Wu2CeuY0m2rtKIQ6
o0AERDQ+gNG9vDEFlnO1tXovsZFDth2sAY6lyAOVvA4h/1iuHAiOYxr+l0nuCSaky670/sjBiZE7
nv3rdT5nGl6A7z7ebwpoBJzlrL/wx6LL/ikPDQAcc+fkfJCP4BijzPd5WQZMdPVv7XJ8BGlEhj/N
W2F0VFZzEbAzsr00HbpC+Gq0UmYB/Qb9+L8JBAwmyPV2cGC0LAmXo6MkyUuWX5GTZyVJwBpt1nQA
OxLR25PeTHeY7yQWEu1KvwNdTp0K9SewmWFMdk4b/U5RCZSeHAxqIEGahHtHOwaeNN/PJE3MtZvt
Ce+cuiQpwqGSYzSIwLF84jdKx84kyFdYXFENBfllPLZsKF3hgem+YmWVa8nGARUNjyU+LjXXwLGV
Aae+Din7piP7ZR+nPtRbfETbXP10AoiNizIL2DSLUKhTZMlhC0AxEGvJS03mbVcZMp2oe9ERVmUd
eohTdBvzPPRRwrF/+txw2IMyhbUkm0dEve7rwopYAAo8Dbc1m5t2Ea7OYmY6MjAbrEl1AM/m89yV
cUrOnb2ufLD1ri3dFJsSKOhtH7CbvMujrr6alwhfKy0xW9dsOdded/fE2yikH/5INZb+enEwgRUL
B4N4C/tkpqHCi8D+3baTUxVNyHgDSKHtX9HKfgskxP7T1Yh6RZI759pCB7snKxBK0tbCTjXoyar2
tQFSXneodA22gNQAZ1aA68dEliVYCcfuzIMu4bSB8O57J1DPkkVw9DYHPoBUY/CgxHf7+smxhLuL
Vm8I8W+bqI+8yiprEag0Z+No63RZmKDS2wrULcnXrTnaqKQ7dUJehigYG2VgjkqMgFff4Hm4KugQ
2w/OLHel4+wkENiJUvJ6wvueJEXAsbJdp4bGylRsGBnqeXRlK5VzO+8vaA587h7TwTot/C65sRWu
CquJ0UV7RPExEFl831lrZZtO2cBTQMc1QmcTH19qjE/MjFe+slzmbNro6zzgb7ge8zskuN5CpYET
WdQslVywkDbKvlXLCvWFV81BJ9eAgm3QbK5kJlBgPoJj3/tKk/G/M85cHJzZdqqfnlfFsIOYS0U+
BX674BG4vUJiujXs9mzuC7qlbajEpzB8kW1EIwOmc8CPh8CsrPP33Vt6U2wMqQitMzAVIDmkhYD3
65TquX5LjjTRdUjplav0R1+v7gjW+nrT5g2gP6BxN3kbjuJTjBGGPectqEPHEGXZkqEEGDm7eara
Hb8PdfYeQLfseEHDL1UmfiJYCYW4i3xDdrXKbVd/7oGKaYLWNZSY2j72Ao0lcFHZOgzeqCE/fYwP
H8+jwTyP3k8MVzQ2T6GET7gW9Je0G1HptvstteLe7Ylc1QEY0MteoHpf+T15Cc+2VuP91pca5WHD
U7EH+OG9g7S6JZoErf/vD3vh4YAtC2KIlT1HMIoooVkQdx5PvNto4d+9Q9FCfwSm8je4bhG++BLx
lgStyamhU2wb4W2kq7nIa+UyAoEYe4g1o/pO1DqUo0ofSAL9EQ77Eilbud23WtR5NROUZ0pc/u/x
YrFVzPkbFwE+XKLZTCTffReb4xcHHSQL7xeClA3Nrz0RNcw/UGMHaAFTVJCvdTPBQviTcXEb2HgL
JSyI/HVjvWDK4yOcx0RrjC54aNJAKHseyh3HEQMIR+XkASBFnDR7VkZhK+JnP06p7NeABM0vpIy/
4PWzWqeELbXpTzBs2Tf5xfBJ4FgDyHg6cilG6x4B9JJ0vzv0rNlfzhARrMJYgG1C0oU5ir3NsluI
D5LbfTZb2A4MErAXO6Oj5Vd0lwy2VM9zZV4BUVdrAmUGKednoOAC7e/lroeMsB90uswz/y1Do/OQ
AEvXNNzZLuksz7lowNd37tNFja27dq8zqwL0NjBK0FELiK06f79mipKMpXW2F1u5wYfn0eovOZqM
PP1CcR0xv2jOgZb2+EqR9u9hFzf5317eLT1W+6BnrHb4uiYHMeLvhZqIMz054JtBdcb/7hHut6lo
3yB7JtMfIdEnc+DjyBwnWGT0nG4ULO/G+pYekzmT8c3I9YU3Mjl9oJPq5QYQK4yaPL8ornFvDnS8
EYCISFYlCoAHgBqPdUswAA7OvA68DPV1c+sVt4W6TdTtGkSKCm7R7YRTO7cd6LZpFlfysAOiYEbl
najp904VcHx+lyJJaa0r5jzayBs/L0+Dn1hGWoQ85DT89WePmVtzbWRsnZ6dUz7dX2Fp3MtS9z3Y
4ssvXMWEYnWRGcDaEwFawYWwudS6oYgmoV4P/0dAkpoblSr0B2dIpWC/3k0gFOxncBvarE9zBAmp
FNNy4s3DscyYalTzTLdZfbPItKpPYZ2/cAHW6BzLtOh7a3btN7WwKwjbGqsZtkzae2p5+qWIDann
T6swHrW9Of/vbzRulMKCCDz6VHYO4zuwvCRbUQCRsof+0A4YC1j0HkuJbV5tOZ4nenAf3cHc3FVX
Npo1BtFPaak2DzH6Oam4+gZy4+IY9q6jrvm8dSVgvBmb4srAKXAul90P3U7OIQ2hGPSvTHGvv6MK
XCS8bEx0B1guY/WNOx2dk0N4bQlPV7hYOAOrANvOLs29GweY5NSmgMapALgyAHrWWwfaSKLf1Gw5
CcXqsqNPV4uGQTj/EEfEis4kAPTiQK15mnDkMtjdU44sBAZJMDVoYBAgf3NUxi5QZHH4OGwdGGyP
jm9nEgFZsJxnDqsmaECbcf4F0CmevZz3dgGyOpkFi0iq7HG/eMS7eZ1xM/qJTSJQdQbxvIedbZ2+
bUr3CNXq8h9A3KZkkfLRV3QWB04jvOY5mTDx/2YjM3Z/gCOt5skKVXbsksWIphjykWEuFf6PzxjR
lPfd0fqsJAQYgFGeQZXUS/CKyWxufVDXxNocEklS0vUqmjxt3/USLSlF2Kl85ZklQ/XFQhURiQDt
ka6WwXpkD0e7Y7ugnuQ+W5FPERZG4+5T6B6XTp+oSuEqy4axYASX9WGJx0GsILVCgDC8KTrl5a+L
eL3o2m8y7W6CJgsnT6Q5ABDRRsI7G9/JGPX0ZGfEx5juLqQcGw3erZbzdRL55HvVrRhDEuRisi/U
q2t2CFvoizvSP5wTaVVYkLOy1j6CRsbLY7cWjXypLHtIgg1canUjXVrzRyBe8WAe6fvdig0r68X2
z1B+qno2M72ddg3HVaeSYI6PqZDSJ7KWjlVzdIVD6WKYc6zwtVuzkaOS/9ssxMnLm7QxWk4ikKPH
NN3Ww4BKMhstHZEpNgJlwNeSV37/db8pmpAcnpZtmFdf1izrmH7UMpmMWmmHWL8YAO1mWrk1Prbe
y9N3ZpI9oDVA57g9PDsJNMT2EqVejGgji09ZYWYBNW3ducPEsxypv0Vw0BzIkL2SO9M2n7AxOBfw
Dyx9XcQcJ3Ety/tgfzq13vRVo831nmXlX3FDS7zk2kG530HFrbUtDsbZYoKkhOeTXZYy55fecD7q
OPTBiEWHX4SZ4su0ThP11KmysiaK7IfttZk7LLM4Zk3kwOk1/zdkeDuZT8IuLAdgC0vJLPmsY0hc
b0A5+b+7TW9EORQHogEjkKZrH6q6YLErj83kxSg8ql1XXQ5K/+eMcr40VxTm8tqW8NzsjcFJ1r9+
8nQkFqtBIgAUuAK3AV6LXIJcLWIptKxbh0EjYeO0QLaywTDpLdlkup612zAGdVSjnF4YXJH/iRfa
3pMT8jRuLMP321lMfm97I/600g7p0iSotjOXJH6IrLw6QAGmSj8XSsdjT4IuqMKzhnet7A5K6TVp
dm1egrlnbhyE+oyZBKbzFd0w0asFOZVvyd8OGUlBGyrGvQCHnN6AGPxw4bOqtXi62bF5OMmPFnMP
Bdy0LWRdyTK6QrVEE+kj3AubUPsuqXpmF4hbx+CAdzEwXkAD5l/WUXKds4EkBRCwLgZf67d3MHUH
4vnyKhpX2Lul9s/s5yNANkcpzsjJnymsVHxK4E3CUFLFa2Z7D2klPIda2+cVB1xvUUJ9JF92GsId
eNkwf1lLl6xqddt2sAMfFPVSikvOhujXcyMx3FSBqmWPHfvCQDR6u2InTQAlCU2dgZNsW5LLRiaw
InYiiVk2t1sgTtWhQNFYqdeFTjgTjZIYueONNN68H9DSQ92z8SFMo1AT+7LFbxKFr22qrUefOIxQ
uhCgHVoQyBn4UeEftVNlUkhOGTuc8Rg4e+qsQ+TmGzu1jHmwG6VN/T4hVTPqiYDyDHxjXWuiPfPH
8uoxFov07gK16O3i3veen9MDKMgxBKw6uwDro10XqXKD0zpJt4bNjyiVapRG7y5kHnpcvAT9rqTy
J5H1boOYOIcrj2xN+X+GJ53eA0eeW9M9/CsxfKF+eTscRWzIeZ/VfK3U/JYmCqvvHra49tMWVYmX
wZi8hbQqLcVJ0zLGQgWqo39kwGRR8PChYXeO6CnenfDqvAw5nTo/XE6PKN/HbuueLhngQaAxfrPG
Vvx0nID92UxJ06BKGeGmOuom6nJphndhb2JYnwNk6CstOMNeXMQlh/KCR6DyMvVe9bsiIFVz2hoC
8iSfVRYsEmhiifCrN+5LeTEyMXcJjg/9UiisOF4599bchcax6I9JpqPE9WDMJKbKs9PXmPLk7i8N
4Wd08VoufseMP/PiaBBFV+eTUqMoQT3EBsAYPO0/N6QgBAevcVWSz0cfPb3H+Fv68sZ8PlCuv8xQ
/riIOUVV3whAPtesxDySFbZVQUhgCcdm3keAn0GCYJwLUQI4ELg9x52ZKqpwaVFWBDRm/LKP8bsd
QxI/rXlhbZkdR4I53yXUUDIoAf2yKSRDdmwrCF1D0YRHcEuWXv1lrrocJ1Fk/0HqDYu9jbgEYXv+
9jS+N2j+1jWyjBRMBR+QPMDvs/03HUEsRsQNsBcDAQoIJ9zh7Y8eUPtQZGinAcalBPsKeO3dYtwK
Ky2V4qBm+Lz4w9xj8D6SLhk8XzVHr00viSmriGaOQWTtW+unJpCe/Kjk396JsQ76MX+AQwMrs5r3
NS4t6/SL3OsgTl5hcck2ll/qTlgbOzfaAuMHPHfRzjBXf2TLSiWguatmObm3YgkZcMnp+xe20lnu
J3iu54ZethmhtW0Fcgsl6TgCpEscfEhYrxBCgyWJoy0E4EBK8CPpUK1tyKV9u+1nTzkOhsuO0awK
onn+BGIIh9YVQgj8q8I4saFWmP457hwmJ0BwQZOHdgr80plyEyA0WZrhW9XTpFuj6ik2hG0dnBkQ
vA2Vhd9LIFI9dTwf4Ub/Kx25yXTs+SoFEn9wGkRaHOE3hfLUIGWDnpvAZeTGY0pa6vL2j6cebN0r
hEGvhBQoj7jdJKcBsg9MaQE9gUPpGIhEIP3jLhQQPZ6TBJ9rEScXISCDM+X/ZU5xJXB+PgJZ7bCM
kfypsZrsfP6NIt6fFneI+1t13ecmApYLFgWZFMm5DHRcYsUf0PaXHe1EOXAztctPL1qdPPkOa7OP
U40uiktg0hO6b1dWfov8xIg3hgFiTcMkh+wlyJJfpPOGEHBVdorhxPaa+JRXct3EBx/r/cLvA1Di
er5Ff/M4duGJh3jG1pPdYHqJL+l7A9jY7RXzQ3HSI31kER+1NiRUd0BR0gd7i6XHlOd+AVUt01Zj
6yZsOtZQSgUu8Ec+RV0xtxe3e+VdMZabymvS02/9Rb4KtdYyBpgqWhhCyWN7pWyeDF1gvaRLuilX
iGhBZbADsTZHuFlqslOBWkINPr8cO7GOtA5GU64BIlw7zYrU0RLHJzI6tiqfOETtGhG37+BqwkX7
7W9kvFyA3exe1YiM8Sx1ASq6nBtoX6mbl5Uw3pAhIdgp0lEuZjHikuz6uH6BGKrCDp8nmO5YMvjg
R0kSXK8Rnf0EMvPxYJurtS+NnjvggRtBO/8ulJbe8dJwVgZS6oxJkkXqJGLOaX1Wud1Kf2b93efl
4h5SIEzi63lQtegbZyNm3qAFLSCi7Gd5kL6haMcHE1uqqRiVxB2P0KyqvGcl/kN/12h5b9l0LSNI
pgXh2jxLXPvyZ49m+pRJZ7VZUKA2PcH3CNIF2ygIBV9rXTzu/Fk8ATaU8rC3RupZIEEh1iehnnrW
3WLNHAL+9FQlKKdWSRbHfMZ74AcU79httOf/L8pRBp/J9/MNir65yyEsN8VW5T7M4Jj4feUR94sG
bVeXk4sSXf7l2wQcmT+ZWKXL7bYDtXQdw9pv2xm3cZ02jdXRHxeJRPvL2dupWv9E7ka5HtTNT/HH
JSrRzIhZw77vlToZCYdr1PwlHkKcL2Kes1hDxMDOjNXML0M/tOTfvMz1p1tHF/sOF1hWK347DTds
a3yj0INF89oGXrqzs6EtDsNWnllD83f2Nf9ceP9vSc22hyIOz3lp4fvgP88mdeUDM6NIP3n56d7n
LP6wWaDCqk6LIeSeVFyLai8cZPQ9uCdM9dpNqbeg8VM+2YyteREnOoUz+wqzSeuRu5AnRB9ZHJYd
yrj58HwbyJjG01GckpkzOuwmU3nf7RfR+/bbOjuzSHJz57kFgcxK2YU/Y9W8EpE1AX/eDI9wAeBx
vxYI4PVjnX9o8R/XxWEbZnsjWYk+17BMod08f8TpOudmXfBJmXHRLJaWmzm1m5nk9B9HEYpjY6Ai
BOVuMDUbCLp9WnWvf2CnNQLmLgcBgLdkd+h0DcnngblbY+kFcMkTPOMUUZvD1zuB7m7F8S9o5Jjy
pEjXGWlMaGtxXVo0lN+5fhJaFO3p3MPW8ytjTEaRu51QjhRtDkcJlq14Cx4KkIM8Vi0W3RYAQKgo
a248m9asj3132IxHYlx8dNZ/Zo4eV3RoCjeY8E13x8Ihe+rXtbimRPF63kPvHHzJ3BILsBTVDtK1
YEs4aEgqUCBxm0hZdrxTDtFB4Rj1UDgMhrgXjAY3MSxEZVr93JDxT5cq8wiDlWy+dMVJl+volMTC
ysWL5GqVWuKpey7JGiBwn3osbsUTRIgazSvM2lt4skiu6L7ooHhK8xZxXe5bInqwuK21H3Gp+ink
Ip3JqNJlUYSOCPsXsp6sTwb5HPqTC7tc6IJnsEqwvZBNC2Bp2KUagmvqu39AYHkdhwTFO4jnC12r
e2Z+YceU3poCHCd5I2cLb4ILCw1eRMBBxb3HFoI9Oyoh5H8ra69gIvhTTqJBZujE0EpSmBafhxGF
Oa16e/f5ZpgG8vCVtUt6zV88wPnM5wrrrMkEHOm8gA+ZheZXZFky/cwkBh9zgnQA4+v1Mswq/klp
PNopm7EdKGc9MdALHYmgNZywaZ/V8VvSSWQ8GY1NrXB2zThErfewYkgaTLM8ipYAb6/l75/oefZ2
n8RNmoPY14hyAaMlXd+dl+Q5QGqtytO3K54StcDIZpIojW9j6rb+R1zYGr7JhGgpysZ1q3pYeyFS
iSb87NEU0yS5eTHrEXcDupIqXHyllQmsbil+TOljjHhidoqAVwtk/dSdInzGzMoSvhkH2etlmFuW
RFluOurCd5r7XzKkFl3ZAmdIrOOQHAAPMwdOL7DLtPIuweTIlpKzcHqCPjLP4bsB62BM45eTpW0z
uNxcZCefB9f6TeDW2TflNdBBr/CSE1zmaZTL8CanpMnaooArNVTe6QSlpIZHtZfl3wtfUUaP37jm
pY6IoAXSdOjG6h5w0iczjNGiBOhN5w4Iih2CjzKAw4wHFGJLfaa4s684XVE8/jDW4lU5JDaI0KwO
EQhyW2VODUJyWOG3Xlt+GtzrynBq9oj0PAvzAdD6y4ygLwoZ6ZU597UkXx6I4PLL15zJd4UyigUi
s7KhgPCoBJRo5ddyDIFdakkEZq9N/imWn4KqH4JoDLzVhKyT5GHyBIZh2Fql4ZiVPtkW7i0vSIAS
fYh+DTfAaVEhXjTyrdYKlaE61rM2BNPT930JuM+x4ycMWGQMEtKuZ8a9G2N17YJ8rRu8LPLaSHYA
4t8QK89iJwdN28/QNg9SdTlnG2W0nfDsO4Bj0Qia+2fNRemOin6skAp5mMtkau5l1rDzWiwBtJFA
Vy2f/l3Qy7dPf8J+gfK61N2RIxjuPT4UoU5c5qvz9dHgBcqH6DsY/pS7UZQDO52XtcjRP6c+HwBs
7gFKwhg2kOsUTKZV2gmYI2K29MdDw/WndSnnMDUXbv4UFTLd3UO/dGH0IP4PujI5c8tW/Fx4BJJG
xfUQ51DuiX048WaUcIDDABdR2NXRKO/05A8KCj6zqreJI53bQ2a+nVEBnPsx0op46dsmmYEmDAHx
fQMnjP6X6iWBgGJuJrZx1EKlh7AmSnKBQuQXxT5WMKqbSJdgmUN/y+JZgjKR04S9rWlYyzW5sZQb
0g4cvhmxhYv6/xXUpnC3x8S6tJqbLvfVPMRMHMWbsQ+VADBwsG7w978uUy3rv7pJM/zZQP5CyT5h
xiiuc4EcK87B9HQDpEmHSr8aNdFm/ZvnZFuR7SRjeB1g55lD3VV9HMiiPF3ewYELG2RKML/6jIZA
u+Hic0sJbJDo0wGxQ7eo65C/b5A+cGYYW+OGkE0P2B2c5U/gAVbFNSwbC8PSXGzPgrYP0tI8K0ck
Zd6vkrD2XUV8S3hxt/dio+2TCKtwV4gTAiYP8oMFE3Jt1Fppfc6w6ZmdG6LE9AfmSZzPMXITurmj
dRdp8qf8W0/PoO8CWZo0gXXQvu0LZPCMFTRNE7DKorEXyj8aiTbq+A676lEuvPDhUDyvh2zUkQZF
CTjkTlUWQf6Ob6aErRR4n0vD97jx3cYoMvP/sE54sh/vRb4V7d67i0gUl+ebpBHuiqObBJpr4hVw
kydjS0pY4BLLgCIjs6cal0CDYmfqckOBQ20KzYP9mF1Dv7TX9Byd0tRr3umzSe1M/ApJ5+VwABjf
nRGbHXl/xa+egddVharQQM1kYMp1KLkyFhxx2p6QFNwOvgTc0BFN1eODNBXploZaAiWN6lv310BN
nOsunQMxRWdf2Czs00Y2lkXyjeeZ1vC4BQSSsH8T3mM6GNU75OBcnZb9gzQyPuR8COTY0ta24iw+
1n3FuC0qyuOFLP2Xxln7ZBmke8+bwtEQgXh1gFY0gsMSqbq6anTGceHycmsM0eWr76tb7so4BfDO
Iti9ksv69ofD2haVIK25oE0ddpgIC9gVg1ApKouD9ckUpi9mzZn16j3BxJWujVqkzmhcKxzsmN6U
hQgAseJvL1hNmx59jRmdUe46quDXvBB+U3QpMcQB2HYxrSy2SMhyTynEnOm8LICsmjUHedpYfdxK
/dbONqyG9VPKXrSphXupK2yIhQnqofSF/d4IXrPmxzFmj8p7zU5HQEPKzV5MwIAWQ/nr3GWIC3B2
XeKStPwmrnn90bK7rMUNXQ+EhsNlpqlC036Ic3P+X5xrp0MDjz6P61H35Gt1JKXIUhDOCzNnFTW2
/USIE2QpeGZH+MT7bUAm3G5T9ooUj6mi33BC6kp5v6xaW6kE4OH8JYJ5C/sSkmJZGiNrHjkdu6bA
1CAq7s+m7YkZi7kKjnV52vKLfCnwF5sBbJ6Mskc/qRnAccLMWC9hBE4MbfwXoIIMyXspB4wVjxZq
+fC0FAUO0ISilgjiJ1RNsCWbYuebKmu1nOwH3x2BNBBgfLtXiNfiflskcRR/pmdLO2wJkm5FPnZi
LlvsV3PY1rCJOoDaGbOJgoTFPveHskykN4EglBf0wlNA8GdvrNDiBUp9vXCEamAxFWLaDxMrVy7p
c8qVI+VxhmoBXKxGHG2zokRHyxZKlMBreKrLNoOChPgISvKqrxq/xfPayhATdavm0OqrIdpkaU1v
1YmkDy5h83S2IX8nL79woq1pGE3ph8My6qi4hW2RO2VZeXxoQjeNVKPuUPQp4lfY1Bk3JTx3VkIC
fO/u5o/6qm91TMLm2W79rA5Eu1jvwnkZ1dDbqX4ORBjauIhEZauEcUpUcFoyNzrqRlZr+UQytqPQ
RerKITqqxba81AqHYgbs+vmqy7B4FtBIo/nhATQO3kpAM+aewXyQn9fRruiR+qmxcaQKG8jQ62w8
5gpZQxKHSULHziWT3WwWDeIXGnDqXtnLNW6jAaDXKWEIYu7pLt9oDnw/xsfC4OWK3NKUZ7aBOVJ9
7LBmzTEOcpxENzFLdvoDs9HistngQIctc11ZPRUJljJlFCzVCa6lEMhqjj21/a5VcvHJ+QJ35x48
qTgQEYknJlqF6HOW405X/J3tfTIR+YWDfUjbwGBD5zLnGHpS6hv1xdcQqXZCMEZae6mDAzHYLJbE
wT2p5Qis/eBHM9nFZKfwdCHHFCMUZJeD3PESP3lQocaHjmIYhbU3Uhv+cthaGJuAmuqT1+eharty
GPiYIbFi7yzDIDM0jpjomW2dGrDSarhiNFxXSQOkmn9B2Yc0cgTEuJ544FG7ELPZZBTAP4AOqNGI
Al/gg2o1nTcp/OSEATAFOvGgJOnKTfdYz2aLzHS/Ib1lJqZNyMMUW5cRCw4TGP6cG7yvCQRygl/5
moIq9zJ/p5kRaPcbDdq611QoMVcrFlaRjW9ckqnwiz1/ShnQ2YUBvGtIxHVKc0k0e4wVCyvcVG6s
1zIIiTEBr+rFZGsYtv8CAvX1dyS8fhRymTcGhEjmrO2IZlIGW4UEJ8v/Qx+cm325y/lyVQxdyGld
itDFNyJIB/wbRBGmEHUJpYUmx0xV2aCxSmLzD0PzTVEBJ71wzRcuUK1abF+gdIAUigmKCX14RZmO
+Dp/tGhf/YzVkaaEevXTcqowG2haMNLAXaQCmrWYrlLkCQreSPVhDrTtRnMAKRkfBhjpDYDmytJe
fSNO06JnDJtds/ZH/EW8+quZ9bWoh2Xb4Sf3lTBRaa8UzONcn8VsDsSAwiKuXaTFhvzq29TbsmKs
464g5xsCIGhIUyPp/1aKzsskeKYVVmsvhZVpXmtIzsgdQlJw5MKXcR/x7kjqnW70X7mM+4Mvba9O
eNarHo14mEuPQrChDQ9msdMlcdY3sW2IEWfPeqbWIQF7jMd0vQ7x4ACLjZmOu6e0QfMvr/xgD6eN
cvJ8Hxv7wqcbrQ2kN3WkArNhzYD2zRYOSq6wx3oJ12XaHgEbhoeqCtUeUMTUaZGBNIaH4lkH9cWI
HsslenpcRKF1MVjY79TIfTnPDSMuIYjEuU0Hram+qDZfWCAJOofQjPb3xbOqjUhkPOVhereBQEUD
GxzUyVQsn1V1l3ZP/216sSCb6XxvN4TlZRohyZAeJL61voPu3usU9xA0IFslokJshFLNrfu4OQg3
V5bvaTY6nLJCPwKW3Wf+XwBicvA0mvXvU1jPZ5s7fXIqJ1Wsua2g0zJpJpLHuFq8I0VDZxwIVPZk
Q6wMCawgewYzaC249CrwBRAh0yF4SR1zr+Q7O55YX/nKb2RBrGVCDQujSavVuocmqLWMdv/KvKaH
kecteea4GwcvZGCC8js+bp+ksT6PMMTlUV8sSr9qjyDDOTQAbiQLtRqndp0x6L+YrdV5K2LUcIwL
pi/ssqn6R2PVorJBh2JQaVOAeki58Xh4kRhvJbCQPRn7yI7eimkO6EAMYfVvo6Mu6x+k2pMks5D/
rNb3pkNwuutSdC7aUiVdS5cAjYIOytN+LWpJVcskcXO+RN0C4TiWVyEFP7AKH90+7LPePGKHvIdB
CPzuMuOiQ1rfnLxg/W6HMcDTEMCuRcTDSL7w2Bs9yNvGJB2ee/vCoKp93ZcPUFWCdr2q3cUcQ/Sb
Uykfon6BJpZFIMW6+D8r3asb+qWVeMGw2iRTKFDP614vi/TIrCmG/SRdC3LThmk1CHiNNnR5Q58H
Mv1rmHx5M1RGdVl3be3y96ZcOLtl3/cuDe8KwL5trb6YeerBvCfH4QoiwvMar+YAngK8IhLnVCeW
EG+XPw83rE5H5K+TbCNV16/XMQm5CoiJUEqlHD3Mv6OG1lXdBxJ+24p29KsqpMw+4XYaFxkUn1D8
HL8V7FW5ETE+vaHR071ILy7kxGQfM4dfSui8ZGfbHo87GkF4XqiMH75bvhPZ5OmuhKUSFM6/HUyb
PDpE7VDbx8d9uZRQ73MMwV+hH/3TIaCHCz0U/pey0SM80bYvW+YooqOQBOTFK2A6DMdRTTyfQpcY
nVteB7jJSmfuTHQPmBx11BRfXLycB4YkbcTCHYpUZ+gAFWMQ8XUJq/iy/NYLT3wPearZkOJZmRxF
6nrGrvYTKvohJ21Blm4rTgIYqeT+cAnfVJ1HBD9RI/BaOKFaGVqq05nWReFEl79To+WmfRtPoRwH
fXzVX+IvUyey85mrrWxrG4ObcIaxh1KwffGiwqlHvx3XEcDqSP2aFvoqEKMc6sy94IXjQutwt/8/
w3yO7dsK7uMoapBtfFzUIINiNMD7Rlwf2DrQyjIgBkmSXf0Ik48YIHQskdU91gkv4qOCCw2iPZM2
pjjPQ2yXQYBvmQ4u5iZ/urNOeUL4oBpRacuEtTXTCfnxMkRYlOEteVWBtTCnhYQ3TtRbDMuUaKTP
z+IzHeXUENhYatfe8CpPVjXjVD5bcPQRZpdMT30X19+LoiSmQDWFKIDwGfz5UwlL5iNqK1qStbxW
hmg/AuNcryf6yXVZ/jk3+0upoV3YDi8XysrDTUkrZ6Ex1vu/w9zomDofgoXbwSkVCkrSseoXG3sE
WvXXBrL9PhSQDp9sB1Uo1caOtWNySHdX9qiXmG8uVjuhDNvRWv/DzotjJYJkuHctNiukxt1FgSon
XAfz0o80ww21RWUY8Zyi+qUFgKH2LkcHti2ELtRDDTpy2vo67VTfIStBedveaOQqs8u8AFM5+3fx
XelEc7auBA3xGGGdmGGXpXPAI+VTf82/r4TrjbsThcIBOMFnJ4Jo7GC3oocCLCUjMeyR9aKkTRUZ
RkCNumb8jUfTIjt03hF28OSYQKDofL8cNKLJ6oNmb+RpbPzBukL6cecTjhSGkT7+0zsDS9+JpbtT
gNngzdpxn575LKczYOpZATF3rXtmH53ji+lRt0mCYQFTcxE3ejPCqLx1rbhhW/cvLHqSZGbJDoOK
/eoUm1rW4E041MdAoIK0+1yiLdfKkT26wpZTOfe+YPAiKLQeU2EAoJmuwRbfDRi43Rr8DjmUVyUr
nF6lEzZk9VDRhusTNMHuIw/QvL9L5sq1jwU058QsYY1HCuUX0D47IrbIlapMS4D0OPj8eJwK+zl2
G9NA1H28vReKPmEyJJa9CIGPgHFvy4LTw9oOkdvJdGcTE5nnOIsFzmKnCk9eUp6F/CRhketeA310
vBTm6MP/eGDMwJnZQIHrXNfLay0BCKiUzIDBt5zQ0mrYBWtsMoceYlyQn682jXToDzuF5ZiDLyH3
LTRBH9kmrJ3bEYIAxAQt6uKH37SUMuR+Sp3piMg8e50BF+RAii+iCADy9iVA0QRLr9Y8gnESL0mN
s+N/aTnpuY1ADHdHmNk4Wt5DMINMCgBFM6nqLdIbLXkxhP8zeftdO6qhKMBYgdhxj7YcNCEvlHRL
aTc1dT5vNE2lBS0SHfu5bFH89QKCu7u2MIIrailFMBjA9EaKtQ7OUXNs1FsVW2TutjAdoFnKWOOL
zDtN1c2HvP94XDhgEE8XHCJ6fLad3SCgHDxyB6RO4dOF2c/+j70Squa4QceMCalkvqrchK0pUNLH
TCk4hRjMZu91jOSU/e5T/NTmYTTY73IiztdkyBxWua0BGlpFxrRdgHHL3EEF7KPE7PVBokuMXn+i
fHIPH1Tq5uwG6IPo3Ft5AnO314fvmUWen8EeX0dabuYJ/AFN9mEMdp94PLs7Tlkz+OS65ssoYjvz
eq3M3D7rb0wZXUW6E3Na/0IFd0pMY5e+W53tnliT1JEnrEsj2DnBtcU0OjJ0giDwutb2+Sx0P3F0
fjOhZ/gjXjBO5yERED81RRpTx+d7N1vQhHMiF8pEVJeUIOBmgWnQR08SbSBStsV2QlcY/9R08u1J
6xO84ls+35L2D/j3ZWKvVUzJ9LghBF+PLTLsf7/UGV4tnzRxwNZ21/zsD/l+zQgrQJIAUxg2kbWn
MkmWzJZCsfSIfEex5+6uHy7H0Jjd6p6Bw6EOZJ0g6wDN14o2b36i+USp9Nt8lh/aVAE1v9CFCl0A
cVx8JbWMSmMhASQMyg8uB6AwuX/l24jk73OQ7r9JB7LkuPJTUVVFAQUfvVHYHuRsBG65q7zLehlz
wuZkRgOU84aCQHrld6B3eLN+kcI/fNUqNWGomaCbcrdumNrr7SB3riD6Gp2o/9VCmX2LR7LiO1pp
GNkNpip72yYNxa+Hw0v5WITx4V+QN6eWoVC4fMg5hhT14iM0PaEujqvJUcgyilP3mRYb4ZgYu3Zl
2tlce2/B42ZHRadAHm00zLSKSXfUylOFAPwTe45ujDdPQi74cDKouulpuNpoFQC7RmPf/pTiITv6
aocHXOLAghra3Hl2Q+VDH+OHmmoij3saPeZ51j1TZN53HxJ6/apVYaSxoLmja0SdmbaVusmLCe1h
y4keO4neuZl4rSv8VlNgxlN2vMN6orGPMB6zJMpYOk6TV+yKEDLwUhe9dK8T3qPFswOfs04TvsEx
TIkqAiT7JcmnG3MxZ9g9sFx3unLml24E2cNE/FfcFSd64ARGiZxftFrk4dGVvLe4FIFU1TYsOugG
8x9aVbidoIOqPPx9c8YTue5zf3Ls6wzd9XwdUkhhX7A4za8zAUeEiVgNuJwuD5mJbWK2Lpx5ezt7
c4lVDbp1B+u9jQ/34rMCJBXM9NyT/mku9tunbNa9bOvAROMbsgjXy6ZOfcGQa2v569+oYojfkMP3
nMnaC7JeITXQTBnMd2PWvONiVNCuvpOR3TcfSaODTDs6uVtuxbt2uVvr1RIQsruMYYQe6RIKRoGv
xnvTHd0CB5SlmhZdlaLoSxPuWInHbBMwM0ebpjIOIOfg2JEjzpV8OP97fYmPwLdunPLofQpxGbMk
F5P2eGb//NGry9aMeKuM3751fOrySwFEJ0HFeQB/PMEc0z5lS8Z7YyZunJTiJNrLvMJUJIB9Mw2e
1mE1+82r3ydB72bx7O2S+zKxzRpojMUx0YnHbdZAWIdnzVSPR7DS19fA/ST44ymsBGmUcZh5whEZ
mi6e29Gm1XpIuisuPp1YaaqO7/zjGcAuT4Nwokqy2CYEoAkK534ACvkT7tAJtoJsVwU18cn7u9aa
X8S7jYn63GaIcgweNiPxIYNzgNCk31Mf0G6b2pFUM8LB6Xfk3ekSXBf5u46XC3+bgfLv+V6bd4ba
5C9bT5dvLQ0epWTMLtgjKRCJfhN19YwxmBg7k8Ialw8p8A9ZcTOLN9OLiyQaG7KEZVTkX6Gqax5P
zwuSQ/+kmjvCnp6CIRUzLOH15vyk+ypR/Yjm1OX4V9EAyMLZEiplQ1JeaFaoqyqJ+lcCyG1/IwXU
XfNbrTowFwSkKoUoRHxjGAy+j3H9WSADghBCGTN9Vtni38Qiq9wIVDg64uOnh7MDpSu6P9iREkAU
0YQRhi5VEhWReU6ZAOsZ4uJBTCtaNkKhuPNA9x8LfvFQhJNJISdHV5f756GqZ5Gx/N2ruNimY2jr
zUuz5t7W9KhjSgE66iXXYV0XN1W+44gRLsQjN86snGpaYwcfGYTuvCaaJwJ/MwNw4nzPj9nm/L7H
/T8YcEqM+22VwK2xNS+peqAnQVRxwA9fq2OFAiSN9pMj23atiexaBEFJ+D1Af6hGz/zE8ln4bQTS
VKT4yWBByIRrW9bpLu9So6Cx96OXA0C24s1DrP7m7tM3iEgZ69JUbElZPdOG0+XpHpiImiJ4RifI
v23WjlLWHnwWsYeTf9BRXbQAj5q+d4W355M8Y32KF9sDWD87wx19s/3UO27SSCwf+Rxk2vogzOtG
VsYvY93R4YKZqG+UilNJpulQBTE1qInrPlyjWPVvw7046yQ/hA7RmHoD3rvogkXfA7gOJ4HHJxR8
cJzitqq6D7IC6eu23ju/b1nD0/Hl31N005l0jSYk/tZfngf2toooYdKDXEvSy1/YNzIh5nqVk4nN
A4zDiZ9PGnsqKu4wktoqf5ZTd8T89TryUGNq/lS7VHlWhZ/+NkCbEPPUgrolexqAZnqK02a5yOfd
x89+Nci4/eMCH0iDMlWccasNgBoXc3V3l4iYstAoE+qKdnCWmUnbEGzYcy9QbESXKqcOEyFG9cLS
B2ayVeHLD3mhRwlmWhJYT2YROIo5Fz3R7U2Kw9reFpA5tEOOblLsBrw07a4OBDLjV7KRuzWgoSx2
tzElxilud/fe79AmE2gy96364mL7ulcuWfngocmbNbvAniieKcLqr1LPdcdGOl3cilX/AyW37Nah
5J9iS7LJLYABwmrq1hbJayVN8zTjavmd55khVFiUE6To5kvDMfUba5EnQLIXSOwbKHbXL3oLdw3B
z1g5xlIDJqmh4HESOZUL68q9JpJHDwNhHWn0RwdN6RipRLcWuuv/m9n77Eh0CsZf6QC1gche/daJ
U3ZUWP4/3oIxH4l2I1BHgoPZOqdk80PLdzaE5pgvjGP5OeMf9eOTY/LAXP1ICfNYyzQd85DxNdPL
naVleSUQW2nwTJkcbFoi8y/YzIrwypD8Y4+SYslAqX/9I2d+hxXRnjMQwPoevUW4XS3XFUCz93Eg
nNlT2z4cImBUIbMAPzptobW+URTx9IajXFRbus5t+UKVh/6NRT/jKhcV1lD4pULN0BtMCDTPFDr+
s3eAtsGfeZO59sCKjPjGUyPYNZdvA/y4lAonrpkl3tBVHgkgugEF+jfpavyjbfAzbxrOr+yh89De
fOGWk3EzSM2H1UyLDm9iQrSLAv9KsEiwJexXeRuieSuZMX2dEVE2YWrCtGKtr3CnllWvHC1V6cD1
lRhXUbwV6+0jnKLBDpGVVtEeAzxOwLW42CS+X06YBvz4HGftpnRaIf++m+JdgJEcmVyaCgrolVIp
WGKzviuB85GpcGSunYafmClfvJq88/qWi6OtYcDxTRvshzoa30wf5qrTbNOC3q0WdCyNI6ndvR81
Hf3H5AUClsz/jESUl8e7oBcbDj/dhRkqfpZhJCXiezofRjUZbCnnpsr1mvQCsHxJny6C/QxrhIne
5GgFC/fhzzKibnP1Wj8toqkPevqjjsV/p0xrzi8bjQ5R9pQOg61icnqWNz8t3NK4LfoWxPAIuqaN
eoQej/mqvg1z27Ur8YEIvAYVwv5NMx5G4GNL3PqfKqyzQZ9aqTvDIOkGqQqxSiqbZXZkhmRUMKnE
xu1TeuSWcQJ8HjKlMYZuwVUc65rGhAv8EDPYQMDi00RNCzWjd07eDv7fG/4EI2GMnF97JQLO9caS
75G+PUws0h0zgx6cTGwJJ4dofgJh/M/9Bz6QAwrQjqzzXH/t6hMRPD95DdP9muH+xxgcpJR/SWbE
rFfwdPtpJGChGwsNavJ/sjOCTduFBs5g/tt/sgnfUA69KVGggLQCNOUmIHyLFn1+VpbHoOk6+k9a
VbhZVQV0YZ74J0ic1DSGUBLkNK3MzVgn6m3v8Q3B8vkwi+xHdLKmd9uULBRbb84ddvpx0/CrSzi0
/QwiY/dF2PAwVsfnhEfXI5p1y4sGTFxj4HjDAVte5yRKdsw/+cmUvgV/Nx7+fBGiQexL7PZXESC/
Eagx56nSWVYhApWHbbx76JBkhuUIYN1baPZDf12dnppIWIN1KIeFM/aXzemt2dt2tyC8UDCjKTcF
+iv6o34prfwRU5ld83Z5Ic/PZnWhAzhBMQyJrTNtbxjOTA9ZefloHwJUlbcDFD4OEYYU3arJ4ha/
8dsCNiZpC9nsRdQYvMvcirgzWA+TQFKziZgi19TyEuGZTRpYJqad4FZO5egPGZOq3XOWllEgGoNb
uMewqoeGIktyP2+IZBwT734EzVPo/mNHin3POLYVmgQTOV33O3ZRj5CoBcMERV0+buObxNHzZAfO
g1TAR6PFLkq7NHnEnw3GC79kfdqRyXYl4mHi7jBpLyH3qZF3qVWCIDO6RdqpPWwn5BGgMHjatwpg
k0QvZ1L496JN12U/HhGvgE1NW8rniPpvsLCy4KnmwqgksuqeNKIam1JNx6rJGAGpFdUbIXKPp6Hj
JfeeKF9Vot3L2OBja3eRsqR8cVo1P2e9FuvNBUCYlwZ5L+hM5PEOt0iaVGH+HDUXWOmssOo6yd7N
CGtm7GsD/gIuKpXvcldrTqMx/cYU9gZXnLvbqp5nP46MEsKx7nx7Q+YmxSMVR5wCuwor/VfVAZba
hQjGw/h1srA9LwddX4ZoWZXTYTSFJ35a1NeHFzCAbB8hbRlkEWQu2IpcaNCMGeX4hAlCtRkW9tYn
Tnf278Z9t6ZBUvrtV+JMhMzbNh+iBI3/rJ+U5Z6UMZO7b+CBucprO5Xhsbm0rFzSUWNzWF8XVIIB
ySsEDK/n4fY16X1DnVLvcjhZ2bSrpcosN/uWd5ZohbJ3PJb12m7XZgbO+lXFP33+odRNG+sQ1dMt
Sas4s7uFWHXl/C/Cy2pPIOiaobGNN7YCzXkqG1jGDeg3gOBV36l7zLAWdvpRPsGOJMwo4rJ+f7hs
nOVSZeknH6IiTlWP1f+7ig0g9bNRfyDGHKZJsdAYzSGWH2Nj6ETy/4Ps87lQJHONh0e48C2ztaM/
V4VXerdku8JD7/6JFf8hnuXLdjfd7PO2g3jchiOJlYUCf+5hgq/SnTSTx00G335v9cN3hMhm9t/X
GYrHOfT3AQLrqHIh4TRzlqK9PprgAQNsPQUNa+s+EGTijvkWaZlDox8MWxDmAjtRRXuS55PHBZmH
y1LUnG4u9+UXSnrwMQ3iRAYwhIbhN+YpTLu2Nxl1oLvmd0KSVyoZJO6iHpDVgMXsYGFHgKOyOemF
o94gauPqln7Kza3UFxH69ad3XXnzTAogCbVN6eGz61QiOays8MxRog5+JspKKQcOmcCOQNIDTiS9
9v3tWJKS5P4oQjToeB86RZbmBc+GIJzFpRd8dBU9vsoFaFRNHR/Qmo9mSWfb484FpCgZapcQ0KQS
5UfDOCLviDi0G40dUYhBGTDClTcjM/O7eezGoJJelCRtajStxK1fOJMqmM8IeNtgaPs/CBQup8sK
/PMU6iz30c/tofJvxx1qP8bHXlKVs764Us/9n7KSWRomc26P0HuvR+ul+f3hZxSL1/7J1xBe8B7i
96DiVyfJr5v7IihgEnoFhXD01t3a+n/LnKRT5d/+eJW86Ulue/9yJqcvbvVmU9Hdx7fPXHKrqjMm
+auW5HmrzWzKwW67Zvo/UgirPRj1+ixDrFbOT/huoCeAxMC6EJwnak376qtrjyrfR5tfOzZrM9yx
UZIpy1Fst+dDbll7uORc6o965/rmURHIulZVUg+y6TRJUhCZqitneDaTVrqDipa7XfZgljyU6jQN
qNe8H0sNv14XenO+70E0ZX+2qhRc2hPAY1wX2S6PHRm1f/b3vueohZALlKTWecsn6UPGOZfKJ8gK
SCLgjEA7xY9yxy9qlC2jl7iOBEU6JXWLEGJHifKYSClng1Lxd6KteP/0plyhNiav824atuS95tAQ
IeJ7hH0GyBDoORwQjLd9pKJy1Dbcw9g/D/oDbNuVM4AK8514SBTtOPChtJMWWLaBffN6jRGdv+Wo
ANgBZdG1yWtO5lN3S16L4jqxdp7xR2whX61aL2t/Alk23cESjNS8hgVr83hM1Gp3GgoOHA2VyYj0
c9+SIhXUC1eo/XjvmPqdGzHEjO2Gx6yKLs00y7lkC1LLoZngaYjcEKkdESig9W4b8CYCP5JhgKJm
4J1WQHEjDN0yS0czXHZ3FuOvd4jK54SZckhb25T9PkLKImiPjEMGw2wZng1YyeqepNqKUwhC292/
xCNK+wAEgDyVOgVxqzJSuxXoBEvbpgGls5ZsRj8w8WBPusFS/x8fhd1NUFO0K7wLZeSXSqpXqWpU
TMQsGTVWm9s1R7B+bQaUAiNbUMlVDVWct+IWDD87gonqCWT1QZuPQeDgkvH9ViC9k58xeLQ3tHxG
DKplsD60CzcJSnFVPLb8uVWMhDK9ksB6m83HMgoGc4dLpkKkZKR3vCsQIk3d5E400spgi15/sweO
cvtOwKp/GlxRSSV6aUK4H63Uydvz1PO0w5Mg2ifp0pgNiwHkRab1YI/dIpUskUtobGswyf6STU5R
vI6nMEt8T0SQ/m1w1U8RdtcbbycGwQmhySaF3WafwXIdfMYEh8UHQXn/B800b9s+BAdTUZWCJVvk
HK69i6E7LtLAqKEu+eqB8qrK8Jek/dpK3cEfgM98H+YGZfjklTTc0r7zYjWvZhexHV8RgouFhl4J
PJGwCWj/m+w9+Eh08tD6w73dnguISBZFs8cVOa0MyxbiKFKKbTJzWNTXc04uw6oABfZLSh87gG8H
VWEhQtRcm1/zRauO5AA5m4CiSmxyojfWH+G/ZW66QVeoyPr+Bq9Q7AL85H+Hurk4HYJr1HMkztiV
2JPBByBfl0SHrraJxtDcll6sZ/lMasm7cN29FFwFe2mxOjZ6Go0lZxnRfaa7wszpJm1sJtC2yQOw
/SJqI6uIMRc1U1mzfaxSVelhAglVtMgRET3gvRVJH14s60voKwXFjxIi2s7Gc/W9TNbbPSzbo2qU
W3xtsc/qvOzylbmLvdARDNu4RPZDfdupKzIZzqqLyrzHhGTiqZhXWZBvJoU2TKaFTaxRie9FWWkZ
booDW2FoCTjfeVxyO5B3TOjqbm2OfjdjzAT0o8y0K1YdpKJ3CPPoBS5Roz/8z5yCODdfjYzFMfPJ
sGpNMgrJK8zCJoQPHJEkf0QJbG8qD1Mc3PJWPuI1IRBfpBnEme22h6OTh1rIbkNucBFLwAdhUuc7
MUIy7nOs31XAu9ioAGXsxQKkGLFcF3k9TfX4mGqt08fgvMTETwiVdEGBzlfC/XdQxAdDlAO3G5X9
0i8JGZpA20zNkvcHD0jz47rUdsYXrN6FCby6fPBNPw34su1+P+/eeqXkx7rF47G2gotQakt35OMT
B/l+2oPDgONnjG2Lm/jEzbEFD7Q0ce0DDusKm2H47vk+AL4t2F6Afca0KfHgyf/Hw9GivpipcE1u
iKyD3ciLq2gCdfH+q3C6+RiniHTa4TSbDyybs7EZat8QYvE+SBocnDRa43H8+jmBJmuWZeye7sW0
rwUbqi0VqleVwPHGmlmnA4mk8x1CGWTTbMha6qJEJLPUEMmtrQXyA9DMOX581/enLl5cittR/n/I
VkXiLqn8FqKNaL7+NgUS9MCJ24YHYk7oMuyhuEQqqOxGJZQGONRN9lVveqCzNyStobqDAosPDwNL
tFm+ukzQNevKKj1pacGX5avz1FMRhrh+q9pAjsG02Su7S5hkSRnf/wbrT/TVqhX3Go4/e/56QTKQ
7C8wFAvEYUbiTWLIBV2MMtAWad2LFezH72q5Hr6VKVeSVUzvKSXvbdpanQc91pnKHGwgJzqKctcQ
nmCDcVVCglKObg8jX9eOQe9zbUogdANurwfMGIP8pzDm80C0WLVF8BkSGU5UQUukHQXjdJSBiwGQ
hNWsLV95P4QZYXuzhECrZEv4zC/84nH+gPmbQWYOe9TfeHtZRLZ7MkEguk31Fvx84ep72B4eXRIG
sFJT61LgaIUaBk7H3pZ116OAGNrMpTXDPwIPfED6JyzSWB/6EzGBjVu+39cq5lqnpBRDGAoUib/m
TxyzzGsd+EqJ2fBwqNeqQqa+saN2XoxRPoDMINE4YNxQWn+TAtXlqmQ8n6mDWhe41+UU1edScG6Y
xwoZTY8O7bhEMP/Dc2MG3Li39ICX4IkE7xpVl2fLyuCFI8DxK5q5jpLmkwGgpPfqEo30VmxUMKO/
eTU5g+49ThQ518pKsi8cMkKhqtXoCfpgwd2dRlmxmS3x9raZPUQtXPFqhN4RF7oB2va4sOOgieew
k/P7HnbN/N/PZMJuaVju14wN/fZm4LHHYzgQh9sUpbb9OJMK3E7F4ZcJv6xvgRTXxNqulI3XprJo
FtZf5b6mCEeDvI6T7b0QezFVdNLf2W7KnWq8DSmGqbYnL795TT6+oIFvfr4BFgKR2npMh0Y3Nk3T
Dof/cr5hQlU3tfm73QqccaII6yF1nV97GCzrHfyICTJic4aGxei7WDw47HxKuT2XKW5M6z2zjQ1X
L8DOmjnN9CjP5lcp40YV2qPQDHQ3m8WJEfOahq0NoiQtwrSdxMsh2e3y8wjRpNqDGfN9n2W4UMdg
LjNPgE6EcUA0JrIV3Li4x95TzmCR4Kiuj0IrSfe5n7B+UrZi5yt113GC+6BnoXX7LI4//UDcrsQi
pv90c415hTg9LGELlulKM2FpiNn5m/mBRxUOKKOrKdwFKNc5BYhFsz4P8yTIkxcCbPo1ZLZXVaO9
jmcI7Ev0izQ1dxZ89abdgaVbVgsw4nW9TwxW73lSilwPVkMyhdGhRYEA+iCeXOWO+txIAQLTcR8b
LM0pOBHMZVHNh/NM6n5OGsLt10PjDGvfj7z6bSX+qZBFaq0F2kDABRHRcgnOtG/AYh2A1b64hv/+
BpmaKD2ICOK2z6ihForkrPBOlSTJmvCkV6utCrc6KXA5k2OHlPiCRUBONHz6RUyY4rzqKOXwPz4r
h3JTrM/a8q0HOlkiYdtCPVkAdYpBHm3lVtrbTzSp/GyTMznOK5g6dTH73W00caTBxee23aFwoKPs
Rog3e6MzzCGopSAxheCEdv2NEVdBirwT5wzHClvIiDfDNUfWLQdfTtS62NeD/XqSRwRfL48qSzdo
p0OpM1PeZDRQZzRvp3q1leUVeMU4NmetSxCFbYGj3c4o16mi6UdrQ8VrAyybm6opsL3UXQw7aE3B
crE9QMQlDmbDrv0B6uujM2RjsnBMVcOCx9Jbvg7xXvmn6LmRjD/yT4KzSognZjhASAiB64uzVIdw
IBSmWMctf2m8HTJWlwHC1RYewvYnaiAr9yTUwk4ImkGn5tORCGU25k5MoUc4fwiqeD2aYATyX7ku
3xjGJOFWKPLQtsjRrGWXjiwPHAHlqM+fbda88Co042WB8aWV2rycjno815k362OWGUN3UIG7eIdN
xaOSOjJHCdchw0TAjGG4FNSCaF+waCba4XjwyZzXr5OVq3fo1z2pRPpAebhnf11TwLLZRs/vQA3J
y9/teANg7Nygf/+e9rnzezwewRhWPYV34cjIQ4ihVdMRL2znEP+eb6YCZQM1BDKs8VXiP+5aeeDb
70amfLv+f1hPUXVqivTaaOzZiZ5XNWK/eU6WXoX3D5Ua3V8BmOJ6nhh5DgcgpLucmnIOjxxom215
n21AOxFJs4+s8N7uqQ9GE0ql+0gIJ86du8qJ1FIGkupEwMRC5+hYXfVR8cko/tkGTAyJxTfExelM
7/+I3KzN+u4xIrgJWlUHkxRcFtxbmp5Z3HCJhEgfGjED0N6g+eUzGb5BOcbS0VAtAecgHP48dJuT
+liM3u7XBit9NNuvcn/ocqQv8mYebxPgmPSYOOwX2usaG5FfjSbIzrQtrOpDJU8T3LfpkRAeA9P9
nZYeNToPiTasSrt8NLrQ7e0kCrSUAkV1ST1PlCDy5keG0/qDygyfnFB3jordEEIkvODL1N1rWFxR
JnclSVBOjxVUoxduAK6p9H/ZdsFB0mAqGD3y1cQuqAjQvONP1HP7D6tA3KwD7R8O/TnkaSo6Nbq8
e6lTa9ditzVphsxbFLL2LK3DDoASJJFay/C94Pmr5nQxQ2i1jqW5SuVn6oAXaU/+68/b6AEWlfVF
tp31dbV7+IR2YQoiZRTlIUw/utMQrBjsGvaaviEpvKlyhVuP8V+TVn8zpdwzqxJaY+z6Qtbzj3WB
kAJOJHS0kl1lrquM2CnFFI+BitBIVRR2IA98zXccs2/deu9DMpBv5oN8KG5hLIeSN1Lg6HKKsrla
MEdGc9daL4AB8lUgDOkmQtHehfSU0y5sv4jhzUmIPkU6eiDobXUzBDfBNg3gH5Nwmnt/UNw2X0S0
tcL6vV2S82nOHh/xA9o2gyqHWkyFg+LQYPp534i5QwJM7jdgWlEqZgfBZEkfnMmII1vzX3D9GWaL
veuXhahMrrBJ/XoBiHDVpOWTFplGGkiFoZV59qNbKGjOzkeZ37zoSNu5JUdlBDNOqf2mIl1ZgdA2
r2pMXYMc2y6ac+aWmW5zrdIEElhkgJCGuntZiDoUpMyvoIX+hTQgFQWgPoQ9R/ShLaZyIj10v7ML
30sdbtcfiHtq3IaoirX3jKi6nwi2BR61kS9+h0MS2tZHZbWNXaw5Qn8PGvYq29VyHa4vW8XmqJA1
8rPw9BPDrJdzw6uzhQcluiQdP5btYuYke8Mj8IIxSgm7iiATITBGkzgWuWr3AD0XHg9JygpeRVNh
yFF0tb7yoffR3L7iSzvqxd4nVZzLyAOrV2HJvg0J5etsCWc9cSeCZtVyWQ2txm51SO3TB5cXF30z
jHZCFmv92cR1mZZIQ5pjbHUx6u0bX0weLZasKAC92JyuU2nmrwWrDM+bhUNdiBfhNvIMXPhJEdE9
1Fcd0J6TF8pH7Uh2XJhGFkR05TCVXklFNFfjl21tGIIbUWwhw6FpGgO+M12SJFfSiUri74lbPly2
ZdiBz4Z6Nag8WJ6kr9qDLHhlsUlPOoeHHm3xlTWr2E3gNO8wLz20Q6lizUgWiIOSzguHWN7/H3Id
yBr/Agt5h379oaPPc6c09Jw0EXh0ATKVoWEmCzfVby3064AHIiK3iTgWv6FzLW1B5Ly6iDC2pZi7
9J7AzGStDMrwsp9cAObtzZlRwmahMRqDZEAUmJbJNxnEdwXF2K+Cn7FtSo7fREoj8p8GFNyrIo2m
RPOuj1HldEHk93UWIzqkkBGC4jdV9LAqXVWSj6KTy7ekM3zf6O1j2NupXduCjrZId04s2GckIbxr
qe333SyrYPrUkFxIqL0a5WTYoq+TZk0/hgU1B34lN+VH4WkVhI8viNus8L2Coxzr6Vmz2igEKhyd
jl+E2mc+Zt1txKHNAmVgjBE/PYUjqffBOCIAA1ORWU/4YPx62hriEhAXQVrfFN+BmaAfJn2wM6z0
Ld0hfMwNdtmok8iDxrqiX6OKw0OzZuWTXQBVDgHkH3cdbC8vGmLqyHZiZkL8Z42zg26dkRebPkNW
fDOJGXXlPLjAF4spVEZnqIgiRfpEdCz13a3iRhN5Qfo5kS8gC0qqH1i8G9Pdhroauo8PoPkwEHTu
LOqaLXuHQ65elmYZ6vYARr5U4PZXLEPlXyUrXRgkUH+SclV9RPMPBP7ql4tTTfQ9zIOsQSvweeMz
IS3a/iqdYscb/y2+4/MCHXh4I6Uy8bJQCHxJiGJELXKBviedFQhzPWDIS+uaq6mrts7LVGmubyzr
KqkRG4k+QaUEyIEv4NFp7fbhQkIv145/layWbMIwmo03jjexl/VDT2UxSBQ1RQXOPW6c2/ynZZNH
tORCnC4UmHsBP/tPYYoeuBiF1yY1k+NVk28wxuBggJxnKjolXTMHM/fABgjQ+ta6SrsCXP9IPfcl
A0+HHYDmg2FRdhD7hxgiEDd2LlE9fHNNUrDkETDrIBhEl8woFnCB1UhHYyVD02M54M14FvyA5ieI
bCWVW75peppLcTcGY2mk5uuP92KcpEbPMt1tXVTOA49Y5RcrUyWnGY68fCRH6GzT8dzecWdLLS5K
4vBUYw5UZ8cZNlPDQaoVtoeKjVeYVombDmN2HbBThxE+SP84tU1HKhYEFP/Pu7m6EtmGjt7/Q4Xe
clLIrk70NX9TDhqD87SQzohMMh0TrFnNQefX10nyN1dZtHuzqpjL6YKpE8wo2x3SJz2jsslVAtou
4xvYvWZrudVyJxyNV3oCPP8zhCr7TyugjCJfQzCQ1uOS3aBngs4+V2iOYOEdzN6mBXzin8kaFgc1
ZnYDhtD10q+FgNkAEcezhXQ8NWv2dmN/YUYNKgIhHQQHNWogAPgePyQrMPQECPf60FblXRhR23HW
17GU/LBBaZAUR70jK1awqTDeeVa/wTClJCN1QQpjFXGKayg0Tz3pxeULiSdsglKwIbjk7orpiD/X
9gSQPpyC4jgYsu9WFCSnNg0Of8VF/M5z6lUWzIi0z8W/pxte4QSpVcmhqWEhH/pG1DSyzcLcDeBa
ckWDSdc/IIoySGILQSsmirBE2NaTAXHA+emEUTnPhV1ihIndX6NcvlbAjx5JKttAUwmqc4E4a/Yh
KS6ncE81PIa3EzHM6j6RYrkyki7KfZxq3RfgIChtAE7MjnirI/jQHQm0Sr3CTipuOryOwzynOSJY
ch3XYw8yw3a4YolNaNPcfzIiXiwnmXXsadxe6JsoC2lvMMIO5EoMXrNL9TrFaN0ZZdYZAsHqmeHd
JIk+c58iL069+fpCvmKJZ7Ev4NJGWzj+J8n0zK7gvMMcGWCOAHNpyp0T0qgGh7jPO+nbmCGIqsU6
WLYnBuh1FYqcp0UFrzEhkaGkhi1HHLI4obzgX/bbA8EsXUBLfvNSaTmIsIv/k3GFRNcbqzngpZVG
gHNha3l5kY+/8rYJe5rL3atcCm7QjPLh/pbLwg5AY3RFy6ZAxLuEXBES/PQcp4vld981VE8rRTrC
OfrBmhOnJh6xhFUKX8fpwqcs1sPFLadJxWPNC2J0+EoxepnYhFiNwoJQNQgmsUyf7ZnPS6VTUBto
0k4CKIdjyqE7EO5NfVGD9O14ZtEJ2U5kmejBjJg1ui/ylKK75EK6g3150H+rVoECh5CS60O6uBQt
PrUW2Ys3e8/DNI/0Vy+T6pichd9Ge5+PwApWM3B6EYTiiP6GxmVXRScgq/PIFTfFf9p0RwPmATM5
kigPH3GFgE03d1xdIn+19dSofVasm1fnSRaigMioLnhv71JPmnyX6rbqL6nGyzEyPM9RwJ9V0Jv+
apja5aF/s6AcxGtGq7BhlLv3fjqMiclY4DB8WEQreGO3eHfgthIQ2N7mmKGnxvG5iliKFBR4+/2d
w0Z24PmxGyiZY8UDCJi1Yx2eAnQ39FHVwJY5CGLm6+KGHihenbbJxFVCLv5ua7zAsWmsRL+vOHxP
SrxTqPjr73zLJh/XfcnaD0Gw0Y2x3GCKCTS5TQtmAX4YDrvoe+wlfrDhwe7A9HJ7fDBi11DQ2BMH
ea3ukGSmHBbJGRtL5HyFtyA1h6et1ebv2OixhIEjxcY1EqGlRorMvt7n7ApPNHfyc7GQeDzYYmP3
yvLTHZ9uzzjHG4e1+zvUuB3zujYOTcmQZSjkJ6d0t9Zz3dI9gFY0p0gTuLOpMziBR752LI9hGKzP
kPpgYD0MXaEDzjZ7aqzW9G6UAv6Rk376XvS3Tzzj2b7ycifIQNJk0kdYmx/veEL8qUpDZ2Hu7ivl
Kz8FYgDFi0PLoRywfPJFtycjZdGzJBjp3fSUu5Ny6nr6TjZ9yGc03IbXmdOTeaMPGfhel1W/rYsC
gHqtSg4i2slw5ylTHhGPajIxy/3Y+GIyRoDX5JtzmePWuKbjr5yeOH+8jW+h+Zlm85eK9Upo0aod
eE2ZiY2ljZl5H8S8JZrQuHOZOkVbU0+WTBK8zKOES8fUo6EJUF9JQgX14Hvhr9X9XVh2gD/dk1Vp
suYzCYc+VWBMN/F/J5WTj6kI8b4MQ9duFZ7o3CUiihBTNUo8SL/WtbzA9zKzhn+558RxF8qUEqIC
pRS8kUCyRXn/e8LrqUOQJJoG9gzHvRRI9NEuhBjHPvuLblBQD8TUFfm8bGgDJRLH6xyKTApKffJD
j1sebnVgGLPO+IWaEVA2zlGmJlk37pJ5Na/g0hzh+5iK+jJKq1sHphzvPJsUXhOguHcxM/zecchT
8c/2TxjYCp9dXaCDwRT12+IKSMsbhWHbifpZ/oRYt4znpfwUSmVha1iAQ6PL2PO1V6y9/KhLpWrE
bDEpy6c6V6JG4HmJzhWF1W54p1aI0t0qhUUBhrFoaUMptBBdEthIRZaHiBkUApmhKhYI9p7Hr/PN
Dt+htNrOGdKQLoqUWG0ArTyZCDfeTEAGtep8sXSCMc333YTD4X0+sNkOB26Nb5vDqzghCRf6BvI/
+8BES6rSmgHHREHb7TW4QQsKdUUJlSzsHxoR/88GJV9UMUsPkuuW41bl5tWMRJuZVWM9NyIaJQYx
nP57xt20Sp5STu+T99rnbaNN2fBkT2hrTYjQ6tAQh8wp3tkFoWgtyf6iI/YYC/UpyxpETkoMHT5w
U32JfDLK65YZ2RTEO6+OOewqsqeOPNlMWOAHiL8q+SynUsCkkbLbdJJboNp23hw0JoWMUtdjmN6y
PREymVfYaDdgsRpgc1fkiFsikTAlrkz3k9D0dElgp2FO3LDjGvgh1Iudd9hVeKdxC/MhEY/F+BKd
pcx3JiKUbQy/VtHaKUOabfW8PX5gnSrH1EglLRgvcqhRPS1QihV+QDuXByxjxXEYpSJqwpA7Fol0
SoXBjLdCglr4gzpR8AC7zOiJ8xeY+3E9gVS0nKD+khJg/N2tKKzhXuaPG+t8yeih7a84/14yOX00
dICIPVDGEzb5DEwsjnHXZKGtfJHvWQhr5T5RlQnee7FKstWTuq+bb2L3DMMcXuF7Coq9qtrlRSrw
oC0wnLuD4rN7tGuT+bXaNpvd1PRt0uCKF14g0QKxSmJRGP3rCku7QqQb6gYxF+HLrruUDnx/bxRz
9Amo63lixLFzAuCl4UbQkKTArPjmSj+wRsx4DzxUe5xj4YNwyFIWD+YnfjXCAWBPTEL1m248ay/6
8tD06o/6A7rHlE/mt/l0NXug0/UODOu5mtezhetRVaODu0sNXzlx6PFx0q9ru94DgZ5pInKTNt5P
V+2CZYENpDueA9/6LMxTL0EDAGSXBwre6y5C9trFBFgiSrD/kUvEF5Q19oVUBWezE+NwxEfQY9mj
X5zz9liUdXuYsSSVPFlFgpBrFybBsXrkMM7wxbCRj6Cmj5TZ4gMAfaJW72fOikN8tQMw9K+XcIcM
5ZuBEObT86mRb6kVHT6XSfmdpiZg5CgSGEiaoJs3h1Q7nRPuSHsW6E9E89ssJjsWnpE5ZC/LWVBr
3C3idw8xJ6cMAm9IgpkafrAuBCu8aea2StVgUk6GwuSSP9Lf0Qn4p6j4/8mA86tKTy40c4idhBvb
6J0eH8SNW0IqnbZtksup46+c2tdsHeT0wZxJ3YurA1zVM5EZGPgmIau8UmtcAbpVTL1r6rq/1u/W
iNuLJcHyOeiuhupM2aHVMOXEOw0DPw+ZGFkzrZ4DJKFA3J/Cjj/M8dpjEdPa08S9Evxcm4U0ffAY
W5zpCbrEYSKHJ9WO6qYZJCR9YMNCtSsHtrqgLDXw/c+uRe5RL51PPeEadBsFwDOdldOzAM6Z1Juu
ArXZZxYjfaBF3mWHRC+SHFqt1E0I1padrTNxMY4m9FHVNnqWFmMam6kDv+EDJ+PTRVWXSt1lT5b4
wIc6l/9rBBhdSpvtLu36thUJhzfQZ1Km+9FSy17TAydEHnNjAdpypC7pWy+mV2pm/0PyfyNxYHxI
J9+oOqQBoPr7j9CtWPAjaSRBNtkp/CdqZoIvrgKypFTVSBT6sgpdFfGhyxLT3FIr8vkQAv57CUeO
kh3uUZvrn3rH1NKytsXksItA/rpx6nEVPlhqqwEx8Ns6CBaWclgS/7t/GTJ7Uj0PmtECu4/gS7Nn
6ZJNJ2vmRtn6GhEab1kK1DjpAHZFDGOPij5sPBQOpDj3/DmFpvZ/eFVqdL35JYVRwWML7ynKYqGH
a4UoKVOKZIGJhe7+SNUsFw0ae13FRXTPz6Y7CNZPNfJgcNsafNCjqU9KT0cEkYxDXyKdwEBjVMmA
/lCYO0prs8EAXBRG3fntelP7oL11ON8XTyXkwzh9a1TWJbYzxtvlagTrJUz3Jy68/J/PfIsyz7pF
islvpAYuFvIPdo6x4vRtDKd0sWAPDvwrp4YOsN8aZGFlwehzNDvf0ocJTcD2ja/tl5sPeeCSmhn8
h5vcu6grfG8JO5GgOldOzIxDf8PEqu0UZiptk8uOvOFB2i7OyG87qsU/AfZrHNAjWoHL+J4cj4L7
Pe3HQl2CM+ocax2dPlnXt7R6ebYOhPhx4kL/tm434meTejwVm9BA5uU9LvN1xNWFNnExhNCXHSc3
YSNa8vJrBItj7cRiWKWCqyw+KVFtYRprvESbePXgUPOuMEG2W8C+2sn2crCl8/MOOtitJlZq845d
MOeGBjslLooSSvdWXG/i4wMKz8vbuXxtuKBfmuRG7RYxhiXEuV+SgFLWktS+yiegaNm3NLgtyFtw
+4onQ0heGj/d0kq03akTIKk86kLkzmahjB04fIDdOVJALm7WWhItihURpmRAwkW21/C7REE9YPrG
6OJdlRblAh0fkb0tpZHX+uacRRbsC3goB9zL4vZK0KO6Yoc+oaqiyjfsnQHnXZwGPQ206uZRey+X
C2mkZXwD2zTOKxsIRptvrPUVn9P9E6wUlp/xYkaWq2D65rZlHhp/8iqg5Y0DGYFiZQ6iS0tqGBmO
NVb0HX+A4qFVDHgZFNQ+g8xGWEG/zgcfzI4eXB7727N8VVokW/LANLv5mi0SK7JZkfBp6zj7riiL
X4hxek0X4SLpMMQd16dO7SCITsY/vzg/Y4H4pYj2gG5LNAzQTb70B1F/kEpCZiRbOrdvD1gx76co
+oCu0Q/y2GXfRYr+KPOvuTgb5BMVuQ75mS1h4GTqqKy3WHrvgsfZWIAao4YP5l0gL1BeT9gwY4hm
DMFxP0abzWwGjJM82Q2dGKdRvFc/6InuNeiD9VtX7I7cfVWfd+irimlmH/Eb+2AdgwwYK6vhekPt
ewp7MqkJqt3/E1npTFwMsxnHEBHC61+dxsxA0XJVf+G0C2EF1qdQm/jswJMvuabSi1gK205QUGoI
f0QFcdlilw3JZEghcxJcYzkNkWuP0nCEIu37xjTP7UnLEk62MKkkVq+Q7f8jpVaHYMPhQzbaB//j
rKC1iXX/5nVjC1DOe1Xji7t14QBxSGgZnZl9fjC5fj6wA1CkM+YBvUZWXR85yTiRBaZ4fFrLNPr1
ghBGL7vsmVP5QZWv6m9ha7Mz2wY/FQ1vXgQjkEoxH2+StltnfjZx1+D4XuaaOJ/HtiF9s5RD/akD
9ylh2a1Bw9AgyJmSl304CU1rufNNQb3G1IBAzGg4ge8NUBSQHFlOCPXClaMIb+1zLeTAdLbZxVHO
qM0e7WtYUG9COgqvAib4COkdodparu6jPz+e6aRakt/KamZar+VKTzf+bDDOBYdQ67yEAgbXHLPB
I7a9IGyARfS5hvzbXwW9N71MlNrqqyjKRfsTu62APCMdRVI1ZV02o/y9ZLuVdjIgywSyNDew+mmk
ABsa212QHYezDjZmt81umljtizArwf8zsdeGNTQVUO/pI/Qo2o19wF7I6GQXqbOKXlF2VQNsbbRb
4BsV595PS4psBVWdFJj5W9sTkCiuSF7nP2qTPQKD1UvfuvDqWL5aABuGUIhGwIWEJ1E55mVj4Hwe
A7Rx4Uy3Bed7tKBMAd/TqydJx2As87LL+BX/pCwYljhVx9ggZ+d+LzFC2blFWQzt6zxq8EuzBOi4
Zl7NKRzqfkrH3cv/hvzMULJ971n7OjHvY5KrQ11LzuloQDdQw8vTrZC+/VDHwg9Btgog1U/iHrcl
lbiyiJ26b0BCTcAww+nMiCXePulcn0Zcq7iR+qHB9BiQLj8rioE2OMv+2/dUsYBCIrI/RyIhunxW
kCOGGNTn96vtplNbEkvmrDaRgKcfuDZ/f6W4eR50yDPgM3tqeDqHkglhIuCGtCU9o63zjQQAdJGo
cYWZBle2Za2SuMqXCOP3h9gdcjYWODb1NpghjiRGHAxfU7sWQ+yK+J1JQRBYA62e5ZW8lehFKEse
RAvE8EikOSkASTrlhGweBAiOsmSHn3SHrPjQ5j7UhiSJMcYIzWqNazpcdniJRC8Ktv3qbGqALVK2
nDFmbW4fdj9Rn/NfSIyod2TtpoEZCddihjrXoXtgipoeaN1R7zpfCb9IqqK8DI+2BMoBAT+WjgUa
E3ycOKHU3+ndlsXOc7i1/UPfqw6hWclyOsuWyDd6Zj23mUIVxxmbzwIYxKlJrjMtecCUcS03pG4n
XRYu5UDZcfVK8BOwMWReMpy1rP+4vu0J3c6xucQUawCab/D4RTHYLQRpp6ekUBTdWnhwz2Ip00VA
iEBLL5vBhu2OGJt+5bUAsq182RcAWekUvIYbBW2hdjMBplMKbirB2PQvu38bSx2JQjnU76+rTdtJ
Fdf803ThhoBS7aS3jPezsViNesKBrnnnalkIXXNRHJxDyIkj7hIfkKQrhHHtEfp+taLg7QJS0v/f
MSMLIywObwYgyzCO9cIfdcFefE7tvMw1Ml70gywSOof8aE2SAYacLFQLjCEjwpEBMRuV4TaCIodO
x2sAqPzWjQdllPH9lykG3R6EfJRvvczS0DFChdvbO8XnnsJWhqRLoax36dHxZ2cQJelsTHq0N5I5
RZid4T4zRn75NQbtOS6DJXmXuFq42AOYPJE1pREW4M5nWs8/ahPhGny7MtfhpIN/hYiGQBtW0y9q
PmnT0at8Xvp520rDn3UUDY3mhp+hU6TBiPB28P2e+Z5vxtSFi3mmh2/b6SOAJkXf+fN127pfUwt/
4RTH2cDIf7NfLNIBlxg9DILhLUgxGGXWhC+bxPLtb9ZEJq+MfQWBHJcogRYEsC9lV1tw5qV/4pyT
ILG4fPtMbm/Az91XkKy8AV9CIeVVSM7etuc+ESBaRlRP+q7iERds0nIVJZKoJojhhB/2R8eqMpE9
4eLc/hMf2mg1Gl2ho4ch/FUfkNsqghGLrQgR3UgmlQYiRNNpxVUZCjsmcIqXZJHEKNmSOz0o6pee
g0XA1NtRh0CtqY1+cgDmdfSP5rgTn8TZInb4Sa79ZTGjpaKwpq8V6N9CzWPuLBr5xkX0fIeQz0CF
1SbtTQVVUo6isTFaf9gKthU9CZTBCtWr9Am8jDtywFAtWxoPboCoWYf67vrbgvvCX7V8yJQeWtzs
oKki8XH2Obw8cTWdkCOVAIAHwoBSaXSpZo8aufdk1THWwy6eKDKP71wYEIWaDgw2Lp+yUhJO7X7v
2fFOU1mWcgThM5iO3IeJDoi5igiEjGdLZ8zgD/HCc/XxdFvH020qoRLuAfSfyemBsxJwpDnD87NY
5pdXD+M1gpsJ5z5DaHpzGszk4GDKEYPVpUElcxGEIu9ujAZDcHYpEEB13VWtGeDLX95fVOAnLNc5
XbhLYkpmsDxBCRBvOroDKjRER0OU0a2oidCr34eY65MXlOrNwMkou3a8FdJmFXitI5OKH1IocuaS
pABcxP7uS8uOBEhGiQRf/PW/Wp/2q7a72kQptloXZo+DaPW95fG5dDrsfV7V8jfIOcs2M1iU7cfu
BugnzcE64IWGdNL0zbGpjmK+1LEvYSEQcx0+f2W0prKSFsv2ibsh+hzFw8vdgTXLTayxjiv5GZih
EsyTJ344bvDbYi89mZJO3TI7ODR912p5LVvqNz/adVNV/qq6FXUmKKqCGHxwcEh8UbEGue6Zryn1
UJsozEuaR5k7J/RKziNH4/LAzznIG5qyltMyg+EYgvYJOIqOaiS0SRyykOnFCVD/TPn1mMjDIPIE
4sLkl2GaBvOo+O0z0AKc+AcLxI7ZRKWzzAnqEis31Ms4d8rqrt/PblBqdFzr9knFRmSBcudycg32
HvoE57ntzTRJ0Ae+2pJZGmjeeqKWzEWKLJLGtgagEZ6DMDG+kC97HkybNq9AYElQFHE8AabaLBYX
M8GKIhgFnN1FJB9F7PuKCA3K38cVpYeTmU4r5u6GiW1hF139g48uP0qAovTRb5Lat53H1feCKyUJ
R0sacQXwCFnwOWlGAWzYWQBKe+TiCwfMIeOOc8wWkc198FOmIG3f2A2l1YmRg9D9tjLXUnZ0fb+g
oBqmRmpmR+wdOAfiUAti51Fc5Xq9n/iskC6Ky5qoBfvKA7lVkFU0kiDL2w0DKXwJ/03diNThh/JF
rLpUsWQpjv+E93DIjkjR1Nn/8E2/WzqL7d37uiix7w2NX1mKK74NyPvYapBTU3igUAwaNxtpg571
z9f+v4iM0uJgHyJFy7jZYPfY+6mOxkiQCOeC59KJI11E6soA55cPycQLEhEmYM5fCSW87rM+D/SZ
mKngC/GoT01n155erjLI5cu/Hjxz5TczoTkYPu4wz0fLIE+Rrl3bk4CBbqWitIy+6VovGRZSm52g
8aCFK+YLQ6Qj3gcJEgn5Q2KHkAhOz6SGHbWSqByE4xms/Iokn8AAzyiUREnarqHnSs6exF0VKiZH
BbJfG9k/RZ8uMiC0Um33uGGS5pp0POjr8Lt/jj8GCbo4j1iIut/o0PdBwfbPL6nux702N4kLG7Lb
xLenHhpurq+NZwBElP0oUgF0D2pc+QRS2Ssb48+1So3++Np6/MQPS5kisXmJq9JzE9ca86xhUkRl
ll8CVKNLOaIFgr1ePI5iCpywEdm/TQuktRjcZrM0E9/H2I/Otgw4M6md4GWxhYuz67megGY/sWQ2
bF2avbMVK9SwnjA8qn6qoPnyNlmhBd4/+MjInzV1+b074Vzo4qHSFh+WsLW7WjtOtmp6A63kOMpw
0gPFTTI4XO+g+o4ksQznDI/q8O260DpbithCk6tnr2Y9BV2eNdrKUSM2BFEzi/ssU84LKsECujPQ
kyuNfWQwDTRu9ly2pgW4k/saIoTQrtybDX3Nb+JX+RvOCg9+S7huP6mwel3N8SxrmNi71NaSWUXd
s6w1yg8bVwIp58Vc8maS8PBeL3ResJTgW+cAz8l/AgJuu8+mHUlOZiF/bhNsjRlpIourRA5S47lW
wpXADqQI+DFEdf9l3ERIlQrI3V0YLO7dAsbGLHBLMbQQPOh0RPmIzIdSI3PQA3WNL0xgyKYpjE/P
/kAhCX5Iwp9dyYFbsxIHEG5wA4T7F8ugQSCNJt7FIiTry0Zn/94QRonUo21GQh/AWROaWFiwyHnK
4c1d7XIutrBXQQ1j8rMZPjXG/J9aO6LrxMBnFSN9iYuqq7xNaFzwyL06o65Aolvq1r0R+qRLwjON
tqRToWsAgFdIUgfIMIjVmNMSN9IUBEAZKovb1DaPlO0Ozj+5m0IQuOE3v/ydc5pvva0IUN+kHog5
c3IZxnTCHzclB2IWDcF5u6i875Xce+bC0l8m+7CCvPRkgt9VoJHai9z/w9c5bemGtcTXjHdw/wX5
cvuL4vlwc7ydEQ0B1ULLtsR202M3xYt4znvhdCRGA9IPrQxqdU5kBlgEfzG02iT0D6U2EtcJgHSd
fCHkaiRCqyDPqbxXi37WTrHJCFpNR1OOgtMlkypScAzkQ855qFKySn4WOF5Bw/KSlvHJ8Oskbo/W
fYfLi+/9FoJBNtWnkAWzJfcFxcOdTqbteYRz2pzIgWDMukof/xwsUSL+LXjOpU92P/z7ez8p9sab
NRhLxVsCYCct7FqdxGp9ZlxodivKpXzUeUJRkb3UZOk3K2t+cjQ05nFmY36j2NI4qkYZb5OqGcNP
w7iSZ3gPm5/HcJad+YkBDN/3Cg0n8wQ/xFNWsEN9mxG5HCjtl+fZwzXap+DWZ4DsBByUoyrA3caG
DhteVHYTXivzVdyUfUbZvQVtr7ZmR9OUMs4yuZDuBR3oaSUNpPbTmctKvKGdOFOHEAEtVTL5wMQR
aOI44WDkE+RQP9lZ5DdiqHLiv/npmi/60NpEcFDwMf9RAMYSxkLMnGBFC/UnLkOkIXW6pPER4qpE
1V9T97l47/jD4Z/rq2mMnkCGgy2S5Fh26/N0st1I+16qcgtGAqoykARdDcNIVeLNqY6miLk0Mg/j
G6fN4DGiJ9p4CgCkKHtK8D3Pev/FEHz1/2mkFqKdFqOPv5lw82LpeobT/0NMbwAaqNKTIEQaicYl
ikP7qumRnBcQGrZtKbae73tPh7ixXM6gwoyrQo9WKngYvLsEtT9YpqUqQht0LMZWMNxZyf/AFQuN
1WUGcWo+8VnVDtMSDw7J+zw9sGmEVUeU/Dx6nyJr0UUi/0p/1TdchIPLtOY4+0ItfXp7G2oi9lyY
TIoqrdBQlWVEDJ8GJrWyiLeK4MmdvB7qyboBOtjecsyND5it3cwF4+SSR8Mn8BWuvNzdH16sRaqO
6Hm0LoPrHWUJsRFDuhhzv2ShYFUa9GhQmJ6C3fdAZrHsdTFmFjriSNiBHG5svx+qkfvU3nb+GBkK
ixX2DLt6nlcYdZVHLyS8YcYDrgW5B+OhyvTNkC8OG3M4aIqO9q7TA5F0E2RTX2NVWvTlS/nMS/r6
K8Ok1kGYvb2K8s/TQPWYEovD6W9NJohX+YNVHuzqjS4tf/kxBGXdfxiIHnKikgE6Cg1B/jBs5E3P
yjxBhimiIOuF0cW7esoZhIB2uOi4UaersT0VwklVjDBxS6NRlQ9YiV5hTRQGtwGt9mBTvPGC0yey
cu289yvbYVE54xLIVXDhh9/2bIMuZlovrUjuGmHVF92bMXp3gd5RMCDXP3CK0dWmnn1bq8PB3nB+
zPzMuTGlEFTdw5lxpYhiSuqQ0p8/JpPmo8wGyf+11yHOaXNsSuwo6zWqZa6kCt217R7KA0Gbclzm
U4aSiXJZwEcsp4ytoxvLu9jENtlLJQUR+DgR2ttE1bUDwZNhFR2Wrt77rKHEblqc+/SlKZ6lpT/c
DeOfMGnQ1fuFqxkzj6GQVWz9t3qhSzbEGGrVjS8kQnyMU3iwMQeWejB8XwShszTRudxWHGyeIKct
sVLpWvdTvIvN31p57AjDOP1ys5blXgV1CN5GQyb1ICeKWIUWaaEz96bMgvx/dOqKovARL4/LPKEr
p7UGZeQNaS9IlnrE7BQlyQoddM4jgxxeQDlA294x/Syx3gTKnG1PtCpqrnbNlOWeSbZAg5ok0VdV
kLJO3fLhpzcpBjUK1OvXf8OjBfgc8hK2vYkg9TgUSA270h8iuNLz86PnKe+qsTIoAssfHLsXX17d
MDx69nskkmgZ6PqC4u6q8PJdlK1kid2gwLFrKd/o6euJw2qOCgZzt1oRvWCvFcX3e1uFI2zl+T7+
FIvF7yq07A0kt277cHJ2t8kEKX2eeb78ayhsqMOymO9szvUNDGZHEePvF1Urua45kMyOMr3r5nPk
77SgzLTdTp7NyjG9kjuKxHXbdRDKcmfTOcOKD6IK/kSUUoYWZVXPyMvsOyqqGK4A43tS2F0gJjbF
IysDbU2ZxqGSl6M7uotdnwU7D4w3yrProl1wd0mwEPPZcean/0hkuM6/exI+Fmp/CJmSXJ86pOKs
3rs9N+J2xeD2xUVWeH3LjrtzvVtA0iv7bPkTvXZ5OflOObCHjsqaolcoQrTsrePqSnuZ+QD/dRs+
iH5J7/PbVxcz27p0CcOlqqvQpVhzLpq1408rjtxz0LXmBHoF/aCfmKRwof/NkbkSjRZDOZqDtceo
vE0EbGmBgBVqtHrHPf2/ufYFK9avyHOV2s9u8+NbvcC1yw31ZEWD5oiJ1Vyy895TOdFHDlCZvG0R
FRK1A9ZcHsy7ERP/2s+dsosmFITHOC+DbZzAgYSJiA7ZcFctmS3B/djMSzuGES6PxqRcVxeo8VH7
32a4nI+Jz1oDpJ2ZtzSL+T0M5S7YWv6YtCGIErQHjHGZkOo4Ti3s+0b+VpzJAe97aXDreJ+nW6Gr
NX8CYWmutVc0BhraKl6peH3R99lKc7f7NQxBgZWfTZLEvgi+IuWWQxzIYgjN31Uiaz/9HI6E+rnY
mnEj+C16ws/dBP3URyIMDsu8BaHh/gkAHKr45kaSiynkXnoM5Qszm3g7rjBwfPVMU5Cz96RDaG8P
4CUrILG/0KnGqKDPRWV8tGkZzGSQ/sHVj/ZjV9nYSffkUB2JhkwqTrB1LnP7ZIqFw9dGrtF5NMCs
RVUuU1zIy/Z2Tyze5V6UUxworc6Joi+3u0Rdn63JKnECx43xXn2UVDbe/CjS7W2GzN3Uy3Seshye
98r62TtQRCOJu5E8RhuvNrG6SfxDj8+sjsLLY7n4vSsKJ6f+Q1lIkToggTUMM00T+hzkOBxLNniU
n1LQGSzu26tgrlRQ66zx2xlQmhZcHFw4CytQHDjKigWkpLtc2JxwNZV7cUwAyddRo/mczY4OJMbp
Ff5QWbZy54GVxSOPV98x5JoRzOgS4m+OjYGwl6yNZybUEzIA7oe6Pvhiw9kOIEJb1SihFkihkMpU
Cc0Q2gVGaDogqRB2kqWEd8ph6RvRiwGHJI7t3N1XnUb2HogjO0FucNzg+P05Bx8FmTf/xqGWci2j
YKpdRji3Un8z+Ja6PDHajSBTW5whyRZS34TDhi6VGl6uOq5rc5L+vwx0aTu1rvR+K8ER+gCQeQuA
wFgknsMohMHQnZxvr30ZMnIQ3ZCj4qgHGR3kupYqtSNaCQfEJwnhMxbjLOji9T9b09HS0UyjFPEq
TGrL/xm2YoLMbNpH2ClhkCEyyyAm9i57PuzUEFi9ZXRMVhcfXsBglNSMVqtCAMGeJTI/SpDQv/TY
V5JdC/t6AkRYu2BG2o4RlMiHa7zC68BjITaueIgdkTRJ+exGUBxvYy+IvqeQXK/O0HxRXvz2bZA5
OpVB4UajHLyrAsgbvAlTxvvUEK99FUNFuD3qzttRPoRZpiT5DqZ/CKxowQoAvif6RflifhcG5d/z
aSV7ryFPochlwK6XXM4zc1S5QXlAPoqtfuW4Shqn1L+KHbnwvcc7ulNhx65Chd3fwDtt4uTKHv5A
duSqfRj1YBuTWw4Eq7bPrhGB0CZQ+5YHTuDQMANpsZIImiNiUP6JcPZrUnJbN2pIAGf/RDBjJcEI
GGKkKptTutjVOgshgI/mD1oGywV2ewjTLjiRl4cB/nVzyQ8vWpIbA2MTfRnX3YAvZdSLlF8oPtNR
4Dik4SdW1c+mShMtK0ZUsAIQDar+MOnPLhwhrGMsrQItEFc+LkauE+/h0X34o8HMs/wyu2mabu8x
grHQWDAzvZGXkQgMMKLDM957kG8I/Q3uIVRpXflLy7YEjAAQ8+UqBRS8Rt/3SIokIbhd9fGh5zE7
J+Qkb30Ufgd+1kpC70ZODBCRhmcyKZUJt3O3yBy2x1r7DsQ718uG26Il8E42zf1LDWVLq+ct4tca
ZW4AVFR8FyhRVAppddk0QnLWKuv89QRKVsgg7i8rPO/v9Dpa/z2dANQfejuwrOc/kYC5Sz9jNfRm
lOqvlPqAWBIZDNNrs8dfpO3xQogTHxkdh4ApDN7diEkCR8VFmLXo+sW4VJxT4SfIn1hGT2dSiAuc
oICwyxDmRa615WMQqTWYzJhA6NC5gHXygVplZWoGu0cagQNP7cN+755Wt4OiS0uKbwCe+yhwT0zX
25bLo0fX6OlEMa64N043O16LLAwTZRuSi7t9gQN6+5cIxuyXYV1TR7WfffGv1qkSq2a0uPnRSh3h
D/T9Ig9kYxHZ0zZ6WuGVL9vtAh1yw9xazcPoLBzm60CyTeypESfRcliSYCRJNiajmMFb5NVCLJct
rB7eb47E79uRnpqzcSGRzS9EcZU7ywpNfslho4Z+HiTxNRrAEX7iXHgUBcVLkJG0DLeH2jyr7rxa
LtZsBGmZNf63IpKlSnwsnqxzjZRu4cYL1UL1ToBpPlizWVVgEmDlhQ8fPYF6RZDGb4bXzmMQOaoH
6ONJEEw85mOo795c4m7R25MxiDKSvWyuBYAg8wcbLgNNX4Yrv2U0K7vuz/juRx4h6u3BvnJk/hVa
pzKGBYe4DVESVQDVsrUzXcFq+7Zppfl3CDNrBj03WAPWzipgnucMw4Y1qfeiD+Ozc6JRZZWFRRpN
khSzultcUnZh44VIqAJqamD3WpHcwXc3KTvuLgCXeqBIdniLRn6sLFtKr6eOXYL5tkF536jSKepa
ygfuYKTjOvj10NgsAVcvUHi4Fdb2s7VyM0Q1G40wpIUaoDvux6RqTjTl2L7yz91c/X2AoMin2x/L
pmVHog+r5r87igf5hhYObFGw1OC/9JLWmEku53WSwDWyDxZpjUJXY6huaEoTmyEcOksnHxYgy/qC
Ehi0XudLNx0t1HUX2RfoY9QoGweZG1PNTy2IU0gej2iOkKaSS3p6j3UVwzgDktIPAt+VMpKNlGy1
iv4DpdUWk1vGO86VdntBC9qz1al2kpGvODqhiQnLy1VOAf6TjUmLXWvQJAk7jzCsKLyysv8Mtu45
sgKFNZR5y3adpl2fsF8LSWVXFHFKDYyvuieO3uw7ZhxrUPNbL4ggWguw/1nIJaJg9bcPrwwQ01X/
WQyjv+uW9TQnnoMKwfdq1LBOfz55U2/HBY1jEIY3PRizqJI0a/yRqi4k7JEOmSiYft44Zn7qaBuH
wCaiA3LwkYfp+kiZd4Tn5/MHgHN5lw6YK/nxgKlmix93/HCpuNzUligOHDf+Jwzdg+AZOUryEvQW
iLYYeNNMpoMcRozOmss6jV/CwZP+xRJfzNM96yr2urm1tWIaxh5fgPu7JmVUQiRngNfFsNZeWUF3
J6kG4jieXtFWHQSG3oEfdPj03TVP/DS0Rmm5wUeL1kf3H9+FUCnXc9pFzyfdk2jmbI0z/FRl20u7
HIpwnuKLOe8eDH1UdsxD723fJWXkQ7zcwQt/TEnsXJFSHLgMwfi1YLnUwJxN3x/6JGIsQSCKBZ44
RxUGCCGJbsQK2euFXKBQLeMm8UJygXakHRWBml2jeAtL7SxsSyhWr2aR4nUS4xygRQLfro64o0h6
QZ0mRVclRcjXHhe9BNAncAaY8NyTRJLK8r4pmM5tPwHpiAB+T+6AEd7JQQ+tVeMHbiDJ2zTBlZR/
Q+oqBKqgfq+lD9+00EfuWYJoHO3h3IbR19gA/Gd05szyy4ykcMmcMbuTwt8DFZ/rEhKmdV35twD7
SRnDT8GnboT5mVXx6W2assforp/E4vSsCRcL6iTGxp1Gx6fUNmP0PN0al7hDGjxiY7CQcrTUlRqp
lzU/8ZMnRZg7+YMkUE5jq+HanzEDSVLztufnGwbw+gh3YrYjFkUSNS0BopkQtMygzZqx+VAXyS08
mcUUTzi4vCfGEqvC2ehXRPwprputi6n76CZUOazKs0ETXXDaJ0yackucsRxo+V9a05DYUwxChsF9
RiQ2EGw/V4tU2/6mXooTB7lzzeCD3eBp07PT3CPDaD/LJkiMTbn7bGYFGnulJxyMdCKoesPgzosC
soUUS09HXztpZqcjvdc0JduefAimTMwpDB/HsE/eI6o5ETJGZXhiwHm5vouOp8xedM4hlpFv/G7J
YrxRz8BTVXVg/XcW9cJj0atN8kxarjHZ2ftZC911uTN0y4+q8dzgai1SMo2KmC6GiMS74AkeT4oT
VJR1mDXLpWoWQgRiVpuEDMB24suoj8nfQ9eQQAR2IJPyrgCX8LjAWdnzb7+1R1Gb1uozUDMzfYl2
fYlpvIQi+j+MJOezS92G3jtp2yntZjGLRl4+hjqVLPGepf1WcndxMFG+oto9mJu3/PE87l9q+sqQ
vxhMypX1vhFzFpgA8PctZYy23fscw4wM536u69XxiXDpv3v2YQfirJD4fN1UOHb9oydMMHEn3/9P
HErKtZln9gi/ldq56Joh3sLD0wC52B7bAXGheeiYVE+ioNDjoUgq2HImdX/bwgwygMS69TAd5Pc+
dvOrNAzu0U4ViGhdFXC641vSSIdWUUKDatHiyGuX1D5HzdJD+1VSChkvBDzlRCbu8rTR/rFLnYlF
e/gbOMA+8CCRViB3+RtDVr6O1SU+p9DbGoflHlO7ut8Xc0CMTF5NlIFa68xGoJ0mUj2WfDO7VKC+
haoWwZCfqZ84VjVn1egQ0Dk+72QHP2vwmaC0v0jZ/23Io77WLXf1CwxPCcZCXxlYdy1r5Ear1QOc
CArwtmjq6cyUe0xiOrn6OVr5BTax2djJzJpgmovD7MIxzoHiUc2H/T4Srbff2tpus10LcVw1L6bl
e0PqNctLNjb7lm6BNckoIdOYlVUUwc8bA24fxsSFVgtS4pmQLFzJj/SebNEDz+xsZn9ptIkGPszy
Eg+sb5/2bW7aj9uy3XcQBBT9E+CEOw0l6cN5wC59MdniGTUjNFMawslGToFhW14FPP70WNDfjMvw
ZChHP4/MoBCWhkL0i/S1nk4rqnNY9xkO9E9Az6yGnYGIJrhenD8L4iaSqTBPAISIMRCbY4dg8R97
dOV6NHjoWwt3YUgMINMBtdA3LxzzaJDojFK/hK6iRlKtozNd0axnKlM0U8AenWiSx3zbX16X1XQM
RK0pS42TdgO1K2bwQhopyrEXICNg+rq5vQ6KfkNBBJcNovEw+WbtdWXg/ORmmSA+nb3weShS0Uj0
sHi7FYvRz5ukKlqqf0GgYlD/hLMxsusLTUl0UEzXaXCN5+daCbkcgXqMGB8V5Yp94OfxqU6IMO9P
0ExDU2uzrIN9azUiDgabTePlJXwSpepuLNF0nLuzi+SvX1cowY1xHqmsKTiRCySdIW20se5q6ZUv
yr3vsFNLr7rXZR5Kk7vn4fTSGDvGQQ/aZSk+SSAo8Za4LferQ1jbyWz4d+rXYycio/fwv7drbU9L
vTeEZiLt9x1EBNprb/0772S+jHY0whvb6h1NP2EUyXdBeyS7wEcee6SYfxNFlgDsA9tGFZbP0KVF
45qwC0AMsS7s2qL1s8f1cHS+MKBIBeZ8DPfpK7geA2wyHL4cBKMFQyGojMGW1A8G0YzchqfDDJhY
IhqZc4tY6zRiAx2cdfw9rEalYgaXUWYzmhgtZRLZ86/3vMYNVLL+ypqleQKTyDe45a7MD0CHWxJy
bEUmJPhwY4K7qpWlVo2o18EVYHXGumVG5LFco4mZ8GG8QG1H8HRApzMnJ8YBjgq/3XoTIVn6c6m6
HE2gngMY8H6i+zUjsTguhFSkTlmu/H/lcoWo8rsyw2Pc0QbjuuPnX/ZwYoRsfwK4IfCmEwFI8Q8W
yq33p43WS0woFNT0tQy3LLhCqRl6BzhR7idH1QU1sW2wzqAw6DVkp7uzDHCc0Hzlgc+AJvmuOuDN
h5pEuZ5+0wIiUTxhZ710soy0lZUguwJneqpuCXv5gWCf1TpYYdyZYIaqQEIQpnDfQ12H5ScelVK1
zysq3IS8llrzOuTuVwfJN1V3Bt7aMuRWD9vLusxoLKjpg9Oyl3WKYEM6Utmab8daGSJa+nLh4KUo
CQYvSlGrM3fdHY8zuCsAW9VpkombBPAfLgxYKRBaQnd6qgQzlWSvCFvbZv6XFNENjoBJHvBCdPl4
ukW37c6NySz2Tqq9knt4NUVL1C67Gune62uoMlIhkTZnU9/oEeXxMQMXeDNbUnAowG1TlNOAqoIi
tcLgQtd8y2EHjltDEcge1meWCs0TWalkwtIG9hEMBsggfn3e2iacxN6W5+9zGd9IW2JLF1iklFmw
DYGkkXV3njkv3z4jyMKK4QLmilh+HquHk9/FbjLWNVhRE06KivXOibWsIc5r7WWyBtey8EDs9Gdu
S4vlcOcXelF/3AUhJvYHdvg4I91+UB4FmGTzVleH9i7mfbX7pzkhIKqa8xy9j0WycI9wVQs9Ybaz
ziCJCau/WMbEhDf7AKTe9SMM55FeXnJuGAPWAJhyWmEw9Xdop8XHYoXVrMD9AlO/RqfxAmtPDb0R
IOUubJQaC71iXzYpYWpS5KEufEP1+i6baHf0VSrij5KeBzhOfNTG6GPqC74uWZMAL9zK4qke+q0W
07vXpP7sVQYHjckmHxRaQ6PtILB6fFOtQjrj+dXc4ZOOdnksLLlDXTcTwVqYUKrGDi5qbseA+vp8
GuleNNIozIpQjSqUzkC7/4FhjDcsA3lXhzMwIG17rx4cvG5k7MBv9NIJfI3I3nwgLXGY94lV6L45
o/gsO8DF5Gwz0fsZPbTCg9mrObzDLPGl8ephP1ixs88spl5cqxkKZTprhpcjXcSwK7PLIAsbXEWH
0qLvm63tiDmd7eqIfEAcgSMngcVyemu58/XGIARKkYSape7Lo996UDQy5UmMX5GcJLYXxzH4b8pg
21hd/BULVQu/+4LQb+toMv2bE0tB0uX5Lp1EBlOlltYcioIuhC4HgsuiwSTBTM1hM5FRGjDY8r09
tTzbGv1bqOuodr6+jMqRtFX9+wfiN1JyhG9JvnPNyrvFuSrUWDYfBQbHiSQhJgF4Zqud4NJTLR2l
baFFXkVPVlYMBJahB6j5sVw8LTj+Bu4xmSNdi3ZwzpDq6GyfB/E/Fx4UgXNHq6w8nkmh3pjr1KRC
paAJe4YoQXdgnGYDBnG4H5ZoQdadt27BFOvklufFJwhVbjojrNZdNo5OLeCSxo8ElyxWaW/IIh+6
O2v6Wk1WbhNRpnRqmqB+TSQT40+tVBRTQN+5/HK7I9NwI2lhycvGKxPsQFoo9AnqRgLdOIDDgnzh
ilsFh0T/sSXu8e60PL3Cz6JeEYFK12OLvxrB9nKE+t1YH9wytXqM+1uGvzaeM3t0vl1W9YK06nxG
zqBAIRplUg/j8BYAb7IRIL6bZROhzxFHa6qJHgULrAWIQCgnzgBqPqn3gdsY3uBEcmSXFRvWX93I
6AoUHVOEKjqSQAd2mL2izg7sEl5NDhJnhslrDIAnBSGps1Hqvv6F4RSNy71bh49crv0WbFVv55pD
N6V+bPIQhKPaqloDUlNNdaU4tImpZbbTib5QDMBfMZD0IrPIKvMC/YUQ5x/gESIBj/owtoGIxR4K
H0pVk3SWWk9nwUTxO95pYioAR9MvM7+gdtdf+A49hs/VGyjjJ1uaO8c0prR9fz4TsRumGkwb1kQX
nszYDoBJcXoK7d5uVTnZ3cr+nAFN6ep37Sm09TIO6Nmr4A/iVhg0Hp76Y6Xv83DNGoNz66HR9zlI
tR/z6Jxy0J2Or1IzU45HgrqGVv2PkPcdZqaAqDr4OCid9E51605ckvcT7fiNnxJ1IHwvt6QSQpV/
vDNeA2dRTzFyU48ZlDRJ9BuMEiBjHRGxM3/5MEUzGVaz/TDJiu3Ixp1lNcxkN5KfO+gKuduAkZ6u
ips5HyyhGLs9QIiHHn8xGSF0iRus5sF953K4BKkiou6ybvOv67yz9W2F3yEAJhzbkhxKnVJ7r9Lu
QUnbImhX5Ywmhj1EcppmrD9GAY15g9LEOO1GzI1cyPYtx+d7q3SeOMutCiFs2X674lrJe+Kuz5/p
ZZDXlqtGqIDby137Ieiqe24fdRbN8Rqj+ef7yCJoLFj4zTn6lDD/44AqmgkSv1anRL/Cm5iyPTWa
G1TSfMgpQygO/5H/ZfQYzc8sZzo6wv/0gXlMQpkOCfhPPymUe/nyLbr0S7e7IBsZNC/b/guu73XL
CKfigdNpCfPSIv5f4KEj/XL7b4vCsudBvvoOwpww8UsLDDC1vOp2EpjsOLszlI+O4mmpYFCGlg3H
ZOpjP3+VoHV6zhuS5GfIOE3R/Sxb6usOqNljdoiyRMJ1ZzBtm5DCGqKXr4w22jakTH+lkgS0CH/S
KCuqXtjsr7aT2Cj7q9haT8qAK67L9Rq+Bd1vBwgTmbnKdhN4Sz6kAB7kgo2ytFbaluI3yigomyoh
CgGsvpKKZmyTurAnNWsqs3Y1T4OsE02h9deG61rQlNkQnrvHJSaaCpd1zH8y9ijpY9+/VgBWcIXq
ABhjv6x67di+1A7oYtNFyjIFYVixDef4BSMWf85qRlC2ISTJE6TtTg+L7tpJ25eBniokHlhbEfi4
3W0u11+vrybVXduSmvLi1qlUKUUGxEox/W0HijzlkKtaLnoOyxCuFWWOc4uBDIWdRb9b6XU5QjmC
c93A8uCjqDKH3BCVNG3Y/bFvtdJZkCP96fCsT85ZIRoduJlS2e6zl473VDYnkwW+NC6jUKfinmMq
PvwZlahSmKjpKHK1P9XIkbwbrIDPuHKXJX6TipHRULZDL1RY9MrUFj5aws9vsSiuzZV+A/bqsp7u
Pk1QokW1Gx60D8FHkddkvcYufi36Ky6M8dmfhsH0d0j77VVJkzjOYHkHBv9iDGq0JUt5/xt/ipSr
RMX3+5wD3/y3MMPIyT4yoQIXlWl8ZS7LG6TSe54yzlRmbxr2QseF2TRYmV/cSDroHXV0OK50SRAR
EgAYGfnDwvxh6GNbTGOD5i5wY8afEl/SYFsYS8pz0HtBP35BhHpikTLdDhv/Yr5i/ELB/3lsiboO
GrggznKCh6EybUT27Sjr9ldw70mhWB1AahgIjHIeMhsRFK/wc+cKoU8bGcEUhv/rUHGz5hL4sgbe
0Q5Dv2rpIOTZo8nXxxpjd68/eSzsehXpTd+gogWpUE/Em7PH6SeidfOoJigG8fluQX3eJdMk42m8
xQDNBtOjNQj0KOK+OYzCfgh2SSwP+JKr+NV5MxVsAMbSpDunR9g5xyQ2nCLEoZm6AjLbQbXhQYj2
TIaRlpgYtj/bbYrurUYEJMDmmo915DGyLXK04pM5FEsAcISOtWNp2NWlF+Pi4UdClMlavG9r99nW
QUON4vhAyRYlAxEpmmr76pFtTHy35Fgk7oLfM9LFb14VHNHycELiIjaOrEPgITHulSO7PfMn+SKB
1ihQKTSl9GEfjFo8Jis9ioy9F55JzJPNmpgKhIpxuCJpYqffNDG3g2caMyFWWpkYP5R2F028mSkH
sLfct28ciY84RlBftMPkisuuUXuo0U4RTaXSYxFYwr+qO3/de6VxqYlh/0KMiFArWwcQllAPpTmC
8Aihf1PA/LWsmUmODen29xhgn5VLrgebn3JOA//y/59pGfG3gP6NLAnr9PGEcTLSiXB0kOysgC5x
LgHz2Gr+8RRDkabyEkQ3EN55aaW8+7WQJP2ET0JXSClrVM2M5n4ggJo2AXx6TqItus9X20sCt1+0
i0iKJNhlOaXvFfhpFN91DVNjHCc54iG0EOVm8cYgscKU8UG6LqJg03mOwxhPqh3oH8kevLQmyAvH
3nM9Kckl/luTPzBkYC+uYsx1MPMovn5wXseeIRjOH6beGDroPE9G180BnlR/vN4kdc4UKkNvZzCh
gMtuZFawFw7XUiE4r6+wweCd+iQn+gnYEk/cFXWMzPC0FrYXlhyRT6CJyxc+NKYbuDA1z5Pwd4lR
UNik/iD/ZErwzTgP4OoOs2hmDmP4wJ+btG2PwaH7mwitVWHyE6TvM7axpaRuvU0HS9NyZXHLOKbM
IPISiBtxLH7KDWtG6WLnuc8QrEhTRjroTGjvkd5kVeOCZqYwGuTvFunGqXaDSbbGWIyqTqsh82Fu
/jSKDx5YWCkp1fUOK5HmGhiqG7FE2H27R9dO/OhM8KX3PwLNB3MU9cZ3OcOJilT8nMOsyDab17TK
Xnp2rpr0WLqt6iU5MQQuuf/sD/luWiNjG14R9QHps3pRnyLdPv/h2GejCD8bOXwFJFBoaVSwJqiz
lTqzKTk9RJHe+s4j7JG5UQnL/KJpjtjd3UGpD0p8LzhMrfieYBEbdpurG87KT4OoZ3U1xj8dEWrA
3XDdHmE//2Qu9OINB9Xrq9x0P96INS6s+RV7R2iNq1NA8u9o60jIV1yzN2Y6a4YXbLLanKmSFgyY
5mIwl7H511oGKe86FnbPsf0gp7RDZLq//xLkVUDRlAhfqTPjbcpVdOzBViCsVT9qknWzXqCLi/OE
K5+2XMLZSNVfnSPB/P3LqzKXXxyhT1VWdkweXSGE1aud0jY2SzGGfsgYDtS/+WkCh7soMuwGMOAw
UD2YoUWWMel6wAqjpqhUqULd0rBZRoexpP4QCEz06zgqgTxnBGn0pFhjj5/20sYPHQuBUjdDkR/K
Horw+cLUFpYOkAmUsbuf/gMtn9ryqqzeoi2eXW4qkrc+Z2DpMP+wY1YeukaHiDkCCeL9pECMAqsv
Zu0tZbQzqX9VtS66Zvvcc19XbJvLw2LXPRc4om5Vk2lCznqnxtFTU4myZ7dZTkCZQiiqCKZd5j+D
v1c41eg0/A0XuXVVH0ycc2l4h7zCX7cgEFCqgbwJbNq+xHFSzL0irdGTLmyPDdCkTqDPqORCycPP
O3TaCjgvhIam0juLkyWhRzkH3wP8oPVmUdx6FFSiq8Kmi4HZ8kGDEuhAQU7cJCtwCox5VR0AL21G
Fxm+3vN9klneFJG21R9ey4bLP3WSVeGPbuZU1fSTw6zOYk8E27kekIAcmsfmtMY4yvJg0SUW/elm
kniGiQXtIJJblUq+2uwPMIMjNG5JXF2tHtH2kVNgqLoki+Gg+d65CQuzm/YASA42dqBaeoIdYiRU
c0LLvWZmDOn9oyFJQ8pQ0WUS9+8pqyKTeSXiFT9BYNalb3z0nDZBrEyQTbrXC9E4D58BxZ2RQsk2
CBUslehNBRGoIYfSvgu8TPWswYM79R6nEufj/xjf7kqXCoKUBR/Lo7kXuy3K9qRPKwgNIKJFt9ZZ
H33JPxZ5LoSqjshzaM1LdQBOg2KANPLg52aSbGvNZVpITp3IC8lGhKH7UlY4OOzANBHQ32QPngg1
sc4w4VMLpKOVWu/r7zyvsL6pp4zpGXDycIMG/IgXz4upKD4qh5wvCOGJvzcTFETiIDsyR4owaE0T
/cMo5FS5JJBglximT2zvdAxwPrPOmw4WpP2Pv0DL9R2ugc6DAJibAbAvseNPLyaAhnQtuH19h+uR
DIdEAMch9BmJJqmAZmcCIXAFD2fLWZqER1ObtcgXTYuNwMtfYpXU/Y00s8zet2L1AKiReYRz5ov8
rLsDJLoB5+RuCQpbWp01dDxF5wehTyJzoN+R25NRGvaX+i96GZuyemi5YRh3mwGtoNFUww77JCUF
i14LpTNQ0jXFSQSF65CZrv7RlwKMuMu9p1rXKpmo9cmHTPJ5KjQBmI3MpP3+tzGaPkNfYLgUYVHx
QzAlXNNjWyWXDnQi+JSpeHY0pv3VaOraAS/tGP547v40tubD/99GaRnJ6fvvGVEsgPCOIGa1Q2G9
v6wtNXF3YWDFBkajn6Ldzm7+khPKPC1a1BqrDDlLk/8/znCLroT5xtjz//p48ugwn0NYmyvHkBem
LxS9jjJ7Jx+IGZF7Wp+nXgWbMXAQmx7gpfO/kTcukL5okcrwF+8Ekh87xgapUz1M3dxb5VABnyRk
UlylOYuDEfwHtKlTuj1Rxc7jv2YwOLfKRZu5suAy0wxonWIbQM48Dvb1u5YnJyRqzclWSnq3NAwa
MY08VxnhTOTu55OFazZEyAguIBarX0ULBBtugLKh4LtXoCLaQ9QpBK1jCecjctq+U1IhqpVsru8t
byB4fNaywgIgSZLSQ/t5VxoRqMolDTv8anQkHCG7osFzOUlRQMN49Kly6GF9y2JJ3fwXSEVLbn8l
0S82Fi+VrSItNvVHd+G7Jmdbvqq2It72H/9FO+tbPNGYOUvpmcUOJ6pyreHVsW7evj0jN58hinIA
Xu+P+al09evt0b9AsKhHr8qqtmhT/LoQEpZr96G2NzdakDu1EQXFSgvELmeY70obA34k6G/QUQ9E
6/MZc9dUK6sz4k4DpdrhZDlpRufb6fDAjJVL+6qHpn3H+Upfej4s9mvpppUeop6VO6MZb+eJfVzm
ORi/oKSKM4uRyxDaOmdt1YxdF8BYDJeGS0/zgDSmR+m+rZBpE9s31W+T6YFZbHp+Ybi6LWC5lGp1
ZjSxKgtgE7cdT1sGhPt1LezUofsb8DpbfB8OH1dIAQX81Ttq3O5YUhTQSCr6APXr0Prh3YWB28Ku
glmfcA5b7pvfk/iOYptyBH8tM1s10YPAXTClxG7ReLAaMbh8+fmCuY6liKQILXf1308f8gLN2mZ0
kQh5ubYGXaUpS525xJvspqrK47P75XtzvBcPMY84R5extOjqngPFgTqiwzfVW2lUrHpnxgTmBNK7
VIU72xNZaCQXG07rsN4XfaezWu8L674yJp1LiJ/cKzoTL3wy5xUoVr2Py1T/s93TnoM8Jv9zfqPl
kwldQ019GEnp+9JSp2XvHRmwOUj4JMqtA+sFmsE08+B/XyptgqH4eazNY3bBiQn0aXLJRDFpmVhA
joCUlGKpY5HZz3879p7MY19M520ue8SI/WLgVQIchElOEkhtcKMSMhbudPu1OrjH10swRv3XD7qo
vYaqtSrjCKbQ3qPviJDT/OSKM6Zlj1KGa4khy6O5bpEdWJgC30flZmClksRHjEcTnyGtUanz+BZu
KoreYPDN1s3WYGTa9h0tmdRys+rg/P4gRK3Hfz2jP8JxOAf1h5589bQzPG9bUUsvDQgQu2k5VMwB
W2Lsjl6sOuI1TwiNLuFyPETsK2g68nCR2mhWgCIUIF8hICmY7unxUz2pCDPDdeA1FuUczMCxPrzm
h4zqJ3iWMoO/c2szXRBp60/Fiqm+iicMQek27cpvBYzQ5G6wW4rGCEJds+yc2DtpFp4SCAkXYrvp
3KAi5Q5+N/KTaz/ovHYDW1Jkz3EjWQhw1hcfhcILO0NyKsrtjrLQVelI2BkVmsa3O2Lu6xjUyI59
ICUikkzY4+HXJ2DESTbYf8ycma13Yr1yjInKl3ByNhm+/eOxlQqvsXyA0lSONQEthcYJoCGpz6VH
SqkKgH4kLDO3GMuHDBs4slMzt0YmTJu4QsJyl2u6WXYV30Nfd1MYz8OS266JZhhjkjuin+gDnLgT
JrQQgywRI6CnjPCbxCmYF9K09PTqNFk9mQlbF7R+UaY59X9MiEhaMyXuXRjfDIX4cSJu+Zjv+1RR
ZGcPIo7wLEZ4lKTtWifZPNQTK+/av1lruPefKjFbR156gLZR/OGqR2oI9rusmMZ9dll0wz3H9ygm
VuGP+nz49+VUpGfa+LX5GxzzWl1ts+3pyqiHWUbrY8S5w2VxhjWRTveo/axDey/tFbX8yk0kEisl
Nn0j1TqFauYWGQht4OvQ+SzPn6nXcZBcyhs/ViInGVt5aEBRPGI2uuzy3mk+g2r7H4sdMdWlLJin
By6BW6qBQuar9ZA1rR+YxLapx2mmUQP2tSpgLIYoZcCivIN/bNbqWq4fpirxw6xQb4iEnLjksdpQ
lrtHEj+KAStTHDkyOX65MAvjV7QVXbIcS6L82EJwYJvtt39QoRWHCaAyayS1U7OgG5ibR6kGlv+4
84lfFZyB/4hFl0JDZ/+/Sp4svFZ+fK3qBksmxSfg3pvGvQrV/0hG/aDBPWfbGyW60c2n3k2OeUKw
ZCmz5JVRcABpPsSRxJWKF6HMWXFd0SXWHhgu5UqvttGdp2PSKvosLQvMV82TUhSmn5+EU4xDhOgl
P5wyxtLLp+c6QNweWL15FvvsYCK4Ek2qIrInyegCVi4ppbi1fjIkEHNE0MDfAbu64HUozCMQC5G8
p16Z3bkX8h/bLsUwnDJoBq/CdBMRGrd9beDYqSEP6ThVYVjvbJZLxSde+SrZhF/aRVJA00N4V8Mq
ICgjAz+k48YAbhQnlxvZZlm2UovfcugjQMoXZEVSHyWyFNrZHvBWfP134OTn6i1qcQc6EBwc7w/i
gI63V91ggLb303rQN/EsPoafydZ0T8Fxh3mnrMxkbRUf5uXPDSEos9rItpqncjGhUxH7YARa7YmD
XaOHqJEII8BwKtLK5S0bT25DcGHJPcXIhFCfVwqjhoumC/t6X0G1vqyAjcRHkL8D7X9obHDh9gLc
7kzd/yLHZN2axlUBz3OvePpxfbRxytokeCBcRg7N6EzWMGbsY+2nfJVOUpEmkMEMObzrjSswh28C
XmBnc+si6Blw7TtIT5eRXzf2pTlmTvwh9KUQ3yco9FZZocjA7vcl3NhOkWFjRb3bbHVwkNQb1kIH
s61TjAfybuJ9c27/UbRV2R42wlUAl53qbTYn0GLtOzLT2Not+mY4ivNU32wNBysUS9seeQQpGXJg
x31RKT2D32Pl3hdbSDDubuu8k5B/0KGPIU5BGYFD/G42k+C46w3ujCr5X9uU+Lhu1gK34oK8aEhW
6z1tT99wNqOGjyU0NEOyA+AjuNIumCYr61BojnoyCOMQeqF8Dcbw7GBFRoPNfzofcwDILg/zoV5R
g8/nOXwlEEwsjEgIeEE3/I9qzN3rWiWDTBgBmrJAazWNLrRXs39tCGKUKW1ICgk/O6MGSEMk42Ed
aSk7HC/ByZGJ2hAh6s9Lb8aN7Rcyw5rRCyfs2XjDKJNVieBvto66m0TsQmKpK9zDvSvs6Gr7MIJZ
kzHem0Oky4XnwTPSLGAYj36ApLDRB727RLghMcK20Ei83u8T788R9H9eXLCwZDWYyerkHCXywvU5
qJepxXI+NYeue374FzCV9oVb3YQzhrCkqlDuzyvDt5UIpPnNldqnxwAUmwIhHEWbGlwBUnXtTsdM
sH3Rs60GcZD/iyl0UfkC8LT7QzFzgb5hfvAEfc75aQl7Bd1n+Wex81tagPVMmyBOjkttlUBD2zuZ
WgipeXHVvpJdCYqg3vKbNNbM6J9M4xzgQACTTlyAYi5OyOG0oyEDkt1zGAE47kh9meqIlxZvwYV6
XJw0EpcVaEZbhclmoPXvbh8dNRIjVnwJvekmBSLB5Im2CT1Dmusr/n4pdyRVtjbA66KZ4Z4fhIuu
ohpXNcbJUQBaWNo5r5IPEY19HEnbcptS0H5fK0iYjlSqvAx+RSv2UP9x57ez/RcROOPm907TGUnz
0MuJwc0vR45u4T/R6ala5VX2OO4uCI0atW4L8cEsNuYt05Kcb3gZ2z+QmjPv1wYlVH66XVnQ1sF/
IH7G448udBPpi+7bP3TlchoyuYRNqV7Oq60GcuamNFdo+FxmdcXMfnDu9Z7iecnMVcWo1Pbfs1DM
5OSUQVJzehi1SB4zYbt/atNzIPpzDOmFwjFbIM81h9zh2CUy+Vv06qw4iVpKbTiN3IB/jxW5a3y/
bWKzsSz0kaOcQLszIOiLE2vfJkZZvNA8E00fC2W/Ibmoy3Taxy4P1KVhT29P76ia9Re6jLnE4VvT
NLIrgRUohiMfJJovfQU9GBYdETrpVkcarSiD/dQZwGeY4efJIvskJH3nLuqmsYqCyL7lVz+Oy9ed
YWH4GUm6WuaB5njK3NYXvsoo2sRCDc1Fs1E9X/1bymBy1gfe7oTCH7p7ECPfEl0D5lXNna6oZlfk
oUQ+o8cSgpAV/P5m4j2GmV/Q3qBW1f0FKIWlHkHzZcw28JkfAYRNllJK2azWLWmd4PWejKxlassF
yaSAD8GO8m2qUWVWN7qOJYo6LeYZjd0/sltNxcWl3o/Ds60C9VWJ6fMJafCcIofTsekuLmGkEOE1
JQoZpm8RMAGCAkQleDoQ9+gMIkwwtw87SsNzzqI9sgMpMGeVxLSog/4hvElApFxB5loCkHya6nac
hIQkcOXWxrdjBruQjik2O0sdDiuBQeSlabP8AxxPdxRQsM9757JdLC1711bw/R+jdjz/Vtt7cJrT
VXVajZ0spv6aDfjqbYRQhPPCDta7iIQZrl10hUCpYeAlBHrTVerTnD5iIDDsRW2vP51Ia2JROIps
8HZ7HPX5LXSE2fLfzhBpHVJV11XSy3tXHHcbcIwCnG81pxaXLajy+0dCPO6do1FFObFlT7Xw+D/X
6WHCvGVd4LroZ1Javfv+u6ySZ8x7M1c6i5gnZHH9eVkInrCJG+Yuy2uMjxWvHALB699tUMUkByTo
79Wcu1+G/6A2OtSSUtxslK9Dwryj9KwVONoVaQPPUHX2D3r+K/4EkFXHYr/fUU8wnDKnn2ymD9oo
OYv09rLCiIaqX3GnDs/i8csqcuZcNYoCpX5HcWkR82Hkn/bOjb0uXE8M54qkjn+PaqCXJ1MqLM7C
5wK6tEz/MdEBr81e/CsejCYOK4MjUhrKJQTCEAUyUH8/AJcu05CcgnuL/YhsWK+Y8TT53JwIkuOc
mh+wLclVZ/nvC3O3TcHSFcOnz1D0ey4ROoSLVh4xQfDW7nHQuTocvyYnsLQ69GVZetSnLFgzHtLJ
62F7+iuuwwv6XCr0OgABDae84b73KXSoV16IYzAWJvxtDDsRxJK4Ucgh/4V8+q13D2waVKoajhA+
QHl+VpVBptAWK6tuOKHaQWwf7xHHY0lnWcfSjpctr21VJz5keHsku6r3l0CkCkyErnsMObnvMMYC
xYqY91EnCECnvypXvtavj2EurUOVSyr9wIyKVfx4/i2WV5P5tXuEqZ9hHui4urn1EBdy1ITFhvsr
xRALnhqYOn4LeHyLWOIIWjPmAp42H3v2ExHwmUGmHGxzE7ZGoGbYAgNdaFhb4bnbv/twXJPSmnJM
3JPgDTdIVfH2gHrPmZ6GniH0QoOIMc1c45y8orfkVNLf4Pn2QXFNb2s8ap2QA2Hf45VFO8N1AyMk
L8TbnVzBZ+cghq71Eahqa5G8dlxHuSLrOh3rf/D7jR0uu5TpLMZgHiK6n38rbx/s3btP36JBObh3
OKIt8Kht6mghI3wBkgZpcXIhJP1ckjbtdUcR4KADz/6zzK2GDK7eKMHA5fxdv+U/9wjstqiP+T/J
fXh4ubxfy3fgkXEbhhJ5cfIH15JiiTHbfOFGxVqiChE1qS6pe/gzmD2EVB336HgVJWjwEnHgzhCE
jgkXcBDFJAD5KYwvK52YnDtbLgef2ckNQN02OhFTsGOINghOg0uT8peUcoSGQ1AfyRzNwSDly+o8
WexZ2y+drVL7lkiMzUH/buNzTI7sYvxKLenqHrzhINgp8SkUa7st8n2nKsIqlWVt1kc5NqaApq9J
tcajMoJRDhBxjtkEA4r1phgKfpKAgXw38Afr0pRao8V1Y2bfLcZAzY14cBaaJjyma97U3m1DkCDf
azG0jUy3crOTAqSpZgTukYw4pgwoHuX0OYU+pCDVWUdl0roM1PACMfJAuKlF+SfwBGE5F2H7TzZS
1OtypHOlT1C2npccDjxm0JuJ5gLDn5WO+37yQNl8IvCK8i3W/vOrcRm8b8dOC12YEM1hbJbAAI2r
2iXO+6Mr4k4Oh5xntUQWMG/WFSHvOGUH4nljxrJ61uaQsd6K38o93VL/oq5WL9QVAB+zcHqOK0Kr
bQr1KPQrWlBSOEqlU1nu3iLypM/+XkZHqCvKsr2lig65dwclioMXc97QFmkgluWhLAk9S8mpSkCW
M3W7SLpD4GjGtR0UD2/mvI5GT1BgI6SjEQNYA99s+8EVpcmqWgQfGndbdDGt3FGMRqpKX5MXrOBo
EuTPDvEES43UyNvvPVNsORiz5mR2ulCu6lNCPuo47Woz1oQoCg/GYtRFduC7ShAfwzenuMmsgNMt
8YnSGxPWPEzpiCovC02PRbUk7JqDt7I7ZxTgJz+wyKDLLA80S41RBBlOKdM3kkl0EnAfly6Zw+Gv
0pNoRPzrVz+Ojd+Ll8mpEd5gR3oX4Id058+MmUcUQ5XumHmviWwCqmWbwzakFIKQHEui+X8napeY
wXT4cy6F1la+OfT+g42N8bfJXxv212vNMZ5Ub1xLTXuLiDGSHP6ObKSRnbz4s9zpaPN7zGg8tuLj
LrZxNwOzGJ5dYMOLH2mIDg8zs1g9eEKR/w3AFS+MlBOaDfpVXATj3pqXa8CesaXzrss60/6r4dDy
Vrt2tOsg+XPGtRTLQBPZ/BpZnJu/I5aEavb5XXeHjy/qtWa+n486mnyKPepmR4SwTFVApHuGXCvw
h+68IsY954MALVbMeAeBB/97qXMLUQfYjBUu9iH0LEuYCJnbJqvu8vSRr/+5qLgUvX8Z7oNu6hpj
QXN2GhqQngq0f5ipv+fS8dkBW53sBcHnXKzKgRkAOXacUXTNNTHvTm7Uos+mZQybtsxpk/UqzxGV
UxMJtsQgVOz00XgsHPQZKy/Zu4Fn2UV6Qam7ecy4Df01iiwGH6V7xsNfulc/gywCl46cosQe0cNH
6kcfdmqX5sxhwhp47TmgU6yFDzrjVM+u1mORk66lCN2mGuM8l0Rjz8BNzrCJftk3PD91xZ7jHprA
dTUtlUhUO3gdTe9i7mniMs+fz6G42bW925zAXsQ7pQScQ4u4h0w4cRvjVeJPJOgHxBbhD0wqBT5l
+wxVT2HkYEwCGXGzpUH0YVn7pHLqFDAt+vGJUDMzc86y5REHH7ccKXauhSwLYqdXizjLNQEDJGne
wuxzaD2xwh+72huMb5W/Pw3HNGZUXHy8J7HEFQNkYcstru8OfLuqtuWPu82CA3p8NRv8EGL7bxCh
lUZSrAEl9IcK3jgi0hycnaeATVjlagwZKFfCJn041KcqpXHEJh8zDKmPnM/hVt2zuvYGKqqcJelV
EOb5ao16L60GtzfuZrKqr8GNGeBqBEHHdP/k64EeTy2DRhiBXy1tPE6gDbAVVEFGnU6pqHQGuF6h
+Oqe7xK/DVgC0HBrRzYBAcj5M9n63bZxN3FFoeABOxo0bsnkpUHbhPKNlFib/IvYPg591/F3T2ZB
wnEloXPM0SVr5dkqVukOm1ezvWffGUfwzl0nuEqSIQdPsjq+iw/7PrvJ2ehJckEV8BHSAbpZwvQk
XdlH3KRP4gXDSzRB3lYuGKVjMpq68snYUly4XfcweeB1A2L/P/zKrCMxZl55j9k7KWVYcJxmkEou
nEew+9j04XMFnF9/xiepOsJC1Khee3/1g8GeXThqSBYhhyjeDMto6RV1hKmED4444w6x6ZjqYzA5
Cv8y85MFh3k+AJ7Agr+IpuPOASZQrBlHzfbOKAjluYlDhsULRqbSPV72UsBuc6cnwtpMlUDf4OJW
lQSmrqmrpGZGIdVneTjgSFFAd6D984Uvsq6c5SeoaHIJCFAq5/TiGVq/70rmW5eKZ6AWPoPvnB8E
uEH1tyQ0MnFWvf1cxP4uxT+FSQTdSlS0xeC2SBr2CsrijsNjMhqYmR7NBP9jFoHbBPIzfNrcV1kz
r7HTogQPQGonRPS+ymsUsFdEJt7kSjvph22E2aJF1QyDWC/XH/ZsgGOQ8z4j9qJtKN/vybHh2UNl
lod4G5An7JLEosiYghavqI1X2KGoeGt3EOHdPLt+drhTqEAbZZoOwOaD5WsQ388q4EDid7iVtXHs
pq/PQs84Wkeu5UltxH/nni3dqZaB5hvlRb4FhzS9DvvzWiX8I2w75CSngVKyvqBawjM+dlpC4Psz
e4FkIY1jLnQ8nl5fcQcIth6Fa6gTevRw9n27Kkb4WCamel2D2DJu5QNGnE6tiYfHisFy/Lvu/ZkE
eYDiYSbGQvcsw1MqxfoHCqh3w0X/U0enz6CDMiiQ3YDDzR5hjC+cZpG7H6Ai37qVLG7bHW7GizDt
1c/uB0sLNTzDpepAHPPTk5lQ2fPXVpziAf3+hGLFm7eSxbmrVFWISoKPJ+rqpnREwePqpaZLy/mB
Aw9Z7+bX5tSRDw7gpxUi9ZB7Je5mySqnjLYOpVQ/EHYVAuUKUJ69yR05IwD/Jf0XrD2bZ47iL8Ys
c8U08MLOA0IH1dIyJvY3zefaNaMSL4Y02AeZ8HvSMhzqb44R/+LqWP/Nl0Irq0Wb2d/+AXz46LFR
Pvwyp9PKOCWwx74/BtPxLiSfF13oPiNi7ogVDxxrKzpxsCR3euurjOmhQ0mRH+rChL+LCNVoOw1R
YCEox2f9oX5ljzczEUoalPD5KkhPWf2Zz6tX4NdJ6v/+vPfwvYswzYeyJQjGASK+v/SRiIgEBtPe
tfiAekr3ZfXDWmvGJO65d3Q5SZPgnmQ17ChNiL8mWFc7Rd3FL72rJsan1FLL5M4L7Tg4dsm3c/tH
sUAUSPTblthaTINSfzY3330jrC99+fiHHDAH+6aNz2BN6iFyLD2lMwdg8ZwL6nzwzaq7MwUbOO4e
fFbJNNxxywguz2jkt+dsilgxng500jGsJW5VCUuKV9lVnXq2brA2C0lku++i2NeMLWFcNQuQzq0Y
UXqAiOkt7oQl15PqpQRS0BI2V2GHclk2dfGM58H1azdbNIf5fsAyXC5luTkgmGwV1t8xqEcz/rsd
EvuXDTSpG1Qqdlu9DECH7goz8TXZ3GHQVlYaou3J8yRpg5YLcj4anw/jBpAbLu4MjKUYkik14OC9
KAVhp1gUk0sLcLfrc7Dr98+RYsNFfptnKNCSius64rA56E7+7kqbXwU3pDq5S5V+mR/KEfJDzU2Y
knMw3auKwTdtfZ2uszgzeb6fJHnuNgTNpOh66h6Ru029W5Xib5oG2tZcizn9Y21IuEVeU9eGlTWE
EoIgzblhaLc5mAudANC6zG6UqnJ2tBWtz73OToA3ElzWcdpcCZAcPo+Y1ph/xse+TkFyv14SbEyl
AQeJtGB1xRDdvym0zAireOtM5dsL6huUnGrsXK2h8FHHXspYR5AnGu+GDrVagHpEVHgSMqRMYHy0
pIf8Jh26wggTomcvp3GwznNj5RsOVt2gNgw61snRm3mAchLlDL1EY4rU2dHqaxkeZWGp2jFi3tNb
S15IA/KQO0FIz4tCCUh8uHWhH4Hw0gxxM12wLA2ozGo4aSxAUgXFEpkVkB0Kb9yK+t7uy/DP3QTJ
cWbapTms+/Li93iPj72K8wo+bSAC8BFsG2hDHIUtcVAH9RjGBm2UsFFRYKNuZlbWzOZfnyZZ7RBR
QniDPBHxj2MScHZSbWCXANIGif4iN1s/eFeVgKyN1zU+NtBx1GNnl3Yngfao0mAYcU0BelG+3WHX
UT1AM2UZxCTfpWfDEKBvA2sJJLpY7hSYKexEezrhuixGmLWFnuksSa7imi1VH2mKBnDQ91t5JkMb
wanZ92mNowhfQQ85/2Kwm51tFBBdrT3BGF63/sxYmnF7o0/0Ufs0nxG4xAeVPoX8iKA31htzvn/q
/HLUGlaLubeVhMCuiBVVz9Rcl54zB4klQictPdx4nuGlYtIlsLD57E4YZAYWmX68vuYEJSQbEmZl
reuFjsBX9bprgVdzcatrb06Xn5LVa7oiAmi6Yw4x0tSWofV2SDcdSDMC2Kr32/i8rCuW+nxYUGqs
NfieSHPs9vmjOCAvtJVb4HsDUK95Ra/lXkpjntdYTPADQ+lBXLeTeDgwwdVoYVaTObjiUlmGQU1t
7ggJLo9dnh4Q2sy/pImZQHJ0tlqauRgIJZA4z96ftmOrDoX3r7QHbXmwHQMywHXMtqJvTRDYERXi
r8SDV6DaDgHqIC8jyO8MppJ2YYMWFu8FuovIuay6rcNFTOr+THXYqGLX99YnOkHvwas2yajXz/JC
hcHuFj02THp5zxiEgcPKu+HSxoyjtzsjrpv6HFJJa5UE5Z4StSgZsUmMC4qmYaE9XAs+yBeP9ASV
S/S0sO8BrxyY8XfR3AH3Jq5b5tm2k9/f1vC+BZ/pl+r8LxVM2P0nU8UlAaoKcB5pI9MLspqpPTwu
VVkx79kj10x4BqhfiG5YoJCmRacaqTz1aRTZWwwMwaiIidDYel7PB77CDk4sx1XSvxUZ1GzkAKBh
NzJVbipn970NBxF03fpUKpeOudA+blQGX3OwYATeoQn56ZUzsih8NlI8Dan0Rft0q1MV2f6tMJG1
Hm8Sa93YxXXbuSUqQCork69/FkFgQgk8/PTl8OtaR4Iw68bcSbb1ot35AsDRyr5IMyz76fIfWCqt
8xPYPs/hwAAbHv7fvRiKhZXBpQyVXwu3cShZKewU3S03niPQyF8EECf1qmIted2ehUvTE+IwdKMe
rDbJFz7MExs6CUlnAb3cyRlK618ZfasXcMpfXiVbh/0VNoNlvo7njQN21tHEERQoBqbEH1vC1Wgh
hxtYPI0JqEe5KmeQoAb3udieZSMN/iGcmLUeanS3Oqcs7mNgy0jP2WvCcekKgYhSsl/B4xSL19po
wfFOmbRrhxTNpu95tlBOTDstf2ECpgeqiBljccnukzAv521ZSUZDawxwu+bXAqH2Ukc7mTX2ZYt0
cgwo+APCueP7UESABS5V2ax5fUoGxWNt+Dmnhw4+0Vkp1Uw4GAuJ7oJwv7P4ed3MzBTP6bvcYLem
6SP0/mW6Q5LDM79bnOJOZastiXVeiUOq3390dGtIua72ljNE+LSznw25gNvWim6ZzRnbDI3Kk+/y
cD9s9C/8uMaR6SXMBlCoO+qiy6jyfsevBWXCKE/uZgGl3JRQ2pxzAo9/qQCVClUilsLoaAseM2Y8
BwBKqABXrMWft1DfDmuyYHLTwq0gxTdHrr4B2mg+VE/k8umKcB9f2+vgRQ5D/CC9ad3hS1j4M+ei
xGLa5PFlf0IAZKt0ZRRLtose0nYPWL8w8GlXXP+suEAyxUzrGS3HOFHTRKc+a0JMico4T8m2TnK5
sfMW57QIUNUa/U2MEq3o6RzSJZ1FiF5qUb/viIdGkpVL/X3qYGzYPBNSgtLBR0ceP7ldtZMrPr1j
Sk3BV0bAlVwqJj2vVTNTvnxVaS9InRrvblvr0LRX98Kw1mMoREg64j5WtgG44E5iNhsAGBVCb/8w
sS8t922hbl6lyrw0O/Uiwtm7jj24gAtr8iE8Eoanapi4iUOLrI8Dmi1uFHhKKZJuM7clT0IYQbwm
t7pRJYDFIQA4qTQx5lb133fBQLBr3lvtVNl+tTnst9OjSszPlhDyHeWGcsce4/pICkO7XsQQ8L7h
q4g3MvvkwQamFOkDbQT4fLDtbtV1y6rtIAn1MT5HzoGCP8iwUnbQz5LTt18babFFHMJbx6MfLvOo
CrFhVKg2p0WpfPH1sDxGeZS/BlkQRFeugIViTTnZHSLvRlIpQiBk6Qv052nCTbHw1X0fN2s5W4b7
mxgEMgVmNPLJx7Z0HzB5WlYTQ/1U5/Y6c64qR9ZsW+Q6nEyovrrjqkGJGA+ywPpIEZNaCx8uZYbw
jYJyo1KNRUOFlyBOg6fofAAbvjo0EgBSb/00thZ5hDCB4D1ApqASKgzyoyTuESzxZ4+BQdRVoEtn
JvhzY14MWlsBGcy3FlF1GuFHjJro6llbCelBYgYqBXGK3mHZpiXHbkZ3xda+5ZJ+tTelZi6mIPVM
i8eAN+qZUYkAV/T6K84tdfTmqChDqV/2FvmvlUv8TEJSo69KHADOwblZfVILw9pV8QkyxhAVo4Oj
jMRGaCowDe2BCFUaHR+ksFMDhFqeKgtg7h7ZeuTCfmM/neTnA87A4q3ih2iKhZfU5C+1LJiNIwmo
a9N/PFPosMJxsz/u5D1TwJXt4JeAFNSO7HQmfTXI8YOw47+DntHPcwAKjVWiyqKysq+1Plp+y1Ul
QqkzyCo7eNmS88H35G8nyCBdT86h2kO7reIO0SJP63PnD6yQWexjPxsHP1WZzq86LEluDyMrmXpR
RhlB1w6hNs/Z4yzjimUeBKj2D0Ks//7YI/mfIDZ3l95e8d7Pi2TaL36IE22Su5qlSjK5A3VqsEMl
+XrIamQ6xWlM/m0l95Dew5KKjtiHvD1XQSc7tXrGe2lHAyNz4KisnVxxs7a/HjbKRMG+zDP0lIkY
IxvrKgWB1I1u0yXyMr5jg7BWuKOzGNVmbfzTlZ711fog6v+hJOVuPokXwk40oaZagh4ij76oqyrG
LtYyyUYGYhtmYliW2j4SiJ63swc33BDzR5CNUO4K6olMNsoxxjUMBJOd9OkLoGWLDGDOU4OUyVgS
5I2CJPcWOvLea5kuKmeAcoKoMGTBz5y0G8qeBQox0sDASWvOr9tK02ZAzZxM9NjRyGBBunr+YHo/
E8LSpcKzDh2X9EK45Gi7W2m+mIwbiuonhOYtRuK/sLBBsTYw9bAqP3JfJIOBxkifly0LITbTzv/S
9Pc4g6ptN7xtmH/anfjTkrr/hDjH0PhtzxzfkVg6T64Y1BmwdRCdrHSWRsvNdjBNdh8/sLCYtIZo
JWn1A0RFsGjRAPvJdjEHUs259nTWBfHWEZGdLaHXkL7O3LAUldes+KpBSUe/SkmEj/oabDB9emgK
X9ivwsFh5YKDJlPuwm6kFMa/Rf9uToBRDrLaJlbFgTeg6v4cfAOwYMAu4o3TWg8tsxhnTTMBveVy
wLP2MFcJcp6WhuynnO2AISFv5BsF88rNeJlBvYOhx9tYtvSMS5tZyT6kmuEokDh/kANHqUU6dnje
ocn35VjBV80YcFloW/+e2iSqUbR/Lf9y7nriInouLpmOhcSu3pkB8+0yqWUjgyKLwNAYgTUESsNO
5fCF97Hr7v9PUFQGp+mcnKwQq0bk397DusHAXwBlNk0kewrkBlv81PJAH/9Vdr7v5phzHcrJkSFA
c1X4Pnv6glct1irlJCwMaNOErZ9RVz5+vv3OgAayhe1vTeTvAwh83F8pc2cgLozeWOzfqKyKeJ23
H+DZwebRgn6o/JUfFtOwwnvJsaPWkoErf35czbUzJpCZBLdFq1xODbvk0yNp5+0Wd/mUHbPwDMKA
bCBa7CcBcuTevZFulo0omHcTMZ9Ug1QTKXKP5LLE7HM949DnCq6hZv8Z4sShrSdEF8kfAEZdBTFw
BSl6stYwECgQ117EOK7Q6Lsi8X09cL9yYthpkgdKaoHFr81daElMgv2QxAQPMd3sThsg2EYxfP+G
LxQDSd46GPpFdA8N16E3EOTDNd91pZ6mZA8xYx3wc0lfuaZ20pYJAKjrVt4KpYnLvx3mWnZwz9Hz
zyxE/ZINhpbVQ9rsQsbKPDYHQ/8jP9+K9oJ+a9RfvuRQ1RceteRI//i7HcFgWh50Ky1lm9ofvRUf
ia65NuRdUTItLnDw2z080Anvt8JRrXEKr1PdytEXD8nw3yQscDHU5yuAvs+aA5PmESZFEkZ4EUVn
E/rWnKW2kxPGo3mEZ12RkLcSL9PCAt/0qfQ/W09w5cRp1SE3qjm8baVeODN0GIChnt3cUvYfY5JR
LWOwEiTuZDml6M586uZ9SyuSgqLvT9z4SkdK7/U8td97gYBeAzPc64U2hGUVQOlqx7oKC5p5fATJ
jEwi62BW70K0Q96vd/cmrDp8kERTeBfgUhQD0RY663bXq7LysBrVh7GqbQ9ChgyfCvkCfyF4aB3u
vMEFQ1wYOwtvpiop6sYVGjsW/VaH6dZtnNxBBarsTW+3n1DUg+6t/CqJUjAOn981Cri1eA6ZaC06
Z1TInmRVszS4zI+TZCT1eRXtQ6Kye/zED1+E3N0YIBfBnChkBFaKIonAS5E8MPQO+UZ+jzukIg7z
yAiDc8qiDc8b2HSyiKmo7bgc0p/SsRqaVZ89Ig+qRHZ47z+G8r2z1Ncy7ExvPuHS6WZzr4FWRoRS
mIwKqcCG+zZ5vafhRPU/86BQ8OWteIz/zLl7cCWRYVLz5hUcjWLtb4HROL2yMwOLv+2HEHcfwTO7
7/nLQLMKSvwy901HT06G0IwEAZzzpmj03tYzWffM+/++SMPSRUtVCfKAAAGuIUFEkr2L2B0hHRBn
I75+NWzah6W7zAKc/UXOrhnutHdgqqWlvCi7v5NMGEhibGWY158kWm1XM54pJfaX+G2CA9TIMQHa
NkNoWsSAJnijfQ+Fq5Ve2x9YGE4svklfXH/ECJ8zZKE0af7P1BkV8eRNunHLEtTllNTc0SKuSmqk
A4jybodfILMVsXPcgbjYjN+n55irv1HisDM+8G5Eh0l+Zu0nByh9bXn+X9gMftYzumEc0ogM9s8M
M0nNB5JX/29Y9BS/kCSED8n1lR71FO/7fIFJaGSDuEGsQgaPAs1rEBIqyE8C1e5UmQJ58OpZVXtd
bdVWzzbZpT54ZW5mNx22CKn+Gp7mvm9T7+opDD1GezENBSWSgrw6NDhCxlAkupX9gXU9FAIBLjOV
Kt+jEooQulPbZKhi+MA9AzwXayhda2jRJTxA0uOv8qufXPo4NYXyPS3Pils16NOwyAGpmHueSRMK
0xABrJZVNQbs9A03YT4rk4EXXckvIqNkBBn/Cl03n5VcyYuzbcYA+vNl0XaQILryutA1QZgGlUIS
cQwPSZP2Dxvol3Ha6rmIztoz8VEaY5kNCRShUUh1pkMMwv0Pfv+n2QLkDYTFDJyA7cTAbc9nQdtg
9xAzwgLb++8eh+gMB9qxilpo2GIr9Py8dBJ2QkC/Mrt7hjJyk54auoJFNl3SY0OReRPSjxVJClBh
FhX/6O4vtYT5Yvaq6VnBx422dsE7sbTT0Cm3A7PKBuCNHmrtrwKYP9Q6oLOzEwTQyyY6PKVCh/QD
jAx+YP8vQzbUwZCLByTWeyBVcz2b8QCm2AjUVpwaC8a0e1lqLRowm7QyJjzkGVf0xzsg+N91UBJx
3WxPwJcuQwXuWQDSaMOR2z2tkhk/NEmTG/0COetuQndCfdLSO2iTLf7fgDubA+YgtFj8xJQJ0sZd
yhSx6oozwUtmhq1AVqjSDMR/com4S07OYiE1yHvmmm5eeB9XBFvNJ69tfEYwDgK2EwNEI+oSczV2
3+5DBu0ymJC9T2aCtyfK40+RP3c530MS4VDvgE51ZP+6i8nK5UTSozHJnZO2mA7MqB5//giYnT84
O/9a2ZmuMZWzlp3r2HmHXcnoe4Hu2A/N+q4BLLCYnOL3wLcexEQgndCrYFD2Cx2TOkGEDgroS1i0
Q7pfe+OcM1pb6ZeRtSiSRZI8UQmAhpfmqJoeq27R6/R01AUPqxon7HrPpxYJJ3ee+RQS8v9onVvY
vOeEcxJAttGEFlV0Ltvrr687yc+7M1d5AxGsNVhup1armYV85XcICqfiRNcqtU2dMo+tJlNgOf0Z
iV9xFXvacE8xb2YRMHxSaWLnUzVcCv13KWhV5uQJkyigMFrKg0UzHTl9k1Qd5wLmbA0sHVHyyhjg
81+SR3FhfrtiQatW78S+jyGuJq0W8YDlBE0ujVTnZa4BN25HUnOzjkUl99yks+4ACwMidCxa1+gn
DRh1VpjpjRWIgbdWIse5V5nITYe/2p7wo+cneENgns89fiI4IltnYoRjEeEYIktanF4qostm6r6M
8dOH8wWHSX14oDUnFy1HIEmnozyetNZ/6b3WRv+3xlvNZKZ4BZUspHp38DaQGixEdsHlGr5ab8ZA
XzPPUZv6Z2PGuiUKmkvAg26H4MmsADMf7Rxaa8ES8MEKmpAgQ9U/GFpKdEqXnU1scvDzWt9S2hsT
jdQeDq2ZraWjwwOz3+1xTxKwgQbVmrlGphd0jqRW+NUbQx1/UMckU/IXGo7pmiorRPUzUqyl7rOP
RJS3ShiWy04N3Xme0IDQUHJlzcqx9cmXClvVJhrcx1pB535mTpVfLSdDuhv9viWCWvn5PDvfHaDL
5yxQpHse2JKCgX3ATiyVSwfvjnv9+Jd7EErnTmkdf/CJlJ3Mx9IA/ZZLYiVQyRbF2Kefrv3DzQm7
xwv11uRtahLhVcLZqOffSOnCVM1K/703nP40O+60y3QS+KLfUx0sQviY+EAeausCiJtXrl+4dKYd
Xj8iSzqgutJsJ8IBJG27D7pfLHFAe36lxp3vSo4rMPI6zLbnbkdA85ps5W2KGOT8RcuuOg6dlkOe
lm6+esspNM56GxK2SHmdIsXGUyJ1NVyO8//GBaw6mIqkEtzfQelgzrJxVdDQpF0xRfjeftTaFf7+
okiCjOqkMdg/kzaLLdTi3OPYk9xAwDOE2Acljsmq3F9f8NIHnd96DFZujk6S6vnplALOnas3VDFr
RVpY/SIbmkZgfvrwwB9BpupA/3zFld3QzhXotSfoXVCz6cyKiYwM94dn30PJNczCQRw7yiMtxCDv
yYpbMKLN5WYkBivQGKET5cWpCzpCu+vQGHjLB8S3LqahX31wZ2RS40YZLpK3xsaXoQ/YWysOHxYt
LJEXRJ4MX+5Qh6wcV2wm7ZJTs4MsBQacwmU5r2bvf0lRtbS8urwbULOs9zGNuKpzznRgKlkqaSGM
/0YAfc90RLPJSta0Ov1jXzZlv5ebmFcfsRl0s4ZjfTZVWaxYj3Vcy71xLKp5GPwMzyOgNG/f7D72
ChD+Q5ET44VZt1fog7/Vb6lN5GtW9kejl7y0cVuZtMyUCy3kgADPVB+dPogv+6ZzWSlZ54gNvihG
552VqVyCBv/+1+RPj7fJh9IN2gQN1nz0Wcg0VZ/wO6BoWRBINiFeMIDJ1JI76yUy5hPi1c9tIfyX
CIev9QnMuJEUbiDIJEVF7iRTiw0CYzaMfip2WIT0jnrrBJk5USu3lOWzWpMdJzFkp+MHO8u7Cew8
wfL7Kli05Cnr/ClGHDlkIHpzFeRJxFMk76bs1oGCpQc9muat3Mcyk6bO7i0smtUU53Neqnopnrws
Bn1SG4yPMPb/4s7Y1697snRtk6pdfkbTtXCvkyC4s4vRteP4if22QIB/oIE/1lofphQFQQUKtBHi
U5pDK7SuFvofU5HJdzrkb/QIhvMrQoSBjvUDjXthiOm48hmDQfVlqu9+Sg6gfPi1LMrCL88/fzxK
MLFyGX3wFxWmK9JSEquOWbIWKamhmWqzu7j0NT4YPoicfEqzMc/9nfOYz6xm3L9McPvjBPN9YPRE
8+9E9zAzb1bo9k9TT6i5Ag14ZFjySvQqGX2cpd53zSwByu4GmAZCVdeH+5jhE9cNmVuOddb1fCFF
jWvi8QnZg4d6N0ffQACP6thy5Ejitact1iWDrolFW1VFk/jnX2w06kusvNR78420zaN93I43gLs0
G6VdW+PnIvTMGJ0H0rXJXdYM7UY+H0suHLMnN1/TYLvqZXmo3l9U5rxNg/0IgOr4snrA3TLcBq2Z
pX7siyeNfeANOONSl5Xa+G8iQzqezMQiSbFqFnGizbsxHnUnFEk+rYFACsZrnKbXmFJaYNr14Ecx
XiVHx7486uWTryiuhWfwkzuBzevmBpRny/sIqoxLax+y9RNvtTXqlkiiiYYbWBWf+MUerXO0j2td
VGrFL+vV81a6IYUsynOKgWE8EO6beyFWytp7ADn8Nu1/PvpAVuASoQJ3FvOr1naqurDOQHCf5WFm
c/TAVf/40wZPqUzTI7pd+4/IyQ6DdA+cNCfd7y7PeFDCAOZoCw0orj25jsMF93pKC9ZGpabXDk60
es6PNAjp3kBFGkHrJZBkMA6tP0Hh1D89dKi2hm9NrG7U4N+FZzicbT6c+NVAAtvhZD4cPBXw1MVu
MGSHBpXJcr3467H5N+AVtj+NzqmJH1t22tu2Z2LX0gwEBZ8160HVzKVseJGZAD5fpbxh/b331gp0
sB+l/ppVMO5W/ZrYn9vHDKZmlCPZ5vfcR9PgIudrFSzCkLeDJUMV3hmiAUOHb7I9HAVT7DPnK5Oh
iZCWzRWcWdU+x0qsGt0Ub4a399HxwxWS0znb6m1tjG9yuvNOTQ/N1r2aNXCBSAiF6IPHqFbLzmWD
hlBzCkeuKNkFwhdOXQpGuVgK7mnr0cvGpGI5od4qbS/82O/k1n+VuibcgSMfHVv2TpH1ZoSVPRXj
eml9CH6MeLWtWjkDYEuC8CgDQvOfbQIUiWyqlUDxAyCmDPIr72ThIQdJc0cwFJ0PYXFhRTliRacJ
UPNkKxzfgEuUqKAQZevh0yexuMYteQdoo6XpGxqJuJDFAgAAoExHNJv2ptIOG0aolR26ZknKl1h8
kJYdCpo3uv6yHtnRABgqvcGMVuBb9xMu7BvJMCncl5otTXLI53YohIGdpN/n3CAWUV3GBC8SZ3RI
mgkNHb5Rz1F8b+CCXCDALIR+zPmImv3TgSLeETTe49QCivwA5J7Ce8GQzQm1gfZVssPRzrKcV4a/
ViYGTE9eOJGF3HIZyWfkXjEMaqKok1pFg1vjQzMborE45kKpIetBWlAbTIgEd5HEvIE/vpctci2G
M0zSepNikdGkMXqldtL9QQQtYqsBtuLvmdzRWUHoMRDGbPJCn1Iug9GgmcbO2QB36N/+sKxeH3g3
5IMlHOjdAJORodfkcGKLUhkGzBKr/3ATyvvqPRPWM9swHTGnX1/fTP3Lg72C4J14k3e2RCGP4Man
4GPASfd/yJ49b+o12G+mxmiK4Ul8nOVnNArXjCGtZEXOZdW+sMbMF3UEMT7naLxCtNXaa7jVJVKp
AbEiBe3MBUJ3FK9kMmughmpxa1CpE7QWDI/3P02JMFoiG3O73vZ3F19yP7+gFoHm/AXY5DsliuDk
tPWDgFEoGU52x3uezT380yayaNP0AXM6oqxEGddl8679BVveXzPZXpMhSwHMvXISRD13szgIvrfl
ZNaFcyDlCiVf62rimFtYYTu3Wzve/I2jXOHmYprIwggiX8dDcAVhO7cf3Z5w2JX4eDs9fyA9Bhr3
wLjskRrpMbOQKcMCng5TcFkjp+wJ1okhvIILHogivDt8Ezyb86SaEvDIMI9ssBwDf6LSl6a7SOAV
uoYHKaflxUcUAKLDXSr4VDhZE8gFpbbLcjqrd3TXsnAVTMLA3rVcRfs+75O7TCURwej4Tt/THCyy
4vpLqsf6ulj+Oh5QYRNPf212cAZRwSjouL8dDxS7CkXars3bsH6ygs8pRGunp3umHSaGKTsxGsN+
7AAQ3msd1xvjLd5IGIOjEdhMnV0LCZNeXixykP5XbuKg1POwKU1od5AdS6wptRagX+GV9JjJAjfg
ZZzSYKO3p4t+yurWjHesi0FONm4G4+SrtEluWG0Fpjx9fuKRJWOaHugsCUhwI23lS/iOs7sqcGdN
842fpp2/VzEwmhYzgLhpeMmec9gUGoOQ0ljoCrd0KdKhgUdq7bpHsceyJ7RmBmMQFMVxTGnErjaG
SePsQFzit6Prmga6FLRVO8NLgkXm7NZfu1c8Zd3QYApS72ROaPpA4IusySli75hQvxa54bnjOVGS
9eq4GykF7NhLnHUm5Yd2I8n1o9ap+GkvNdl0dnWsENmIAyGj9cs3JB51Ooq85simcA/ro5tF4qiY
yU0vuHBGkuGGxFdHpCvbPkLxCBeCAGjoFyn0xJXcL7pS8Pw1JNMWP/RZXiHrUMpUudFq46dnKueq
Jhu5atoiiHuCw+dN1AT7wBrDa2xGuMZYEfrZwqlDMaHHvDZz8DgzDUB2JMFxVLblJjzqbLn6jifJ
SqFTYv1SW9vrsf4DLfyi7csUfu82wKihtrGcUK1/bYNslIWm+t44fbOOqlXHHPc5V9cyDz6vbdrB
oTxwM3kbIEv/AsYQDp0iser26/u/uFSf3JGKVOEsFM3vjkV1grc/bqXeGFyAhSB7C5cWAJO6KYnb
bNnlefjrwg1kVZz/zLWSPIQBV3Aw/rCnhDqEkLhB7S3YKB4JLVIchGYR3vqk0sG+g5PwweAXz9Qv
w4XYJBoSjt/fJmlyMGOjHQzVU4now2PBOt0nXX2C2sFo5dbkj2F/K+BfLmbufFHtBw9Lgt0/AbIP
Z75rVdy4+wFHmr/G8GxjBHmQWxYIiAm+JGONC02Pzu8Lxy3rx+baA+Ry8BERI4AungwwXeHO6Y1m
s80AeJpwSctNkBbkCvJ6Bv4ocC21zxl4Pt9AUKXidqYscw4w721aD4MQyphKfi7U0+VmcdZBcHIP
fiIlP3rKkd0yrmh/WOqeOjVptIYfZTUlNzjwFJzQ9ZRO6cUlvEab/OwVzjzQkCTS/qvEVKYPm288
/48GH1ZDbiJeeUH32zjSIFXBFWTLYwdQaLR9LqgN/CEfaugjCC54iTABo0P334hJ9cWnyGTUba9d
M37sEDjdxwa5d9kMdTCeBE3E+KKqhn76Qv/ysqv2VXJ5LAmAxr5Ihl53Xodmtn2ZiXJajP/WLC/9
wWxtHho6CuywZrroLEADJvw4UvuIMZvnl36N1498sErGNtsmFKOSPGwpxqbenLCPD13lfliOUJGP
6aikGPUjwp7N8yoMyy479Xs4klsz376Hd1o7+/uJU/YSmBPWm/PRM7Uyzlsk+1Qus0e0XWM+fEtV
Ru+EIjmNPBEWOEX9zPhTXkciv1bbQxktyH0DxjUFpa1ZTyzDoc8fzqnb4HtNH/xbd1sIIyyOy+21
4LkST3kLj7PkVC6syRHBGSNzRpT90PdiEAlOzefyTNR7m8UrZjbVWk4arKTtFQsAfJBmY58RiPWA
kW1D+GQk3rkIoLfV92v3vu/FFM/Ni0lgUQOxSEx96B/rUgjaNfPcobHH4/KY1Qa+0oMHukEUT/JZ
tuRT/+2VXFtHXOPf2CpzZQ9FSuwxh9Z/yCwpjitOAMMO6DQJ8I8kIetqne6I+TQ0nVYOmUwn97Hu
aDFhIkVsFqVdgsHiBtDq33/H79d2Y/yJYCEZ6rFVbW66foFmGbsmQL+v0Vz1PPVb5r8GiUmhab6D
rniLjlZ8rSICxApxd2yxveo3enoTv1vR+s2HLlCa3/XKPvQYxYvqGix46Yf7tbC3AkOA0vQ2tR/P
OT1/va9+ORE14Ebh0YlsLkDRVXb3IlruPHZ/2XeqpYqE6oGWXUS75iXLddvffl1iTuEt3vO/c6O4
ovQ22R9BIgH63pIg/9PYqvggEeuklsCvnyjr59To0StwdsxYc2JDOXTWFbfK6I4mzCPnttBdE/TT
VC6XJn7qcozM4e8P5F4q5fK1iW13e9Gm6XwejJSuu825drw3a8T7/si8t4qWDXbAkMKjc9Mr7/Bt
HIhUGukqzwEkM41vFKF93Gvu4AbvR42+EnGfAMk6uIkLFWR0z16KsDe1lVP/VBrWKbmF+gn1+yGH
029ppkxrpb+2NR9Uq66EmrUN7JjiU3B2os9m15DQehDYTqavwsfFt4LmsMm6OgeIQYRBAnTYd9v/
jb2WNF8nPq+oRLV/XH/RCLCh9Un2kP/cbUoAMNHwk31v1BhQaLLvrfT+Gs+wHYPshvhu1J0L1eHD
NLqaI9RH74xlj8hSENC3APpBQ4YRiRaFeBnPw3T32mkBhKgnXNtBoGn+RheqIuAhmv6mXU1IAUB/
aGsujOQ+p/HnjakUZ+tqkVK96hx3x+3keqrDqSvrYAC1XHRrPEy/JNIcAWt1l2aDyZlt7IpZwOyF
kIfF+wNChTuxZbIYLGWBo3QqXoe7ds+gk934c3a+TaKySZdR2oFc+xb0ec6V3n3ofuZrX7hOB1Pt
3n/+IMv3ZonJeVX3AJAT3Kx157QoMGao+qFbCc2IEqHaQjlMk8oVySCc+CuSfamWDFL4pPfAifSu
uhagOV0v5aZ5M0FDSfsUR9gTwnUerrw41CB1/tWteAM7vQ2YOOc7nu8qbuPXcDVpEkAjtVCLUV1Z
UMSa7A7oTSfs21qYtUpyL3L71szFCwaggIDhdh3Pf+Jput5QX4hf4Z5D0iK2GEN4Ei4Bblfwc3wD
Q2wwnnkgCYilJNALYqFOVH9k75DkdTLgawdxDYr14+vB7WiXUWGTSEWQcRLilabIpFuJKTdbfNfV
uvMIcYh7QTLVi13nRQYzUMVImyBtVPF7c0swCBqqJDkA12W5g4xoRmSbi1O0NahS3YF80LomRBnb
yS54byI6YNnWs1Ct/7jwC915DqNYYrKcrdOMoY0fl8ppet3FPjnw/XPxFVP0T0aqkzvA6D7npgEy
jXlBjGkJIybwJeYyU3aystRHbguL/HIG2hJnQ4UMdcy3DqVAUMOWJ93Raa+CmgcsyMmwXpJvCtVO
1pf2RScS1uLsp0H/lSohH9DZcch5FPUWUwfGUeXv+o2vqLPnAMXor6wO1vOeq7rgLCICCcIoQpL3
j7+1TksqYlRCMXF9RMm4gxmt1B7xmsYIhvkEnAFZjb7GORSTfVX2+ko87eJfJ7NpygGXCpZqosdB
uYmRCCDRxIMVUsM60zKK11dFZtIW3N6SoHvVqwN2dL2PWtthiSSJ33FWpcpu8OOKJo8dbbolNcMx
CYcBvfIedeY4S+Yhlh76175W/mMrT9imA98G/UTNHrKgjU/NwRrsaWFeTlyvkZqprwG8zaACWCMF
qvzyTThSXGtVRcpJLoUK9QFPiHr4FY/zd4x8u/B1VsKMViBImmAMAz+z4bL9AQptpOJ8mYW5IUUV
PyxjOcvqkPdpcyzwONn7JCRP4Yu6HTRXvrUY2jY6SQyawbi1xJBfGBXfZluAvhcX1S5Cwxr2ul7+
MN7V9p8iUStsG4u4f7OZNxdHB2AD51WNc6i/25+jlBxZi+eluLrtfdZM0EheCFaB81JOvCd9kSvC
4MzrrzceJn4rScw1ojDASnyz9XjlMXpwYhp1W51cHvACdK8gQFUQHTHrAVd7XzCR7mL+QPzGtS33
+gRYsdFkefQX61Gn6OSeR3PkpcBbAoBlm9gFjFAofEhv6mb2HpR42Fakw4XIQf0FLj4k+XYWMwFi
7t/cG06qLanPFhym/vr5eHFnDzbbQLF6gyNH53edTqnsYnL9Bglwhr0ShyXVvvvlTnKQC5RRM7On
TWEQ1L5vAZCZVK1IQzDnAxC3Pt12FPKPZz+CMamdwb9fHxhzZDj+JUw256t0vlQWwbzOpxaeu0Gb
WqRsHtT6i4WvFiHIa/tXMKTQdKPP5sOSZrmeQn+8Id3Hubt5Icz59qKNYePGSDTej5TIk+1PIT4t
tTXQ1QgBqSyfbfEOxCnxnIgstzX4jBZDeovBGIO0h4fpkAuV4SIt5G18fDiEJQ7d562mb2OAgFwz
gCqynGcJ6TrYoFY0O5oqPIiqpGIegu/4SUTzQ+JjHYFuIqp+XKVVvikakvhYRsKuNm3dyJfzfF2g
YryCUXtNZHWUgnF6wYiQ/mM5gaoFxQTjeSCblWTmnRMxQKPA0WG6lqZt52FUCNlvkKderJjMunQw
Ac28Cp6ZdqwGkxDwFLouTsRHF8rtfrrKW12eQUC/xotDGmPKX7jH6bgZTizUjPXGfW6uNIrW0MJ/
l244hPiWdiCZtWDgqXOjajhGEJu11yW1m8SgfSajYVYRcvVUlBu/mI1RD12P/NVsIEj3A3HpLe18
prJ/8w0cH9Tqj7OVoPfCHdUYlEFg+hp2Hvo0WyxkI74F91QVcTtmmw6ybIcwpsqc4KzOgNBW/1dn
gtKdjjwjwiph0YqX3W9UgPB//l+GSZPB/LhPMMTk3hXmXHn/z8wv0ovSlrlDY6/B1V13gg3RDJ36
mx+84gPoffD5Zb3puuFrGxxhTWNrYwkojRqZhznCeX6zlD46uF3SqatVCzgGJ+Sk8Ai5Go4vdt5r
ywePrWy9U4JMwdkQNUy0OQO9ccf6l6Kze/tuBqSW2GMTz5UZWBl0mzZNo8rx0dxlgu8a4V1kp0qU
4qWFJsHqwr0jViD2hdbdBJxsTnkeHDyzyMmc6RNOj5lx3V3CN0bLHp41v6E2oVPrz38qwfXPrnhD
I5z4BurvMVDiPJYyzho1AsRUGhfO0n6hwgOUnQHzF3P+EaziSOjBg0zaNeI2YMBSo7IBEM5eiDR3
S+AaK6FBf3LnPHfw2YEbmnhHbWUgtsR3E/jh2iOCHofb11xylQbN0zDzC2o/DAH3UxU2REVcRFxv
rqD5pU3Zp8a8RMUL1qAfkc8D63R47EFDIebksszHoRJ82US9JORv2T1T9I5ENiVAyvMRxUJLBcqt
RB+u4mYXH3ku85Y8Wk3Eb/PjUZvSZ2aM+ih6XCN977PACDvN4gOYL93lo5zsTdXX6uaewx9G6TS3
FRQSFUXko+fpiQinv2ADLZXJTL+pe5IT0EuTAaMDQt24hDHt/UEqvqMRMk4VHTKwdsO56hvmTSJH
kzYAVynzj+e4VU+3wRI9eRayCB0MVsRIU/LgDcF9SdjVBjIUHRO6i3AnSkZQvxP0dlnMRrB5akyh
gXY+gKwBOXT4/SnFnmm4yRc9foZZOlW+W5WGx+8uW/bMbQMTNFHKF0BvCh9FWVQkKt4qEZHtoZZZ
EhH531X+ZMWTry1nVZhTZbRzUh+AoNIJR78PblYLKkCNx1kUDyZ/Vd4v76LDjMQewvzmgHTx1O4W
zti0K1MprzrkTRvA6+rWJs5WF6b9mZTTYppMRM/FGFTLcsYlOpH4F7HBmKWatVjn+yc1RsD+j6JF
wr6Dn+d1PCpJsYgFRDDSegWMwcofu+iUZaZMfBflms2/6wuqwrPWuFZXQBvOTnXZu0As3qbVMdBl
a44RqFEshfYH0AElgl379yVwAbYfqDEYt2iUjE2uB4+RcGCSyAlC35Cr8J0P3WzuPJtbK4jCagPv
laMWLlfzzvcPLs344I2kJERD8bceGwsLbRhq8QTOQVQWAvubD+XQ9Vkia1RXk+uTtb1UPsiUKFW8
czq5FFck8IRGqVqiNmb6MLM8FN6RQEIBGpUdzRx1aYtEhUGa7WLh54oV1E+9xWU//jDmxtAm0dhK
CzqIfKiWufMiWEYsJELcPl2VUtOzWkOd6UMNklF9bMC0hbM+pNgggjoe1DjjDkF0NNyzo3nOYiGH
dvu24Xl0kj6Fe3zpPS+NhmVyxQ+lolxkAzZvmzvCEkFSQSuktB8wMklRy6qztKj/9eix2/Xcxsgy
Hqr/9NqGldcvBuQSPc3bRAIp3cc9XmfI63P7MjG75QP3iyCHzSbrgfdYX/10iK8ZBtKkitA3GedH
tcB/UOeIFkWH0kh+mk5ZXyh0q3lIZw1k69wNxW/72oai15mLR+RZJ1gIGIFw8OZdvhJIGYJkzi25
zJmH9Qn4wCslmctMeM+tecCwd1uffqRJGtmrlY2P0vxKtX5k9jo7MCfFJE8Wrae6Be+FQ7Jssq0V
mZaXec/IYKfnKivCNu135o+6pBRidCBhmRxoE0u/R24pgz7tUuesuBnK+gYJIM8HPEA0v3l+XQVW
uwoin0dQxo6qo/j1bx1aa3F/NFXVXn6qloCkHQOIJDRWpkykJ145slDAjKCiLPy8XpFO7yvQyOOR
mDf0T2d14V5e+WkbB+XTmQKplSBFRYYBRvgwTaWqeKQ6IuFW6NxkycUaeCpm/+Z7vjdO32kmEgEC
xxT/u3uJkvR1fhvg1q6MbhGNBhZ6wHUz7ebfRa1o1SiKrpI4fdg7F1XHLqQk2toOzD/557CGZF28
NAGyNPN4M7q9bYNwkNd3q2vifFTTC6boVtREvPLIDIImra3a75qdQxgc8lHKswxOFtlI1vJf7RXe
+iI5XtC+Jk3bOFzjKywbcSPZ3ygfmojheWksdhOXSwfBwqp0AnHqpsOluKuBArAbP8kz6wpTx+PR
lm2pV1mvnhGffid1CaCNztIFR/n2amyr2ZBSaQdIQcJaXEsGAP4Risz/hR9YFv8HxHqi3bpeyTmZ
qyciSWR0aGWBThPb8fgsav04wSCcTzov5294GcS6qap9h1BcOUkSfctgrJFbHVkzyTW4fISeOav9
/Ig5bVyZM3zQOAn2napTDyzSQXMcSbfwUthtsUWVytV0QGxZSWjjv9S7ny3eV/sxSukisVaNcMUg
7UfbOEkRUniIEA1q7lWo/wdTjBYybyJ2NZ2H5bkPhsW/Jy6tHFtLDtud7JNeY351Ph8OCd2JpTwv
aXM7s2F9RRUnuP5gnQHDeomiMetUVMe/cEQ05xwsW/UMIngxtu7kVfnYuoPgogFF4uKtJLjCqjD+
F2hyd1j9thv+Fzh7uIUPmn3Hlliydb5xjb29/pJY6XjUokpMvOXajrzaqamgeF/nHmDo+J6iykmp
KFt+VHkDwDWGF/5naCEAUuCyrQ2YKSpnA0U06CTCgRWltW50OVXfHeP5hAjPqB7pxzItDbktXDVB
StOL/yjEGlWbqZ98eKHj5gZbExf7fGo5fIz42fibhmejaxb5dCX3/wwVYgo+b8mi9F2ttUX8dXGW
7GHqhzTDxVIKJfsbtC+hTvb9vZcfSb+RynfVVykrFAW6ZeYcxEbYe6IQjYoR+rxx9Ndl3wlm9Hzr
u4DLc8/7gm40Cu5gEtC2RGKbBelkQzVjvKIvw/wNUpoVFVlfPxzJs/zeXQuUxlMvS9rnBNRcezWH
pVpUbO9TN1JL72fzCUksO7d/WKNVOWhYbUJCmBo/0mJeN6ly7QxjQIhKeA7Uo2P4tYOB0pveec1y
qvNq4AsDi1YGOpoMMegESb6b3B42oJdtJufvdwEW5itqg7wnjU+nGVn6BGb0EoTN+kxyKJak5tGO
nRNTwmKRS1NyeaCafcdPuSwEoCgDQM0HQsJ6d7iR8RRbseKpITIv0dhr/B21iPeFn73p8XFQpUkv
WVam4Mbz2nAaNTtwAGm/Obu0En9tHdzaNYqWpPZSpSfkF9DiYQfWGcvGkZldc2vl4r7BvBcZhx51
uCbaJ1t3Z8GYoVa+4CDWk+T5AITBnfZfHXd3SYG7+jaWiI0MhBAvsu4QjMxT51BUFrVnuyoZN1bB
fgTJyc325d/f8S/X14rag1KELa35G5hkJTnA+QefqvfZ1ijVRglGzb/oX019hbYYBWNZxoJY053C
mro4IQecprHMHKiqIjGlA50R8FD1YW9FNkNiX1+JBP88Nh820Udh/QQMVDumbSWIbeZS4IXXd20h
1cwV/kIOY69deTS5XDiaY5XoFwOi2djS1GaOBH1AvSsTiRJBMRkzla4VzDDjkukQcUlH//R/KHPp
vZ4Z/5YVgobB1WVb6mJFYwsmJEutTHLnrzHvhPBf4SEPdKzHbxymdF6QtyWdREMiv6It5l4QzdZR
RLADVFBxWtvfALJ4CMUA4SUjaIwCUhBBdpcVqqE1V2ZiB12Ixh2OamzE8OZmTxWsyYaf3K11H+Na
LOwj7lU7yQa+GRX0ozjsQEeYaAKOnHtrq/1OBV+4Ca00lVMlYf3Xf1zfRoiFGvoNbf4WSnsFJEwH
ymZqgyt/TalLdTskjuLrx7SQxypZIrpCe5XYoPW2HKB/7dHEBOIeImWUck/2nt3t+8NsqyIFAw7u
O+6qoJ6c0NbsaqHOp8cEWKNSaQWiwuVOS9kawVw6zQkPCXrlDBGw/lfAWNNUlVOrdotczrJg3hrS
8PGh+EdTnKgyMYw/rD/U/eFaKjxM+an53NgwLnQaLjg+pu75BN/84W1+Zy/60tlXgXGbTWvnE/py
tp/xd1jH7J0C/U3Os6e8wIlpFUvVWEA9pa6/6mp/aVsngvfyl13zHIDdZtG/nl1H9/SQ+yj7SJmU
DBQjI+ATygh5QM2lwlEeUH0woUk7UNsfl9Yj3qBUpwoFrE6eRsVgPIfjHXE4kHP0q/n/w6cdEBqu
eq5+hGTVW1cOCuHMfh5qqv21rbthDttH6SxHWX4IpIpo9as855SXqRWj7WgYKT1SKkSAzPi+HsKP
LQslVo6HDVUxk97IL9ydem9TZD9YMJTMhx6Yqkw0K0fzKlj5R8g00ihzq+pgD5HhaGbnp+Qfr6KE
n/4Ny7gdlTELXBZxUpBUFi/kkApqULXwthyPup5PjOsnX8oFiPHAzKGAF0ox4Hw+j5EX0/vPWMkp
B/KbvvPueNSzgUDnyH7nABdEm/bVoKsz3FxXmk3MLgSTxAU40A+LfkKdy0Q4MCB91+PH8ddEpMoA
EDK/P9Dn7CHtY7JxeO2xCBhYIjcgYFInFECOifO+AuAHktmfBbwHV9tRH209Oe9z+3DGYtc50fR0
RHT4gLTDwFl19IkAjmzmdBMKYkym77x7mlYmzV37VDoNV8/27ry/L9fJdqaU0n7NUqLzxTyNFDzF
FAHSnLJ7+2viC+xDxaBP0rfD6TzEmXS0u9+BRqpvNI8sMojFjBAJ0unXYkqXpfVJplZypoyWJDI4
qvCMso+wOO19/v4oNieQzOvymjoausUHRTQ4+Tb80q7ijPIF629teE180nx9JLsDr3Fj8w0NrNlz
y7tO1+tUb5YYiJOTRpbpzBsGBvKWCSal04jUGOI6IvyA87b5wVlt8Sa8Z270/CW0vS0eDC8N8hxd
2+isRvrzBGAQjw3Hf+M8Tzr6Qha2nuTB7ADHJOyMr9XeYc7c0SvwokatN9eDtTXkmkFjprRJYSCW
j9fYuhc8HlXEj5y5uUZFkv5qbTyps1VJ9ujLxA4e7cnB5vqbn+gHNeF7gyuvfIOH7yL+KXj8H0E2
m751WNeXYFcLeaLgXwDvUrVMfZ0bPS0znLZ3YkCPSJXUeWku52E7xFUO6n4iGKUz+EAuopu40OS8
TLf7VXeRE2R0EVJDyCqdVLSYezznEdgtN1I9of0dnexUz2WlD8cyIyoSGBEyYHeBOAVCk3Q+CYxW
0S88UrMR4u6Ix+o5EejelsPceTn6tpIQNZo5uhFoxF3PUyA04Y8b55GMRKG9QIa3kR+V2ROHUIKM
R2FQjVFZd5PxlhUne8ojSzAz9OPrkn9TiV4IzepIuPndXynWSSJ9AJIRDWaSsUglQRdNxESdIzhW
Cc+B6BfPyXxXOeW53aHvq0F0aHNMijlaRDAmEL77+2PRHw5ZNJ9AwZpHqR/Uc3Hw57jm0ZZCl81L
Op37rs4319k1LEkKy7FwKoP0veXnPgn/h8Gghtymkn6uq3EHbsCO7Y/n2o0+iEVC+Cccyfsx1Kb0
rhtG51B+IT6WB2bsaaKk+Z3Th+5jM2MaV4PlsMNcmGahyEsqgutLqvVrj7FaSVfGNG5/K/amW/M+
L9iESJBb5kv0FXid7rq5//Mqm3Gq803zr8knruSKdGXX5iQG3RoiddTuGcQXS0Ir51Yonqk5woJe
Fb1RzDuiy3goSEy7U4P+6R2RUUz7kzzCR8TTPU6AaMBmg7565KNI9orGcGHMf79tRpgx5kOF2hT2
iv7YdvpZMnHx1dEFWDZVpSlhciVUI/UusGW65dGdeTqGm8ZlV11CSUWkLY+UaR4pdnusbLHZ/ytn
etjDoLcNXEh+AggkAA1aPBLeAqYeyOKSntAtcf/s4dyk6inC/UKNVeGY2mQpvg/yEKSQHDzPiiU8
xsq/V9K9RKl7TGttHJovWuhBMRahntcfdS8Q5CEZgkSc/634w5hW6s4oILJl5Xm09sFnEhKrVd8T
7d6py8h1dr0ACc4MscLf2lDhEdzrPd5e557gTtGdAt7zvwjI1xNi6DBabaR/0R9qdoUdTrtMfwsH
vd8/5SqTa8cLVCQ0oeBDDGvBSAf8wkGuzHPtlZVtY52NBUCq9Loa5issrBMSxgUKk19RnUFMANzA
Cas8MQRXqYJJhQmuvBNFjh1bIaWqEaSdkcuVLca5vUljxBLKX9hfRsJoERskmMOlwOToypu2kmKS
oTZMyo//KUp6xbaCsAODRQVVTdNJ1jlpTPnuwszlu+HaLR5Jy2C4mZXbktALQKDcewCXChu0O0ZC
KdhErtmEW+ykfVfqYEl7zrngNj7dv2DAqkoYykpquyjRKUx/GEhLlrdQ+QlWpSRi1QAcJVa+JnFL
yqIQUgETeqHXG0NQfJ4UGbGY4w0xUx4mSuN8rrOcOPxlvYL2zfLl80xFtry1MjURWgto76RH7MQ8
EAWdYS6u3E16X96sZFNjNwS3sdtwEZgJQG8wOlJYJbUuWfF/t11v9arnosa3b2mXzdycOR4OT1Cy
umuisMn3Ddka+sxXjgYv0Cisadxr5eK+KADlJPlb04elXL7bL55BgaFd6uDNG5xSOFEjk6iCprHs
1dWB/IFNH72vFRxDhmqgey0oo9b83T00744vsECTsfY1fsHmOurOkHQMf+9p+0kUi3OuN3yNRGHj
Lmej/0tIO3b965U4u/RpNNDBPSVY+k0Npc3HplOHDo+9Lc+TWkbDkFLBJF1FQ9ToyRCMVvjLDTOa
1nW5M8qroU95+UsGb12cvTN9EKzNuQS9SkOhkv7Sha0c2urmtfIZJcG0yKPGfd3ap7QCo5wnsdDD
zHwNIMK+ht7yvivXF0Yxntnu7O5lfqf7anfX6Gc501wy1h1T90n4xLqSh1XgpfUyLoQ3JjooG/r8
k1HLnQWAKe12e/pivn2n/NuufXMf1lgXrGjW2eQWNwALFVgz8TdpnRvEm0SvjEgZcCGxe/w9CyNT
Ljns6oRxi3c61cJ/it33b2CYTnml/dh1jg/nwRSzL22x1ybdOGkZy8OwG+Mo6MsAPhwWa9mlj5cS
clLmwEboXvohbj8ZdKXRkCJ8qwc1O3+kbsQVuFiEVbZqxIwDmRM8AiwCNyeSrFNxdlR3VBvG/vFx
UmMYY9DePMO+kqqups545fa5c63ueUc8tcWe7nx2AZt8oWO/HCN26X51ig5oafI766Y88qo7iPr9
6KhAZYTpLThV+4RKXbxN889qghg+dbrEPw8WHgihJNgH8UQfGYzkpl28jck2A4D0ozPkDgM2oYcW
B/b3iRotB9I7Vau0a9AvqOJzhJA+a81cvwb4pApGZkGabvFIHOwx2gEp6bJcnwD4wX47eXDpTUcR
DVMJ5CUD+sZY18k7it3Ln6VxwiWvALb5RUYZcdYAFen+6CZLmsL7g+BYApViUCSlzHx488/5R1Ck
B3v99PtoZnPrHrmZsnZHJQXs8l6XsJWGveCK0f3aI8+tFN1Hz/elKX+tK5dgoCCxOCVa9AJaL/SX
XHZJIfoo6PLHCMKYuDX97Lhj0cjyIHwrjs9dvn8Zy5Nnx8G54jK9uifpx8lGmMfvLE+GTCInnXBz
URCgQLAaGkywpMkNx0SJP18mWcAGMp6oH1o0gunIt5c1JKX+sUnMSRrGRjbGfHoMgiNq3SKnNHOm
0A36iDHY68dYys0yIsOE34U0XKa+uMC7bjGjI/vUgAoQue8095sfXL1JRh7ZYnhDjTBGXXIclQzM
SO/jHokxbX7sOec/jKzcvZoHrpZimaNv5aWnFDp1vG32KqBJpNbI/2NBY9Srl7ZYrPWzpfRPJg4Q
mFUHhvMe/6zMxs+vY0oFjY/6UrCBTNWL7LffC/tsti6xk09DWZ7mN2ALlKGwYUeN30Uc+2BvGQ+I
vNeGlkG/ert4jq8Doj4xmBLHqLuadeqITym50P/kaI2y7MSO1Me+7NXxh5gYtHnTaoVu08oR2i6X
LICHwkkssQDlTAMRABqz0DHXcZrMdF3BrIv4u9AeurJcYybB1oZHygOaLdFVFO96FpVSZ6mC+CvM
SqSfTHMVufmU2l/6N+fiJDPYAMWPC722cW8s8WMSCVflppM5ksOEVxRL979HVTUQZrLJAzlITcOF
iqGuqPA7F6t4nHkNFrXcl+gx3I7Gti+rFZjHIsUPT3Gg8AbMQ9lr5iTLwwcEZBFthmdeuC2/gLUq
FLwkDRju7XDDEKAKAKaJwiLnVClXA3cnQQPILKGqDCjcdHgHCqlYx7gM66L6A/pOF/uZSwOMduTD
F5NUZqNJ2SJ+Ds1h4U/Kl61cNjN829wQTwktyY6RM0Ac3wFmNvrQRSLicV+x00UZDAEgnXWqI3B+
KXosR40FkBq4UoqYtNJR3MZJiFn2HxjSybwWCmPasl7iH0gSYhbyXZMWKy3EGCHJG8alzwAWvmsM
0nhJaRcEYG9AHZqzQa9njh5NRvtrzSUvrdJOpcpfpw9j3ZHuZOgRM6qOoy4mE/gcGSt+rVuO6qlh
7viTnyaCxFaPlvNRfhSq7iXfuOcSdmYaVte3cVXQUJvFljDTMzvb3BiIiCdx0AK5d2XOFSB2UAU0
kJy5dfDEa0SNMPKm+NIWZHdpLmhpf8pi2Lh8paJqnUZAJlyeJB/x0pL9/kuwJsE/a2hmXwx8iJBW
TCYsgq5Kt6kOZsMOGht7U/jfqCMv2G9DvMPLb15ezriaF5nMxiPMp+ORLtH/s1rLQb1phiWYOUv5
ElMJFep2pqAMVW5PdaWaqDIhqgq5nEXb/bgSq7D7wayiYyD/rx7vAfklLhlBZTRlQMqf4wZlaGpQ
gwMSzQqpZkQIZFz8nHeMuGn6HtfOTDazJqWYnCoOwCtGR21ndD491xHZq1BvVfcKW4qf+shpaX3r
95Wf/Ibr9swdXPp0uQYbEYBZs4fx7QvxConDsOq73s9xGiqBSvhZI2zhlbvlo/57Fc8D/AS7rkuq
gPfcFu5sXKS86At3op/jxCwKhK2U/4OxRr/B0rlf1/erXtZXBALTOHmR/8bRwHkml4OzvhnFoWD+
K+E93xFWdez91dY7T9xI7SBngKTkKTtK6gIAiDPI0XOhKRGM2oMyM1o3UJleUDEP6F5piS5X8xSr
cZNXeIFCQCJYObIhKG9KxlPPwlJ7uPpxo7o7XRE++egAHjVEIogQoDFwXcEa4Lebx8XLdNW7126C
zDKtnPsxeYIviNuQNMVrlUHUld5x9ttpe8XBw9vot9dNJauJSgOofM0w5P41IHXb2OhsilYiz6cm
/NyVBtu5nKuBPtIA0+99Df3la+XbbXnyQEizzLlH3jWT5PSZScwpXQFy7vUwtekNRdZjaoVUqRb2
FjVWn8RDf3VwO9VFPNog9pfzpqXf8mqpQoRefjJ0pWM8E3lBitup8AucYxR3cp3ma+cTHBMGuOoq
YQ0nEhre/f2wUljDasLzBxuJAkojmTVv0ivLqxKmOLKliQ+wzs+SI1mnA/t9pUpLbTUFXeZFPGMG
kGVcQgUYYYzMNWw1vDXR/qkKgMMz4eEzWAkdM9e+7J10/ubzCr6WDF9g2ScdH3CDJ9OaFGnYkq78
lC82wWyLXmD4HTwtP+wOd/qAx8Ft8U5z0Z3/IVLSdDZzdzuVBOOtNMicWHkq+TGbKZAWRsRdMC4k
juuq+rs2uTZ5tlcWcwPm+nyZRlX9p6oBgrSz0FDoBP6ws4DaHKKWce4DWdglg1mldtAihpeibPVf
B8hI04p4OMXpy4E0ENeUQ8EM1GmQ7ATa6+E/hUE2TVrrpLDME0V83rreIimh0Jn4ukeBurwSzYdB
wVUrf58/xyWqNWLkPgq9V8DEs6ZWkfEgQcchKXB3xBRfRRCrzEfUq50ItpapU45OqM1ST+o+VGh8
+jzwz4bfnmdbbzPovZd5jw4sPK6///pAByMpxUdvn5HkginxHrS/HsSL01NNWxmwOYX/6rTCRUZH
oDutfvw1+TqvYcT06ETIrXbHRhkJfyeB88x8X+5eaZaEr2gAFIiuCl513nUlyaTafKV2264BmOuC
GGtq3+Wyay9Fgki254R5IZPR7aj5m+yS+gSKuukAMXiesmi5TqSJaPTXBawg7161pZsfzZw1X5nN
ri3/COTLFDXtriotn096s7GQb38Y1W/POKb1xGE9jwk6+wtTnixlT6WvAqKTDl7EaIr8tHW2wkHT
26Im+IFC775lV1KlVgG1XcZOfkg9fA67vRx5V6eWvvu1tW/jvxTGTqLznJKL05+L+CIYfcR/SQz3
1yTt6wG3UYWToOBfWRKBpVE6v3R4/AGTSq1AmT2LaPPOrj+YRwBiRijpk0dT3m9KVg+EGiTU+aV0
XTzrUUOL392X290HDPpZi0Iw8YkinA5tJBWSy1NL+2MCp6Se7fYNZYVrSOaPF9tIJ+jNEjwCambI
edJNx4297wPmfxji+3FV6wjV0fcpYnw2VePQFOZzVWDFk8Nn7wTQZkz5LZ2M5eLKB/4TNzslIMb8
XwGphgumQpNKMle18SV9VdmEh73nAsFwxt7bfIR1JV4ZJ2h5OuHcGxU3zCRhuPCZmYlOHzuxxcgz
aYw+36sTQNrVm9NCRc7OXqLoeQ56TnmAYZACe5LaZVzdx+WMlQiRQu7/Jgr5PN1s7G5lfmNPVy+4
EhnyNlMWRytdq/DDoAdMywz5TBg1bI76NRZdHSxuD9CmlLUHW6cRuUnF9uqzhr4kyrUay4oFV2bx
Na+F/4VtIc0ykIz7juQwFiaP4ONhX79xLj7MAMrPJ9xhLswHPjUE3N2WCzvGQjBbp/5hFAA0yTXG
+t2gm/NzUhVi8HaSDzbwPsWCDTv2Jbn0RmEMO8uMglKZ8XTdGHCWokzpVYIJSDo5K/J3t4BIbM3C
w3/2E3LAQ27119Y2nuplj33Z1XoMMBppYKW08HdMeGR1e9zDxRGdYQB0p8wM/xeP9Eg7P5CUqHdz
Di9S1/De4EvAPUvISDOTf2B/wL/Pa+80XbJw6ULIFzG6Lna5/OQCDAcS6TODCAYT04nJ2aNj8H8h
zNNemSQkdsFwoQVdjTgkwE2LPCeUuumdtjzbJrNYwEMMqvRmbiGCXrTT88uguTnMCRZEQ9vF/P+m
5uswvi0qPdy+Qtd8O65kJc6WRcFjFU+y98Zdmm4PyJ5WcFurQ6smpyeShYNNhajh88XFscy1+zEj
OmPNFgRP0uSUd1pIGGrAeFEgxiaDJBHjmzdqP5cXNsg7u82BfLRxEj7YHgj/bi/O7RtOJArb4m0D
9s7Ubms/veE0K5WaBrtyICbU9XpL1zp4xOIiy+zNMstEcstDp3OhIFMZwWZoi7zhdaxGoefkxy5Q
pfNGe+broek0LkCE44br50D9LKaaNhBH9UbSvJP98W+X7Io77XlYMgzFuy3fB7euOEHFp7KWHXRd
YWhb9BbNUodlgDfa5MqPThZ0HwB1r7EbN+6HhvnctfamL4r/ZZyD5Z9w0Dj6PDN+1qKWGgyRBpcQ
9c0D1Su7iXwIzIst7f1kdiv3MAnzA0JZU5xTO5BTUdb64M+4BdqQbY86rmOwIqW09xyUPFmxMpuW
MgpUKMDY37g9dhkk5gedDPVqDt2NggA521RBX8aOyqorLU7mdxQHpdhjN7CZ1ploJCdJEHPjL3Wv
5Up9xeR/7NdKJdduBBbY198iDfUlOS86TYsloGYm7c5/MZkQwFCA5iRsLKF8w3xjiBQVyuosXsMy
oVqRg9ff5eGr8pwZwLxxTXt4z7SDvSZTGam6GAQN30Ypj27SL/7ALCIQ6hpwWccaU99zhmv4t3yJ
XGzYQi0UttBLkz9dDHSqxnZiPQ2Rr9Hk1ffzgzT6Vixeqx/AMUqd4ejvbtlUBz8gdUjr3EBOE6FM
+yZiV87aWIbaG3fhOvthp3qjE6uG5901ylr+P1XK/VsnmGXChaNKWxlNa5au3K9onntTIRbBQHx7
wvvPunJ+r9r5PedwdeQ05f0zESAwpT4cBQ8VPkA0MpQHgn1bYvX5jsun+2PJM8cw/YUbQ7bK5pJb
QmWfQCHmJAn91T9XzxC/R1v63JhrXxU2N2iGyiEKZXeBxS1j125SeRxY3Z7RKAqLWx8PiarBwSVi
AZ0PKBr+tuuJXb0YaLc2Jb5YBv+fUco/8d+20qIByygw+oQSE6Y8ewWph1nzK5BJzWn2RXXV66m7
OZnKncK8afNJDNtbRP6Vghq/eC97OGHXMZil+HWP1q6Kq+UCJ8tYGhNDOkzLp8SZOU9QhEmWaOph
X8E1g0tBceRfHfzkLQYNmqIkFWSdQVXJJKsC2jaZG6geXcsY+sRkoEAdjYU8mpTjGaICrlLVb8vO
/9IcPyXrW8QkwkGfLWn73TT43zw/Hf6MLio+oMz2ycDIgWvG2ZDUe9SpG6Bj773l8o+eHTX98+Up
ENrHzQMIkf/nDyLPLgA1HKFjIDK93WD0UEChcbfrgYfBJ2GckFLk28mL7IAkEya6EOf9xCRuT3J7
ilUaXKDTNnkoyDFN7Y1G3euH59FRetdeyzLy76eJTDN+uI48Ai/SYoJy7F6HIy9GDUgMJm5R2bYQ
NIZWWZfTTqV8vvlyWgMfPVlquM0YFpjIO9lNxgk+jpcGXqoIjiIGJj+aj2q3EgPBtkcWmkCBBMjc
Kh4zhCdiDtMmlhWlwQQG6jeZhHIjf4BmKnimJLczLR2toCS1EQfeg0ddb2jqEt1z42nx7dIEMe14
e9C+MTOpDtj08GIuvNzzyl0tqfV9LoOsEw7D6/Hwo838FNCIxnluoENbl1072TI73UctGcwOYHJ+
XEvLCG1AA2wmuBERMNekvr17vRkKEPFE+2N3g96LfLTvU/p5pPgMWUlQnvSxtb8h7RkoTno2GOvr
m/AbUlIGMjuOtV9Ah/emHO7NzUJeZvcc36yNyslL5FM8uhYApM4+yQP4hk21SLkbvq9dI5Yhh0E3
h4BH33TnqhNpG9HAJyuKlszU3Adk7w9JACwMgT5py/3fQPALSbMUPAz3AFxJ2OyYHmPWXbf+k+wq
kq/7sGcFtRo6HYxNceE1i+/rZpIU3QmpaTAsXh9kDDCkU57ZbISLmMrksi3h7iushgNUiwcF7par
/gpfzxXnUwUwyZYqdo0UJopG2cGY4kMtJCKoRRNbTsI8NcK2CT7fwPFPh/FdcBsEzVqkVg+dNQ/F
J4VPW/ML0tIJdfnjDjXc70t+XcR41fJxOAT8jfEpkiGum29/EzfZcv6JWZeCbgRtnO9Qbk3ryN8B
paI6Arwb4s6TYAjQbaq3pY9iOgQ6fbRds0njXSvuNB7jcOo4VJ90Vld8BGShxhAOpW+cyxiOfAE4
jvuqcY4guMRQfUdIL/4kCI1JLH6pVnzvP13nlzvlCrPeNKf8NeJIpQ+RLgKPJriOIqmcwskUOVxm
4WORHw50FPtVLAJwaD3ZaoUjDMaxUf76d/vXBvI7WCrxRBjycN7kH4LPXY2qtBcUtKYA4TkxXzd2
iN9KWJ3BTrIIWMiBTeAC+Ao6EddT9Rr3amDCMh6HOMaKBrNbg/Jru/AqTMduIxcKSMztV8hDMnc+
BWiSbCt59aa5v/+DAgt3Z0TLc9BsTByfXoUDHBayA/MKRb7N8kNuAbbiLucx1LNBPtSmaMs/q4bk
uKCPrA+OxnPjIZy7YWqCrv50lpxiCUPMuDqeBOGX3bX2wYS9w2KnedNk5yZFrK4yfxfJUHTo1YUV
aXfeFCvr6hyiA0k50iELYtuWH8TRjoJuDsiNT5aeu7W0PDK6XPDfYd33BhAtfr4N56MhKCEjM4cl
JOafJSb3s0LVeF9uUFExGgQvA6YB1DP6uA0VM5bobJ0SqZcVSRc4ckc2imB5cDnK4GyH0djf7Kww
sSaamhWBCBTGNNj+wIJgQOB0QcCC4ChPXU0ntgsptnO4j36Uj1YzTrdL0TCLvsDlWUZaUU1h8X0j
NRDfv21HKQPJYOt3qQSp13aadHq9nee+6wfOH+wOFeUBUn5gV40PJfRNQY7Ahd1QqpG1vMLX8GiZ
5co8DI0X47J68kINePbqRopPE+ZZqbjYDOTxBajOjAaeKqa6tjD/q3iV0ArhSD9NgLMTcv1FfMaO
2McQhMQX8N1PDPtYMi6C8xZpeaXuN2Y7M7+xqYiHi9dQ5QCq27f8cfAvNOU61/Y0JuWDUH6Fa/d3
o/S6sPZ03YJC37b1bDF/DCPNiz+fyeTu/18imHmWwX5mp5Qp/voXv9SasDZpEA0G4SmUIuds+2vQ
zgX8eatjXB+0AWsU6PB9rE5m41EixmN60PJh23sFhWyFdivkaAENdEPLgxaq4AVPSns3qdrY5sJG
jKWVEENvQf8qd1bzMvaV8FjXs4RvewRiwMLlMgv/nVnsbImQJDg1IrDOmepe9EibS3RP+e8wj5LY
duUBrRrSMZOI9XhxD/ivUEk3nfLv+Tn9/WMqKe5145qeA6bn5c1vT2tXaNYWjaDsd0K8I5kx7lBG
tmJ6VLdW31CidAtoQDHEtz7m884QrEi3vc7XrMsg3R96wpbeSp50v4rmrheBStzanvy20BOECKXA
qA+s9XvG3cfMN+sn7v6x2VyIG9aBXFoJlRHoWTWTlf7E1gNJAzGwUJXunSxxlSwfxyh35Q+1rnfF
J8+Ko19yJvTBZz/kQ2KsNo58qxr26oIVdRHG8dICQvayDglJV24OgHsiqi4hsrrinOVmAikl7Jh9
znsW/inNzERHFC1nBm+un+XGdZ+Lec9aQOwkNEjySZub704FkmTRskR08pvs3u6vwlstlSgxQLOW
4KXEY4pFiekoCu92u9RkqeT2CracuuXChs5metXsv/QBtyfu9lBC4n3cYGcm6hwN8J0mq/kWxlQY
aGF7BvQd2FQOJHnIK9Vo/2xPN1/Sabeuxc2sFnCniKYmoM3c04cubKKZ7v9P9I7yEDZ1Pw8FtSHy
98m1frTiU3Vk9Qte30gcdIwcPrFFl7bThm2anwEpIgPxDvS8LkJL8qrGwcLsWxYOO5fDSbtLDVVD
YmTXOVwD/NdzpViKp/mSYW11VBzigIO2ACie01/1vhJ36vb+B/wI+P4iaU8BVQ9QZ+d9sFnQ8vam
8Et7bJnWJwMq4yF0gT4EGGcxwIzjotuDk3Uo3q+17B+OPXNKoYsTtjW54tlE5sESb2aKQ+DUggV8
EX6z3JAVuFR4MK7+A8cQemVNwMTgRr8fcWo6GxAr0r1SWq+tGq4FCM23i3+Baxo2iEP474fw/Fxb
wL9KV4k3k+wTBS3TroAJaYW+o9jxhWi6Rl9OO0yQJy5POkgbgA2mL4rlfolAKQfYSlZ5bFdUe8xq
+21u+A+3M5VRP7WAYUznemjHFL8eS+ej3v2wz8sZ1EC5On6REY9QLwDefGPQ1Pa4nkJ4J9/oZjCW
Trs/HtYyTh6HE409Wo+9XsYzUWc5DxOhz/KFjI+jZfB5S4NSpdDDfEx/796iFD5zpasjMr91RvwY
EO01O075rB/KwzNElMIJziRYFlFxDqfMn0Eh6swW/Vm/piCL8YfsMYrgSaTZBLBYfFAfWtYiOLa5
sHHF+/sIF3U5N0Qmsw+l9GhFbiDK4QM8L3dh03dS2YUxflMlTPqZAv1N0DhR1sLUj67gCiQZzzXF
exC3wq8ArbvRsO+FTvxS2sPemDggIE6UwWOMGISjw68AyyesgfZQLjybpp3q1EHS55irxDdSLTEI
4kyX66G1vk8O4I4e2uJaBr1w90Lh9gQ74L20Eo7GecHxzHNBzYm/CvSNAc0ONrkFxA+zpzQS6fF7
5jaei+akUy4MIjKiRusyObvKomZcegz6/BCzD2vEv6iKcdl+2Mlkx0ECVvRjbV/GRmNBWgkPQ+LZ
pu4s+9/8o+rzYzEYVZiULYrTaCK5Sg6uDjjWGxBpHY2adnUbRy4TijR9ukCs0Pa41EqbtCHmScY7
s7hXp1Uy+kmAJw9pgPmEHi4AQRzNHq7tSpU1PHGqzzDjAZl6PbU2pvHVv6cWfPR1HrHunZG2kyTZ
SwI+1BctsMY6YLw3V5PVpYroa60cYMU9gOEnNgNStNiDmj8FELbHY15kXLT5MoR4+zZrpedN5A/0
klgttwY6PxSiAWvT8j2vJiUixZkrfcInFFFlXFlPXQT0dCn6IPHPQP5hpqML4l/U5zsuNanhqiMg
rcBj8ZRev83R4zijwlc4I3ZUdm4OAOBGVpeeoRN96H3zyo/uLCM0YEhZEVGtJxcynVqM1PpGNAb0
I4CfFeNrBZqlrxCr/84CwVYNhjsxNtT6jMgI9SGJcHASDc+J1LoDbu24NzuY9nKBxTEg2t1u6hgQ
Od5GPAL3vxgqvanokHrkbJo9677BzUaP0dPl/Oz7MRFdMJyLUVzUOp3dPLsf7D7S8wGNUTI0rCPj
C/Xjv1cJEvk6owPULaTZlpT8/HqyP3aIhqca6fRxk05RcHww/hB5kAZNbSnExyZFCfd2+YUKA6hB
q9f+WQhQFhYlXxaAXTPd40UY3ry4Mh5qSNQQN7q4XtFXjmptRVaQSI8SFbqYzL/I9+82y56RV7+g
tz20HnIe4F/PKDwOHTMH3mrrZXYuknTEbqmUn+C49QdV6qV3QqHzX0FECdv05tfICFFaC06LFsFh
yeEvJdLLK/MIG6qzQZ4pr3NVFSssChLmARSXW99956P7CvOpSxsY9yPrCDHXcivPFwVgI465leat
w9wQnw3mLxBJtxw3diRlOYTuFrs8ugd5dpgPji8+vkiMxJvrA0Sw7UkK5MZdcuOrkhSz7ItXbhte
lWe2ggA3f6SwM1Rf31F3uLsW6jQ7ClRP3hccHUpwOzPvqY2I9uho9nSB2keqnx8nu3MnJyinCmko
DstNXRaM3ZfhKyxBqjJVORVDrtDy7aMbD/bRSKotPEoZJMdc4/PByoZn0UkwnP0OP3YmELyK8kRT
jsRB+JsfO4yf2aNTaaEOcryqTfv1KUrfM/srV4y6q/UxMRBQCHrIUmaS6XiMAsYUBXYuHLKs84Ax
tN4FH767PGlGPovzkGedXOJ0vmm/nk7731S6eTSKIS9sf9AsjnvD1mNx52Vo5yf8kyU7cmmGlbD9
Td8KeXYFLBlSwLcbthlvySjapeLk1x+j92cw/TRc9x78TVbFpbWTQ6k5WKYdMNxJBuMrnReINwxu
DLp/xb1LVd/dyBZ2r7IFrGGJT7WZ2aRt6ZEVgq5RndmtsmYZX7AXzTyi0PVs46JeZaQexK7ZeNOK
4vzpl8luIOCjicKepKkAh0/jqbcxcpK1b0jpH5XpisAZu46cocT1ZVI2ZUfLcCltV5oy7t600Yuv
H36WG06qp2ZlNI4+v1ke06mwEsIhmYoyb19ldszaClmx5nmfcs3P+pdb3IxXDuh2Q5X2SKdk8U4N
AfQWvIzHgDiK5qci/m4OiXZ68fmDwptjsf4yoPqMXycRKdQlpKLxCYWWCHnZg/h2950JIG9awt6y
tZ2swJdNdydR9J8O6pezMHj33OdnHHuK3mhP1WduZ2iRcJ9aDYxhsu1DkV5ed3CjtTeqBajOJZhg
0Br5650VS6SuwC7EL9VRT3jogoXCgMTcqbA+AxgG3tT4x4RmUR/DZuHunHjvq3mzOgrOpLWgapKb
rlHO3Q0ueB+zgaN6vSxgyLv/eyhKrFXTHUNavYY+fEqmQAiaZOJ9dNiJKAj9RUKsbFYBw8iObYio
oLdBnEUGIdh+SC+fQ9Yfp4P/dzST7mEoZ83aOx84eTVarrcpeokV8d0aqI5E5b5lXnntZHq/ppNY
6UGxYmKYPL18GkVvXrevqw1wXEBcOhBvB7iDMX+VZTJnApGxQCg1IPCs174toaIbsrJ9gy6TaI7S
eobjWKRaqd5xJ9awXWtbrAxKC03oMJArRA+A26twBRxXFLxJKCet229OkszN5zOUzE5ZsKshbaN4
EB6ZYAvagfxOfDyg8V8vVhaR/xa44dCuU/oeN65+jkWXaNK5yvRx7nmJp2Y4mfODc3vPYoGFX0Y2
9YWMGH7efZgzVmezojd0JCY0ocLEfLFxJ4fkAzGQpbmU9JD92jgAyFTP7DYMhBhEW33X/2unUe6a
uSO/DVybQVO9/gIS9rr9B5wnYDMNLD1aUm6eyH81077pekaaLeg7Sq7+64BwQ5tMJR9TnSUwnSWt
5WJDIAwkyrYnV8pDmO/UY3HI4FkQKpR7Ly0vQFZ1eR/Tu8gjKZeUlCFrIy8e6S44Oi6CWwxGA12I
jU2rhr3KLpwS4B4oA7u7ibsJsRtzCZgX70EpX3mSUb6QGIHtESxUbjUDkASq1nX8uznzfoqUl/qZ
+2q+SxBPmHcH1htiIMF7KGgXfx2D0cPa4EkF6v8tQmRfxLET3eCj75AM3Xgf2ckNjuyrSqWdEW7m
s67FiMaxl965gk1eN7K7NIR+93tHEtwwDL23mwWNSffY5EJf93XlwqKoy6vqa4bJ3qrTBI589EqS
vpFrGM9ggltf6YStH+0p+tNt/c59Fgv5nNznh9Gh4E7uuSG8wPE4ZNmaCt3z86p+smWzG7+MkY3T
Fp5zpAQLJH7eaC3D96o6Bu2EABOxWiCcX49bpICT1KbwEwHR1bKNnZ+euUaoCo3O5tPvpzBMO0mu
DIwOhk98B2zMvElRjBa9R80bx4lWYV7kewo8cYHeakY0LIYzJG+hd6utvRU10cDfbCKtTV8J+/4H
y6+T0Gf8gqEHyhzQoRa8f9f3m85k5NJBeya+zsw9RO6IEmiYRNJ85wFu7C7BapcD+BdofvAiF8vP
s9nk2PvMdlVSbHUnoqQvY2VKIQER1lYzhe1SLoh+dOG8N3yvl2AAqpUs+XVOC2iieFPXBK99cPL8
3XEDaw1FG8uEtQRhfKIytpYBbJS6bqNnRKogqyCbGxqyjutJoWX3CrL9PwT+08AMWz5ro3xvDRi1
zW5szRuGCzfx2uJpUVeeJtmbcfK8QltVJg/RHnQprEwpJ3D+6iuLMqqqjkqtRkdXSDEisusYlIpQ
kuc6/1/KE64pj4EK+91n6MQxpLQZgaLFXOXWnEjnl/bPi+rxMAe/odTz23N+r0ZSNnr+YyO4byuF
eEH3n2x1WhQqSEC3Hd4RDz1SCbKEjo1YfmqmulJDywdC/hsDKs4pW80+XXT7kK3ygmY5UxXxnLvR
P8GjDkW9JYBBEgOn99k3HlkiNDZUGYrGRn1ovQ5JKBw4ePG9HniYXBVS7v1fpIbOHZbUFs0e/Rdy
F5246LdYo05C+/prSOMSpLweV7ePY0geGSDgu6knRi7uBwEWw5ykzCl9b/gLOp+OrjwPkU+gureJ
5VaqxLpB/e/vLsKRVx55x+V4kWnBhSu6KnuSGzc5pEwkKsdvOCe5QqpzT3StHkQXbv3QjfXtXNxW
+a7itIopb8/j+MJqComhPgkkis/ooWOwzflltKJ/HYwV00cIMAttvKUDjRB6R+9AXjAFQcKH+Vby
oJTaipfA6gXLihnciGett/pSrf68B+9Q1diFhCqo1akybcF1XbU+JrzxXoMI2KmEXhK3XCX6dZkq
1xHu5g12CrtuO1Sh13FH4fZFQlZlA5n07TjkE9UEZlkcnYPdyPj5HloiELxPxBjL/uCtn5uPbPPb
HCuPIp/iiaByd6Q1HR5V6UApi7YSunG81KPxv/S+fr26P98lDmYymiu6LFc8Z5w5PJHjST23/Dxk
rVVDE9gGt2UO6z6cuLYL9gVgwPmvldNYvZpyiXoJGRHZBPXmobP3IkHu6hNeB0SfUAj0hIU8nAVm
mdjJP+sRg+tCkx6gPyIu5ZzoxSQfp7nrPzlBsSi5uaFHLlK8UCaKeXrmdaeuYt2dyQ6uCqiPwBOE
o16lLmWbQpWtMS/CuGzpZwffT3/z3eoLso9cThnX1Z5O4lLDHjcjULGGg6YqwW+kVXddMZjUFfwF
820/3hNUnztvMVpP3WfnlspDrO+OpSvyQCJ5WYYcNwQqkXIHxIZ5TBASr5BloAwwH4TR7JLMsMku
/hBCsnjb+G+oRRC9kJHUd3afxXJi6WYgqxpttjh+9bvWg0OHInV7uRRfm8uXdGzRNXxVAGkqSZJF
ANX/9VQig9kXi7rzsWoEtUZpJEXPYJssnL0XnjdxFlF6TJIDzdtn2+SfFfy4mIr1pjrW5zQ9wC+x
711Z2nLiV6kfrhfETXfI2BL97jTYlYrxIw4Eg3Hkigx3wd60O1K4pMpb8RuMTFDdPaj49mIPg+NC
Nwmdc8zcgJYGbFSkBK9ytef6/zTyW2i1i9lHE2fPmK7ZZyouwVfROFJmLvUBbunfL0hz/ji1p045
ccLOt9CWoMx69Zg7/SkKuC2cp0vkCp+onjvOE74jqaKGjRSlQO7vlYLelmrfkg2nTzuEJrKdtf8z
AgpvHTWZoSNE4LZ7s2+khLYkBCPVUdgHP5d71EnDVx2R6t0R6cpIXMD/hylo1a1hLdA39ShtETkE
letoCbw/MUy0u1ieELVcVKlit7/W+Dug6yAXPkPxlvn1Dbd7Z+3yySycVW46wQU5T1OEEFFI2SQq
bOJp2gkBnxi0M4UYR/LiA3zbs74xcX2m6z24Lm5rRDthkuAbNAEjFVp+BE0QI1ETEJR0CSWUrsMS
1cYHIb/XXnSHoQ7NrWCWvuPp0HALedj3ileG8ofjOcbnK6RR1cn1ykDlZq9cltZ+fwhsYohDkwXI
vVrtSavbH1pZffAbuHJkjp43qIZvYO07uSVOlDxNfDv53eTf3/jef6pZmhMMKpojisB4sAXVH2mY
wH7OQ/yunIaGsscEiIuqDgpEmo1McaCqh9fLPH80I/0IlwhfGTuI8klOUs8cP4AUeWKeTr0tW1Uf
0NQ2GL1OJ+U9DTCmLUBYuTyUBngCq8B934kL3x5fRzCEgHFeqTY1pedqfF+nGSbD/Vaksu0QwdTi
8Hw+65qOiG3iz0qybjEQ6GusIpUEfA8sbBVAKNXcAR93EKSYyFCRoDvKVJlt3fw3/b+UrIcWP5iH
CnuMeNieH/A1ORkvjGoAUmf8XxoqrzYhNtKqU6x6XTNqjmIG9rDDTEaE+SzzSUVKF7wCWnYJ+pkD
gwSxYUxHtTcVYKk8kkBA0ODfWYuGSSKmrwqxRWPLscTAQ2KHVTuojwq8DW5ZvgSqEUrpPgGJKcyK
3sgePR5bpDxUTnUdegdbDK1iApsRzSqGvPgZwMoo7fEyixUj3DhDta0c4Oii4nzqBlaAO+0Bit+F
+U7YGq6xF+URKxcpDmhlfa7nURM9qzlDy9eUdaxXcPsUEkdib7NneGmy4fbpS4g5WK10rpxXuNon
+a7K2sZUeBw5cHvsb/T3OTfKa7XMK8QsN1j0cVT4MnMTg4KhBERfWreIyTwhfZJbTpAYev5o2NNz
axWWhvKedNCQFAZEIdJAPPzbIVywcqhdYHDPhIqmmks9k90gvddOFbMR1436cfL207VumpTA+T1D
JGuQTBt8LuK30j40v+7IRwacGTkJC9jFyZgtnI65e0Y6GNMSlSsZvAoRRswmiVAJOmjVN2Ig60wm
KW1/OJVzPLXy0tShyrZi5TTiUeckMS3MYWGx8LqIFs9+vB0eNDq0D8KeSzUpwWrERNlRse3FnORy
nVuKPiyPUjpRIJGHSCPBuZRUivwbAKRY5Jv3pTO6z//ufuyThnLy3ziiFaMgEVmNK67jBGAjCjkS
esQKVy6UfNzgwol/RwFSsHgPXMS6EQNgLZ/1PjnG+0KHvuXCW5m36Ffx5q5hCjEFVmfxvK9u9lSE
C3k2s/iPhW2B7pkMDoGqe5t92MqW6qxNs4s/cNwDh9nIVQFvTfgEQM1r7xcf0CTCw81gvKPsd179
M1UzZUHXncV70GiOQaJhaq7HZfpwoZ6EyR7OAkEXU5cHUcshwUzcCaDtV401IrGudehWHHPk/Siv
pXKy42QGgUSWrQ3o/JIPyy+UhdlPzNRCDYZh9/Rv4vt1EYk+BHVCXWNyYJANOesKZe2bnt6dL2qL
xJP21PHhbcC2aX78nAWz8nXtdyT3V2DnmCSPvBiQUY71XcOCNhsB5nSk02B8B2AWGkvoCCNlXhWb
G0Ux/UVrMJ+Mi49yQXIsLHSejMquKfWgFA1bKvQ64GFgfYQad+evttcCsiGHvlXvRIUH37F61v7A
FjsEF97ye1VwG0tFOHCo9BxTz/EpctVlx0rcUJ+UcpN2riC5TvEaSRYU+fhZ9tKrVnSvZCb87Gj6
cb3ZgVyz/42kZEf3YvOtI/zyPtMxBP21HucCL0upPB4omOSxxFbDKee+V4Y288Yr4hG7zDTppXS/
e0WKBBs5iTEw1yVvDabxXmuf4md6yd9V3TqHQqqWj45XJlirhRl9GguYS2mwgRG2HlhkQMKK2t9W
U6ehb2TTHL2dVhRovh2dpkfS1cMLYYJHQzq7flnxwaVRPyUsCuDSu1zHSq8YZNAX4WyiSK6lLfs1
QaRjUX410S5iqJYHYwVjtgnVTqw5rSHGCcEP5A7oFnz8ZNouga/lE8VzsaxVbbZ3pqyiVksJIJDo
RsHRVm1fpoxXFjDQEOf2HueKYGhIMLZ+SyGixJIj0vSaT87DNrH9+AHUUSzLBv9dChx3mtGBl3Un
Xrx84cMMh8TlgWrpX1H+xwRxfnKB6KAq9Gihlf9juDEysadZmRLGkAP3Cm/T123LjvA79dOsuonC
e4Ov6LS8tO3LmF+vIZduvPQiEb7F99f5X2bmfRjKHiU4WEDOlgM/VOEmoFhm/5922fBjHht5+c4M
BuZUtHg/TXwOrLDh39vAqg2l/zfUnlXVLKqdrHFSZLUh+UBvB7QeEPjud00Ni7Jhz5S8lswaEQi2
txzyE4GuR/wE5Ak7jgPp2Zx+RTEA5F1C1w/a0oZf2fkp//4sxx8Ux+WlKtIpncUm4IonN/Cti5zU
xNp+xGuVwI/lGNOJbgtGpOJa+UFzad+HJ/AkT28YinCUlZ6vqQqEdD60K+E/KYJjj6a3QFkfJaid
zCzKkLQvQHqM7TVn2hC5gRPI39ISNQNSaR7GXtPM+Y06CDoJQQFPUpufQPDZuwmER/BkyRjBfz6D
MRHC/YTh8hGUleKb9Sqtr2Rddzl2mPaVAJ3rgzP8nhCchvIH8lz+T0Z49WycBsCG7sCoSr/Q5NSQ
YmsoyO7ZSPd0tEb/VRuQjs7vX9YyN9YdVFCLtNnWpfgBJ31nDBomefAjUbzCy7SR1JRc2hwFxI2M
kjO5FFCbCINdzRRwYGnKuxoPKzfPBBYUBXysV6sjyn4tyBWdIB9+0T95KC+vbiZNgqw5JkvWh1ne
0LfamwOVmHF6Dx9voewO/CWdOLYAD5K6nafNXBPCQQxi05VhXYxn6d+WyBsyf7DRPB2H5zsL0vd7
92kiQAoy0QewonqVz5i6xYlB8uFCjiMP9jYEWs9vDIx0ZUA6nPYg8orGBzXsmK3SfUKF0NT1Mctw
InmZouRFGBVKWPDttrNLAmo6Wj7FqpM0ChsjLARnJgj3480U+mKvfxzkpYLcToWUw8thF2Mi3Eoe
jY1GDSlyhfy1AoVtLZWGagORrNpmcYPoIDJZIaCVj3x7xneOzslEQl0UISei2cAJ6P9uYCULdFFC
PJUThF8K3kbAUKViNkyIZqiAPtdnuMNUE4xMjbE1KchaSn2bwkKpSvAwDXbiPulVoPp7yVX8mP95
fAKcA+dR3M7L0I+TpOHCAbkNrpomIhMHfxBTnmH8ty0hNcaWS5FI+ZIjThC3NNsluH0tVaf9kK91
fzzEQmeBbBY/InGQJ7GRWzY74pp4oNUngkvagzQ9sO33OWuhN8uAt0SdwM3+rdAnTBmG1eJYsxtW
ofPxqKeXXh5t7j5XFz1pTg5uxC7Zw/Gw3II7hUC2qBOAUa4sA9NDzaquobDYxMNX9+CEkxt15par
QMkh8rpsQon6HgmngcaGARBLUqvlhZHvMytxix0jzXL8sA+MRzT2elX2IRU/X1p+OUBtdEqe6e/n
dctIfRp/MfhZ7WTOl3wcoDAEHURFVOrDEOcVnuFJF3Z10hKWEQqVin5tEUn40jlDU1V4bDeHW73S
ROvOmU9uwX/ga5K1ehOm3A9PzLR+wGtH40n4Nu95LSbvYHYH/tFJz2G7tALo3/X6QHWiHHqLJirv
esUgL2JwwDEV8j6i61atSU2iU1Ajg++kTR/sCtGSZyN3uSRyCaOTeqn1iTVdOHGXsnXZptI8PsUO
W3KEXAJoVVwO4DgMWYSoWCTHyhVxUvrjoMsV6XxJcNR1YWZg/1lHP0kNPNKoGU0aehqYJ/l1DdXx
DO+vyVNyxreitbKETQG0gFhHKivH3HUCNi6OL5TQaBw/gltK2c5BX5S9c5at1j8Du2rH19IoAEuV
7v3UQxv5xXFdPd2ulIskDgXuav/WQvGwNuPQevACtn5+qsynwF0MX7NmUhxA58zi00MyzcKrIMKL
2KWi0njhxfSF7OpwtSm3SfDfNJcqNyWu0Fg/g1Nv24PH1AdsDI476zcDfk3K5uDWnD9oNVKAv+kA
P9qOoCUTD5Yf2YYfHkpnOEDce+8Rdw7fZ/OmEvMLknIy3j+h7Z5c+emNGhDLRNRs+MMRUrT7NwFP
nUAp5ElC0kfUydfw3UH60sSMTtkEOpOx3PQJe3tthaYr1PihseTbEi/O6OYaJ13UmM1OzoLvXA5T
Lnte3YkaW3QkzZJuXaGWYgs0y/HgbFRt8YXmw0xiAiBnUtXuQvh+I4TCbQi7C1a5/EXMpgBinxxj
P/Ynyw9FAYhoU4+SjR02srNDIppBng26aiwRvJom5HR/HyRzd+m7uwyF+7P1ewffRKbNqkI+ge5m
YeTxEEN1MDfhrpJ/aaLihglt2d9Y5iFHP9OD6pX0VbiO8USKGOnBqqYPNuT/0MVSrOV5DCSbK/oL
rZdtbKaGeQUIX7FWovwkbF6eJPT3pZ2zQ5YeO/th8Fp5DXy+mg==
`pragma protect end_protected
