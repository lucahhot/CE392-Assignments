// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
fw95B5NgA2b0Pk7KL50kV1xtAyOHKCh24kelyG2hYL3mWLo3IGwRJgHNxG4V5H7jT+F6xRoT5kjN
Nq8AiL18UOdb/oqzAsDoAQODJ7ri+K1fnpIQH0Noy4/wOZvM8LCS3+GbhQHLiC/Jyfo8fVtzXxbV
AFGF4Q2vBZNMi5SS9gCqE3XmoD/rAbibjTsKin7K4cTzzm4HBOsJ4j7bedPeKuANfVcpjDmU9pm1
5yI7uQAGydIOdM1usPmAIxk7viHLlOXJc2M78cWZZen9gdOi9HODu11n0IwYcorbClppAHGXQQ0p
wWq6F7ef9y+2G9M1VBZDU8ReCMCj80saCbwLdA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8304)
oZ8fDsimcaA/v58dxfRtH86K2QfIbK4QZW2FXQy95JUAREOTnr/Ow84tLtD1E7b+gm9pVClAdiXN
8vwgAy2RjQXfnAbzqn3rc34MlrAq37kxwR3Cf0LDlfOMiuY4XaBMZ6zFb9JFpuf76gnLUx+ru/Dm
neVCs+ErzjA4cAJHujgRyU91Y3QgkV2Y23IYHCME85aprH2ib6oK1qHt+Q8suROYGP58+nSBci2N
hIFR5Zjfz6I6ZUQ1Pra2oY/Ruub+1MFLAkLquGJbiSkkCh+m8amdxEIPXfDKFacrBQDbRxFU4Ktw
bzH3QijJ7G38gUfPzsujiKoBptWUCd4Zlkqn85Rm8WOSnZ/CrhJD8OMSzuPl0ON/At3n2JXQhctW
1T23b5P29VGVmeM+BSenwoFb57HnWRmR62fEcB4Td6oBd2CSIRpVvY5v25JCIw3d+KuYoJYJxLOU
fXr/ngf43UlxLkA4HdRXszENtHYdEy/6gE2W7asJ6iAlpRnhiOAzQGmnQoLqdbh8JUN2nXxYPJS8
PVQlR2KDJlohjzXv94N00GS34fUmNIZ/385uSteAx22grArN6TrvyWxTviIUPKDx+7Pvrpk6gI/c
VmS+T58VoUt67CuoutN2HVdDiosmh1xKFKbV1gZVRNI6a8zfxtccjgEfH7P047xx4QqStS4DG2Nf
4i9Qcl9dzjXXHRXIiuxT975+vDqv2v9ojFT41RegoAbS7ELBYhtrFjDITGYE0/0ttUMAll3+yGKN
x+pJCXJOmvD49NS1JgjjNZoq0yqEXHGjjyfXr2baOwBvnsGB8FUyTT4UZzM8RvcW2OW3bbW4jklT
Qooua1CdIR7XPzSMo36H2RF/dWlLZZqTI5rteF9PSBpCPQHzckvS4ZU8k2ZodXS+nE1dhW14Gxvx
kh58VJ9SwAbCfAv58vXggM+QZ/B+/jr7fAbMWNrQG3jx0C5bSpbj/ITMrLHsUVl5geFbBg8BzW0w
3RU79h3xSYVSphlTRAk1MPO0wmyq5E/1lWmwjbYxq37F7mEdb2sYrIb6iecWvyXLqohtqyvUOx+K
HpekZStc45KCwx8mr4IhwAbhhghGoZn2dYi8vDmjpj0zzu6+F8SijKULAK+gzjvPCMR4BuWEAgNw
PhpTpGkEv3zt0Q65O9KYD5E7SCESgJ5uj2SKxHBDva2UZqnO2XE5MPZS7mF5UQCExQP8fI4MMgdR
tqdJQVFl2lvLHIkWVVeIElKqpPzoXj59BcdsP486eMrlWkY778rb8RU7CDsYbzwsX9R0aFj+yalf
pOcTOu1Z9NL+G/uJIT0ojIqLPu4Ivkb+WIlrxTMOES0uD4vROB55z8I63TDmKkkzsTzJ98LKCkd2
oXAXgcButMC/hs86Ay5b0nTkOinbV9Mmj+Cv0LZu5xNRv7kY+I6MgLVi119K4K5m/LlsHjN0tm3z
buRFCrcu2v713xiDzdqkwybW2Xd16ERdSAdiZwt7StrOfoSDEquZPNfxIHrVySYVHucAjZNpmDI3
K3fvM9yQJZMRlG9jR3etMsf0oFeROi0Qjm6LnNvN/InRpzuROHSUgi8s0iOoOnRKqMwEsU4MboqM
0q9/hJgfxeOFieg9KHc7xwrPmekHPTqKOp3nIGHEOl8DwJzHrv+6pPH4c21TMthIpbJVGzG1IHqG
Tm1maz3bgiFDpEh1RUWyYtRSGYlpfBvVzk5W1iK5s/wVPCUmuGa82hjFdJ2cqxb1X2di8qnCbBo1
LEgus6vRt+iVd6xsN4k2aN42uQcFVm8Js6kIdWXH/6/rRJTnK69q89x55C8uwlS9KJPrTsmZPO2F
rSvrmEUmE0DYdS5LgK3Jz3ECKzdEMQIAZI/pN77VlouOYKL9LwilHHNN+MhJ6n0tWnzqdaUNyaHX
jQga7HOf1MjyD9OEvHgo/CCgf+FHgErU+D3GJRqU4pdShgH8bBETBR/D+glvy1GhYQJxw/R+G79z
miyFWKQeqIAPWuUacCEm0ECOz5CQtaRVRpf2GUOhnXx+PFC+K1BRVx2zfOXRgF6KBXpigaUbUGDo
xCM2qltKpHxA9SAE2sHdS2mjmweLqFxaS9UJZ9nMljGQB1w5Dmg21LPOOC2W7X7LrUvhi60gucvt
iZmZLxv/fI3D4K1siwqM/W9MV/UZmvmUIU763kaXoiDFBh9zKYDMFMIH/+WIcNzyr0ajcVHFPplj
V6lc6VBige1FErpEHRxfBtgUvWvxBU+BVS1NGnZNYVb+O1G4XjfwYlMeUssj9r9urrNeVqkZIkOP
drBhDueV0cK6598V8X94dqrwmN1PgAiFOCswFOoHwidrJ974swJSHG9VU3yZV/0R4Qgz1fm5NjXd
IrHggRcSteHkBARU2kwLqy2nOckvO+TacfLkEmiqcTqkSS78wEt+Xdow2Rjbp/G9SuKcUM6nNiyN
0e+KYftSSd/V7z1OGleWq5cF3/T0XCo6ddhtS00L1cSjHREJCPGh+RsdGj5j7a33ytIXF9bPAZyD
592niuwrFyhtzCSWjLKe7IraPZYsThOSxgAWcgv9kWp/9rpO/EQFaDuOI612iAzo0ds3nmA8UEer
8Zv98RL48I7xPgqys594UA6h/g8wz6nTYeATNFfMf8evze/dKoWrpPjvCsl5LRTtvQZaCzld27t3
5mus7esHo7qvWgAIut2ddCpHSfO9U3TgZTgYGpmfWSU80BAGY+PQi7fzO5shP+kDh0GVjIaihfpV
3iUwAnPnaQIEeQtCAWd0NZl/BMo7/Q3dbKrbz57rT0KlCj8EFI5CjaC8+bVm3W0tDZAJ4a2LdL1P
lyVe1D957/1kbt5Miz5sNk9BOEDOZiPqvnCMFiC8ScF6dM/Md1g6YTDn3Hksvc4hbQcauRlFZMP4
y6kgZemsLnRV9IVNLzJ6h9sexCoS6aHpTUbKUvCDzCxA2OPXMfRGMyAdHXzrqbNqEKH8fqhpR4sS
8qduzEDP1+F+Luq+9RIWOfEhAgwy6vl9E8bF/bY8LK6JkOfrHHKuRTY9xAGa3I/f3+sxELFzQMii
TMh6KIvHBTBDa6BafSSztWZ8B/13ANtVv/hKE6tCSxliuVido9QEbvqCbsBBfO7Qns2aBVHiLc71
8QuGi5zj4IbdwVz9ZnU2xmkdoJvaZ6PaI6vjxbdfDWu3fUqtKpsuGNZ/iCdx5IEjkuEB2ZKoBX/e
9YYiZlfuX2nEsO23OqJVWR72KXfubXoMs0TUvVZJqfyMJFEKT/7QwRhG7/jDHfPuDZolXiPUUqrJ
Cr0KPKLQy8N8I54j6uuZtFtSGHleoSVIdP67tpUMgqd8dubL3MQrZVaMnH+plfcglXV71gGZnfbc
uyHJjnti3YlgOoxHXhYWJ74Os4cYlpyjtre67ehYUL0ibILlNoP1q+eI+ZNrgZhI5Kj2zlMUZCBR
f2rowbnW27wjlQ78Eugg3bGPJUASWRbkSlXcTTq3NetKNXx9txmvJD0OU+7oZJ3Jv3rQlEDY6r71
h4Y6LgaK4zQ/i1giYaP/VqXVQGQc+1Fu5x4n3ZYSEXBeoyT4A5/19DkevdR91X5z/dtfjBHwzQ78
dIUPCm363o4uhPFHDH0XWzduKjUWuutAogkSYwd8zmKNMOyr48pb6CwChjTcucKbyEOrl8C91wFy
UqBy/IWF7V5zpmBTgv5GrNNCKFXudUMswUpHVyMAD6W1HBIDwe8++wD/Ba3J+KqIgkhpQjnLDHu+
TOQkWJfev003IWC9j1p06IFulQoAl7reqO3wpxj5IUVPWc196SHJmUyh8a5/Fr9AxhAs/iFCTBjY
yRmIqMVQNklu69bTGAyUat7Gxf3ttBDJ+M0fjNhlgEZYAQ/42aQZh2RYHwVxz1GwhNOIknj8y+2Q
N/sFf9bulvByIuQy9F0dqwtS9yPMYjF4sAReeUkHJAAhRPGAwffMQFDzpkp7tt6iFlOqnGxTyYAo
mlXmuPZIu4r1jr0sq0qsVhGXMrvF/eNG0NA+5UGgvtBObZNF0um1ls+AEOx7oLeD4/4VclJCkK8d
3ODgrqRlZL3yOo29VQOPo+LhGZnkMyTekgUEqcaw7Ff8nyHxBwmxaMw3BEzLQPr8ZCfz9tedJQa6
DkDC7yPh5nTgJ7jlc5Z4CflA+t2+SDsfGep4rZL3xIHFUR1A1EwuEtB6LV5qNVgbn5w9ARE/CYPR
32ki8xLNjlzV5P0y4LvWcqXTszzSFjVt+KvUg6FpN36kw3XvBZRkilhdzG5lFQ9YzwErw3mQ1sNA
nrCriN9rKN1T5mjXmduJzQ7GGUOJ3OMFqZDKIOFeUr42dgSeHvB546PDZN3FpsaXe3MHgtxrPCc9
UIyaH/l8LSyLjVx1BhVGTuyrQIyz1f/8AKxnah64Uj6hEriVwMmbZHExScW7onNHGN7/qlYfH51f
hHOwzMEZj57JuVRRHkjDMg+iDMYXjF4LDyFX4V9LcQNhTH6Vli4pfZXfj38Wt5KJVtF2FVz69QoB
UTQlZjceU7kldnI1KkjNsR+U5AIDgp9CTHxy/O2Lwo3E79S9d3TsqlMIjD8Jt5fWDyFV7AP6+TnK
HL0sCssM2uGnL9Uhl3L4k/79AYcnsaO+SH93udeFI7B2EPM7eFK5egLdkXUIRFwGCQpu2qFWxrla
swA4+FIA93m8sCOlwKy9u9U3gft2dZedTf83MkxSBCX6Kb8An9Kb3obSKIXTIzifK42PJLmn85MA
38EDGrEblJF/sqmqSx1oaXm1s4msTVgryCp+Zccwj4ip77IXqrHv0AECEEt7ZWFRDyNGkaUNswj1
LypWTOWV6dnSezKXIxcJGs45h+pl8MRX0Qneb9gH2EF6yVvHUIkvU0b+jpKX4c9epC6PfPNpBfmR
09BPdcCdq+t2BXAmJDaZxal6c/AY4VnFk17Pi6IXjVcUofSxCSeZTDFfAqiB/juO46fcXPD0zl22
3kNdYOeCbqT/LQBKTZIhDMQUSiy9HHgg/C+ZihOPww9qBiDVd5+uC1R2TISYNMaTsFc1plzAmHui
Zs5zDEmXXT7krT/PYtEu52UmKSf5pOArg1BeOZlfLXqypsbZhPB4VXqwxOZcK5KtacJ/I4eDEMhc
HeroWyRbl6sx8VGTpyaYdzpwpLqxbrtfqp2mf4tDkuKfESK3fVwhZOCFs4YxhtTTBEdIrPWOiasG
IvgwRTe4TnbzMBLtx5OuqTJ2woO7aOZvhq2mlnv1CsecFZ/96Kfa+1FafXEwdrPIoJpIWrGU9eFX
JYBScbvkmOE1ev2gtJBem873a7FG0Ws4jTgU9bmRLnAJWqF3QVFlqw4Q4DVRhp3W9ZxiGcF6SQPj
uS4N6dGvme0XZ8TnlZ/NutCtbA/o9HbOGEVeQ7y7kposCdgx0cQdMh3Xh2nBYrXV+zlQZhDEhqSK
UUvWsPNky+IBAL9V3VvH7TCWlseNk/TrI2pL9adnndoPoizSjYSdwWkxJnDmKojnc7Z3363l4xSO
C9H059+WyLtHDmVLny5/nJz9QvKmdOLZUHoNA1IvRV46QVW5H6Jd7CyVlma9C8l/SpVeKjtDguGM
+SVo3dXSj7vt9h7EThukLSX02B7iC5OPfRXra7byu/8xd1qquja1iJxqSZAGDwqbmzjG+QwmS6co
QFjdST8MI77j5mU6l7F8opLlC4UDM8CxXwPEOncOEWg0Jk59OB5M+cGSGVktWHM0q/OXomvHIBv6
eUs3GJfSjFBxT89rPJChEOOzevfbxsKAz5W1RNfwwYeBIb7JWasfoWJwwTnQgWRnCF6RWJ7RPLGj
02kXDB/KK+KY9HJqEn1CG0CC6QnAreU2z/+/YkKvUdDgfnic91MshFELcMifI10lUtPgFhhKI1RN
4bp+CaYydx5JtF4M1xbk/BoejdMUNOYzmeHZ/mfHjPUeDIU0+ttNuyros0Q65K9fTzjvVQN2NYiP
qRg/e9iDrdoUaeNpRGcy4mykRbJy3yU3412UgQ0oHop2Ayk7FUwSuwNqEHzjLhBqtq+vAgpwOFGT
PshNQHYHmSjHKwuBRBLlsyZTnObDSZPeupqIg/DPs/AViuMRaUOfQvrCgz+JCl2148xd9S2gAB4U
sd7oRllE6MDWGrr0SOvGkFy+3PbKgTUvc4vtD/Lz0SrOphk2a09GG0UL65OA6NZuey1ZwiNQhc/a
TYtyuFNcqVtFsCbw+JIR9p0d99k6Wxl6UK+DaGxd7xoY2xKjXbeEr2tsxlzoAS9N85HTXAwgk9SY
KDruil80w8HdZ1WpOyX05KvMHlAk9PUawK7lTKWDtBNkgq5rT2XHh/lKR6WraegSygrX8fGN7CNA
35QMYYnW4d2OBsYNWL04iMUED+ubBeAX9iMwX1EvMRAUHBWvKmgLr7Gm/yXUqD0S4HU4FVZA64Hw
CxLa8Upr0iqrRsD1psbs8qtQAsbzaWsvzehIuZzKcI0Bh0kptXEPsWIDgFxQbdKbcgN15S6RYBGd
0YXw5ebwvpFdPhpos9vdU8RPA+6+7ByPmXNkj3iauUFDeQmeNmS9Jh4oVism05Cb4RDO4cgJBlTU
UFwabpQomKS5CLdNlxwhzn3q40zYGW5CvLiiNInQkHKAgkeGMrC8GD6fNhssBeUAMaHp5gD0vWJr
+U7+BWCko4UWX0Rr0U3W1MJK5HnXg/uLc96fv0OYtMAAKGUgFvIgXo3rtcp8yWntGMMLBPGgYJ3s
YqMUyac5JT1TpIEqIbq3X8qtjLKwKPgX7WGA2x330NuWX5W2pT8PsL3qsxVE+UiNwA6vB3tO0KPz
MrodMBjNDJI/2UrVENsJxRZXjzNbyncHJWsm3HdiJGJs+XQBzmftjaHG7TsB9TJQbjmJ/9g3H6Eo
J6vaYZhk9elvRR1wPzMwE9tb9OhE9Sm8hTM3Qg6yyVJob4qy/rOqld5cAFOkSIvBU3vUHvXBJs4Q
qU/Vp6JVKkjqwvXHnDQrltkZ3VJKkzzB2v5WaBjno/KQioS/A5SVbmi8iOALxYcUb86H10yQEhVt
uC4kExSa0KcDoYeMEDpuFj2NNq0KTFbs3JaeSn9eu/ln11k35qlVXcuQLgj3k1Ay++Y5F6MmnKpz
Kao57c9mDP14hfQzQ7TxbaWlLTxFn/sAmVUrOYuGnd7rMJZQ8eSdULNh4F8spRLvb3gs8azT1jxG
rw9Tw3AK0eUkVXCXPWgae3tJilzNjxnHdjNsabCyDWmcbtS1rA0hCMohWjc3mglw1zKYxAHCmzRe
GDlhH/ozPvSuIB39NQ5eoVBhxl+rCEXNrMB7qfg8K8MRION0z4QQK3jXDMRLPgzpJc6oigMOPlST
sjRkDJsi5hN5n/iefaiv9F1MhhRbsKnot0HUCV0YCeiq8pwH7/JWVWbVT0Ezi2mHVrM3xYFsKMYZ
iVvG+dsYgMyZkGa4qhXfwgFsMROTW1wta6K4BEZN02mYCb7QWB1G09kOowAsKdxD5QXQm+ZCVdTr
xS9/YwbdMGHvpy4z05zGYTK5I1XN5+9eyH7oCIFMsmm9ddzNwmWVT8Z0IVLrCrrmevY4MoqVMjto
trdbxCKONdZJlr36ixPzS83/rP4AKgi3HejnXt7vPKz04Cg6S9eQ5bESEIDl9tAL+kFCUrzSusTa
eKViTS4/Cuhl1NFzyKAv4UiQeHNDCWTsnQSmNOmPblyUgAyGadnRc3spgyQ9CgVwOFkxpmbABDth
bGKbWJQn2vBFAwDFnZReRbass5Zo+UDfkuvPhONC3+KJuBMYI7rpswmM2DNskc0mII3CNw8VFe/a
trLPAlj9lk1RFFfzCqdP63j8Jp8lNvHygol2ThsXlbfvVGSLwzcBsBXAhNtRLxyXvxiKDdaQW6vD
sDlFHz/gVEU1POXpAcsKYyg+jxIUaq/+ILFJTUOb43FVy8AugDpLPT1kpjjHTLGKE42reHb+wyal
zcvi2XR2Dvw0OIfYibk47T8gdk6nQNk8XpkVUrkBC4FDJAAd6HSu7JaJqHyqNFusvIl/jUFCQseE
CxZapeOA1GPKvq5OkgityB5DN/ZjU3QSnUXk0CmgsjinRGkmn++0/DmjJjj0SAOkUr/ALZPREJvS
Hvgwjjz3ZySFaDXLQ8H41Ci8aa5+s9NbOtL+FD5k50UGLNq4JSgWQw1Tr/U8lZyilivSnJcjjNCe
FyK39rjxqfVou1HL0iwKp9ZoNnKOda7qEEBfWDs8+1ZLTD7RBjHbkpP34qU9PESUoiCkaAKdeqsv
BE3Z6gQGV61fDJF3CpWuYMkVO9SaDDhPy4pFXyn+3jfa7siJ7QJ+SvG60eCAtl/kfGPi+FYph3uc
EG0GNz4b9tlcndbBAgZUqcDUnshzHU4qqEo5HPgmxHd00kDDRnulCId7K/1UNrUKViMmiloJK7py
5MxmyhN5k8+ExueZmeYGTz/wa4lkJ3dRoUYRkfJp0sOhVKbCaKumdJSFqjHwfk5EIoRT/0zewf+q
AamTvkppVeIL/772AQh+upeDlQW3EenVskU1BASAzf/f61tB6mNg3bu0IvQ4NdMTBbE6xtMFbEG3
5n4UFPFbE0mhPJMhZmCrqlLswlU1dW4ne3jKYiEAuZa8z1s716zRAigo6/HOYMPTeby1Lecd1L00
tZtdJq7Oc1rewSxNxqz/8ZBZN+5Myt6oUFkV5tlzEpYXQemMXuTmlIfQ+8leXwwtsBnyunefzqMa
30IHJ8wjCsPXYtuVm8k2nnPU/1Vk3Xb6v7CAqIDWum5rczOeunbDGTIC7IRyljauVXCEMUJgamDg
0uTKXxAfqUkhKJ0v3TXafJaE5tGh3p+5QReZXGf1aZuc0SQB3AoKn9XFxNMzfRiHHldawXrnFySa
79sTY63mHUMMHflO4l9uPKOmZlUGuNdw3UJYuaPgOYVE+Bfstoedn6ml8g9d3rbDY/sgc2XBRAC0
/8kcxrYLkt48yl4o4jFpiBZARTMW7Eumvanrcp9kiTrl3dwir43u9byy/OcMULJQAMh1Lp7MHJkh
eZ4NI4ajRO5UlF4f171IZJG1/6Tdkudim/o2i9AYJLjYDrCwXIrtsq/ZQTI6ITNXjS2sZ5BgHX4c
4AN8Y1uX2ASRIS3j80AMmWqNEZHvKwOSlyLsYUzBhHBpE8WURj+PJu89oL6rjy6iPe9l3MuUSe1/
q29r6USIui7OXSGSRAkAankIoXjqDyz1CzJbJgusQwl1JPjYiOQ6VXWJosAz5sF2BAAkeU6gTcJ4
Ndl6I/6qSCG2O03NEJ3kr83GU/kMWCYjv7QkpUbPL/9gx7XlQllJC6modUYqurbCs3ByrPtp4TTt
kow6uiQxdE4+Dxxo3pD6yoDNoIpAJjnFUCuqqkAOlzr7aZqKjeYHqqbzpV6WJNvkeMpvCpvbSDw4
DP1BS0F5HpNAUBGUiNmUkuxYPTTxaR8P/MblV1dys4J32gZZWQhHeG1OCWzALJCs4iYMpgvFPL6Y
ompypurJgIBat53+kjJGquET/rk50oX1RRFaG2Yo4st4jnCn3t8Vhr1BuyGb/xoIPhO4Rwyn6Ak/
N8hr1NLyFRS0abSOqMmpb8FmNM2lNtfje9hkVrFaumRXrupYrV5GasKgJn/qz/SFrVhGdSOGQrcu
BJfm9092VeaqQmFrthj8PJmXjbc/Gd/iwQLiQwRtLTe/bdnHE3seLSSwnPeyIex7q65KPD7fwiRK
CrukA+nbGyFL+SeXLMdBMwfxZiDadzAhIHn1WPsZfnF/7tfm/YDOsuOWrOfahp4mm5VDiWXP+GWe
A5+nQ0Mp9n9BPW+4aENVKsLTwqXaXJ9iUGoJ2jSM7HLy0mN3eHSCyXPUURlozG8SSCjpZ79tlPqM
EcDKUzf2TsLOFyTxR3ik8sqypkCAvtyI/tUU/XgtW1ZkOTUzZPjnHpGuLLse1Jo9Wpt/nET+RrST
2K3OhRW9FZAfyFYXncy5ONQVrH95b5xF8TNpdiC/J44z6P87XwQGPwd9zB2vyKhQ//TFCX3Uc/a8
kUdQ17I4eZxa+70RrfcIOSDyoZr0uEDGVHfFlAym0Nm9cHv7EzOy9YztQ5ivxfFy4FTdTV8UaRKR
/lASltBbgMKa/jVUIjaKssPr1uF8iYkKxji4WTeLJ5I0kZqCRepsqiZqnktZpNCwP0J7IN2BKuDo
jItaMiBuE7coen7r3K6KcGca+hNrVU1spizLFaGBM2wFJAQgw6V7bsrX98vz1hs009OkNgoWIune
QQUWRBIbXm9grbFdRAGVkor586zr/LG1VpdyN3y13P8z6mYnCs78JL3ZNIYCYmh/+E3mqIc7eqWW
EpWHmsfNzD48IQcMyIUfWfOUzyuyg66LvtX0BwRxhxbnHGfPOqmYsJRRaTZQRkV6y29h7+wBYzAv
jsb1f0F6bM80Sj6fuUqEYWEuT565rCzrvAvAtChF47oSgTgobWU4ZFNmdZPDe0JNa1newqxs4U2r
DeX9GlqQtVzFGVRyHhMGZ1CUTuSmwjTVNIzp9c+/td0ye5T2agOF33j8S0LNYtGLPm6BiEmCF3Bh
pgr++22NRDzKI/WMgWvw7CfPAtsjJR7nuAOSE/YeKgMmLS/u9vFauUD5+VKQWTYg+aapciT07IDH
ReR/Rd9EQBHNst8HSBu9t1eckTMiHCRTriSgWkPbm7QgsY56O1knz6/hmwpBYlyUKIyUDL+ykeqR
heBSAVsKiTHTGWwdVRid3dP8cxTXwcK919xt64X8vwC+RpJAsZ074F4h7E91tPlaoDNwZE0hFozp
+DhXTfoEBwTqA4wYEpmp2aR+4+Pp0AOQTWeOK0eUscmySt5UhQlo2cJwconnQrrZsfDbG/Q0cFyU
HKarEUdB1RnKmdHscdySRUA2NnT8qjHkEVWVXhralrmpE9X58n9MgcK1VV9K8fw2HqVKrPv7c13o
E+1yOqM/u9pU4Of3Rf4DpZclyRhwd1zEKuSM9+dBgwDJmEPHGEsjyD/1vRa67zpc7VEiP5M3jNgq
jGNBELRofno/uR7j7DJP2W8w6RcAauueociHjziWafdnsSLSqq9c5HLpHihVBoy5hbrOMoSYp8Bq
O/4pz8fVLi7HUk9V2unOL4E1c5XajpedNnjd/G/Bxmekv/SgY6hK
`pragma protect end_protected
