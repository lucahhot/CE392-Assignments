`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lE9V58aBbvAKPa2aeMgmQ6PBjjufZUla8UAPUD86ei/C3uRp322z1FSz8PxU3XWW
wb8/1vt5c1VS5egoST7u0YuCYzGnLSMSmtl7LKgxMEg/ZIHdnieekiO4GWZt+mkA
u/YzZt12ER43mZdaKipj4gtWuFr1KXBu1CwmsMVPe+o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 91424)
jQ4YyOWconVlIo5r66TwPLEfzOXG26xNAEheWGKq9YtgxQz6zbeQoeHv5eWqFemo
Du7QRt1PaPrAZQwKDJFhedUEk9XM5khZs+SYie0Q068CjsX6Xpa2oYl9syqvSpDV
euWOlrIwEZKLRPnDOSh8F+02l40VyYbSI6VS0nM0PkresqtliVJ08dgP5+1XVHBD
VM3KlPqC1SNG7CiRwH+BVCn08pg0AjI0JpbYbDdev4G+rPAGVfqcOWrIiswCqILk
XZ3aBcIoO+74crEUrg+uDSMJB3l/sYNsmUKXLWdcHQzbff4RrByqEZsK5MqPLY8L
AY5BR/6dquep3bJ6AN6VG9AI8f6Jc/LxkelJo/qTNOk1ScokcQ3oMul0U6ArXZ13
N0Oo3YhAxc2FT5zlWUkN3lWqj8SnZ59+QCN7IV0wXglRFmdhRffp/0kUTtHtEiKf
2uBNouJQH4OLw3UjwjEoF3Dn50kMNa+9ZrJdxePToRB2gCG64htYas/fc2WIXDjZ
3giyvPu8FdRAfwut1xAHdElcsNfdVgEZ4qhFV7ElABy+9uvQP4Cp5kiwmHOvTKDo
lSAUlzu4z1g9QBY5GP4JIoRAr/+qKeCt53TkRXUTq88WN6yyq7eKD2//vpCpbtHD
5fxoYLX1YVVKmy+UWHHVXXLvhAa3ccpW6oCSS0XBlPLRPPt35G49YwWSwJXA5xOY
3VMf6hFqigUW0MdDgH1j1abors//u8PJyBgifnKMDozdG50jpXxDuQ4bu7tYgl+t
GYA4tXS3S9btuS4BLzeTbta+/yOhcrsXSFPLRRj2MCd0sPt0OkRz7gRMvAJsMoB2
ZCz1MaB66wy5ac/m+QHYKfQhJkksPTX9oiEolh1kGhccnzEO6KvQb20Wxa7PsEQj
uQOAQfoy/7of/ta2V5n5LjezLQrbf4FoixHuO35On6ArveZ795H+lck9QnQuCoD0
VfclfwVcOFiTV4InxFM/ajCqMvV1Go2Z8HlFICYhef4+A7vzHbTbmlNIQyVNBv4p
ZY9hNATqkGPNgX6S9ubCZCjUfo6kBj0EZXqnutyvFNPLZk2D0rkWn9V6fwyID3N3
rPNKYOhLW+wlpTyJkygA+JdSJGJFHX+TPHINm9os5Ez5mVlpwFEY4m/IG78+4bkq
cnIJ2U8maeAQkvabjGjfjj+9O8aCV1v9f9JRJset/aDDwHHVySZDL4UJr19b+Tso
7jara/P+xvy3iuHiALETqwBkK8dy6Yj1Cbppvryw6VXjsh76alVZuXr1C2SB6kqJ
9TiFmJrOu4srRslPnx5pKvOLPI7nPDDT1LgOZ20NgpAOr5Z9q+inrVWHvSJXZA0w
vo6r8UxjrP7AMvF7Z6ZgcxZvLURLNXbGoyVX3IMO6UYO758mm6wpe75KtpL8oVz1
Z6rKZsxabe5YVxyixADJH7jtpc+FcX/r4jR5qfCrxpDeAkL9Knf2FYNXI/mMWjhn
CiYG9ahTRDQTAMfbVj4TekMKzDEK63OmuChqiNRWBR71PI+A8ER+hOhAFrG/PyCg
yRxGXCU+RU5RtLecMgHMoIL2xWbGB9xtdnS2E1vstzOn9pfM2OxFd2pRCAycS+ks
l3kS2/bfXISKhErLB3VN0WziEwdUCgCifn+TSBhpvIgmP+g/G3QpBV4iBiNnaz9x
N/m4TOciZ7NdSwU185vMgM0D7/qUVoc8mA/RcBIIYDE1OlzFB4oCCXr/Rtt2hbLG
Kkml3/ioF4Jakyx7FaeE9BIiXE0GWJSM5scHuNC+eNrthPVUg6mRPLuXodc69ZK0
mCVGaBgcAeJx4VwURXAD8tLSx0CUdg1uQDsYXOFMwWz0caBvcbz3mLa8u5JTzToR
T0xTDuECInQ8zToT+ki2Ot5aR20DUJ+3AC/KciNinHK5ifEhoVUeY4ChIVXG/xHT
R6NskE3A6ZiiG6UT10S2juZ+Znpzb09Io2/Xv60ClCRq0uGq5+z9UAPaUpt3gUMT
c5DCAupDj5akjPL0wHevYMiUqwbcd17ivHOOtq1pWCxkxISy6PrBsBWw62uanbs3
tEzTYb0R3gyvpoB0E+8jT3RLzdVSTMNmeN00S9+4d8Z5Nwj4xKZD7dA7tgGSBYm2
2r3B1nSmFgYTopseC/3F5ZRob12S/DWy2Rf8qp5SIlmbzwsmop1OaW7aL+JvNgb6
pwd8lMa1Avf8jk2tekxODVUuDXATu7rCwiKJyrB+fpPG1xtIeKbjwCu4hElEEv5w
00lyOb61Jrjm8EtK7thVHiMEGRwZcuHKnyh1/Om3FQIdYLSXd+X0MyZ27ap4OAhe
3RcIFbpxtNwolUmtiUq6fxzfsS5NIh0Jk7Ugx/wzD8OpFHTjC9zI3jT8VLSKRCpf
syIb4XqKFLhxuOfPMIrm4bHuPcLodwHoudWKd7kBk3I1vv/catN1YnYU+mWeJZ95
W/F3ONXAaOw+DnuO1WvPitaCk7M/gNteu28ZCc6LLLV3GiMZ2mGzQH1PR/gWLpl8
yzr3+c05GK3CyB14pFROmXyCVd+FaRNiRaDNwpPSeIE0h198lS2LT/1x9Slocd1x
gxSBimAj5o7hNMCpClMy1WjCwDU//PXTbuie9FKGSg+0EAljVq7Ju5exCrU/w7nC
Iukep4SJJB9iIhMXyBN6QFlwnYjElO7Mj/oODfuzfHsvIP/okhLFWU5kciDQwixm
xWBeHE1YXuz+Kjrg1qD8E5aHg3eNHhIfJlFclZolHfQztxDdWtkhgsV4YDDL6/Th
0+VSMPcmdwB+weMptBwCVjIyCIM9rRoMoTM3EKslJUuWCKYdyh/JZAd9KEcMjDFC
VXDQZafn8+3J9yrFU9XB+MXrkOpflKMvp2ZQMSNOXjufi4rsv7k1HznHDQU2JJyx
CAy/TDB8Y+hcjGuH8ZfOVwxNAbZ+U1j66cHtG8pD5B2KtroEBpkagmDP2fVT6783
3eP6QC5O2ZoA9ql/VEdQyqyevN1scuTI9yjaAdBFAX2Vo0noD4+GFo+p1clIQK8m
63zSR5Te0dBjkfyHhBOkTsgRIJnflgP5DjYMQvwevkuwSKfVUbIqh5R6unWipp9a
5Gzi8bYaedwlzb5EI/zy6Xkv5Rk1bXyPZDJfZcR0EoiCA1j8XLCcgaPgt7/7aFVb
TonoVefL3m/IJCYhXKOBi2vceFm+4UxIUfyc5zycVPncG5A26NbIpoUGc1p6GHCK
1PCBBC43kXnj6Y94xHIA69L6ospKadqij6MeJK5d/jfSSV5q1cGKAt5el9uDXcgM
85gPQD+ndZWtfk8iMLBmplzLAs5mnTCXwt7d2SE+3f7VHUH1f6blOSWgzDh96N/4
MPetENIXeTtuOg3yjzvsbiFbThUJ9PAR1JM1InNLm9M2hmiSWr8lJb7eQSDZlAKC
DhUcZahlc9zykC5dfNLV74txQpZt5y6qBG6sIoMQi739QovdTgALTfeqkmYzyuKx
x+DKS3F5G/ct7fkuxj8y5pZpENOqcX+xOBE6uH3Xure3haYpbl+SRuySnmDW5S5j
z8nx4DQFLT39/ZoR4/PPj8/bBhCGz+4NQrFzKNQ3G1wEDRNxrcMVI0p9rGOytQpw
jaxmtVFabVSVa1p6frpKYAu3WCb8mNmHsMhHFjVts2MxNgHkj/aZYN1NNJlJ7TcF
ES9sw6T3c6w5bxNqurPlZh65l6C3AParPEI47LJjdm28PaGYAq7OWuvGpY1paSqi
22HJDweAX1DudHj6jFcBqRRBpYeDEhu4ni5xuVy5wnPbNKY2egOSgHeygD4pYT87
HE9INCUyz9dEKSEO/4UetgGPXviIEDWtgit4ozJ1uSeuUijmNR3hjf82mRMfhcEU
y6CoZ4a2lnzurAT9QFt8oAq/5hTD/TTy2pg+88KL7Pp7j7MtxgIeRd1tnqh7MPU/
dGYBPKrPzFikBlz8Q9FzMPRRyGff+xm8/qRaCD0OSTkGtmuxH56tzGwsDiGKmXq7
rAoU310nIW4NNRhJ104IwrsD+SoHjz9YzaPkr7YbxKthSYfXHfu9ojYFOSedWZcY
P1aqqf281/79iW12tQWA57DX+WFLd/ZqvhsPV2ExbpPDiS1ojmN4GTAmv2ouGiDw
pPXT5WniqR64l/yerfEix9pM09D9hL7capQuP3XudzB22v3ROEB3kNGMGN3vaGna
Ma5n9BaTmVv9eOiqUHTVh20tS61wbarlC+QnCKBn0jFru26eivwXH832r2v8PjR4
M0o6AzSMD3yE53mMC1Cl0fm5y0/DBUnZw6DPjfdEePm5yZIT1lvojbqK1zHBpsVK
Fu6qv4ZrLMwy3IvYXN97jNpjDPbMfedVQLGOMLjHaCtk1Wp1KbgpKYmJTdrMFsKN
6ZqxuKlXNGKOKhS4eQMuDngJf7Z3dq0N3HY9La876AgU40I0qyOu51Bc2uvRAJ00
V2/mM33t2Jd0kjc3sZLxhffSlbEVScnwu/e1UDN+7xHGbiAsxDI003vtFJBEIMzj
U4XGmj4tO2YlsefPwnqGuVHbtKBeVVyYolxy+hACN2P8CYuafjA3xs4QgJOmSEqT
/jMjZ6lZ36v4KKZNyy7O+4CEWZEsfP1+NzgOkftt3Z19sMjE1GB1epJZI/bNOQjD
xudz7a6SAN0NF88Iq3Kaf/HVrmdODlcM55ORu0LFCtBL1Ljwg8iPXCfMTIDzRwfP
xuBphzEQj7rBeKTk48OittnXov3EIg74Vo2qaYPtaQ1g5dtuVpN7qWwCxSXRQxl6
iNZRw6F+1bYLMtqWmq6kPXPWJy44afLsPubOLNFn0vkDLIKrGtloA9i95Dy4zens
qj2dg43S8Pb4ZJ7JYzzgSIY2Dr/esymlfnAHg8WhqPd7nC/o7287X6wd5mMxghAP
odV9p1OuO+h96NOYKCNPAaRRy3mmLbhqd6olkQEhswr3XT9j64pdnY2CseMLqEIO
xHM/51THN7r440CSbhnr6jUxmQb9MweJAqnLpNnFsDdweVUBV9hTE9wSw+rm+HQG
VL3dWdkoIZwkWgAGPaHkRLHq3kbHyPX78sbbK0uhU4hnF3R9nwzmi0W+sN86rF5H
K7nXmaG/GTYi2JRkcPtUEJjXudzFQ47RTmqjdO7TADvLbN3ewCrmW5+3D4UPHzmN
L1MJY1j1hnKALYjxA1W95sWAKr5+qIMf++aIhRVuw8R6MDlLSNEEk4wjEj+yrVfg
unxM8VpEPXT5MjET46yYR6TQ5jHY4WeuQTOM9ZATl6vixFgvFgFes6G/qGiG4P8T
0U0R3+ZqyGcpXsdDbSETxKEH3hdBs45wDN2kS21+6wX2FgiLe7BrarIXkDvv3jGs
B7ahkBOr7kUzHOF0S0ViAbVtsbFxlX3WqHkEB+fwKfRRuz5xRtGZQEdNqgQeYet1
7oJ5LoXw6bj32FQ08EFp6y4F0rnTkfzVM+r8d4i6soV+u5jTACFzf37Augtk9cxO
gpWhLOMYTTGUkD0m3F076Ga+//Ie/wME9/5hTbWU4odPBm2GSLTAfHRiPYMVT0FP
ESuWxwmoLsDvetGI4AIuYPsl2wXu/Y9nF+hd6eRuhz1t4Yy9CJCIT+NrC7BANtzY
TiGFT7l+PogYiw0UeIYbHbuf9PEwQHbk2YNXhsY/T56ZKkEBD7QLBtYaJ51dC9Qv
umlJE0WDSGur2mri2E3K3h+bW2ugOaAZpTaXzd5sySahofESIpmFW6Os8dv2GuFL
UMtHNLbbyEfrdUlPW3C1Ltu5dhSQ5yE3nohSqnvCKUxBDM2FfUfcM4DsS2p5SdH2
BRg2Ugx9vxx8U4UyFUlD9OczJaf/gPU6GRnUDlUWSNtDN3agcvPdnl+gKP3gc1lm
/d6K0z5sx5SO6qE2DVpLwXxaAQIJ/KLcekOdn1wAVpFIlRPKPbMe+MSrBCR6tAaf
Eza0VXkruy5QAa+/im4OHScd6nrYmGxNICSCRJTIgBRNI+RfkDjP66hLqNinLpZg
0qFVJh9+bwnz1/2I/0xZbq6Ye+DxnX2tH+17F+0dkSBNSmG/zXBX2fIoDE4brW4R
6jwB1yePUFR2zMWXjAedxWMh6BLZZrZyjpcKmFNLp1Y2liF2s5NMOJPURvCiOvZo
qIEdvwt2BlZLj7n/98VAOxuDrq/6ePPmzlbjosDY9VZwrKP6GCq3yghTh8dW42A9
MQa0w3+LPaihs9Au4tsKiekBoLqzsCi5VY0ppo80BHL0DAio53xEfzG8ySFXg0yw
L4Je/NaTci08N/O9vZwIjyT9QNQUU91pjk86ND6z91B3+chEJ6+aV7XqdidVmOm+
0oMtUwprhxciUNvw0fcQCUvM3Y0HncJoeZg0qwC6qotwA2qfo78ais7OLNNF3tvs
a3gW6gA8xDvx3enVkzrs5AbQ+q9BjICkB3nJpSylk3O8PO6aWpLXivrcGNHO6Js5
EM4500Dw0ADj5hvM5kwky5/NQ6JIi+5p0eGQHp2gLQ/gdLM+KF3UL79g1BbqL5Lz
kW+2TYqQ9wjo7nCfkevBbTchesSqMCDnb1mRUFc2or9PvXMri9xRYjVfKdulAhh6
p1gYUZVEgi9SrNFO42wX+zD0NLZ6GtHvyezbMhWjblYG0WKaGvUFE7v5lobEtacC
20vdYkCjmYPYHW/zwxiSy0NozND7HyuRPu8+pY+D924KnZKSZyFQIZB4LU2w9sgU
lNyqkFpuPdNWyThGhJriSuE3WaQB6tVLCUkppi4262+rhvBD2OtmWxtGNitf0Xy9
BTvw6YAMsuWGfTv86qhzt5WmgvMlPV1NG1U8ppEzijU3efE5mK8uKKDmI9wACt3N
ayEvqdII5vT4MJdwUbg82rsLpN0j04VYRH1b4rRlmcgTYPhdyPjaFeBQOlIF8vUa
mUNSeQyk+KB+6BIIUi2xtLF7PqrL1K83WG84CfaT/JpQ6P1YI932+Vim8Edg1erY
Yo/DLR7lxJVqMfyjwiGPTplDMU7MgOTzDU/kH6PV5jZg5X53uS+0z0lCtcUOU0Mz
/cbu4y6ksnb0NU7anbpIodrX/bGPNwv/nPxSxcIKvd1PEobxS+GsvIkMngUAd0IL
DlbcodMUxCrCdmkejVKkh39ue1qrd5Ksbmh2yqkxDborRoQlMTT2vlguOhHULQjz
0MPmfbKlhPmh3EKUkWgYe9tyialtzPnNGtXi8E1YornYUSmHnUyU5WyEX5vEME5g
l8vEJELNq+JKBR7Cs96B3jRoxVgUuSEQs4gw7IZDwSumAkP3+8cOKzN6VSS8jDyG
FO7vRzVXIiKALkhTQkELx1c28LLuemks8Op+owTsBvxrMJM1N7CRLornurpBpt0S
YU8dokaRXdePrnS/RxOWBwtR+xTt630LK+anU/wtJMDfRJZNa8uDalIRDBAdXVk2
g1MOoNG5COlth6wZlOTM4u17tStrgblO40GMy/Fbu+Q4kkzSiE+EiyF9OEyFXpU3
drU723FhVyGi07wfL6/oVo7mWwUYV2Gy3lZJxc34mGb9rGTzfeDEEBf2mgB0etZk
5tMD7ZDF+ak8WdaSOi6yRkLTxKq7gnHnXM1XgZT+LTwGxkVT1KljErERoKTOHkne
6oejY5lrEf6MBg/6ue2CugO0EJK9Jz9ompt6mr6ehWb2tGcbCEN8K73GOqTTtAkC
XQG/Uh41hJBH2Q/ek12pN9w6snjwAjj88st5rbPBlm9VB7AjSOaH5xicJr0YHQs5
rom1qH8R6oVj5cEs/QDOsO44ZW0ETaNDh1KA9gmL/I98DecbQNANEnGMM933SEEz
GhUMwWuSpsxNoaWcZAbD2aqD3R2nmM62dmyFJY8oM2wicarRCaZbjotDNrQVuNlq
QTKkcUvhMopiQt0UM3HjYK5PAvOBo0jshRGKyVBrZLwniUONs5yRObz1G1ELadNj
A3iKOS97/r/CSDd28fqGiWxnj08nAPMM63/ItIOkda6bktESWusjh99ta5Rqyr0h
ycsLB3ivsV2X700tnrgmgO59n81M3OdmlmFtj6IBXpYy5Dun1E6Yt2smD+hei5nF
yfpJ5F0A9ZbSDFsXnlMCG3Pan0+SK/WIhmM3Zt4CQ4tR17allek8R/+iZ8/IPufy
Jpy/MHTFyru9joHmxwVl/QrndsI2Cl/KJDgBbFb2fkjmy3Bp65cbRKHC4jP9qYax
zBdZVyvdTkK6uKvHbgrncST20iMdViPRVzVaWL1IjL4azWtL3uecjm5raCTruvSR
tGmeOEkLlRoh7ebY/Y9PjMJ8CAdV2DuNWpkrOogkQJHyrrf2ike46xH+WtKyQ5uK
281OAZa1ug/PcbBV+nEYaaJhg6UT2+X+p6DtNNNqxeNy2MBkVi3RKI7FwjtisIqZ
kpp68VQGPzJaegHnXqXGUl7JzMX2jlzX4SOKKdP2307+tSXEJlBq6yMGXwITcObc
cRFZ02IRw65d9UK/5/DhvATnDt+7H0R05bxbVrHi63sR4zjrhKoztDyIq287ceX0
fRrARbmoOmFOInl1AgVhZ56QdiTpgipu7ApFGiMntHBXdqyvVwdvw9eKANmqWHpE
pe+ad8D+ZK+irnG0EfKTB1WEG+EpdEa9h1byOZCTsUkE3z3XKutPuSk5K0KeTYsH
YNok8lFL4KDW6nMfwVc4QCovqQGwM7PXSCl2Nca2jwcFe3oxxkwOsEKvMSoBP4UV
tv2o0UkXuIF/HXKSDHuvzMLKea7yBNPlWuyo1RxxolPEJh/xH58fTJ5SAXntks2G
6YH/fFrymye9/8Zf0TV5+hvDYV9zLaPGNrTXYpWDfacTtnQHJVUgXogXLK1tLZ0R
eE8h4fEYy0JA8ZPK3QoYvGZO4GhQSYOPI7JBW30w5ZKlGcY4JGUka5Cxh9DiR297
/gh8tdYoMUGcX93WwT0N3kNFdQa6IGroKt/OlS/mG5iWGe0wq6L+ry85oDYt3oAh
S+n/OUw7JRSeVHjNhfJRs7LiKEMwh0pgoDaBlEhvGcWy/S2qxDQcczK1TVAIYkfW
OJ+5wjSmmzvae+VaeSVke4iISpj3yTlcyQWm75BcVwaudPLC3S+dDYxUR7piCSKB
LqgErQ12AzzIo850P221T+xItscEDID4hxPCS0Sv+uUwDTcyDLMtRW1HHtRwsx56
aF09cQeiGiUSNBkniuHhHx/y4Sp1wvuarTP8gD3A3p7UVVTYDu8vg0OnGKNRUdwM
dZ2vwT/E3qhGFBptpCzPtedq+ixBNSMi5EjFxqJ2UqWriIs9NDsX+X/YfxqvT3Ab
8B2T4egq+t5BqLcZZPJWHQ6uILr4Arblx6Eb7k2aqJ0AtiG9+dWTSiJ3P+9LZTsY
g5f6QkHCqlM+JXsPN7Da3dHXpnxCmIYU541FVv9BCaAbgJy2+ApZSRzarSZQV8UQ
KISk7kGY2D/y+RlV4jUrDwzKQASVVFS9Ys0Xrn5kYzRRzYCxb8gLewXu1s4PQgZN
yiD1Y0ic8W0Tzov7eVzPUzIvQR6Ydd14D2j9v2OKKye+3c0NuXdv5vqToAHoBQD+
Dj+mh8w/MLuokef54cz5g5J2+ScYYS520yE3Xwp5HUGOKcjuWQnL+Cvup84VYZfe
VmaD+8zdasyUnjBeq4MQ2TI8fMfVTDE34GmNidTFo3e/ciGcRIxp0R26YnwTdqNQ
R3+EwsyTSHES9r044NfCpXEXXkrTyIbqIYNNcryLUbziGERGnpEroxvQBfL3ell7
sPsZbs6aKcnBBu75SS9g7Z3vpHanX2rkz7/LsmIFeplg7lb3n18molHYxaywjG1M
66MLxpJnbSm33dlawhOsOF+43YRitH2bnWjIEVOxlhaCjtiTEt6fof60Os1fwTPt
pzhD/kIKx8G+KpiD7Z+e4G0mZwFaHcVyNWA22Pl0fE5/RAMnK4ciOOK0tRaqKoRM
W87TE7ZMIA8ocmcru/iinSBdkmEj8WhivU0vaK3gEWuAcuHp+m0RXrXsMTFr/GH3
WClMbrBT+YH6v4e+ynon/9mNObtPGwe5FXZRUDttmF+axAs5IIXR7sMiF3Udn0u9
ho+hEKH5qBw3FXuEnpYVWKCIoCKll2V3VIaDFOr7BFYwBau/aPZZMFpeFkHqfiG9
oq1nQE2xS9yLoPqCMZjTCpVQpbcOQfZErUZST6NRlG9ez/up00JGgr/5nRJuxjNV
o25u+bYNxcwLMTLYPstXvbHybIWCk2pDEQ6fdf+olYN+htmu4zyVCy04R9NIx3xn
JYyt0TC9gjecxoDNnSmaeku9dHoXMIxKgsTBOztVjdbdqulkika7In0xKGWX7tJX
a8vSGZdRObihz78XGbNJ16Qcb5wSMGpepm7ULwOBhC4W3Wf9BMTeR3mt2CMBN/Rz
JM4ua1NZUf/NvJa6mBV1BKCmnTedpACyqJAPuGAVlUCXOxRQbAMglsyxbd7qOU5W
vryk4KY7qYA63FG+SLr6hqEOzXu32JoZi3JXRUmf0WunjoYiHowZywj/9UxVoDu5
tX21IgMDtJbo9UJhgcEu/xO3003x/naTxT9s0dS4RQg0gAH645x0YIF7LeH82tbk
ygB6Fk0nEcOOpECTh7X7c4swHBkh4OCem6znHrPhwJynKa6EHzG3EFC69YcJy3pe
na6/ILkh5r7JnGRdDx9V5as4vL/47LXrbxRPYcdasvkTLkKvLIZIRXY51o4fxLZc
4BkSElCcWlrQnQnRyFjPclErGfN4tXBNGe/HMcRnAqeub678QyLYJ19hNzZZe6DB
qW76W6zImKXyMmy/bvvj8/An8ed2DOtun58GA8rsGX0BTCCkhy6u1Hy5nnlCPdKU
LuxOJeEV31Lax6rKFE/lEWyN9I+eMsZh4SQaxBVYhKEhb821Iv2laI+91Hz0qJms
Kmcu1nLvOYIKLk8YWp0b54lquJRHe8HIh4WROMSWXo8gdFoUCkKCmfH9xnWO3aDT
2w4Yff5elf266ZsJD8CCRa/kI78w7+9gOOz5Qnl245HrUIjv5lHYR78VeQSU0Mqx
SaMFOG3CqWkFl/a28cwCbyQDokOz1lyclsthC87OmeFP4KEkiEXq3/a2+sh7MWhi
Atvsac4p9+8OSfmKApTyM0xjvwH4zsZW8arzDCavkU/X+ypnIeHC9TcIp/utRWNe
oadAfJvb0no+z+WE2XmE+jVLdOKyI/HYEm8hoU3blyqJDx4Hh6YXbHxFJnxOeR8q
4m5hJJYVfCmer0HiYCqn8qUumCw1efZF/oKF0FmfHMSpP6x/9ATa1BiH8k++/e40
6RhbaO8Y/LgarmJfNKZH/b4vpwL4eTZzQO6r6uNjZGp43+eI0ygJh2HxGYMJkFYc
3WM/xI580uZ5rTADheJQAPQdcqbOYrLajkqpfjnSl0bNoZ0FBt2w+BYwsQ0TVFDl
ejLCgGoNy9cLOWOofGY6o37LJv7EK4kpuu4IxJPxx1LedImFBBQylpTXaQwx6IeT
fLcO5Wec/ywTvEjPuaTTpz0mEX5RsOFq3pwLrQHmNxNhsht52V3j0LexuIUCzruS
vl6vHW27oJ3tiKhmRcRB8GjHBWnaRNEMb5lmEVbTF53q9XimgTaunwHoXeJ9CKMg
GkK3MwfgAGFhiArwNjmnzEVPSD/xynZHX+Z+F7OEYTSAWB72AkO/Rs8WNpUE3cCI
PcKc9anBFnoCUsv0576CJExhGLZU+B+1qP3iWPTrYrgN68BwS/CpW+ADYOKkKOcb
gTRBkp+zmb0Ehwjwa8KDS8g8wrYksAt6gGAuzC2a1ElmqM3QRQM/zcpFuApV1/pa
neG+pk2fRYHC8ExYYs9HT6mcfpFtBUhO8TbOBOqlSF+TlVwHuYMD3DufHdUkqk4V
zJ9q4ipONxVWGkMy6YAUREF95q0Msct+xV4ou1ATqakySTER8hWUaOatXk4w4r2N
AiixE0LKk55bbb0SgQKv9UuyjK0s7cygLN5H1+2pYT4MBYLFo0V5hAlQk64YOTRw
2/waMP1Mlsdh2OuU2hYuREK55x4uU2hcZ8+kQCl4U2iIkzYd9kZUfKph0fvVARbv
MsNKTRgDAXibDka9qo6bSFx1xkPd/BTyhdrp1KJm6Y23WwF8fYcPfprYfXvPR6S2
NSUXW1eB2Hsok7HvgvTgBog94NAOYtw//GXD06D8FFSPeV8x5hJ6QoWAaajLlOCK
o7PvEKJATCwy7wsynOGAqlFRk4z8VK3BmJH25lfM9pNlmCXULfyEOnzW3RaG5hrs
gKUqE0FSLIJVf9oMU3Sth2nd6mLYTD4Zp+S6VhflWgQ5yv/YNdrkj/xqJYkVWMus
pN+Yeh04kve5aQrPtDkJ0t1KqL0SlX7TmDGweHMVy195eIP+KtWF0HIHBn48cVwm
YKGM6mqQEw4I22GFB22l5O5tkHaMCoiDccM+J6dYd7T/B/zpby7GamToJb/CUTgO
d8w69ZI291v+UUCmIjfQN0OLu7KPAESHL2Nhn9tm8hun3KNOfk/Y5rbixY0LW38A
ov0kc+twc8+2pfBDQSk5n7XATZIwoFK2y/eHs54Hr/dv0sGXDPzONDxMjeUpD1Ab
zobPDX4nLo1RkvnA9wMA/ejiROzBjiz399vF5mVQnqiL+wpXUgQGfcdDBzZPgVdG
6h2upgkolMft0LFnaVD28MrLnVJpKi9LwYzgHWYbUHNjlrsTZ3LnxoAwL/9VYQy/
KASAS119Yq2UyNH/ggyvGk5KwCXn7DtCITJw6TzloPpeGqrsljgSYRxGRFZvBkgt
gH0l3lQPZVOw7BjSbw3/erC1wpAPILadGGN5DQb1fF+DsZtzMXzt+dSM78Z0GwzV
85tJEZNeKVVbLOy0zmQmoAoOaW7Aa1DUsZC0683CFuNR6+MJlaw1WzCQkowR53ta
a1CpOGfI6f5cKZ3GyrQwZ/WGvQ7t+Mw31QjNStoPabUrvX7rfL6h5WqJmj4cwFDi
b9wKFO6zdx8DEAcZgCkJ6VILIdJTZ1iU+OjC8DzQ+qn1V5NjexaTCSeuU5UzjGhH
qn2hyiqSyhRuI1TXTLMYAxcMJAT+Tmh/ZgMyeOXH1KCgFWl1Vz15kGSXHEhiW8Lj
5jSDKlQ5LXrV4dyymGPhIhaLhc2qweJrqLq2m5AlbjnkTuGE1Lt5AiUKIac7mnCx
4EvDgjR2hcR/VxMjG4SDJbw8y6W05JLIy4qcg1/gXBfkgKmOo9T+huQ+FZn0gDea
dN7Ywx2dkITSwHe3hJ5/U6EzLxJIdoL52bijvMSF0IeMXCMc2SG+dSQFo80dm3Rz
zijEbtJZcJf5anQnX41fUaL2CnNsU5edcVSSz8fpV+LsJR7dzZusdMEErvyI5wPK
iwZXgHMlxX6ftHAxMABfNcv7Uzz++8mpotKW8uuBjKmYklrkWJCPkc4sUWvELGEC
lLaJ2E179kYhHRoZwmaUwasy8NTfFn7U6kYoUulZZ6wBzA6Pu/BinkNtaNN+8e6I
nH1vWRYSsSgKwFxzwr5zpGtXh1XyB7G0VwtWyqB6U1P2a7VmffQlHmIhaiINBPv3
lA0o43qagh/JIHvx75DauE6juYnvRdxffgtMZBekgUa2+7qWYVivVQKmWUR/hmXm
FTuJ8DBB8NOQILFpA30EscQyF05D8XCWpXyiOD7qPw9HRbCmS3eR8zm7b8i6V2CY
Ldlmpowi9Wl4BPOkLU52xySFun6lpIoGsP3A1zQFobAVDtihaEaVPFD4hSBOBnan
8AXrcINNVezh1TUoPTgEqFwyD1pv0oBreps8B1F4OtuYq56IiMW9s5VyIdrXoNuL
p6foDO0pvT1FR3icKf1jc+/00guTs6ggd43DTvy3gl0uZedGjjebzma3dRS9Y7/j
4tVHfwpThnERcuLirq9apt8/+umE6v6IExIc6nruFBPTgquu/daS72ve77MXARtu
2pnCuqN99w9viNIgsbBhqmkvpXs1soXQ8rtyq5HAP3XyGyXA9E/9Kabt2u9UukfO
1He425yC2H2MMcGq3+s6v3jL3YV1ILaHN7AC6XYbLmMkWBiI2q5b4BJC/iK02VNS
w8JbwqkUkWBoSMin/C5ebKXkb4tIN1c1uOnTZjXrilN2TYimIO3i8ZDh01giCQhJ
SpG2v1dpy7GSJvDhEpc6eQkFTPdutz1dSZihztQ/6w3tZNpqQ3CiwF2PHUKm8arQ
zuOqCj4VUG4FH3KUsTd+eCQXkQrnGWoMluTtxGuFmr2ch1wMAZkgEB1ier68fpxE
tYILmE/TxZoTdpBZ5tjzQ2AmoN3LRXuwi0BxDon0OGTy+TqJhkwFZ1p93noC7X3f
K39Njez2JBbGYVIps0/g7tq3ZdKi3d95iYExmHLN3vIS4ltGvEHR8kK/MOtAvqhM
Oc3Xj/qyWWu5kceIej/OIwFxh7trCP2BuYtvA8g6o/t/DxIuJnG3yr2SFMy2vnK7
3plwuohBXnCk88AilPIaeMyGcUbyY35DASv6ErUqlG20XXYf5zx9PDjo3/wqdqWi
kwpS5ShHuVI21voaVBL8wPcSBmHKF8HTvfHbQDeeb9QHfj6tWjcZ+Up0AXgXA+3u
zm9E52VGFR/nGzYGVSrt8ExzZQzGh8DSI3QR1nYaTyph66hmfFtVtjHkQO7/djjl
12a355c6KPdMOqqsPQNGdbUf7ux4A33jwup4e2dVLmLBYYF34EHaCL4Oa+92xwhH
i0ZErcvKIy4HfizZ32bNFcqfv2vk9qjzHnGRIV3vTMVGIJRAjPU2kkb8lgCFk8cC
akOS5IGR52Ti323dHowUDabRC1lhNNBeJ/db/xSIEEvkac6FY8q5cp7prz4m0Jeo
PyzRBC7raczPoeaZtGK8YhDq9obk5xOFWC9+JmiK5yhZBjBMXeot69du/2YRdNml
jqiVWQb5Y1X09R8pn17nQKOoJ1kv704IFdmjH1X49eGPKVu4cCspcRwrySK6UvBg
S8BeTq0EeAtcskBIXmst/+7SSXVDzxW34m1OiTqxcFXZAlCknsT4nhoBOvbx1UZY
lEoPfb5MbD+YKdmkKD+2kFM/uDp0TbY0a+OVS3dBvV39Ra14jmCk4i46Oe46Yvzw
Cs6K3dGCLPmV/3OLvx7WHuU/Jpl3YkHqCiXIe4sre/9SdBSPs/+Nr54VJbl6SHXy
eN0gCvawUV0q/PM3k+9ApUEjNrqKjOP1Cx3NOo9o1W3fgYlG9fpGKsBcDPWvOGIW
Mp3cYK75nM3qDycUlrVzwgs+MxVfaCZntwDucmagiC3N3cBGkauesj0nbUwpSFx8
g9KDLEQSaSWUkBFatSKOgxeD7TZTu5QTv+tYpCKlZa/6vs6S021rgqPHdZinsXRx
bQXRz0CwpxIOZFADBAATDEHIFI78rh14tmAgi3Vatk0PymiEc/410W6EbzrPX2Fv
SAbNd3JQsyzEo+JEoChvFjh9D0TLjlJZieNeoBriW79qia8PQAXuPlHwvZxVVzrb
wnvqiVZlypvX0/ND3uNnux/yYULczp8AjjImOG9TpMEoPQ8GEVakQKc+Zhq1A0/B
PEkWC+bZjJQh4uDOEqfunWhRK8U/qcEjsAoxG9Z2V5V1c8w6SQlTzzB7NXdmELp+
JMH/QJ0TKkWTUiA8iNtCPNoepvZPgWI4MshplAqVsF3p+nf+V1jggdenMZknn4s6
jJOHXlHQoLjZwOS7WUae42JJgyuX8221HInxiZ4EJPsD0v60kD4VHPfIn44LFPqH
WG+sdWr/IKlw4w1jQV5bugZU/SvY+NHKK1VcXlcqJIvMdQNUyHX3qo/3gIuQ2sZF
dq5LYQSrp8LbY2sPhbRJy9yfys8JHHenzDd3NQS6JO5byq06a6TFtfHaSbhaX1RE
5+GolmkQntmoSkc0x0zXWBp4Jscb1poh9nPV1MKEf1GaJ+YyQKu6YFh+rlqRlz5x
5t5Do2BkOkKHrOweVXgySHM/OwXZKr92UjWKSggBPnfD/F1pVVuGYnEhNY9XVcK8
tb2IIo/tdGhj/jJIwrMhrVDNryX11zy9FYgwmPvmaNcBTKp6CuPWWKhpNX5aCQ8K
GqQ1oraaUKAjuSmUViHJFUeSwe7SG/O4VEUIlP107KH7xHC2FhtuuVQeouNRoHNg
p3f4tV+t7AXxYx6uTFAx3YRJKWsYVR5zbTrfPhHZfy5d4/zF1Iyo38atpmMuE7LS
JTFDg+gETJzMIXwdCYi0/MBJNds9BU7P8mdLDYwGWBfMQxYPD1HTno8M4qw526fg
msq9zf7eaM7yvlNNaR/LlLcGWXJYZHYb+ZAl+BBEehGoA5FSeU23nNCfDIh8Au1d
XFtaN+W/fziTqdYrJLIJ/7VOlEyl8wH0kGsLC3ZFHzlN36ddU/xAU7OCuJ7manFx
BkaRLX4SnKGssLNdL8i7Pf8uGyfL3ZBlc6+psv/NKKU7CKR6RH3EEHkuJayvuFYO
oSp4yzkS726qF0q6iPc/otysu5ns42VkBUM64bXp+eT+MO58kvQJm6iU23zEhQjL
1QkLiHpmL7SC5TjUD1pnRjkfhgs5vNMKKm5BLsxWD4vzcTRb++9VoJ+V2GhPWVFV
eAxcHzBAtMUPl6PlZ1YD4/kZZG4jL6Nh/qHjXVy+cR2i8055ZH2FaW2E6UcI2lKS
bIwkX76/CdmsQihRo/9c5fupTviPC2bne4JL+/xM9njz1etavLeGKRiO/gIed4/1
DWGDT2+Wdm9tmXrN1zX9yQSwvXfKCXkT3wKus+MTtLySVP+MnZ54pOzNPqtR2iO+
RKscZnZUwjPRtZjzUgmSbbw0NtopOSuadT8E9dYOCD7d8HHf8tVNVvrEY99JXq1P
LbV5lABtqhO/dfWEyxAxuamIVDOQBtI+pg2dCAGD8R98pJHV0yVA1Fl9NPGNhhi6
ARlk0H9AORmpmudNvSR9An7nB1R+fSfgpz/oKaJFpWFk6aT6wTMM3TO4cO8VD6qR
pJHAN8sNBMFxqkM4o/lzVRlI+IQP6bB1sRizhwXse+iXYfgwqW63jsRsUlgDvXoj
4IfiTfotTjusRL91okCmMmUxwQPRutCOHz06YzlfbmPx4qj3BTUNJP3vFQPHm4G4
TVFnB26aYOV7+bFu7blC9hSmzaplhbYVRpttIjeDfIX2d4pQphgC82UvSBQUvjN/
dCHHfuOY0xaB3/S+BQBJ2lKq26ZrRXPD7ilzDMZgjUczTT1rxeLnllmypejaOAEy
7irUosOdWPSGw6qmR9nyN1QbGHmbDsv8qLD4R9InQd5aUhrdFIKu8+8VcndyzIYx
H9PucTAAPt4I6KzeALUMCEp+j3by4f3ujwrP7UjjHi477+zJF+ODJEhfb5rLdWYM
LaS/G/BdrwkEhd087A86m5lxp9a21iSFwoXYEF6sTRcjqK0JWcO0ij6314+kYuFU
prrq4LLEeVw5sfbPjlS+S7v52afC8GXfegVmzJ9xY2dRboW+uKltLbGyNdblF5mP
ISmYwmSlFX5wV9UWCrc5rvf1sZoYI2jlGwWwZYfih7IUk4GbUy1m9QHA6rdvu4Oi
JgCbdSy+/2z63YUOHwMLybU8o+jy8Ml4IP+PY/t4qMDY1sEegRw5pId7cv2byYmB
mofR0vFWexyl5tFqXk91o6/8Bev1K1Z96rEDN1n2mVKDZK9Pto1ntY58zdGw8WFu
D1hzFKlQno3/OPwyQ98Keshn8MrqYpAfm2+ayxSg/tGF4tiNSs9dVEj3nm7o/6zT
jRcBX7OpsvuV1OOJgLJwRoxoqw05s3iK7Ne8DBFmij5YJAFR0cZP9R4Y5WUZWR8j
/xgj73tVH0ccvxAj9/gHi2knpojsse12t1n6Y+LnDybpDCix5iMNbvj9MMYz18vX
rPb9o2jw+WVB3eYdEMCi38DflIKK3LqimeCarv6j9+5oVLIvU4Lne4YLBrQQrodF
D9rxmuVEVZryj/Y0IBAfWA6FR01qiyx1mGNTTgF6LSV8O66Jda3G5fBs9zy6+LmK
UE2hmFDvYHc6wGi3ZSCHYKU0PhtzV8scsV+L5GVEZGmPkI5CqKQZ9JT5T1WNTtym
HvEFtbaR9NljMhRfOLWJSxQx223qT8jV8kS1KMGX+t6VvVZyNKHrq9r48b5ihUKc
epWL0bhXcJSTchMXG+xFrudmqMd6hrYIWIPtYSbdmuN0b8XXk3t5+0w+ZfshyDyU
ALEp1hxGFIf023mnFKpDyRntRwLBC1q5TqC3Jp6E1pIQLF/qHnhK9TdXJa4vgphK
5e2hz1B9XrP7lKp6u3SUdYaj/kDIaAhIpn+Vv8EnN6iCLyCCbWGj3tV3fGiPaESH
T4An4PyzbtJXnfPQRUWhssJ6xYl2MLHbvEyN0kGf0mL6MTI61r0oOzFK56UMci3a
rffpk5QVq9WNGIXQupgwiSTg0jf5CVnGIStLiFPdeNet4xPnbRtyBYsaQDnSlJTy
Wcub431zcjFzMc1etChk+rguS0TmZsCQl9QQh2UxrxwKLieQqF4zFsOFJdQlk8yl
77OXdPWU7uF9hykV4W6P3hwBbx5KNorZYI4aUtfJdr3BvXTzPPB6GtWxoh+N2/6O
xbZqMF0ltMHCfRSwZvTQ8V+4Dl8V1N8Drv0To7TJ4pv5uFUui2qsn46zTTSMSv/k
gwUy1lB1ppLP8qTQ8WadWi3SzwwHXKqf8K/mBZu0s0r0e8Vq5l3cjlggfUEfO+9d
QB7OnDaHP7CANgVbrUQ7hAEDxT86ifGATvEOTjkRlAhKSAiH+bmslCiQEwdixUnz
Uv9k/0JnAJftcxpyffd8iYGK8XNR5fKfECIDDr1hnkycpE+MFBXLcqQSkZgRqa/t
dFbViBzEVWp/gIrmM+ca1HpxEKkB9PF9MnMGrpwJV6QUmDbmatNJvSIfE6bUT39p
Ny9c5Lv7ARmu/l9mvf2kx2180SUlArD3KXkWIdBuYHjQX+k+WZY+BSc46cPAwJhm
dbn8hlwRJd3qgvL+1pv7Ytug2Moc1+NrN+7zRhyrBGztpBfb0LF6j8UrTGUNcYnS
Je2Z5wsZhJ6iSN9XGwcQHyLn2rxgxQn+dvT1AEwPvnfeA3JcT0TuFO8HdjexqLFu
+J1zJJv9frRCskJI0UDl+9g6v7Rl3tN2lXj1+RHnvrEX4Fhm0Ht9a2RxxjRSUybc
nZUYAikjTyN0BWtbux+iznjlEymuZbCV6A8GFNAz9dS5bg5HyrUXiP0vjJ6QZdVS
ldkvkMwt7ULKytclhoXNQ3BQq2rId+amv8XswR5E2NcLAXH8qrH5Ybj8DRNuIc/V
TygFVyNG3edoX51JHvt6HSRj8aFmYqDS2Y98SDl7r+hJSWqiw/UkiPBpXcaHtBQt
qz9Uoi6CAuqX3QqSAChOBDNGIRct+8Lhkp8PkejX/oUQRlQTB1Ye18+GucQEdBU6
CD7QW41PUTIRWcOW0AUHh91uLXB7yyHBhzDzo5VsCwh1oKykmOriJIAxUdkPXHuR
WLpfW8TV/4i2hzUnhhbBeHI4CX4/fAZKHdwM3tx8IWqM5kV6IEK+ZyIyAH8Vc0hQ
FHAuYQFcNaKooEWWHKuPH6yqGygFTYbZH/1xB6v/2RiNFumYCzJTVnbzdA2sSubl
eqwSpB2dmXzqHBVe7EaGGMST2Eq1wLai3V3VG3kIGUPoFV2Nvu/lPyV1RD92MeZz
GsKgi2WUj1JCWh7urn6T/nVhRjVqgyAu3Cqm88Sw/SmRq6PHRPlFQNNwVGkJr2Gh
v6Y+Df+8a5I2JLmrqc9cc48NQjGZpIMl1pfRc7RqMAcZe4CdpZZEV0m0uafs9pgq
fH65kHx6K6E2nn9Y4eZLNS3LWFmWrUHqcVrYaHNZhzPAvUU8sd3n2/xl9TqRYEKg
6nvYJYL9lMl71arWJxUCLYXBl0bJuUA/quwMQF7F3gUoWFI1X+Bu077J+EeYqucg
bLJUD4ZjlwywmCudjYfZ3rtzbYksGRS5TAydY2iEk90QSWhVUmTz/BszL/2V364q
+CxS3BflRmCQ/yGiN+SOkVqd9gcEZKlBC+g48YpW8UtQbBWDiXTHCpZgQYjt8MMU
wm0xRCbfjqYsnOQ/LCcwI4AsSBp77Fge8KndusqQIjErfyY9gBkXhKqNQayxsxWq
aAs4crQK/vXWWKEJF+cDvmEG0c16RQAHo/y3X/CxgYhVLR430gw72pDPveVPlj2t
ODF/f1g+wQLejJNt3d+EqDm/vhtbT30VGslVj+50AJRTKsrXZCJjwJxS9Au0hFOR
7TWvbbX6Z7V0pU5Aj5GIdsxUsXqMp///cQF6PlmNO3kl9JKnO3HNOoJgqjQeO+eb
XaatKyguw0Ubh4BnL/cwoivXZOpDQfeIsEBGizlgz1b7nxhS68BMQ1jOGiP0Lbqp
ZJ5cKM+y0ihxJExo0G/hf9txFYwVbYeSDBAV1AwfyrVOAAMhZVfwWEcgxd1otifN
p3Wl3fEQreHvD8MKtmVfMjiz+2GfxHI9w/tgyYEF/tH8drXe55vNHD6iDrKQeBIu
B+9tWIduKZFU0t+F5Ha+KQBKAgbRwojXTi9AJjUGKiocr3L5SdNMhsQg3hk+FA4Q
cTaKN0BjkaRJ7kTABkiIyZc5YVzSATr1+A2G2jHrjJtis11uz+DyABNcMVQygW9s
SfhuKiE6dtzEUDQnk6Q5TyX4oeWRv8YnpE+7NyMb9lDatF/ESa6UU3t1jF3EM1qE
zG0NVaatJjEFW810Zm8yF4Vr2uDxKX0ljUD2zmqHj1sxb1Ueacn8nqK8Zb5Oki5/
/6zSZBnwOv6S1M/hrOwhEboF38Env7yK/X+GtOjsJMvPMm2Y1qt5imoV0HVE9yf/
P8EeB//pXFhdHHXHI4PScSbdccO7eFXFTA3llHRBVGU63OEGg/cKahmoxMT7aOr9
L1ApfYkQfDAN6wr0e3Sarl6nepuNsk1NKzhVRo0HKSwGfpP++fVbbrw4MvIB+/8H
A5fHvm5TvourgTgaRp7Bg+Pa/NAMD+J5o+84aqSSpFiGlrWM98gqntk3Vue49Bcb
rj3nz9TlKDuvmZCgVIa9GJoeaUhqBv+sns+4+tL0LRJKUdHPBVJl2EJxqLysA71w
YQQYgoQXnyCEefohuxMl3sVhqTNhminJOJTxi4rCexKaZQyNk9SsQVFg0h26P25V
a+8so4ka2UN8Qlagl9NRQv6Zt9hfl16bhRqrvN7wI2SyMrhRwIK7lrJa0sPIPbPJ
JGfhniBQhCHyWdCwYOma+/Kzeo5yOFRLmCkXwHmSMLO4p1kCGD73RhJPw8eVfTVa
fUfKFFo5pTF1xhipjT0u46e7lLpQrEkJeZFkiaT1GiJ36i23A4/QCRjbYUgeiUC+
fiYMy/963ekjDhK+T+5ZB6c7RluGUWtkz/0c+ZJI5d8OPXBtJ3y4KJ430bhiF98m
pW/4NMWxdq2ZsQTKdAtu4Mg7I1FnxxdoEMB2Sd2vmTpgY5KViCItFXemCaX20y9w
D61oyuDQZiR2efnJzNHAWMMJ8qqt89AJ+Dnzg2jLbZ2zhH6He3hJ/gK+YOged7FU
LR2fL7YNEW2zLBxYXmc3i+970C9l9JYwKMISalqaqNBdr+ADvwaZ8GCDV+nt9a+h
0eQLNlK3NU1CIrBKNm0jKXj0iiEEHeAruUrqW5iPfhCh8unn5CpmPmi8IPAKG30p
7WF7ZTLip7KP5PKbbkIJ61vug4J0mYBQTKyKqXdrxNZjQXTnhYNY3H8S9UKks2sI
mGalPjI2bOOaVediPslxfAvYGss5NnR1zArzaJNSiuoG+pKLVJVe/ug/tR8jqmeM
V5v6FGSHk9vr6fmrPrRco2BDtBTr4gtzbCdUlUnSmxADt75aaI8AxZxMnVQX8suF
h4Jh7b0jsPQd+vqhYxOHpuI0IKhCwHb1cTloAoZWu3VKMNJBJ435pantsbNgecVl
Lo7HOEeg+CLTMkUxCBx6/CHaZi+PKXdcCUkDu1NZq4oPRVDY99ZMse24QG+XOXdN
1bPkLgHvW8XLs0yKelQZEaMjXy78onHXZ+jSO1jx9adJwBhvps1qZWwpSLBJdRMp
/3zotbH2pQNb/8tHL6VqB/Y8+alIWPodrAYkIugaZ7XPN6kcnl7055fvo3HuTj6U
wckzeEaOrVENyyksY07TZ9iFci+ZiBb/T2GOVuKPn54C9G6ifNAwqEfPX6GqNLLf
jdfpw6PYY9TV/y3OmozLlhVjshmryAO/cmL/U0DGdtlzKhk3DS37050mGhq6Z692
0vK2hYPSSHVNKpzQcvFKT+DvmxWArmw7C9olBs1ut9aTybRWX4TjvrOQZ+4qfuwb
bYFlSE7+MsebZJ0a9tyIa9dK6oXhP3N0N9skRsMuFXUa0VC4IUxn4Ecw3HpwE/Nu
FoYFGamBsUbMjgcvIYVXljmyeRpatGaPWklitl0PYqAVEt7T+Kq4mZB5Yz6UwXRV
qD9/c1ebBmERQVbQaIRGerT4rnHIPpNmI5XJud87bo1cFSv7Hmc7ROZLua5YSYOd
ANa0C6rvibxvxRLXCDICRTCF06euk2gJbXC8N+zalKRNr1UTvbx6abGhqzfmq1CU
WbCMYImu9JuywZFw015opF111h8cE6ftKPxuHCZQCguw2yrF2WhUoQurr1aHRfYA
UMreAqrAiMsHZaEwCNx8KeP/QvKe2GNW3fQnzZGE3WuhRYvsHTq9SnaAx7xACo8H
lKgKE25oAdLonFA0yZhyd0q6USp3zXekleD5qfcUb7KV1nUxWmqdw5N8fmz5dlS3
zhw7rAJrxr2lqcMrbGikIjV/PGcY3mKUTe8mOh+F3Xu4PhVrTdJ9MRPTeIlIme+a
TF6/F/5SJDHVv9hKnZrNdhHxcN4/cGFFIxyCTuHLurhUZZJSuF2/MPmNiCtmkkc+
riMwHU98Y1GoyDE1fCQwnVaga0s1z/U5HpJrYqp/GAcDiC50tg9oeflpVmR6q9BN
TX72H9cVOEsrZmZ5i3H3iXbs1rB3GTcWj/gaSD3rWvXpeCq+ASYZJQvY8ICgP5y7
HXLhdTRx63P4HEdOnfL+DtmRlLPIe3ispbHmQ2/oYuHUg858GWRLNVIkDTS2diNF
4CTp/ouXFFg6hDRciMGYOnqsWP5hmUgKu/FXnct8wD4fRKnsxcT50XhtmTBm7DrY
pWXjWOnKpEk+vQ5u2bvzbeQeLc3zl9HXQkvHRwabg3gusNg4+xw52v97ilao656f
jI4QW/O90/AHVk4rTsSI1t9Vupom3QjBNHz9w32WNiTix7gdSFkwZHR5SDMwnQ+H
RoyIVvs7/OiQmvZeIyvGEAkT5L/dD5nzD7s59bFnS3khTTdjV+PZEmOe/KFhqceK
qBveCXZ/GnED9uWtUH1w7NnOXg/5tnt8gxERCWHMYWZ7yuqJa4WlfQk+k6l3+59w
XfetPznQG4x7wCYJ4C6ka+seabLuPvf51/0zKUMRFyYMam/PodZY8/FZMZqFl4/i
GfKCEAq9j4sS26+M+70xDT863bwsadmQTArB0Pff0QII89mr3kX5pNVyNqMFx/88
EyymPH0H590/luR1QBTGnAUBqm+rSV7shatZQJaHOAhJmUG9XxaSJlVBovNq48Uf
8tN3voFMtf+odMzNNScstrt1vSIVpFLyeFRb5JRuyNAX8HTx2MZ9/a/CN1oQOQWF
cd9FdDTgsQR3EPpqI68cQF0Tg0qrASU4t6mwm/IY0prLhA8EHYaz20Eb9D0Vnlpo
2gO8mrDAbj7ozyRU6zuGdNWXGVb1BJVTpf2ctjviG9bQprtD+kKFFmnzVuR1cfyY
lWre2LKfqkWEmBrigXa4E2ELp+ziSOUYFBYwxEXOacXtHYWNHbb5og45IPakBHhq
MK2tj31Mo/PrgBLz+OPpXeqKuz5MIA9nRyjqkmPx5RvADWZdUijTipTXszv+22VG
6/zrR7w8oVrbp8c6Kf5Qx2HMYNEydJv2rQfGyTtqVpRwhx+Jo5uQBq+bWo0+subH
pi5BWY3v0Y8Ek/nu6JjmaIL8x1WSQ3UrPDUKtFk0zFl4Bu3/tsVuolnVnz1fX1ad
7bN1UY9Vt7zyHEtJY7yV99ifl0RkxqpaKk6Lg9Xkyip2yYO5cKBZcqDisX1gY9sZ
NXjEjJxgeajjdRrpAzEsnRqFLAp8W5GOw6ybSy4heraOz/xA9YjBX4aIe+b1qdiT
k8Arnvy5Z0JIm/5OSB6YPN4+MIFAt6Nzsn4Ll4lKNwe0xBRyOV7P7fxh1SWk1dws
9AX+LSaAaoytQF8uSpV5FnU9rO7J7A0klUVmTttWiOrPdeF0fdL93A0Aa1bhh/Vu
HI3/yolB1AvUTRJZwFT/S/itUJaUvhK3htmouc74To13vrOVNplNeKQ9W9Kxj07J
RLUr5kUpIOULvD9J7MB7NdOc6o0dX/bq61Eryp5JzQpltA6j0wc76V9rDgIvCX+U
/bVxmJ/02MXECpAuYJFHGg38NsFsjnyCYoDy1wcPsCnL/dulRJWhF99wSaEfgZhi
UUj7Ap60d8Sa7P71mECh+cQu+mvy4xsNIL+5ZMlLEd0AifGBYO4SjtbpeK9WMeFN
w3FdUzpGaBvnTjx32t8yy5kpj/MJ4qXwYv3ZlcLL1B/kZkfI4siWNpJ99EOITRnd
ZDnKRPjhI1oJASZoWVV6LfdtoaipOWQRo8p8Nq4QnxaxG/rbmCCSF8iaWAfbr2nE
d20uwz8MCeY4LB8cxoREpQX9r0TY5IlCNDCUpv4GJPBNi3JwWwpt+dCB6tk1jDIu
UFuX7qiO5YGg/Z5pCZ81xL0dneh58YvHk9Gmf2JbazrgUaS6hvlexu5nv19aw5ZA
SwVoK3ia6QTcEnXv6ES0IwPUTG9OKjbJnguGwLJWbTFUn3O5uBJt9ck7cGGornxp
4jo3dPtxTDwweHZL/VPfyrcV0qC+HpCUMh1uSLUkNPbywtBl/ulBmfJRUWlXK9rb
30mL49/kt06AnDaDPrFu6hJmkG76fioUl76l/+VZ03WmOWROxdtX8oWaGfI3AMRR
tprmHhX/1uYqW1dAyirAw1ybCBGQPjOJ4cS6LbWtXHHAE/kjpanXBHj2DhDXaMGY
h+XFC/KG8iRgzChTgL/556hm3fIEblci569amS/avW+2BO3w60cIKbg7bCeIpn2B
QcTNsj0qDCD5wzoTSaSKwouq6sGHpbPi+cWd6ZZBZz0gC03fWLGjiDRkU/eVCvuZ
cVLZ8pdNODXUL6KGH+o4GXkJ871PMeZmEx1Gc9qy8PClFBmH/1dpL4D1vPJNd88d
tLeBlFIqnNd0oW3+8a6tVlm+Gk90Lwflk3vRjXTLMRZLqq9IEGDybm1z+YwccSL2
49445OmkHIHDXIbrF8PBDfR1Lx+oVk9E4JY1v4nT1bf+7qaCWCEq0gZXOPYtmlcv
Xbkp5dnp+oo+SIclApkAzDlDhKNGvOB4svf8Ob5SUFarY7LERpHsy1uCep9ZlFF2
wQvIix/y6R+JDqmZA5KN/nTMOveXVwJQNBE2IBHuteaYsnbvN8ssxejv5/V6KSaA
hZsKVD7MUlv5zgZN33X1vSDNuiSmgsdlJGbIHxWwfqE7fqDJqXbmWZjWs7XIfHoF
EF+erJKtsNkmK6MqKaMPkYpCF+WWEqYwBzx+H9yHvx98roTZaQZjtCaNRBQfdb+n
ITDDKIPvMgY89feu3pw9OBF7QNoKba2leqtAMwj5kJ8MQimgZ/5td3F5rqU8UYwf
4CAJVtRsammXLRdEmKkyEAXygydB73wep2DBThT54LCb3xbdAmjPQqcUUErAkbst
Kt97UPwKABfrdFd5JMF4tV0Vmd0qR34BSV9Kd8VkgnHLzo6JrgrxypL15HOXWAZ2
hya39Kd1E2qAh+kRApp67YE/gpIDkZwMXRjFC4DRwSFoBCCjro2yXWE8NsVOP6sn
GD9grcdOe1r0Yxt5HL+pYu4yuAS52oYqyJwXB0EXKsmrF7G2qD7wozkBT0tvb+VC
UXYjDZSBqRYSRgKylV9M6+DfTj/Z1kQhJL3blSZ8whEjmfpTGieMuRR0QY3g45Q9
62w5tAhoDFDiUz0EeWnRWuhl3lAYYZ0K7MzzXAw7Qd/RPDJkOY1XZeHbRay8hhrl
Z9d743ykydKINmAW4sG4LCYZ/XjODR+TE4nQ46ch4cKait1FUC/sIaL958lv7/Is
Xj2kWGRB/C6aaHT3feXA+BAT40aYPxUGn882UqyAjYYP/GQvWSF3PptfNRMFf0fD
OBoWHLM/i6WRB2n3U8WNp409hgUepYG7FkhUQBBWSCKsBglmUlAGt8TRwOpaw+D2
24KpqODS0Ywg4MWOFnIty4enW6SO3rHd9XbAQCsoVAmeUBPvl+McfznAEsmxoiS6
dme3McoIU8UBcEhFcApou8goTWCfwTr5/u7G1aRqlMWqprY13C6UU2WQCLXKiDRH
V05PbLBx7CFQJ4fICYPrztZG/xBQMBk1f3LMRLzjze8kpth0WCLSfIWCAJVzt8K+
x/cDK+jQtZpf6pSRnGLwSN0aZKfrTbFuGPZu5Jeg9RB4wlmmcQZjg2X52nC3cbHl
SoDwqmKD9MH8og4J2JessMb8ODkPeaSpexSlnjsgziGzgXnXX0k0pNkQlPHpq0CS
pmCweKsPVSPOTUez6DsFrwTjY6JaUm37sLsQMOEHAJ3mdu+cv/iE7EGHsHnwm+/i
V8f70fKZpKjIcyuu+olkAohxTPBPzZncgKawFHf8sNJjiQWHYrhBpM+um59e8bKs
y/xVWets/LYdWbVlZCFSsfM/0lSwM5jDOnksA72+r9ye+v0o83OVE3nhkB2UD4ng
Q4kPztb8qI7KLdvHXG0KbUoG8fKY/BHfPujV4UBC96eX1WcVccorNRz39n3ShaIi
zZ+hSOJ+h90kxuNQ0DHjGU0sy920DvIhHadJ2pnodJz6fn+OHRQEzrd53XdYg/BN
hHKaXH7dN8NqlPW171TTZh2aGDdeAkpZ6nQgFoueCZ2F36aasSh9PLFJ5GzmM/26
D4yDO77xl8ihKQH5Wy2ZUc9q3SU1SkWnaCD3dVRCMgL9zOqg6i3Sa4GKRmW5qH5b
kZmOVU5D93RyW/t/Qu94ebYjFeCppv4GkNPOBRWLmyMx6HQCllBd6nV9LkfHzzqE
ugXBB0888WSC0waCy8uPvWyfwhouoGzZJCyFryTU3Z5qUtODxML7I2IgXGi4yL25
I0rZ767aZTOlnpWHjT3KwbEvxkOrYD0sZm8D65+9o+YRQOlZbU+rFcRXgG+1kkYx
IupwHvkvCFCTf81taSMdGBNMgJJBCGIbeDHkHCZCgC2WwgbyJQM8rrIlkc66mf4h
9Qml8H6U98qJgzinOoMP0r4RMFs1KNny+p/BdFrpwJDIxVRxY4t23jrpJhutHZvm
qmn5WSV5bygTc14R/w0NP/2/HAVNDAsMmaQuxlV+kFCRgQijX6gWgoc661R+Uxna
zxsqFE3f23cLRdBJC7p6pu6f6Navw1/jXl8z+26em1HlFalYiZOIhlcbYdzWuu0J
8xX17IptfjhijKf5yI2BgcMGhOy+UUsBR5oWrzRtImlhizOtNEH1vfs12pgTWW2n
h90aDVGBx+ostZI0ApXZVgu1xLedO9KVMH11Ez1NE1L5s6qnO8SqIYvXF1YUtM66
LzpC4NlTKb6PlSigHyMDBlLSzks1EB8NEEdq9WxOeO5SoW5zfu7PgQfjct1QE5bM
e6u5Zms2QYapkKYyxkp1KuTZWhRcTWR8hP4cgA4K1axXukAcBjj1AeuV9aCwjGsK
owpT303fThV30WHdySTQ7wGqpLkHvdEYoYfp8UZD/ZCvPbTBz880QE+bslrCJxbw
Cf4do5UonIQNn84grCjW0DzdipGrDMgjttEZyfGco7gR/cl+7mv980UI7/g8Zpfr
dxqJUyTMoKgzJFiqe7eZWyzwkIpp5xs2KMRzvTPvAhrVaMhxeCxgs6m+Gox2bupR
ITXOyxFe6N6qbB9gx4VXSpyW5EhoYZo4bTMQslHDm8J1pU8ZjDFzniNOs/QQq7aU
8oA8FLfXs2Qhxk1NYY1I6H/1IEgWsYbZKIWjl+q5TisRtEVaPT4Y9BAIUsHQo5Ys
w6ZohD+9az7f/p8GE0qBPFub2AtI2RFUn9BKu58Z5fe+fsINRpXardQMQN+Axrk3
ujbYavWJxl80qgdRrXwIdrwArEqPt+PbFJ92bqrgt8ML8yNDAQF1AXfN1/c0fTeq
2WOGhgTwca30MQ0XLq7ORCn/6Q5yT46NUzPJ3kH5N+9IhpjqY3uMIUW5IBEXcy0y
zjmxQbPykSe7eNRY/DHXSqPE+vOO3y2a7POPP0nPU5S+YDK7S9w/LkWy32RsVpU0
WDOQN7eUKcuvtk9fjwyZJupduNpH20pCRvB0g3Vsirr9Nlgfg9GCHZS0NltjzdZt
rioOZbcEvbbP9o+dad3cypf/wH0Kbl4W01Lt1JepFrdEjPmOyojbCVZtbXUGmHOl
0GbKjThfridO9IF7H1MkJzbJ8Qs8WOL+A7iHs4+m+t9GYIM1FSADmnncoXaWZlY4
wToXu081hOCBkOlkh8PYLDKQ0OMMl8fUuauu9NabqDOKmmLNG+8MDI/wSLfdP1pT
i/Nl9Z1OegzgxVvoc5ZPIuWbIU/mbKkL+sxw1K786wgHMU3LH1nZpqI/urcotLEs
1W1OM2dXURf5dQobYPDLD1+URYgWfKc7m7r6Vtr8YnGNUUxhDTJRj6Xl1ZWAg95m
bcgeDzso1S73D3Z5y7GEDpqXGeNcQvm+yRQ90UE4rIsYhLyolIwc2rKDGDq/NGLM
7SGwXOvkCR4j0vQXf0aiaZD05pC5cP+dvNhbh/aup3QWNISOCFYU291XGuSPBcXd
QhQlh64UQcfjdBmraMTrnoRfXa8tEJH6h22kPU3ttWToXOZMG3Qg3ez9zpWyfTQN
gOegyd+PCvb/oNHdgTQF7p732nJyt89V33vFVEZwk9d1qMo5SaQ4izWDDPb0MHOG
RbFzRtPn2AfBGCk1R4DBg7sjfGuMEhdxGL/ovPhcUE5VXqLOOTrXPHoSL0xuTRPs
3TngzUOtgomDxc+AIwdTfiGvr80GlCHqZyYYfDE5CIj7Zo3tnMZ9P7woa+8P6fnp
6XiZSt5jiLeDUdDU15vfmPMim6A9yR7QtxLL+OuYQTgu7vROzgiOG/WFpq79cpnQ
bqen1L7XsYz4S2MatUrXacvHMs76+PH1il9TN8mDnSQ/A2FD891fKJH4XZ99w9Ak
kqAv4OG9LuS1MxDEprtAS1rlxlxeKtBUmHUvdRYEVKk0JlT5GYbj28upEMz8MO51
1mPU+2SQAA6De7ID/PRAG/M0t4pT7+lq8LtmuIHEesGzRnrsBVscX9g/SG+6VxdK
UMTG5Dk+VAJQgstU3FnXjDT6UJqJvmsScmeNCMPdd6ZD7UtwhWiNuFA5k94FmoCv
opchMsr5ihHzxzuBNXeujpguKDxoNPcK3tsbdAqZz2TeNY6+3+YkF08QmEZq3QNa
k0wUalTKfP7sIOn5RRSeHCxnxfceV70lMzL4JkjUsrtWHekWA0jBJT7tEaYGt8VH
IWSi5w82ufONImF+sffzvvwfxc+7M/mzUuENztCxg6o2bB0nU9Ksu97rA7+HZkX+
8Y2jU8xqiY6cI0PTSEcuHUk7DUhlUNNMmgUQum6TY0HpafdRzb8ubmNA+fjVKejj
26MmRhKgV/Mgvr0qP//aV19RIuYigo6IcrJMKvwMQ4hvFuK043le2Ighc3ryyD84
su5zKDHpmIUE+Kg6pinPqgvO5EYVRUMJaC7wb2e9KgGZvjszLAdcuRFlzWV6VM7z
mMPorSpMX86JTYjZ2wlWKNQoqcUlZy76ZkwdoNavY4dl+CXqWAdYRgK78iwi1xBs
Ky1N4aU5L2IVSnDyZWjiO9r7Vs3vnk2qBj/osANvNvDV0jRLctQNHL3UHBngucD7
R+dbI/R3DZXMl8eRFAK+tpZ6JDZLsuuJWpJfnbOIR/0phKK0O8h9NQq4Cm6UdovD
31pg0bEEGKDNTyAncL3w9GQdrupuFcoAuHGXGmc5sCVbFbTM4dcatsXLipw46EEJ
Lxo8TtV+VMfr8xuMwnYgGPQ2ckswzjPHFlyegOiCG7+C0SKdh7z9oVArChh7v2Xb
mRIfXRSyh1u8AKsOS4W40aqIlpDqmXvUN5yn1Ljna4rNpU+TFBOf3kp3nfjjyrNR
eh6dwdpPgW3iPiV9CDkH7pSJyAV4hZZRuxat6LOAzVVow8aPl55of3v1udxqTGcM
oNUBddNXNnIrB4L+lg2I5tz9Oqc3CZx9B6mACJgkcplGvBw74CvL3jN4MzAutYaH
fWXRT8uK2CqSLhoD+XeJOMtqL1ZItO5VWctbixZkun8VyT7diVx8mFy2rTCDXgcU
XaYal12XJL4rMfAs2j1rBW1n8Ox7SO75S10tq8xVNHrMTePMAYQUp/jgiSSg7Rpp
szbiyd1msqn2rzOWGmLJj2NRZ1cg2x+CQvXdyckfyYo7u/Uq9HrmuhyYrmfw6orz
iKTU++0vAMXvA57xsioL3jyFIG4imQE2xS0lfK2Bb7XvUmZcBxdGjNzDMOVBfobI
seG/SBuxt+jpXc9DRLQswSl1Tk4bWtEEZqrqtoHN5eW+iry0e0wtosWhjym/4rdr
Lsws0wPTQob7bSn92unXgoKN++hmTCA+2FCUVwZQSaNT6+P3WembPsBeGzO00yDj
xdhHnwa945kkc4gCj69xzfYB6bYoI0XiHnD1j8tpRu9Gkq4RMuPfFfoHCEcKVzFU
e6g3UV+zbMNLJ2si4qorPs4PupR9/6DSNUfdkfi2mAfLd+AIdIymuZ2t53pwda59
vRwf/y7Detp3FVYLMMapQldI8k2bGUTKjPsS1ci9GBl/uVNIYXInq2I6WdFsHxdK
xhl6AMCj7SXrfAdU3MkBvZHHTfppJIu87BmPo3Bp4FXxWHuCi7CqDIdDUbuBZGE4
BFAWuSa3RhpdHuIiD6sOttX4QeqAIt1YN0BMNLxk2r8x9RcSW/C/Ll7sUPSakh/W
jiF39/P295JHT/FeWSoKZyja+jx1zlQC0D7fyLaPMAtDNVgTSYupiODIQnZqVnEP
zbzxyNaYeV7/y+hVBZeB/6CE0USDUQIT783u0+2U9yVnmArfZ35r2aPVOwfh4sq/
wcpl7xYPaGhEKpB3JNpuZjIBZBrq0ZPdMvtaj6nhGMA05HFSCcCqbL19Hi9RuSMl
b1GEcc70+G+5g/B7RIHCyq0BHWuIh6pJWalpfCWh5QGs/6H1QiPdkVbiM3TxC8si
GmX1stFhN6kQoq+A9EWF5USGBkCnPcL8Q8cMLIyyfHf6Hkyip6ntr7tD6hAfs8ca
hxLekH2IbfUpzceHSJLXTdbWpCQhP3B3xASPQGCR5GmABM7mc1LVXuMp3XuXzD10
YWpo600wQnOI6n8JcOdyhyZ41fV3+c6cYRpC7gHkgbyJxtQJCyf37TZDpBndDqjr
7kEZ6q4H8rhq2HH7dBR1OfIo7n6IZlMiOzJLmb+CR3uROGYygsPwQ7VL1U3Gz2Uo
I7Wbd2G1EmjbzUSkRF3C1WSvY5e2V+d8BPHFm4hyrhpTVJuF6/848MGYN/Vd6bIl
1+KEDi7jydKu9a5bwiVQ/G8acai/PdwdLJ73lBDntWlaQCtMKbzaAmvhOrQWj9+T
btwxxoQUb48fblCetdQivAUjCX5JK8AMrBzfAfQ0pfiTM/ZqUBSTzd1ogVl/pOOq
PGahOtKUK3hu8mkOtFmvuy8gEnW05pi8AYamQlUndOSwQ9rX+oLJ4l+jCGB2Xi3r
arNIy4TUPUrcfGiPt+wjIQQ7q7fA48iBXCfuwk+Wb61nsoHUt9mpmgd0r4FrBTM7
yzy/HzRoYnqmsjzRFoOO6oxqd559SnJK2SSJ7HKq8NbHetTgsJ5I3OG+ROhqnBXh
/W9Em8YfqTn5I7NYIeHiW8ZzFu7Xu//98U0IkjjhZvi1ISfQGXeNV+D5/caT4v1R
AvOGwfe6XkPqO1G9jDWPz6MHtBOC7hZXtVxvoR7XOa0PpdMAgdwsSQieXp34aJq8
xqf3j/NsL6nEQIpn8CHwb2eVxpZy4iZ6lL7vy3KGxjFl36Jdx8hjvyNFNl5bQRHU
kYkIiCQkmENhRYuTGSkWbZPjKgj2dD0Kk7nh6ziU9sdGy76R8bhtK0OFdRl7ufCd
Xvs7ZMLcoQ/1ScjBh010AVchfZqBUEgnTetYGtK8p50yriK7s6TfJUE+mxP1QoBK
dEalycsyyajNdeDAPlQ5xAs6EEkUBTJ6YXzT4hSnshx05dlFzIxz1t07zw1/153k
Oh4eayK6j1qsJ3hrazykLFSskyZ0fn0VkgZEAqckznSd01JdpzPHrB/GZKS/5XVV
elmk7/HTMvpZ97njQapyiSs2M2AfX64WeYiYV32s7hENOC17tx/GdEZIqta1kqMj
Pmn4C6lmlLASGU6lOIr/vwdY0xraIr67OUtciGZYHFSJAJfK2sreCnv3jffchwpJ
xuWFyr+S2UyutvtrWA7/iYitMTwTVVzjr0ucWCVnrLhoba14kEXZrduLIPkVP0PX
PvN7lEnwstcVjT9QnCVjAQuegw8bOdj9v+uY9hJbSLsMtoU95kxXpSXHI9aqIp8V
H/7Q/JdqqrChymeCNw9aMsXCRzIJjKT8WdzqWdnlby7HxtEMG+g6ztXHsrsmMCNe
d7J5KabNnXhThUivPoo7K0PqQyB7cstDF7639OaqiBYvBHJwhrjU+Y0DqLD6Y1Vt
CYptCRMPfG7LReGHxcR124jP4gXvLE3ir5ojK6ofI0Npj8hZd0VDo2hE0B4NbLj3
4LrS7pKSwy2C1eCOQFFjc0HQALlNLrQveInR4wVIY/thYcCjxfPE0Zg+rl0zhI6b
KXc+KWPomkPwv79z7CUyQ2tJegLI96Zj5oUSlQsAuNMeVREpXEJrrCDctVkyoH+u
gZd3y3b9TEr5wR1cKxXl64srO0ShyALAMA/P2bw3IWBDvW2noFEcwM2Xn1xLMX7k
wsEZp5V+rqEfTKDw0SP9V+iaPfjldVcKQgs0ev4Gz/dunJ3t0OIk1fdTgq2ES9Gd
mSdgI1VqD+aRnh8hVMAczaESbhkiAN8Vv9WqduiMh5UodirJuLQgTxfAVvS76Mgf
VLhPWHe6hczXJe0kp5kFLqrK3WFVDnEJx5UFf4paZVLhG3HfRxLRSgnUw/SyijaZ
gG4BQVi4dSxYIh0I2PCL+Ts9jRscTkw6df3L3jj7Kg/742YBLqrc1T0dwdGnfh9C
jWZ/fGVXQOLt5yMrmUuEKhCehe9ouK2GBMY7x0xMMM9cwi/16rJEN6MNp1vEJGPg
57uduq0tN9TVNvaooVHBRVvLhfbr6bKK95wNRf856TBhp/C9SYcPXCLmkr9x7EM/
fLUorUGsXSvlXGp2qF2omU0EA6vOZiqKHgpMLfSWv6ecMEg4syTUQ4VCXt5FmwOo
7i190icGsugIgcjV4EXUuQFFGNmzzAWlSzwAi5hdUkpyuP1aZG0KXC3p0FvTYSVA
MjuUNSDkShOeF1EJpDLAi2Zv0fHziE/KOcvkMIGAs7x4MUW+gv7DkHxJ1iMvZDqK
f0QUM1iy46uI5dyFM2oRzZPGYD2aLry9LfTcP44NpP8OJuufGLf8LOHeKhT1XxVQ
cFUZOQ+NWq2AbFH9FzDfHugdqsGJA2R9laszznHKlTlgFdvqDKz0akL+Xjzh7o3O
rqQHfAWqHaRKt8VsmBHUDHDd+fuEYE9YufTSCpvdBXUKgGWBeJk3ZEkjbTgLSFjc
4hPRk8CzAlBAisorhTv3xsnVD0s9l/yvrtyoABXx5fV6/1O4WgbYl6KPp3eC4laT
6vrbRh9ucF5YdkoR41+PfpJRzMODKTuDtVPKt4fQu6lDylyy31ynbDjTra+5G+Mb
fvgpymuiluq3iQ54V4vv9u1W9GMHXtKd4p7Df4idiZq0c7vDsHEzLDkayxyFZy8o
CbmfVitHIaVsjcQxavzqDg5J6vsEOdJPBcvP2B+1yr0v01XF299ra5Au5UfFuWEw
Kk8XRUSs3DX99+Whkxzdg01IJPiaK391RbMf4QPtiQ4CI2Wy2JMNQkzAkvl4gVxR
YME0HXZsFkY/Qa/mDIdzK7S1hXWi6fGt3v4Dki8lS3wcyaEsIdlRgvadbDKEMOTt
NjxC8pIvu7v8JzCnXfgIem/VIhyDhzbe7k76Jbc51Y0MxqzP+wq4yIJ9+mRZI283
k4NdkChgwpxecAvI+vk29JFAaPfSp+x5ujmS0V0mradxRR0FlmBQNWSljHS4BUTW
uIfRudrLDNmnPmQ7Q+BYpICtGtbJwn/bOdzfql4xEIevnbLZqmZmssYr8W/tkmqw
Ds+UEqBrxMomaSA4GkkESKZmvT1C71+16Z2hJguD9zGQDdN+IJKymtcqixxgCBMo
LhZ3c0XNv3uIvWJHYc4uvn1xbJnhRZ+KhOZ4od8OzeeO4bY292sNtiIbvDPTtWfi
SSqv6QloxZ04q6CF1N5TnsYHVnO1uUVTl7Ec4XK2r2CQR/dL9IEsioV3UTYXpwR+
5jEI4WtF/LR2k7kAGx7SaQxX4ZNaKNtHh8lM0VfhEtWth9ol5JoGcyiVNwmHBH7p
mohWU3lFQThq/dUdN8g44c0QW5bCLncOIoVUeMy39PDHsLjC18yS95HvFvwWpVY/
1LQmL+1uysAkhzCHeynHki8DrCnyv/OAp+1TJhcJB6V+V4lbg6IPtBdr9n1+zKIm
gGnpgxQu0DSryfqKLlbfpjvUqMjSTBXG9URDJRxcUSnHzl+vO3qaBvyxAukV76E/
jBz7wD8sHvZmaXNVfOlKlichFHTsezAoGwk3WXeCSX7MMayfLE1pgTbhkp1oi1B2
rDCxNdcE8das/v12jsan2wp4QrNVmMuutHTyUWtYYxIjm6QrrEL9lI+FScJCSB1Z
YNgKOU4L/ccgqEC6dGyZYrcRQ9VX4dJz4iaMHm56b/0YWRb+7IVE9fS0xXHF1DaH
K7UmSbCaE2I+WTgInjkTO2hW/wqos+7i3ua0OYKSM4H1ySjeVswUxnpb8LAUDMGw
6tzBKurisukOTV6TCeqqToJhW9DoRCMb9lGxPSTKTegsXc0E4prI6MC6pUUfNjw8
3vocQt5WiaCDqV3KMg9HIKsQINyyKpaoLVr00Nr9Aw5H/eqIIGyaKnpncVGjV77f
nNtyBFA4+Lo9b73S1OqGt88np4UgtxqCU14LodLbCDH8oHhwhCMKWtEv+Mk4sfTo
KZPH5HhTLxEtfMvmfWek1zSaH3km9S0wp27TGthFtDZgCFmdy3/1E9POmAJ3Awv6
B2C48JYGq9VyWAOYUXanerucvJ3MXEyup6gSm50JC6+sAJnzBWXmGLmLBDOFf9GL
Bna/Z2u0AK5oCNN2pBgfipi3rggc9JaXrGexY7SAgvu/hWVxw0AgbTpK3dz0hxSq
jI6XAZn1CF+eLTzfuPS4nxjIj5Osc/RSEXbN6WeDcIDm9k3eQlDk8yI4WuTB+kSW
1uTsCC25oVPJsPA1pL1ZPnnroqEI+FlWgGc+mQS8t1fAzaxnbU7jQ3i5ahemZlbh
Rzw9fo7SGg6zeCE7VJXgTBMoGed0kBrE83LZ0JzVtu8e5jX4ggL/9Emg5HG1wohK
jfKHPlcIuZhODuCd5Z29HHx7UsSo3QbzYYkhJZ9F7860nh4vjYeFs1HIpVlr59Wj
nYx9PpM4P7qkvQC8galfLJLEqbi8cAlRKE+7rbyHarhia+WABmY8Ju/fFefkdWse
8QxY913ptvQakZRwvRL6TtFD0UTkQWdPB/ST/By0mqp+jXo76yccYhYNBhNF8e+a
ZlLZjASA5go77kRFTjqZV7YIrTwutRIpQg79V3cs+foGwJWpYa8igjUONHZn4W7m
GZAr1SYA9Y2FdUONj4h2gX2OtQg66BmQkknDpRQbyly3mQz6Mw+q//8ktB7HFckU
w6Q0pxSP17EcuZC7+Nr9DgKIKOYwoPerZmb+rEAm4TKkuwpFqDiU9C4Db65GMG94
lJOrgJywGesJQPTrzs3VGPXF3b5W4Dt/zQmadwPu9NwMkvdqbtRZKopMKTn0eWPT
TYJj7tLHpVe052rA/NaI12Yuhd4fC67UB0zlBvUfXQpOm8/Qu7b2uC33497k1wPK
NBZtARlxmOA7kPpcoKeMo7Hz1FWwox+qU352hjmhhRWXR5Zvqn0RgRMj6Ud2seph
C1LIpca1sMyuLca7iY8zPIgk8/9Myp9UHRxJyq519emUM9/cemS/ZVtmtxRqDB4p
MFY52MvnQJSEcp4QuU9N/fI/HmVqAbhw4KMtO6Vdo+oUuOvm2PqEuaZwYHpxAgmo
bLYpF/mfMnaR1buzm7g9lCysWLdGBSPj2vj1sCaA3uC1OR6rLG+oaVOV8U7l/64d
A+FPcsEqehiqS3wpW68UxZTzDcxbXVj4GPnNbIxyxPug5Rj+tyrvzibnzYi1LajN
VnSxuiVB5PJG2pHOssKtqcUVBKA51ku79WdyNsQWAaWSFXqzs+PGXHWol7zSqZON
wFce+ZQTPGUVPkn+FXT1Uv2poJ3pM+UwUGLCzYVJqKV02HheSXR4TMMyE8GD/lrz
Pv7oYBOPHNIq7TCK5ePVgv9iPTGzx5H/rzex72AoTdyiP493xz52Ou1XpBry9Bsu
EzsPTbtANQ3AodA/09Rk7hPbKf3eS35/WKI3EmeU9dawxXWSKzzC8RBhohlSmjSX
oUmTu0Qg5Ct3IP0klOrcpFW3kpIatCTFaw2CdmhJCf3BYNj1U/9JBE30/4QeCzD5
3v2NoKUPx0nStHBo57e3TYfY5pzDPduLavVAf8ynNUzI41KRGUNDe0xcEOkqs+oJ
JX70/JOTPSXINCdm5QYNiVlxJJRfMrzFgwwdUwmvjU5gJPnST0NboxLvB3CMu/vg
98h+ohZpZ9366gwqaXq0lM4pF4hhBwF05ve0mZh+5SZnFSPJHFPOs8i1T50Y7xAM
q4B0pbHGfu6VUHWND6u0tUeGQ+d9UEsCY6xS8cAuMqSZ2P0ufUeTlQQKtKfUOyqW
AqO67ZAERvkbCeauA6pqF4ABeitBthOzSijO+SSMdPS85dtzphElUowXn4jbMpx4
/U/2tYUdMl3emHGRwV9c34AtutHnI3habj1bawkBuGQj53vAtmmsaOeer1Sgu425
1AjQ5tabBP1EzhP24XNq+T5kW/7axcYB0AI1EChb9pqUZPthrS7ImXJE9JexGsAb
xyfK+AnSRsWlHrYg4gNFQOTsc4ezBKFBYxUwb/9XNWxh+fK6faZp6eE0TO9vwyLp
yryRSODRWDWFltjjgv56bWdCq7iD5LfL9hZiQTgGtKMdhZ2BEaZq0gk2AAbnP5f1
VOThKjxDWbqrC41rODUAB4q81/6utDfZigVZ3hmqvPeNpNupv/EMMuL47GcyPOQA
MsJgI+58EsfknLIfsdumqQUc8I3CYhBYpLpyoPbx1QBFTWkgZM4ww9n+N3nW/b1l
ChLVGILvkjIo37hC/3Z2QVvOoo33krlSWMyQm6R7LrTfKAM/LD+xvFqM6TEBpJvq
AroeHu6gSfH3SlAdQ96jV0JbrtwCKHdbfB/w5t8gpLAcF2s0m+sBXoEr7cKtLqdc
cqHpwavsPzG/VtHhpPaYy7c31noAGGNG6P6BQphpGXmEOyDs3MN0wIW1w39bICDJ
ysEPxcL7CJ1oz9X034U/vzgjcOMM39Jvjc35jDoIDASOMvSIYikQcrTyT/xxEj97
CbjVPfbHiwE/w0TxvqAJQcQx6+3SYL2WZQ0OY3g8RbhukOcmi7TnXH0dIBr3OnfG
k8/o83p4ETh+HpCSz3DJY3JYDumKhBGwUQhXkbGGaqEasI6qXi1BP0bzPyWMdNS7
oeFOB3TpGSG5DdiV8t4ptuciObuJ+rujaB687RSeLRWVZoL52k09WuQri0E53cDy
DhVk7i13b5ZdH+wDMuD/S4NPFbwo3Csvw16W6NXPDQ87ybYPYa8jzP6pD0tC8Eky
A0TcHVuxU4ibj4tPIt/NHN04fYkSLik8SqXXLOUGwTeLi+DLxI87qLDM8Slq+4F3
+pU7ObsdtvSlCWRQiA4eNDJB8dDNUPDgkjOgf7vmGqO3uG/jmq6OlXqiJesy5xiw
oO4wkin3hlemAGjxunId3rgPpv5FzYVPJWQu7gRmM6EvUot3Gd5e7IOXtCu3aBk/
lwV0vFNvYfxka3o1BZuvOXCc4ZtCDdn5wIopC/vj5OKIZ8/QLu74XuOfUtHhRalJ
AFLwyD0A1+TNfHNQQTRRQUfGXwJD0DrWNqtDdSb+CjAf6Ktzf7+LWHPpclZQIQjY
U0MrTsFYayZzVFAf7FGbjzgqlnJwh044JmJKXgmuf5uaExUqf24RF0y0IEF93piD
A7dIHq3M5TdDWevGH1ywAKVVN21KIynyKMyC9prxkWmMBfAi6vcGdR9ea5aDrHkM
1UyK05Dg91yeuPXxs91pXLFxy3iAJitIRAZU1PxCPCwvjoeQTgJXeyCskPgJibu5
xT9aHeApaVu+SITeVNyNBvlRCHyXBSvMuz/P2IMOSgDVYpRFuqultLqKVzy//1HH
2x4UxQ0hMxhx5awi+4bPahc25N8diFyI52ZNOYD3M5DNisXX7E9o0Uj8FOo4/Ytn
Jq+qi9LszCGE0B0xEgYdC3lPyvFR7HnVDxKWuXc57ddUQyOtpU/XmXuIVqaWghvS
tCZ+4Xyaa0mWlxAW8A+542Odn7iJuuAIAKap+FiFPcnf7S86R1xi/NEMQ97KNIZK
HR+2WIiL2DTSq+muU+JzgAhHH5+wYhkR9vREQli4GR5XZTARHK8JTM+SifTXjsv8
tZ0I8fOvZjJh/SFBaCB6JnxfQgoGODV2qASPzpLp6fKB0j6nCOeeTAs+puh2y/j+
2f+/DUYgLDbz7s1/+W/x0NCNrtrr2+yWQU0zJ+usf+Sbq/vD8EmREcJThXPZ96t6
fLWqRRGhYwnaZ71yEnW2+XPncXvhIuTh9NLOOq7Ent9NWolk9oncPcn3l1kJPCkN
7Omk2YhgOWB4GSfuBqtvPeWw3tu8TpJO0p01CjJux3pvw3D/xfdGz9YiMvmXBp9G
z8DhSVpqt6tIXtufEOxrvPPxritfS0PFOfejkeRCeLXtsn9M1D5dtY2atfCrjEgu
NTzitG2L8UAJYYPxEW52YtUubn6/Jmp/CUuLl1BenTGcN8/gLlyqowelTcCxfPL9
/G/R9qdETeTUfywnzz8O4JIzyRNb5AaqCRjgJBwIJ+2AcPmLwDxIsiDG0kE5BN4j
pRuaQbqSeEONoyKIMsiHg3nRy0S0uQRTP6YumPOhn4qyRaO/skCCvNPg7NF0P6b8
372/scDN5miPZJ8egj9Z1jGyVvLchgTOp99E9PrW6ESRj6T6x8+I6Gxq6XUjGSxG
MnB4iy41r43+0yYApnsU7cp0KAvoiMgfMOsxxbXWkPs+R1H1A8eRKAGs69qfN/gs
2aalGkRYAs7iESV3YeHFIrtBhTZsRIEtbCXrHH8ghv07pZQyXAvzlXCANFWvd5rN
D5CbBYMLXZ06vQ2fwL2bESIrO4H88D8OgwwYeYskrnqQDl09fLXVo6LXBh7yoh1k
fYkgRLhHMG8Q8xiZVH44/GFvYGHpB32YGsuW2nnBd5ISK2NEP5u4K1QesVL39+pK
ObN9hYgf80hAWNX7Y8PlXB+UnZ3S60xlD1WYDTfQIBF2NYVRJynpODeMKv/SxHm/
XR0f82xulBVC1dsFTg0awESCA3CSoBe0MWLsuRiBwrjwJY7zPMJ7tv0GuZXiSuc6
NTBIXpF1RP8gzE8t7SiVNUiw2P0tPKYPrcLE2ZCjIbBicSRvMo/UDZ74PEbdh5ie
EG4kEDcArJ1RAXCmDZbV/TuoKujqUXF4TC85KJFq4eBjZKAEmyMEJOGw3d1Yj+Tb
qz8RaZEYxE7hdodvPfXPMsXrXXP2x188ahZWTFQcb7o74TuNN36pJ17zzarsUDAb
+zETzBCZg/hwyd8TtyEc3nXOy9RjoGZ9y7JeIDKruIaoOXIIIHGY4FEO9L7+uiv2
XBM7k/Qm+Ya4BstuDc+gpfhmSCOqwVVJZ/sGIAOT2aJAwHZcTPYU9/uBMGcex0JQ
/LY/AdGLM62IGi3LbRjt9SYJXQ/fIKCkOMEZ4yPqEKV89rqPcpk3PAtsCATGzd/M
OMiJlSgOmkk0oW0EqN4uPRDZICMicrvrhDTGxm8H9SrAHdqQFQcgj95Se5svwBYU
OcD9UuALAmxSwm0lVbjVROJ5dPLQ4RKUiF79kg80m6YP3JGEMkaTJHRJmuxNGrcW
OtXIy5d/JIyMeFbMpHHKBF71ecc2gUkUxfe6igASy3H1mxTaTnkdH5PaJrVYlSCZ
oo8QKnCiaMW83haIfq9wvG0lH/Ve5jw385aiBMjCbn0hZkE++y9DfEfakcGoUvCn
mciUBzr0Emv/rTcDBT0NgltkKJrFkfwO5EJBok3d3cdVDJ6OPqrfn7ZNEWRB06j3
Oe98jxrEjva87WC63kJ/WJUMDJHEw87DSTvQLLfYrUaUNAkfWL7tM23Fll3j/+T2
h5qfjTfi80kQHhotYvLLHzXwT3bD17yzAAfidcs99slIsUQCucx/hxSm/+vApANt
/3Gz3SkYj9EEx/fSCiJmkIkXZpnLkWky6kXoUPV798AqRaPLmPKGk6GwgqKaPGYt
vnsSHMb4AGlqYXueamRlLvoE8BRlMD1Yd7fmZUCNpQlHT6D3Ramx4UaobhTR4R/6
ZmplJ1sq7RpJykgmUMn03ckvy0erFSE1lVtxGRRoYoKMg22a/epONvVpR7m2y2yx
goOwsGtI5APW2fCZkHwEdCzOHuH7wd/uPA0GOLiUV2xhWFmTChrzx/t4EVleSkhc
t6CYcQZJkMxRtu6PH7DNnY8hYnFQfBCV5EI+e2bS2ZYIFuvOxRUroEp8gaw4FfZz
rSJ3bWkCx5rNkhJyGT7fseI6NyPqw/Of3bXURM9u49celYJKmRhhFdldYgFnwFrG
EHR7SZrZSbuzVW+12+IwpTcylA5KfdLA5yMdSlK6l9d6SuQwSZ1ygXcjO17p0fEg
dCLXYcqlJtfp0rIbKZmD8R3dzG+IVbv16CgZXj1sJLJo3bVXNlDhOsBkkeTIQXxN
DjpJpxHSOvBN7qMG41XclPCk28bftDgsbv4c4HyjRxka6szvTkSXN425+wBPVDf8
q2Br2L6ZkVCvj/TEJNwL6V7rkeR6Jrn2pSr25qd7pv5dx4cHsnx6OHHD57BPs4Zs
lwDmP7Jk3rL8ZZrsDwOqlACz9p6deIhavV0LFXrnbYEz8dvH/X/DeJa0E2xPZntH
WcVqGzgxsoHjfWox+YwBnyp09QrSXeK5bSWK5ythgECA3Klj2piAhXgZI1GVVz8s
W6UEmCmTHoEZwnhIHqXzLL9vmyWiL98qALA1m+Lc7zdc5wPxtyWcEQqoes2XGWkv
Az1gGY0LPuKoc2vfRWkpBHsUeWhYvD5no9Po+437lvOILuWD1JBCgT9QivYWwKVI
POph3BkL19bz5IfJZMF32OEMu6GHFz6G25u38TCEWVCfQNKK0AZv5xDfEVe6aESJ
nBtjWivROD1eO81EToiMLChB7Zmghdl2Y+Qgj2vfGJdiAXlx01wPLOkrX5NuVObJ
FZdcrcrhzVPD8oceCG06kqE7zSy3Q06fJRaIYfeUQV3pAK6jL73438ZRxZFANeoN
LkupiMBxYEq6kAiS37DPpKianECgK2/iFA83oMA86qP9QHsYBp8xX/VlSo+u908X
SRCwsaFspvsNagIekwjrtaLzostowHcsCbIAYadnUvSs2jAV2EHVfXekCA0WszAq
hd6Dc3hF+jnWKT1nQGbL7YHpnBNltxry6cghSYevJyHyCpe0pOEusURCWpA6a4jT
YagAlb+mPQe7MZAwitb5+mtqKv0Q46mVLkzcSqYHU9mfzfTnqcEMqgVTpnmFKj/c
zoeDzkitTE6OIyqRAJ+rBuAqZlNnUp8Aq/EbV4XTMUWK1jUL66jLDragqH9gKlQZ
Ti+23lpjJH2bq/dPFDyihnSsYZRyoaN1CYZmlS4oayyTHvvaI1trj89paZ5L5IVS
AZFcdwyCk9zfY/yceWubO5kr7RSY56vIY4cmopPd/l/6YCUt6Ji5WUzhBHBAXkJU
HHrui4uqmXX/nvPMsBL6gPlBcRcwo1/GIubV05SPt16MCf4278lrvaOkd/4FNypG
Si7jWNZGha/C3Cyxmd3zAcXnD0+OUzRZWpaJiAK+0DskzX6Kf/IQhdMHWOKgA0x+
EKQoxIiINLSbgh5IDGG81gI+QWcnPDuGnTqi6WIHjX7Vk8BMD9wcP2rrftW3dXhG
PjWNdCOVJ7WAzTLFwSygp6RVwyb+VR1w03nivW6fKMaeSzpSIZbl8msIzJpo/i0q
WG4i/QWHfD2hmmMTRKE6VMJjcIz69lF1YowgbaeSgwS+Wjd38P4EHIQfKsvLwJQ+
SI5zQ9l4ECBrADKIlLr2Np7/NeYx6pQ8e5c+807xMBG51MzJrWCXkQYkQuICL/PW
5Hf2bE7IDUndexep2nTa/dDNsSyAsaHyZxBCZqI9a3IOQiTs8rAA8RExraZte6FZ
YxxmUy2Hxz/jWDDOu+D7QF8N6rHB2zAzqjwvHrMlWWCWCT73RXUYgsYVZpAKP9RP
En7pJtko9LF5Qk3uXZQu0eXzMdkrBTnj3dQqQ80iDQRc+oVPm00Xs8vnDIV9TTmp
QyQOOlKtOlAfpZrQaYjMARucc+dnshzOL2QGKKUSghj3dWiThfVr7W855hl9J9Cx
1vh+c871TSDBBQJ5UGKVQJYIlt/9zMWPnGdjmdyeHzy2sKKLlzjTCI+W4LLEO6NY
vthTcyZ89/Dw8Ekas65vJtUPYz8sIkE0fsw8WA3PEY/wZxkV63DDIq4WJCKwFrcq
a32UDo93OPrjhEOorbC/Rn2EsAWHDb1L0Gy9D6CCHVVg5EL1vi/e6YgjZU9xTVi/
k4JRzvvaUtH34M3NEHbmoTLqZvFG+75WwDTNSW1boPApr5AvWafBKZO1H+Zfrdn4
Jstf8B4e0MvYJ1YjP4yeqE3KgHOpDXCpXbT9J34ZsAHwUtY1qYlY0+IRXTwgCW2S
PavWJlpHiWiYnJ6tFdV/MgVChZpO+Q6OUoxZQbscFbQ/oc5C1rsArESuNerPtxCS
iziebSbEnUzFA2+ZQbZnRSYRP7oAaaSHaDb8rmjGKoQLC28yoNZdAie1siDVz/RM
9C3b7SJ6ssQovLLBZV0s1Cp3XBqwmw+sdd2jTLptvxhcS/x7rRrg+k3rmlE9Vc9d
/kM7t93u4v+JicayvW2ftKjTIHPwkas23n5wuvJ84tnAD9SZ+Ijp2Qbe/5bwsTOg
pyAIgPSrD97jLYl8CCqbuUx5UgMT3EBpyBdGlnnjmw33cjkFIqU7tiElJozKjRA/
yfMAPuoqWoRgoITTcaGMIFmjQ5AQcE2m5nw1334U695pOBqQtcotPg/cBSR9Y2B3
7lqVo2/DGMwrh9AXovU+l+ApHDIq6r0p69ZXyZYr+6GOq6hSJsM4zXy//Yz969Uy
2I+1MO4HCgvZVCskkgUcHjm1qkmlw3PtMexKDHBlWMAtCo+BKJIOhePnCWI1HXrY
ahcF+WZQMOar6Ob3hiu5daJBccU8g33Op2nBT6gNB/QhcGrDPC1dlGi+WBRs1rSc
DLC400/97BR0uucq2vdFg10fWJ+kbjkSNa8OMV2HMKsZcF8AI2RQY2jVHz/4JpcB
U6LbzIMlkN/l1ETbLUtCC2WAhwSFvucdMMviYxvzTK6P80t0pjbvY+zHyOwgEHye
jESrlR/PrE6CMxkjXonFJp2uyTLr2IuKj+foDD7iRh0dfd5BJmgSX2B7o8O+IApV
i2Z+cPU11Np0209dP7x8LJFk1BJ5QH5qKtf8jRaQ1ao9GduGj5FYkcetVdPSq+dE
rZ0PfbS0kiPZHuZNgnDHwkY77UjnMBwuIMY1W/1cW26dj506A1gDUonqbSPzJib6
Wwwo0eDBazJ95TyjoqkeAMdC3mardrQ3SwSpRmpMwrCOzTX+n4gbllFB+iRLmTkZ
J+zxLRMmJr78pSpqjGk/ThU1iNIgF1yI0hhE/Jao9XmLg+W+ydD8bvJv968W/6Ie
27n8zqtEYfk44ml+n25Rwi5I9T7u7dbX90PoJGTFOLSzGq98n9jMEfGO2KVvQy5I
c2qJRAg5AeZMq4spqts5qRDKpENWxuG8HS2jo37NfRf2/X8N9ttdYsiadqZRk8/s
sKQlAHIkB+J49ZvNdC3Xgcg1iU8cL41an70v926cu1UY7ViJtGCWCpXAUl3tcfGZ
vtGcKeNAtwA7EnGNhanNGKlV41mnmqLC+E8yXU/QzuNesRKwP9uIVjOfm3mlKBxe
LzxHBtwrk5GIAZocdzxBnkm/sFdXSubZ+5RTnHnbyWqWKcooGqcdnz50AR9lMLD6
535ASwZJTcz14nqIPoAF8h/a6vyPdVBMXxr3IDBwcxpEMW8bDWbPlEUbSJJ2qMIE
QGagNshQT1w0kygHqAsVcuTp3A8efhnt3mB6GQbwN6DfrJEzEyqJLEgnsCt707wb
vneIDxwlm1d8T9CYyiUwu0I1pC6UTqUDyVn3jcpeNLe0zCnEjc5wsehCj2zwohT7
tKDVmJm6Gm4f0EyzGuNpars6iZjks7XtfBcRFI4Q2lxRpR2xEszbEjWijboehlTG
E4lb5fpRLA43HXUdjLkE/w0EE5Qmk+E0usWfYq/I6Osqa4Ly1IbZl/Sy0RK/per5
7X/aBWAu/8xSeLpSqP9IhWsXJu50I0dNPhOXS6JvPsgqcKuM0M+J3PLl+Y6KDHmG
r+4Sm9uF1tlZNa06uiWDjunwBtqjsKwlBUMzeiinK7qpukMmsSeBGYqRGbRtDyEV
t/jp9uiDrTb1HwGAnyNhStchMc5rtxdRDuFBOkDe+7tcKQrPWcC5ajS3XuuJwBBB
H5LYwBYEkX3VfxJh3Y0yOe8TORtuMwB2OJTMK26L5YsYAYEUJsATCV/oeOvq3POv
h6cJPw3e7ITrHSEzZVc+TMOazKJ/5lskqP4qoeQCEhp/vMey2GdzFjOI9OM84QDC
3kkRt+24yEMPhWrRQk7qhQIXFJ2B6U9Ci8cqKM+NuhpTK4q/4mZQJGrAmyVB3RyG
nIMi96yVUjllePbzIBzNFw7tNBWSsUbTYvBJH4yEIZ4QWjnd1kHCAVYcFjdfbaQr
AMREtShbzgOGDxDTy6HNYA1ahnhIEw1SYyGZW9RIVimcq6ogNmzSrX72i+IwE+ku
GAlYtjwjWpmezeTXQRY/YnUHmlxc8pPCfzCfrCbR3nx4e7S0T3rPmQYiNvC4qrlX
LQxFH8wy2dLSkZw59n1VkrgaeTzkNNMWO+gGnv1+YGLZgjubPr5+9laxofFUiJDR
cjtEIRF3xY1ErU98/70//3JMaNtDhl82R5ipqe4shL6Ecgkz/hd471NSnpsaPYmg
WRdL31QGHC+a4yiV0gVnKLVFmmCIeNJL8wf4GyFX+Pc+Fm9kBd4Kfp46Fz0EY0Wq
zLcDy8ZriYKzfpLbR8ZaggfFy/wYymoJjThZIQ2FmegPxJidhd6kHgUsHknMS2H8
EhnpLlI37h7n/eZgXoC81bobQ4QGqnX1UmNXZSKYPxCfSCh8CZT5b6ustaMMi3p0
BgqKXlvzrhIWX1+D3+x/mLNDjRuLNoQxWhSoYOHNhj0SViDcxueF/Hh4EjJj97VF
QyNtMcgqV2RvRGuXND/YQaQTIX10uoE//6t4BPyWxrferaBLpOrOUftvWh6VGDGA
ePg6Sy/Y+gm8PLqqDYxS3PdyHs1qSNiHF8feiPGHqOlXQBLEsevaqDeteVceKMCs
OWVRkE/mfQgn2oR/UMwz9KpHDKVaDWc4d0+LLDOCm4c/Qmqszq/SjRiTycNbAty/
eCKjHf5CalO17e5Q2OVdbbBENuGYAHSxKEaMVAZ6jGFPtpYZ0EBQTFKwBredrHuS
Bx+/5mZMxvBrXKBunu/xcXmT2frBe3oxZirAltLyOyPcomcT88ondXlR6kynYEEB
faR+Q0HUtXjL+XzzAkRO+L1OdRlsLiHwv5t8tta41vhYnCB0qkliTNSc3iB+P8hV
ZLBlXu7Kvs+gW3F+M3mQP4a0AKrIyU/7SBspKGLq4WRSGEALIMYgaQPYp+T1qu/l
08INOSJoXW2y5iV/NbWkwwLDGylRVkI/bKQtTPrsjc2PhbBmoeAdMEluPulJErDA
CbOPQOCuva10TL7+lhSauchO9XI8qJDCpq/Fok2h58J09Z86Eczgi/PBgBMTTqWc
YrQ9nRo/i0t3wknPKfIvCAbMOTRf356pjgjwDbPVCeJSoAyU/ZzBkw+vxTKrsTpK
VYfoUbpNpaz/bUPm9c2jvaqMmlMDKor2+adm6EdbN0DsO/zfUe3igFPhmzbFT7ss
UmSpMA16OVTsWzgyMH4VrLDGLuEM2+wAKNFB9q7SRW9Rk4NybQp06Gy1yLNY9Fva
3WhiHMYEgH55QK27Befzj5eBaMeCp81N0w+BHwHMB+Q2O/+2KmEQF6tIVStTUmhF
8PImCcH/7oqwbdk2MAmSn4W2SaMU/FKuCML4WbULt9QUl9N65XMq/uesKDTfTfiN
ncL7bWvIHihbo1NnK34hnugMLMo036dy9foeTQqNjGCs+VpC2pJX0RPbVfAwgQdo
H5EmxomVVEHFmFdgKIa+2ZLsIXbyCKlCHA76FzCJ014AQbjAX7vBGqifeNT/1oCv
2J1o/8abYe3DF765Xv5sWIgqi4TlyZ52zbwlxwe6XU9Ymaj5S/vAyplvZjQgNbZZ
hnsC/CpXdWmbSH3n/oJxmDOi8bFq2SCuY0tgsKSucb+LEbzDDyLuYRqedzcOeEPw
RIvXsWuskJucQqb/B3gCZCAr2VqDmruZf+PNkR27+rqI5PcrMXwgoAMx+tuqAUTu
hhlxXXadb6fYlTxtS8dyXzXpmcI4WwKhqyAUE3E39ogrYauko8ST8Hj5OF6hJ9W5
wRlo5jTVx0lukmyBHb0M7Tfqla0wYCMlBANw7nNRARqazsiLtSZ8BrsRaC+J48FW
knn49M7CzWzxQPnyPt76/GZ3ybneDdB0FOqVE9jo/Snmq+n9e9Q9n6O2c2WFFcHv
ysBA3o7ata5hdhAUoPUnGR3cQKuxYJ4TrQ17P6l4mpEgOtTh4DBW1mLl6Z9aqPfl
cY0RYYP8rjZknWrhi5OrACjcvvf9hPrkfosHwgHXgOqq2z2elT0p3EkDbUB+8ATy
JI8tnEeWCrlVnGk4Q76rZfwqQL2y8ycEJ9j8i0MMeFYV3tTdU6SmNxeRPWSDyaLb
79V+p2UnlzCHFGgn8pZcfVNDeX80GKrActfkQYrzBRrRzEbQVd0sbmfFre9yOxgd
Jj73m5zgbV6OBjU/ccAfBoa3EY/An+nVPhM3SqAJhzsp/aq2mc2YSSoINhb1siSm
+cwsLjNMHfuhpMuV0y9NUNdwBDtKkouF5+ArhA5vsgLD+/owxzO4otE3kL/8S8Yc
jgEbbI+roayWg8eWCzTpnI29lYLRYKlO/ocNg+Elf8BmTuo4zha++Y968QWl0qEY
Wj/TpKWbOqtrRnT6wuvGwMPAad77lHpw3hjZ+WBFywjnLauEos10zQpaLrq8OGau
QZRLDP7tc7UeRzc3CC20y9O7r9OWBbIBijEyon+XJbMpWvGvi8Uzy7x+QSedlif3
1oVbjUUI7LIq4Esa+iIA8Te2C2OADmC9/sNKsu88R2JEGVt7fWvPtWRzLTdfnlrJ
ZR06P3RjSHejicgqdI2LvCAqp6UmdgAL+6vLcGZNNbHuMZv9qYcomEGC4l3GM57/
g/4/yq9Qasm5xaO0iQvgWsvmusynFZ4/BYhsW0iK5Nhr6GlXBVIuj5Tv4vqwfJmn
9nHsFEKLPSME2uDdiCuVuVDGpp+2Fy1HKyz8HR+XKTgZS7QZFHXqZBVU1+ofO5P0
W+kdwapT8fEOeTGBHHlVsjTQ8MI4OZDqWv36z/4lS0JrLDhmDb1nF6dCysTWm7mO
gYNU1EAaU1xLFzhP3fmVTBP4/TnMS0iD02SvJCOuPdav88c8/bhZ39IC7cJwVdDk
f8DtJNCAgY3b8QBiHRpTuNVR3ue5+wOAgVX22+pMFyU1DJgne6HM2+rjV7QlxkkJ
vlVxxTwiURjFRzlnZSUMLjwb1fcMhzs9RNj+Z7uwZ8m5c5hrR2y0mXDHIQcFq+9i
OcdsXFGte/JGOE3L8axUO9WcRlK/2slExYhm+zHWjaBG4Cr4+D7AcH+8Ijy6jphA
RlhMmfRvN5ZlgfoA5YgI8LBNNYGDPoXuFLapJjvrD9IUaPAFA46Y3nE0nnUq/dxk
BNdVrmIKNw5p5QFqciFmEE9FAoyhaK3CjS3yURX35bP6ow5EfU7FWqC3nHgdOPKM
ddDGp7P4vgh8/rdb5BJnx8ZflX1nnd5ci8Jy39GzXVpAW2wSLlcYXkEylTsUTEVx
4aFMvDyFzFU3YIpq+h30e+m8Zhpa0f8fakn/BYUI08bvhQw9Oi43SZo2rmOaaq5Z
oXuXD6HiEVlgHFVwHLiXRsdxIctWd/xwGDPm1PU+AX4DvUZC4aozi0qUJTYrJsSg
oZhfU3ZKIoBZg6qUhXGvnMQAo3BOCNLCUmlFaXGCaIE6eAdyyhSxryfcX6nrS5Ep
oFIDz+pNbFLJv1bOk6qrrhxI/UVrfewTo2Rdq7NUM+yXJukp2WrBm1HQJejp5yVf
1hLwaekL/1MenUSCLDZ2x9GRi6m51CjXSyBIpx9MaQSSS2H9TDVLp0H4HiuLWNQn
M3IW2nYAHPOoWI5ypH17w2eeMrnw1jwK0AvjTAPtoZhBp5so9vpMAD6TTfPTuHu+
gae9LX9mRkgYAvkg5L1PXtXCPcFpKXu3ytqvdVgBWaiGG7z0VkVi4RsJyzJIFqEU
DrEdJYVYCbrufQxalJen7zeX0WigO6MZtddo7xDQ4ejOzx9kjGlJsgGtBcEzMWhr
ZSYqTxZ8eOqoE8cQdlE5XngZaOd/apqi6QVXG6Y/dVbr0ZXIwTpF1sokj4zBSYwF
+j5TgUVBjT9mHGdxiWvPPSuvjLvo/BfqP3zDBPD36JyUkYc2YLYIeUTCKhYguO0x
pE/BVHEMa1fS32zE6SYexlyrWtFI5uIfD7mK8mocjSSaGBcHgnesFI0VzseMbXmi
nTgtMTI9C7qSWIdhohZ0oRcP7dizDbBbw3J8xJHan0leaJopfZXN6pSv9KnxXddb
iEcD527Ei0tpuaxmwALb8HN5Y8LQ7+FEVPF3E3cy+5mZTa0LQpkCc8CPkrvfxXuz
FceCgkwnZLo7RtDjtFmIbl6VVVDUJvwiI+75HU8V1HwtRcSRsimrb2+BNV6rZEP/
/siUkSdS6sbgiq4CGzwFv7DOLupKJbXaI+z3ChLlB4PYZlXX6vqqNG+goKKJkuTv
TW/QAJIXbsudr46gIlObGNdJMTPL2PGCPTNekUL8k9vDzUre7XxyRZlRDDQXpsdW
ajuc/6CvbSnjtNiH4OyrstMsQx2z0Oa6oGhtppJTDpuIh7rcFSWHH9kNW+lHx7u6
LiOvSc6MrnGJWrMnsM3u7yl/3V9RxpYOnuKAGL4Oi2nHDAqcfasRq1RMK4KqeMrR
OMVRpBATYAv9JyM1DgwT/d0fl2geU6+MNUFK8zFN1lzYLN1WkA1+H7lLnoyx1H1h
lKVvWCs2VKdv51Hs/gjlmpabnSX6HvDmyG4cmz8qkY1VPNHVs8ISTdPIzYzKXvk+
xrL8BkDelnVtBB9Ldaaj9nVh0pZha8Dmw11FhCFUzN7Jayu6P0ZvDSN3Q/Y4dPTk
qQNfxnIkrsGJCgcHY75DmYoPbg9TNZAF4pwHyaWNtRNZEBUjpAu5KWpcrFWhCl6h
/7JXQpNq0/6ZMmBQpez3tHriWqyYg9Biq90uCGPM7hipO2ZfVOydy4MWhtG3SINu
/nOxfa0W1VDlqLIVB/ZFzUhaM5mjSqFclG5iooenT2SW0/l24qHxpAmD6aifKBog
+Zqf9oekfjn/JorfjjF1jkHSSUc+XjkeRGBMtGdSxyY/FGRSTJzreR/ggaTlTwxN
73VL1RxpHLqkPe2vj5t8L4WWhZrWhP2EJELd6KNvNCcfYPlQinH0SVPKZO5Pb/yb
9qHNgHuBjmkiiX39mvNuYpH6zvv9AdZ8OknBAFgWy8NM5CKUwKk1QfHQey7bCgQj
Vkmy+bL0UrbDn85H0v9MME5nowFD/FgG6OKAR0aNtrEIrcA4w3Yhp5doMuUqOmLO
C1K592VTiJ9b7T+FzHlkhlI/UXvJdKlmyS58l9/h4uUQOFgWz9ooq6bbQNn8ATB+
0PnImrjKDDFiEfwujDdpRZuJpoaDhFSNxRXuwOzIQrscacnjph3L4cBy2LC50FYE
2lr9+5SWPVwa1l8jSG/cl+Heg4e+8HQ1D78bpQt4INUrN6f00HWEWdWuQuDUtZO9
1elFzU/PoH6+d56ri2+wOIC/Nl4EH9VsPLaJ+lddFXKA7sKYdZPFqfe6X70pjvJf
qwjQB+k9w7WwKSvBwB7ioTHlqINLgGZm2CXCJSM/K52ZNETE7QuLFsaRCKGD/w3w
pxYS9iyZEI9z+Yfi9hIDtegQkqlukwdodojJoM3uNtxL0DaF2d6A0hgoj9Z6kOle
NxbYc6Pk1jikXytStc6Sn5pIm4/QfOGFGJObDjLyordzqDAAaJb4uvikoJkaF0BY
NTatkVodd8zOt5LZ/FimvC8NsjNEgRDHVAE9BxggBsIzKeioUdviFb9l7Dn3XStM
mdkVRp2jBo0SKk6PuEKffGV9074TBqKPWEoqbjO/Lkh44supC50WMf2CXaqZQFjD
vOiDModv9w6DFQNIcfN2PS/D2AWY1bmLaHR1rHG/z6cJrMKIVsvhv8SFoSkN+EFM
famfc9z/yr5DqIa+Dtp85hWVGhIjpUC/0G+HvB934iFJldCojqUvKQl/6WPlf6hb
X7Vg1dog/paQKTM9DO63MuUw+kipvJCF11vsHBwqI/2JCPrg3AwiuETKTrqWZ/bL
K07xlXfqcR6jaGVByArlne+XDAdIqhxvI/WPlLAldNXVyVh6kFeAG0c2iaKBS8Ek
gT/O+TrSgr74vVk6RQ1kJLhj2HhjxLD1e+CI3NUelh5oh4iMXkJ9iypbBmG3iN7d
c+m1b2SNodFmLMyxxSf78hGxsWSzoLrRjYJcpYErL8NhcytehTjwqxUCB140R6Z0
7NbFtUL4d1drbP8+8Ryf4o+xklNVw2kg3Rq9CWgrjZl2f9j2cxhd7Qu0SioAHr59
RGSZ89w77TTYnXA0AWKril2PHZjDHCccBmqeTfFuCfSguNBkLY1OHDk45dyEiMDn
AHJJHCdQuJBpNXAop0VI68KZUwLSdHxUKQpU52lAutYmo8uy1VVmWJGO1uxvlMwn
UBfPjrttbGggtdlGn/HJO57Oirxg5oGpab11MnpxFN2nlbJ7G9UFxr0uhJ+BMook
WxFbWR9r8hU38Nc/Aie1lrup/tbYFtThpDEudLNGliFxObqtLy7KJNBfdJw+gC3Q
FlhY6UbTpURl8Jw87a2sYyOLQqlRXxjICGNP0lQa70Al7vPDkKNr+kihzvQ4fL+I
RrnZ4EZI/ca7dXEHfjNuFPWTGqe/cKeGtKwQfzRlo8Ju3md4RigWbFZvMMUKANuC
8o4osDairU+/78Re8bQaSIEagQYy+Au+B7y4g2oRxlDi/aPsI5VTyIti9ElwAagX
or306FqJ7SxPryft1ApOZ/j+3FFmgfFm/YXKWOa1T+DJ3LYjeIM4Dg3nXtpv70lp
OpKbINmYHG+aJ30UPxhDorg+/kNKcPwnaCQCKPTL81jhrDEhMuFWvjL3mbYFizhy
edcOOvDJwBxwJDGzHgd7jSe96d+3G/s95Gw3w7qdG5zhavuPqLGl5qz2TuHdGn++
A+A69RRnuqn9aBjFsitgn/ZyJtUInXkAK6l5HLb9bJlckG96CQPy5H3KpjgJg8Xx
U6gLHZBZpZTmEE+TJ3n/JIBCnvq/andicPQxc5dGxGcHdwRsH3Ak4xfEInuBMQlW
POeYhpLePu9YtAljt/GvQeqlgvgBtfxPuVWBrpbkkHa22pa8fgz22Lt/XZ+Geo0b
c0YJlRXJj5aJStWD4qypCmgg+D7pBHvA6HmJUpUg5qZSoAcHltpYOIOhp0aO5+f4
q0TNzRlWkNAjgJ/N13SgsQyGABHen6lQeVwAGlDyNkGq+FjtdoqAVQkvWlLbckI9
lek9273R4YSFmEbVmX+VSA0u5Tj1D16jfMYlo9x9t21TTnXYuOHetY9x7wG0r+FD
ieQS417dj+BNyBgCO2ObkLs2FI8ocNWGL3jjTXwKvljjfMX3WgLJ74cvLIcmmgc7
9lbpoRvOAD5qEjsUfKm3JD7Z9OmQiOd6yq/+hZbkHXAyD0FJDSylBx9UVW3+SoMT
czRWpEJwi84rM41O21/ZLwCqA9Th60+SS7HIgXRNtLTm05Xlw/fsWOq4v8mX86Ni
6t+R+qimc7djFPAYpLY2RC/ygqvzASB3vsjOWs5fu7RQcoPW93wrwnPcUT8IcpNM
Xih8CiGUhxkTqLnZ39tV74c7Pfn5/c9D9mFWxH6fwAgWQ7cBJuloDOvNXx+FPJGI
x/V3vOT6Z4o6kqXOjuHWW9S1PvBidBpFosbGNrxykcbkgwXSxORcgfiw3hEf98ue
qOmwM/TTZk/uK8kLLqKKc7yS5l20sWxu4Oru3vYkGTbPMLoJMjdlbnaHQenYr5yB
SE0tK5uTw4XPJ8ZFm5Llm/A/myiyh8XZdtZ3yarg0fSOAnb2idCAQfmQyhnH+VZr
9BiRNwxKekeJlufqA8d2Z0NBNnWebp0JHxLtcoS/hxXgnPnqeOtroFdxkwCvr7w6
fADCuuDiGOc0+fdlZUfmL5lqR778v9WiLlx/D37jjGH039bXVrEbXs39ei9KxfkC
bH33L43bqFyRLnBG7hPEtwqX4NV3fkHEtoV7Yngj37ybhZPtsOJUS26SSvF8PSQ8
3tAiiQTgv3ut3xAefwWK4rJ1cphZMLnZAjF5g0h33lGvncBi8YJNG1y1yJ58Kkfp
1/Pml5wnVsfVrIC+St4WTuDqp8f1IGW0dxsqdc+SNEKnkoQy/uz9d44e7yRcwUO+
L8jIKdJzmRnm/Kh5R+HENjik4vFSxwRLHfZ3MfUTUIags6fvoHcj/CIhW9KSmesp
/RJ2i2DDjuDls/98Pph5p5JQZmCJVK/epPhmirBcZU+hgpdSMDEqjQuCP5afESfg
AkZcEiVpruyUlB7sjRmZATbnyvxAddijOiKwmPdHvnPkVAKwCWjxwPJdzRVGEjIE
xJ16iooJCYNzcfjB77egPpTSkvKdIrbWJadHPlBLzFZADWCYrU6E7EbvikcINeF+
j7PruBpcknKNWmLW3dDqdamHgfPskZ7dmIBOT8iSNFTCaCOjv2p40v0VwiNpG6+t
4+zF25yQ8Xby6Nzi/q7r6FMdd+Z7CYY49mImm6VFgBcyJ+AxY1gAo+2xfzLiBy8N
iS94LJGRtJTrWkKoBQ1O5ltBG151MEeYDeaQWphbl2/IWT6+P0oVn7Wo/355W7GM
o4EI38DqguH8zEBZDZ6slCnzj92Rg1DdqZ0C47znhRRxWY5x5ZhXT+O2UrsjF9pG
7vrHzRs7OhWCpGoXWzNPfwtUxW4cxAW/vjI53eOzkikeek5Loq/0MerHPtQiy8Bl
HYyUMaTJ3mPR2E2fYdXweMbhYIFzCXo3RrhWzs2YpvmhupnfnYXoPNUhDT3SrivD
u6HLc/Ftyp6K6Q7pDjXhQ65hds419uRYWKqnPXOrLUz2S28EIGAD8yOUNtc7uEr1
a0FH1f0hlG+7GiHofrtQQt/TRUM5GZFwZydcKWIQjc06wxAKd17I4V7goIuYLzpr
CFl90CIdgAI9Mye5JLptXVcbkPrjsmNgAJU+OcWPw3auewzuqVuQAq7k12ShmZ5N
nWqlzF6y6vA71fOjImrl3YXtU5OaleLyqz3Qvep5HkM2hc/0VbJWplVCTH+lC0Tg
o/gtQd4x/yzENkXS9IUNYVa0zFOjBM4URln9QZp6Mpv2k44Zc0M7TUtJwpeJbhbB
rjVbYilsnIRZXkzNvQHNBNX7rxfP8mRdfT5rBMCjBnK/LfjsZfYJYAbkq07YaxZT
HQfCPNbup3lCdFeYmU4YJUWuuueiOqL/fZHDVYBYjwYyh3RmMjQwVU1o0pLuB+sb
4dtIGW9AN8IiYO5Rv3/CA9m3wlycSgpG9DaZgLb3dhfhpM2pCd+yWUdFeFwGhDHG
ppcj9BGTj2rFLaop3aQuaNHTWGRUGdrRbajMar+F1ji8lC701PWVLz/nt1QTxtdd
Yryz14bina0esD0JYLHgbiGs4UhKy9iLHQ8IEbx+uYUz8+lDQ1ND1p8MIGT+hr6z
GZsaomxkp+m94thc6DgvWwtHojTp41LLfI3JiPPcH6Oidrdwb1BIiWEvq4FKsunH
F5DjH9iwLEr8Dw7U0Mpnf6SYrS9izPlygblOjfvZE8ngRmNZCKEXTVLqLAxChQuO
APcaG1EcgAJA5XnSYcR0LNCgH0OQTXfpJ//pAy9Eh1Gz30PWVg53y3NVCJlcQuP3
PvrXldGdwC6WLxUDB2FHBBtXJJBZeIaSmjPDdN9nMUZDULGMYet1ieGXxgj0/38i
VEMhumdiDUgt6NBmuRVt/QiPfQwh8RdSf6xbZxiLqxFKmYkJZ81tO83NFxvVoUY1
IKTAiI5mU+Y2PqFayUK6AuBVizeR97E5rW0pC+fPAzBlOnOPHWT0yCR+mKmXTUYp
xavoBQleE6IniGOKS/b9umn0i3T3HYrwD+MlUTKmFG62eFsApl/f9nP6jvnfAPIx
ORBL9Fb7ZNJb0MFpFDR2dUawD9dqtfkIPZ4Bv7BE5G6aDjuDqTuD85YmcsDn36EW
NLo8KW6dUSu18k4jY9jfF34BqDjW+SPTtCLzGy4O6OvjL6+C2hAYydC+rA8Eur8D
jXTY5PI4/AV8jXVFWqdGi+SxrTTAcfWGaouEyH/fal8rTZdoOEYEid7cYkd56tnd
EPleMzoi8BBoeenG1cDbGYK4YFWiXR9yyJGYmyjylixyHt8ceRp2Bl3D1Vqoc3wp
JvJIDNq8gsoKnuidNxxeno/3oHdHpWyH0lNaxbgK8xJ0J/xjP6d9KxzHEZqtP0qS
C+SYrHWQJcW1K/GBUtnhjQUlcv7M7mJ45YecBdYWtA8EjWj2Tj2FoyjyWRCqGto7
b4xQ61AHgN4bKY4ADxCVAiB9UhDEPhygyNk6UtNG9w1ooXTNyNEkAVjKXBjJqfK/
WqYrh9Po21UJ+BV1jOMtJ0xiS9R3ES90Mlpnnk3xNakl0npwCsd8ottLjeZr22TL
iUlVR+x822M6rU1++mIzNgzGQiUKpGlfa0lMkpRG22+IzL2QgfOg0k7rAM35F/EV
3BxslUrijtR2pL7tEhmneo4OU5IfMFTLExe2XHEay7010ztsJa8D4KGo46KCvdzb
Za+t6ooR/vOwLZCZckChQjhKMMth076ANn51NvnGioLxcyQEUPwzWFKqeZgBFDw7
kFF5vQq8vjYbpQBtX9Z2J4aAMtPCpFVYxFMPhPnQUR957dBddA56x4zk57Pl48Li
L5p4/V/v2Afb3IXLv4P+Wx0AJJ2183UuWIqIsQGPTJOqsxM6GneQzF/NuIzTh0Dw
goxWyySBZBnioXmkYWb19fuy4Di7Gyhlka++JFlL+QoRJKBde/OVSEpeuEsbEKli
1VvUMG7BeiqLcDpJF/BnWrF8mJY9StfrBzFYNJtLtQJe9Aplgb8tEJ6zsOJBbCmT
tB2g0NjgE4NxAflMffLlGp6CM3ba5mo6U7DzRaXaIQfCzwHIodSTaNvmNz4+IqSn
HVM6VrDhDSq5+tMxwVIdfsGiCdMyPApkMuE70ZmfYFBOKMYdsP6XEiwt5RV7C5r5
iNXXrG8VousstCVpPIrenpBzuYSsRXzOKRhM2uhWLjprq0jA5f4i3O5XX6EJ7gpV
nThB4XKbbl2117mHN6iwr4FCo+7Dlsmxp0f8wWTJu2Pncvf4sT9DwAEJSSiuG8LQ
RCLjQpEC+xTfqxScWNhYWYPUjCVg/wKdegCbVsNCL5pW98/48lAR9r1u9XtFaSSV
MU3XYAIa2JOAk1DslOeoOnWBOd4qyoOCfEM2dSIH5te8LsVs7Bwda5TcncFMtkhq
a35rtxCOnKjJJjqvUcWCq8sz1kk9wVm42ysQIDVa/g9qvWxBcoNBW4gyJ+E8KutQ
2EzgwZCj2uCawLVytDMJqOIV/81/rqjpoCh/lG/cxGu8dZ1E97nIdbxXEjm0BTLT
qKAyoTQJXZpvzGTFavY7C3IsNTTBEzERE1Rgx7Jyr7gzfkXRdVt13Zs2vr9YWyqy
AOXs0u3xCX/zCJlN+kT64t/9C76XWf6P4AP23RQQpB3UPXV0QbL2mIk8vWAp3+KT
lrLUmCbkxNXTUoD17urE4GXgDlKK0fBO2I3/sWfpWI3ss8sXea4M3WWU35cStWSb
k5Z+L3ugDGzfilg9a1fwunjyyVY4yNxmPdKovSPs9LE4Qn/s+x00WUFd29k/2eqv
nx66bJCgpW2DFkET0joOd5Ccg8usFVxFj7U5s89bK4P+BdSurPlBIb1aYP+dgKoh
m8Ogd8D50SrM1ZT0zscsy9hLHajgD6FnfoUoXNRXEP0ulkQRFhGMpttUsUKUrzwI
bZv+xanR0QogNlXMJ8KAFLVZdVTioRNc3viiMrmhHhBDY/fnDhUHFi8qsJuM715V
tFPgC9rgkVY9yzw+VH7zny00cfF7b8o+X9c08mfv4dyc0JY+0pARclWOzCzejo1u
mVHaLqoCy0PfW/9v4i3d2hxRM2NaSezkgbsc0OP9rDKLZ7H+0l4CkdVkt9+vwimU
L6IMJURNSDvqprt3Zap7S0xXpNYE3LJAN/oei/omSYMZD3HCked/rO0GiMobujaF
NnHlaSyu9GjrMOK33B8zHL/Z5Vsz88XYmbw9hNsFsNYLmHUAfS6Y+OkQQCg42wgj
HPJI66eSjEZcTUxcvsKK+wYYu2EU099J1SThpO/KdOjCJ2O7F7pBVlgKhBkrfAaY
/H/541SWZ6bgjC5XDTzslmOfiAtwzB7JjoHiX5Tkvnxz5jmQ6zOD4HrMrUQq1869
CGho5zgaELiMkvtiRX40YECW6zFpzXPGF0fwzHr/ZBzl2xePF7lc8kgxu5Mf/Li6
Gkw6NKIzc1ZnCPDLnaZDrSGtb/2/QlHC1wILuI84HhAGfR9YIZ/whZkPlllEkvd2
HN2NpGebR0+LsgDmU9mpWN60rDk0oE42UOXXQiLg9g5XX45cQUiGeAlx1YvnQhrN
uqr/RIK1IqdGasmHo04in9bqVMs1mONVTFM++Q++r1n/twFBk4OL3zEW7d0+ZZ8G
Z5TC24drByMsCiqfcBO0PP2zKzVogIy8NgGQ9HRjdJpczuXHnKpfOG6FyeusXcft
dPCL9oZhwMwDpTHioafhPxBSpIHWAJa2ncgsZjFVo18EdTcbOlx9Ui3KYa5nvr0t
0cWohIrJbryI0ELktRgqeM0kSqXnHBhQnHO/lx6R03uJM8DfZueH+bBg7y8mMvTk
jzFOkuAZy55b1j5/9Fo1u45XAuzg7s4ljisfYUILbI0rUKsG39nz7OIqWszItclu
shLEONN5IoHiK/8CjNlf2mGowDncGmTTkYVNnTL8WAYFKHAfhE1YSrDRHsLs/rhH
PUA7B344GPlL6xm2LqEA2NOu7H4nkEfq7pzFkBxalouA5FlL5XM1cP6+WmoqbBCS
Q8XZ6OCK1GK5qOiKs46HfgR+Wjgh83eNh0QcITQAytO3Rh9Kr1X53km4MuvVH965
0idJQLHiWvAjENbzz4gSDogN7541mLXam3JZ2aIG68zJz7zT15ZrnDqb3qgwcW/e
ToiF9R1j2k9LhXqHKyeJmVAHDpwQmPw8sVCnP0xHhXCovncVxQy9ri0iGOAuzZXa
X2wjAU5RnfgBAwrJg8N4DppgTskGzcacRSl9cjkAQfDW5nZned5KFvoDk4E6a0d+
KDPe/4n0TQoktXI0buT/0J+c5x8gAnGUIy5B6A0wvoFCdtVZkRzRgCseFd0oP+pb
4rL2AdP0Bwb0TfKKxqzH7Wcslx1MJ/HoM5DnfsxzMU5jeV/SaPiTqDp1p0UEQWkl
Fz17x+c5Svq21n2hUdr/LaFKK/oIt8AuIojGgx4eT0HYFwUFRHZ2tYwt4elgKMNI
4L6fw+0zu5y5EberXXDya/SQmeSlPYFzs23n9r+I09ej3TnE5QDkaGnagb8txVWs
UnF8h4TxfF5+9btRFbKTKfY9R2oTKAxPNJYUrMfE0st2mPka/nKh47zqc3nLLdTg
HckCtxMga6WoN3HwVqi6l+D+Z/ZIkLWRQ+3wC89C9zUpQ1+mZJJs9t9adRRCIK0c
S8967LLWwDug1hhMDZ/cPM9U/GRQ3xilgDAo8EH94kyH4gGXcJm5MyfCgf02m7KR
Ls9HAV2PJ/FaghA7LN5v3DSSVjVyD1wChMMpYKYvrGVCNaELnVGiQ3FdczkaBLL3
XwrCRWsLvSvzcsHZaQe5JmMyDaitEhXRr4NV8/5eTGIsHPn381nLSinPwiFQ5vCr
y6tRgptPNoz9gN/6twXKKc+vttaS8VYqVsl5tr7y6P/AlrvTaTL9DLVtCXh78U6Z
Mwt3H3RjL/lFqQllmhf6wcRdzfDpc6ZRvBYUh9W2WptehD6ATW+yUcJH/xvBSvXq
WGS7G9okKiCWY9UvycqIHFWD6gm6j8N3teN8qkzzvD5wMFoZ8QYV6iZ8O/UYWMht
l2m97jKICRIpT8uin8jYjbjJ9hOwWzM+nwfGQrDTbarvJaWPQicLDOARKZPiMJdY
SW1K5cbWKQw+GXeDhs0g1vOZs79CsOQsBA8JiOsOAC+CVV54079GipXHUxJMfh/x
A1pEeMJivbcCg3dDD0UXfazD/N0aHXQrTJ3s2ZG7uTcfqoyQobSGQfQUTg+1Ng+Q
TRIb/PhUWspULVEPg00pyEohrjTFWpyNZeQAI5PFOkGLz1b4ENPHVfzPCjMUlTuS
KixxhFZkOpEnnhaVlzasTW47peTN68svYtO2qurZhsFYuwNeJRF73Pvr7kGmhIGl
wLo+bOAUeZbHpHt9VZ/Ui/VzZvslV5z0pYL/nbvNR7FD9LiBAYx3mRyc19jRuwZT
ywNC8+z3kxvMae8b6ywOWkuEl9awubha7VxSYuNdzQ6GNyd1G8oFZcLjOjDLZuKb
u9Y39FhGrMAkxBl0SXzKmchF5CTme2ssih8eg1uC1/3o5Twlwiu2cFuWVnqwKuQr
IYDoiElHAdoKvZBQVyF1ORXZWeYUs+111jmb2cRK704KVXeTjohPStonLITfo+B0
BuE3FhGtnIhd/D2a00F7t82lezveOvFKy4OdGZcrsvlcXeUB5/TL9qeHIc2N+QJo
SHQ/zNWinU4aS5dMXtjVqnALkv1cgf/qMiLUxNznX1oxhbIf+z5rk0/R2o/mLJnb
tSSyG13hMjhYs727UaRArpikpXkRo8r76mmaRCmVpjAtacrjXP0ZdNzEAFsFVw9x
pJgcgRipMgS1BM4ZEsIV/QrQS8lJ11bnmmFm78qVTlRS0i8Sau++24W/+sXbFdU/
ZxnB5UOeRJOe666IINQI8u1FaH8v5Cu0DwQ6daZ71d7YbCa30wI9UXnQt3xvwNU3
ZY6Ts+ctcvqPeCfmHJ3M5UL/lvFED76SvEPJIVCwujL+ZoymFfAT0tYOhcTabdUS
cyG+8s2iL28Cph0Y6zSEHjM4qGOWu0cu0J6O22yAeBwpPrQECGIb2ctK5joKZ0o4
QDSDg3IyxFuz5J6Li0CZY31hvASvtPcHSqWsYfOCm2umueYclJYGBqO9Mb8Pak1Z
GVwfRyD6RxS5HXkJfm/eJjEL/5VDRjXYnBgemHNkbmtrnuprk7g8Z8iEZ6ZNdqIy
EEG6KjWCU7StoXHAxscsFJsi+TeztsIAOiuTIlauMycaitFtN67gBr/hEnARAa8H
nYg9U2Us8RcvBL7TzcUTx60+EaurdFohn389aQrwIDFOgxRX0pSV4VUZGhOaSC0k
1yWmX3ZEcLjZmXcZr8cAEvZ5KPWwkuoTWssb69HgT8j4YXYwcVbeL/9Rf95PA12L
VlEQahKRsFibsqQ3u29FayRP6X/YxYRZE9SBK2joqW7hCfcYcyUuBvM6+MYEnK9L
HuuTc8drz9EjrrZZAd5Jc504chkfx7vKZuQYJs3qH4gE+/sK0jEy+/hQ9OdIZVmQ
knEm7F4IIpVSECXFnIVM4wLICLX2WadJ38/MitnDU8yZkk+QwFQszu4KMFOHLHTG
3gllczgQqhkvMsCa6m3CQhCXCCqk6xd10KuVhYSt5c6Bv40jk/Z4FG+2qN7lak54
hsCj0JEz4/3xC0GnFcF1HY3gpLcDpqAG2zjaB5a/Spred0PEeG2Dn4XlLCUTMf/+
l40DWunW8bS0E2QJWTY/VB3S87YTqqZ4x9KgTaBhY7enfvIvD+brt/KX5Dz+hX6G
yzOLSIfFLoCCPlgPVClJgEXqt5ZtTyRqE6oJFMHJsptO+QEWgpCV1mji7Hilrpft
Lyu0qbEw0QnF/HTItQ6CD/TynxnnFQh9REqPsJgm4TU/1Yobs8kovx1Y6LqdYI0f
vd3ziAQsIROnDgqw6kXevfFYZue68TwdNa7Q2XjcdHTGVbuvMVTV2PokSRkzwltr
EY4274TAqSuzzLruLUEMDaLkNeKK8VD5rgfS/9T9bjMdD5iMAHCwKHFzzcmYzlM6
0bUsIPDamxhZG/sLRLzZ4a7tRkEseEE/G8T/8y3/msmry/qWFQt06MgfUxiPy4+L
u3u1ub2gNpoHFjsEw4YYklXywqiFWt9WIkQcVDb7ibzaS1QJnj5FXrW5DA1rmYl7
mpaEid12qVyBsUciKwR4I30lXDdE+jdDrjAxLdjmvfgHI9YHTvpjkuxQTbh2IKJp
HuESWp9TZKI/LrTvBSEKh8RCatEXuuNiK8l6TSXP/+cF4ho6GdyIr0Aqm+/smoFg
qnRlwCndQya4ZTAH4uwjmg+oWbwPtG8d6Zexw3gUkbxbK7JUbpmjg8FUsheOcAmx
//lCXBEAZMuC4q/D1KuJtWVSEY1duQGP1VtfqPiko9GE/wiMhubuB1QfVOOnTrO7
k7B3DX8PvBFX2yxLEBI58AejNULmoGUnDte0XfkOWdHKOPtqB/FHQmdWrH1/Bkyy
7NVTm8W9zOnJUOzNX6ScdOhmROPm+2Nt2iMpTq5o+HjWwnPQdycyQIKV6PcCWwJ2
ZmbWHFw48BrI+wYz6/EFGqZpo82A+y9G+MG7QL4UMB+LMvvi6bwnW+DvU7iacFq0
Gm0174Gka3AKuvoVMaYzMi1XQeWgiwTvfDZXPBCdxe951bXyJZwgFUvnK9cPfrl9
UXI0MJkG8WbpJIBt57MZBNcvsXIWAZOxVjk8RkUVV9BOyOh2103pTwRjEEbsJSNI
FImAsasMJmVPlREDiOSPgslcLO63QfkQyWx+DZ96kyjIDEk2Z/AXNTv4gXTlInTr
dz/8IZObAiaHLTH4Q5o5naAoxOW0pboiz5K8wWXiXQOoZR5FRZ+kxk8cpnlV7TDu
RsyiaKN8B1IuQaSesM1iin7S+dhCzuXFIlDeQexuH+k9e1gOm+hMOHqHZpmT+g1o
7fjFW+UGj3PcMalrHBoPsfpHRyZOWNvDDTZLlBYDTKElXYOZmLxbBYdzPyZ9ku7G
UcKEl6PlOC/0AvapBCND6T4iG+fPXQ1mXqI0/q+bY8NZkTkAasCNKqQm4mPqtgRr
dpg9K0YOiIUtnkbV6foD7PPg0fuq+yw7an5NJlnm6VRRuihRn2MysiU/4AgdNDfB
npV3VnNDENVjfzC4hXXj87LAKeUljwjcpvJsnAOnhR3rGbmGAys5Eiz5VWgtaXM4
XcuiX9ZchTp+sQgvT58lIVlTcnHA8/THSbAlDhxrj656WPF1vgoGYQPWq0nmgORc
0wsRj+PBaBuhKaVELKQiarVpnJiGyRHal17t4K6yVm5UgbFNwwqBLijVl514NBwt
eAWCxN+sOgXcab6cbSlj+04Ffvwv+MR/vz2OgeFl1el6FYqsLOHoKs4djGcISOGx
aunyPW8fjKxIdTyZ7KBA19bwsKkndGRCEVeAkaay3jA+pYM5rlLdNjH5HjSWeXSG
tAGkuMEuZNcwVTaBJcNa+LB+LsV/T0IEF319JHhfz9FOQMsMafR37K+vEb7q1rz2
70hSDCNgIay1AAlVG7xMuWekk59Lup9K/cVaF5VaMxHZ/j8CBeSsRioWSbU5T0Ti
qITwxJ+T9AQjvJP0ml+Km1b4vIL/KPZXQ6tAE2aD28KItqITcw7mG+1VQkOVTluz
nbmGkZMH4J0ZrCy9Me8ItpTJ63ag5W3K4j1182oTzRZp6KNBUVsUWzVlhDDdiyNL
HlUZotlYD9mGK6xZnvIAOdliq1IZl3Y9k+hPPweGcjlZpn+Lz7LoFes3H+TCt329
1+hkA0xC0txxTpidK81gjC3vio8lCpZqsUu70/5IcMZu6xCJlBNWDuPPRESJp7Fv
wEfksQnfqBp7ApSbd9B8aEpMXIlLyJa3pm1Ocwnczeb+1FuGTZpv95SwOZs4Jcli
jlf8PiB5N1gmAr/FyupeBfQHrZr1k4kdUaJqTL/BUKRb+Gya/799xDdju7CRI/t3
cZn8/IgQuzEAZYhrwrCsMV/JF7fTcdpr7hk1oyFUa7YS+mEPTh+0HrQ17l82qzVN
TP8hbP2y3UZQ9ZqBEOWOvI/kpX8x44JFJ/TEbvTvZrZE3loEXa/Jhe2YpFjJL3rC
iDHVE9FfY2cxEfGAm4PQ9q+Ob8zhiYhq4+NmN27/Fgo53txrzhpdEI6kDKSZfLlj
voqBuw8ByJfj4/F4tPtgh+Rx6MhsdhpFff6bO/G4v5CvAF2WVlku9/s8Stpet5JM
BohuIdHnPDTJLV5cn6X2fw+A68V6X+VsMXKY0UAgvLlCj/AwS4sq4Go0rfUE9jYb
UwAq4hQTrFlqd3NWPD5yOveIm+mOqr0thjFERFgVE28wYm54OKP29Fdq1zO3b0rG
Ln4bY7J9XrgA2BfawCHtgLg+Wtz2pbzrxX0jh+HXJvyXlQh7K0Ju8Fx9Uhbt/GvK
ef3x0LmYKbBPthCwE+NdbUcCgJygeQaz+ojDoAUccPHnpk38CnWyOZEsNKechf3d
AuqwaR+vvmpyu2ZlZxNiwd30BT2hfgWqKPL2nbcuKpYI+yag0LTn6w5XHUvPp8vt
6LXTy3mUHU6hGmxbixbkzpHx8RXrUN5kMoQNriq3YXJUo0kQ4uwl7tqJugnm7uXn
/WDEodxM7crBzz84bjvdtgm+rs+NINHfXuCCXWwEQhLpNwfm624oFc9zk29dtqsj
3Y+zQ86K+d/bmcsnzXhJN3HXACr8tMElfNMXQ5zHKeH0uYoEhlITwHLqVWNyavU0
94fo2e2Gv3BG3ZNtspIMy1hR+JH99v0JjaDDbs6Ovjh5MRn5uU8nJJ79PtI4TCke
q6aCGf+OyAArExh74teiHmqoNye0C6f+fk2WpO2CRWcPqJ9BAB3iMUA+/ZVkVoQt
xDoaSQXUNSrOawuFxnCB0S3mznjZ0OxAhAbP+N2HJHjdLy6l1Q7QUFPf1WOyAEwE
/dHdQXDqodAYkMQknVuRQzCV5AsQymOWSmbazKRhmv2UoAVoRKw1CAQDTJLLgzII
gkfGYmHARpwXk7RWOOPoV5r6l3KvYyxjuE7myB0M5cvKhvS8H6cGPv1zxxC7K/p9
q4bQKmecAC4/zZflhbXaBddekY2u4YkGJEEl182Z7fl7rqYwPL/jP55lrKuwfJmt
b7G/6VlJ/tXukbajwTQhLHpnQ/SniBsbg8kWzi3LrFIIgxQOYWN0ro3CzkkERnLf
JzKp7uBYGkjKlBjj1wA3q/I3X1ZCALpM2getVpc3zfV7xbPXZDLvb2e0I7ErCN6f
+GFDHua6S5PtQMNSGf+wxQWX2+mhfLnY6sjfHztGUjRJwhv2BT4LSlZ5AV80s3t7
SEhwhWE35Wm3mLSzlH7MTGKlz63HFLuyoXBsGZs4tAACC5rhodCj4Vw32eLDQqDf
n5tlGtN0nemTGOhWlSTHMdzwysLnfghKFl3F7brgDRIMhGM2iiJ6Or07xlh7Mgew
ImDfBcV7TwN3yXqvPxfn55lSrNBaNb+HwtICsL2/zPx+/vxTCZ0ROC0M3oT1Jmvy
daCjh4r3arwFWw7eHM/zRHEgmpJnEDPDhMGQfUWYw9qrZfb2z8MHSUuDVt6I68+2
0o31EUrZNjbbJNfqWlgXYZZct39d3mYZHDRbNwriiwMMYHUaW7czflXDFo5HEnI8
SgBb+HzS3xE6iV964ZzEE/YT9F91KAVLJngV3kT3Q2iaXnWRP9qpOIlDX8JeSIdU
gjEJ0LAhPba/fLjceH55x9p9hh4lfqxf+raMUeU9zv4Tf4LAK/cwUkHUo8Ev2PVo
HUEyZz8oichKLZuupgYR/MhAag6D+UHV0dd2LdLilYMSAhryjrGN2/SrlEHyxWOv
9quT+AM8PoxYkMh4yFA+zTxehI+V/QgpDmIvEGrhkfQp7ozrXAm4bu+oKZCPaVkE
38nYn3YLTPG+fG/tqRi14OrKRRDDTHA84jNEZok3ujarov+/+ha7C+a3EAzFul68
4NEOIAeuPjd9bphzxJtU7s4MO71Ig96Vz5HwEbH+b6UsRQ8mkT1OjwFPTel4uE4V
0wPqwNvkFrespx3iafvfttu2lUs9Zefu9blBio41ux5OWOH9mjT688/E24ussrWa
DPLHxCJ8twJzEQ4r+REv88DSR3KByw9qu+t7bhR2nQoCtNRdd5lpk44q/k15l/QW
/i05kesiISFIhdHo6jVE4yCs28zrcwCFEaLERDbzF4gqjCn554CLQibKHlzTbZir
MMXq2NXKB3noIcK3xicLWKmLkawAuq1wvH3ie7x6FuYatlLxF84wau1UKp9VJeE0
JFDnYcyC1/4IBK/VT2h7L8MsI6TAzc6kugYJ9hju5NUGTx+SWZ0YtCzIjkDqjV2N
ShXFQLNIY8aKvCYTYhNs9qIJw2K+IAkmbi2j0FkMQgWw3C7TQbduPmBy2+6h2RlD
QqX/U7YZ3LaW9rb0h2PcEf/RQ9l5g/3WMK1VzMCswX4NMmOmLyVd5EyE4dL/aUPB
8zh8CsUzfjYAZUgwSC6QYoMacdH/4e92hxNSUPCGn43L7bJeXV5kzZt/x7S5XRUG
cDngGauOyxL5ZkX7QLQV7e+Xj3vUlmzj/B+tHUhaJKa8hCKVPxjrIDdRmm6z5dvx
RD1KOLuZ4FcZG0ERK5szX+hccwtJxOz/NOOGF3KnF6sYlcWTwP2QOclkznZaQdf5
Nr09Ak4+eiWf9y1ZA8ORvnvVnA7B0nZfGkjQURBbLVo92sdQBTeoyp8pX7eCk2uf
Nw4+0YtkA1tCVgFOysq08G+drtQSBafO9RGu+XievgTXi6HNLwhGZFL+0oYwW9SJ
lyWAyzxG4KPZxrLP9jLMm5JaTm7qTTpwK7jcRAW4YjpkFxzmg38gAz2/+YnLGXqA
o/S+68/QxwEkQmkIViOsZCZ5jBEyF1ke2gW5+S3XBit4t351mGhmeRVnj7ty/Ny+
HbJh35HvOSyrlOse4MDnd04TavbfcQXkQeZupdDJ1CLfi10mMQhR4Fj06ExTLVxY
EgbZkSSUK2n3QqBgNs/YNBp2U1YmCC3g9PQ63I5yln6tKtXIoqA8AijUeT0lnlk7
RNbDPibRZfeiyZ3R+m43fbLdU1ePqqDwj9p1T2lF/xliJWSLcv5+bLtq8nUTQXwW
oYdNx0tGFwC9vZniUVrizaYCi8lkjlT3L7l3lO1SwURKCqehsgzfj46ulL80fYzT
tkFZM736BukqaAHrSKtpOzIfVBVebGLk76pdaVBynaoibKtREWqlCIsTZAVRe6nz
dHGIvLTM3DMytQ+BQ288k4wwPoRtscfqD2u1Yn8N10V7fy8tne8prkzq7tekrUoG
evRabmsAIE6vpyEcrzXWx/5lY94aoTVZ0qWghzxq5Q3cx/csFBX8fKdnCtFXSZ7M
7MpNle9C04La5gDrBw3zsy+K8zH5KL/WcX/WViq3BzVQ/Sv5xTJqmWLmOneCRjYY
PlDTKI4HMxn0hF7Exm5xcctFXMrVZyzuEatsfD671EA3LyykKpKjPcDt2UQVtING
KaOIXdVhgpxYW+ZUfH7ccCZvvIw/DhnqaAdJI/2+XXyuE7rZAmNkxsnrbyLPIJyR
E3FYRgfuW0/gbPY7b5O79KM7Q4Uhw1Eo7xNL67D6dSlFF/r8Zu5lWCXlqNKkKWZw
/JM9Jt5T8DHNGJeFPlgoLzix+0JmV02/fsnA64UAS83bBPXewFUG1LWIA1zBaVjl
L7h+dXeJ+px1Dv3ZRP4vT0TEr+MzKwsuA9cVkd0S1NTObOcjdP5e+laZTSq9LRmT
5O40zvT7/HOB85/iYyvE4gZnsk5QI/7HvKn3SCkzKuQlQGITUNXKLEuDx3r+YaOs
urn4IMzxizfcRqMmKj+K37XoXIq2+7za0UJnQIWhQWCxBoJXHnQbU1Yrbh7cNpfV
25zt2oWlnzH9lwXeAefX4AF2ccnfY5pL/2Lmd8LsE2M0GWuhfcBdpOzm7u5yRApP
ejsaZpw3TurALE0QfsW+M+/CXKQ0Y2CwNEjuX6HfJ525AsaUj9xlA+GHFf3Uzy3w
ZwBR1nklSM/O7R5KDNGH5Vvz/u9CGaw2fQ9FvZbxWUjhvO7sBnRhqqDlmBNhHTgF
6F/BilhMiev36W02Kwka3JF48SI37fOsConUqe1bI0bJ0kULPrYE0/r4WtztTN0X
XXoqQXdGWMuK3rYemk6bmHDNcyrVRdyZZKwi9kWtJlL9dpjiJn2x6dXQaX2AIHBh
LBCnFPV9T0Aoprxai1V3Ah0wm6tmZ88Udn3Du7bk+/pJBbk0cyQTWhPWg0juiURG
trDe5O6RNP3Dwgf76c4aW9UfbnjrUjfeYjHfAx0Yh0m/VmrPxyhT6GGGKaRHiS4G
FecUtOk2UzuC5DVXiO5tnXC4qOUzBcYUS3F3WA8O32pc3X7MhQR8TiYihJSMnlx0
EUyyWs2T9rdmeCQW/YUnR2k3PGc2CGn63hZwHN2eifEEQNhOY313rwtAObmiXp4i
q/biz2MV788ID4Bljt8+hrLMpc6lP5H3YVMLEnw3C6PkgNfMIJ7Q2D3oRegZKxg7
RQJmiwzQBGyPnnb9GSzP+6Y5g1vt+cCr4ZV0gi+qdnSWKQWsbCDMkGldzKjuHnQL
lNLNgdbykLFmXM7khArelYObwnLPfVxaxNNKzZMnr/O/cs/GGvTby8vnUgvGnOed
L8zJYmvXzXwjcB5XCGUBHB9373LCQkL21IDAMqeRcodFY0aqYuB6FNjO2RpPC4Yw
S/FhwrzAjUDBTgE4LuyQVGlZg4crq/F2gG+d8ApRntIyMBDj1D2g8T3Z/cN+UsXP
fumFHxezuBfQ13F3ZLE9Ls1NmyZNmgh3q4wvv/3BKv2bPHA/CbFqmSOXq/YyAJjC
UWn60/Vqfki25t56qK2kS0Hvr1Dmf1KCyF5kJR7iJu7AUzvsYfj88wf8IwNPGmyz
qfkydNv6q67hKFU/+7ssBUSurh+S5X3VsqqSgESxxOJrlZs2iok+hah1yLd4yxpB
0OXjzTaERrYOKUtmz2hIERFDIMNODHRHDJQYqtigxhQ2si2Vd5uo+1GQQcbkyS5g
lCcKXPIyxFpgxWX1cRaNLPEUR5bTPBkDDpV6aN3wj1wad/Fzfqse7V2/BVC+kuKV
25bAjdxPnWHV1BoCiWzQAMRI57Vs/L3x4wkGZwMsGU5YKvdBqTTIlWbw5qWOnE9X
SX9avrMNU/zLJ0CRo82qJlkeuoeJB9bGii8NvGAY88f+i/2bSef/JrjTCDh0b+aE
RzgSTVasQrCER/ZMta8aVPiQj/uPGd/8q6NdEtZggCBOwKv422lBBBAN8osELuOu
VYhezWtxVSqSizYenIfGYszYkX/tpQjgIXHH9oTb+dIbG2XNdqw7iGQEIgo7CCsb
N7llnB4xJPNXRWDu7gy6ZtUqDIVnezUXJ9It7KCahCljJXFhuAGyqgZEuBREc91A
WBwnr1Sw1x+lXIbT8q8bHprNJdT+08Jrgf5gWzsEwzBdTas8i1WrukmhXyAbfYNH
j+E7Bf9YxQVLhI28NTHeWH/FUjUBNxWFa18kr4MZ5KgDvgy9ARpkzLEt5Qx9ZpcK
zTQ94rCTEyQPEV2cGEJ/+J1ycW9eS5W5rV85IWH3bDLPBEAUF6ujiCc8nIGlQt7z
M2Fxoy7PPiZvef3aBADV+IEBt1DuOZyPQQS15WJLfmVgKjUMD7VGwygbGolEJ3h+
qq19pnlMs37j7zqDzmkthqP5pZ65hy/53Dq+LJmfoGEBE8zEjCwAe98dXvC9Diou
4PKZTKbD5IzgMYOSOouJbphudeQg/Kp6JCG6x9pJ5eU19a8Y28Kx3Pf8DoDrePC8
Vy0wowrByeqMtlTdo7SKdj3/1aFsacblCOv8QU9vUnH9bLyUmMp9t/fOX8yIRCrG
vvXSMZogjd5JmGj9OeEPpGeEWwBAEtm3DqS1oZRxzxRmsulDBhkGoGdv58oVS8R+
IlpzrtnAnEKaWzX5b9wXCo/pMA4zTK1yQJVo0+p9TmKUVITNCw4sl2MLX3z2MFTC
emznrru8dAoAaMiHuzgiYXhy+K86eFrgn4bWUAgNlwmHYpfYwK7mOeB2JWOxsIlc
uYFt75ppdkb1e30PwW/iTKjC6eCy/Sq6A+6Gw8495cOMMk4Ch7Gn12PscbCs2xys
+O3zpgsxqqKtqmL6GZ2YkA4mUo46+McF5VQQMbcj1QNpI1Za44/GehVCMUVg5Hif
tAZA2MOeJIrKtdVseymWElXn+fpzEztyYsP196fbRpGc7DUCUXvssFvK887Kit9L
A1ulZElhvSJyjGBaY5fJAWjc6dedaR/9+oTOcoExHdHPKUxZbDjIs0Hsj/E9UvBG
TRXQ07/TqCQb8n3ERBISBzuBAftRw4vhYwKTSRqkFtz2sFa3RpbQrEKIPi61KUDf
sjVuchD9c1E+rUGV9sx9Z5Dy0uOXVmJCi+xjtExhAa+wg2QqmmIKSxKdxBkXasl5
3I9vQrKgWTDGZWweWfdjElFtBOmkX/kbfRQfEC9YutcMddf4uSc7tTcMJ7NJUbxm
HteGM7mWawljUiiR3Ezoo2L+t16goSZr38vVZxJ4GG4iwIkuYbk63WJN349iDLAf
wP6Wz6ELraLAK5TLsm6BBLDNA6nXrJchOYARixhinjSdw5B1Ixyj6b1A5bJNqXJH
tzhPg1pNzr/ZM9cNuB1fZDKFbZ6pLUuFP7Qvw3qYni0r9l5mGZlIc3kEY/38g21H
Z67km2VYkzbDvnjV5LXUk1tS/lvBTFMQltHLU0PDWv++Hwd/R1RjCDyHtT9h7kPv
GR2YsGhxTCwKgRPtMy2XXBoGtBRgzC8ZgBddKOLjcj3e0jJkMqQ46MawIS5sIbln
zRjkGu8/imcRWNbZKvbtHxPwWo1roViwGRfbRqn9asd8Kwmju0TDTCFGFQ/JWuBr
SQo/x0SI7xYT7y5Rmy9lkwbPipauQuk6XfI4ChzrKslW66PJEk78trNVZO9e38Bn
DD3b6FzWHPFagdkUETEkqiVQjpvFSEBsGqZsBdtW74YCZ5fcnTMBP5IEA9eDPVy9
WCFFmeIBcBG8PF1kF8oIl2G12wOfXaDLzDatD1vMv+pHpEkWW5eDxHVWXZ5ZT3bJ
SoL9qE4P48CHz+uhKpf/4RrFYUkPQ4SAopQvuiJ8L57Ce6o6E0y8dfs71HY/rdjs
lw7zyPw3vqmSzuDK3ui1PPdvWpCQw5fYhJ7CTZcW4a0PTCRLq1JdlYVzfhnRHuDz
gHHZTU/twKDBONJbAHlwzKhiTvWxhU8YirVNtV1NJFeT7XGCi7RK6q1Gm2OmK618
ZRDn7jKg4Un2CdbGhmT32m0xBrs/XtHj1Zwd+PvssKKB47lB4oK5XGbT8iv4v9V6
3noXZ/jQ43o5AvJ78ZGuiNew3ve5v/AOksM02jmZ4w/npkqwllW+8ZeAcPwzBOQD
otjOx4e3cfPXL3qyIBviX1yRWv/jROlw7wdDclJ5Md8XD8PLD6cTD1OJt8hs0zdg
Uskmx43d/E/tb26+GsKD03RmlsV2SHHPVebw9q5KrhzaQg62BaOIAgx8UVOBwjIe
HBobVRS4fXn2DfO9kfl62PPk0pC7ASLxA/pUpKfZ1DPqst/DCzFexCkA10CWwcZh
6mN0efdAT3iur2KeYekLqMLN9NLlOALOBtdX/be2Ov/FNLqCSTAjcGQeDOpFll+A
IQMchxin7kW0gIlyYuUYt5PssfmQxfzZaiT7GQ3PjfbO2l71Fqv234oE+dsY+Zwh
y8T7OiO6bTZqz9p46eupqOCmG6cLXQjdxZhOLD44SEPXnOZ6PxkjH4Ku1Y9EmkMY
1Lbkqy1IaRNDVoPAqT3WgJRi6byiBMSSbkd2JjCnSSBYfZsCmeKo4lUDp9UItkN6
Jbcb6o8Yp80FKjPRCpSD3BJhq7Z+je8zKCsBQ9jRgE8nJd5GCoLoj32deWNDc/vI
ojxH2S1WXHQgEIhe3exIxPm/dkMr63Q6WrZ+eUGt1tSjKygCuw2tR5DNOR06ivXS
EQExjmAuRshXzuolCSRC8qucp22B+ddhy7vt9YCq5H7WU3myelXDElj3LHmYBfgd
2lvTiWD6Spd5XoDaN3GHPKCrBwjxy6/JGK1GzO6OICkvQUdgHb4bzoZIFCETFW04
qFMd4RmdFjefgBPh/kXyLgnhuSvpyr54z1gjum9M8YVVsrCku4xZZg+MgnhQ4bjo
1bmQ2BYeodGn4Dc0tTQ0PSQ9d7Fxg7miSjOmZfHo5Cqw3SdicbNCb++NoxXl64un
mDc9BSUpnHPpZFp5dZYfxyEq7LKvoRoldKn2NWJVXKXZkJPiSDwNn4s6GuA4kAxa
TzefZ2+TDNb0NyiyqytdR13iwc1yWSajXeZD7IlGOYtYfwtd+BZaOfLGiM7TB+rk
hiQLoCOwJJGd5H+0BP7xLC8K3usfI6daV7GfYTxPu6y/dw2l0P+AIc1ss44XhtHu
WScZjo3ZKd7pgRKqhOUIyI+D2tM1vGuDYxdZkBv8LX0aCJxqoM3YUcmGIY5VhCm/
DM25naFJrA7QmmDsaxsivS7rJutZiMwy+PapFVvKvYrCVCrEGGTGkD9hicp4431F
g6yBexmYnGgFQg1qa2XfPFN2ep+wuXkpQpd/JVzjmwreOe+mCHLAQpVCOATllOOY
IgMIkKOUO2kJITQfJ+8y3C5LOo4sR0tMSkVf161pFscqU5m/SpCvxuxyFn71OyaI
XGTsCEFj2NS/8ZDKCz8qVZtw0K/fIlmJNqDf8q35fzYzwVVGji/BMk4cadzyF6FN
lTFLFZVSA0NjCl+p57kISeNDmgH7MIBgEo90FL4lB7IOFJh74T0GsYagUtv2SCKB
yVPp6NLftNBBo2UbsEYerbrzVad18mL1NUo0P2+vseOdiKb29ZZ9+ZCnhPq7rvE1
OUKB1LDQMf4r4eJEgo/j+U6xTHnXQeMl3PVpL1VeSzaN8v2NADUmfCoMW9ikYkFF
+kegSxlNBbuELwHZZh84kd2hHwwZOLTogxiHkhH+MwdvAve7j+TmQgSSx3p+rKyS
MutALng7+1XUCQnrXP9enJx9DVjyWhZ4i79PfLCo4DGsuQqSs9LahDigfUkAcVde
RrL71UNt2SC1xxLVHyIQJ7/VF2+gXKvPbU1ibx8o0lB1vMAXtUdU6rUhcCEx40ie
S6wR9ciCEtIOlu72XnZEFb6sqgoNdd503obx/va1PTNzQ95AX3TsGX366WW00vSP
G1JPiSKnoFevjt3U3KV0awUcELyLwG2vu2uzyk/woyCN35Hx28WPoRpTGqtkXCET
ZNRm0BvKcCwdgIFCKXW8TMLvrueIGGet2kQyCOHpbyIQsabtnouHSQblIshf4xN1
m8z1tPN+u4aOQafv00T94Wn9xYX6zqckiM2ZGvDgpjfCB/bpLFhycyXGF1kvWFMc
SVnQ+cRR1gxOLDg8wh6mnMtNIFxVX65rFUdYttrAfPnS/Bt8A2VCvkpMTTpVWjpF
6OVv0XzoEy8ncuAQe9IUfLnnUykGoVDElBRfFhWOaEz0RHy6HXytKI51gjhC/nYB
8Ma1g0VDsDVdLWHcz9H4nI6zRP4T/PVSSpJsvDvL6RYf/gw4Ri13TgFVO4OYodRM
fToCiY8L5MOfsmKDhYIoiYwDk9x4ZTkLYLOigWrReUszO6Unq0ig7xooqVOAirOk
U4Ss80KFhrBAxU2650apJKpFcZ722gwB0KHzjYp2o9lKsgDEEUPNq0eTIe0kkvap
bOerhTK2UTcjh9KJhe0uR+px8fQUMKvNG2QgoaIP4DzwmvFV4xbYX3k3aZo+7MqW
qE0+oAwL4KREWC3yvXQExw7oECyzXIbK1xaQ+JqtGPtBGx1M9wEGWIsBCihbIZTs
llUdNULniQobiWAbyRuy+6xZB1Z2iogD03HGlcfaGHrwRptfPCHOspK3O5XLsWG3
9ZOqvENFsRZKkC02iMdwuA4oBYfHyB893eead+Ko5KRxcbnEkxIZ7W5JLvo7FvNu
HjZvT6HiZ0gl6dcxQNjPizoY+O4oh6I9bYsCAbpRPXqgzyheriSsU5RbEAv0965d
OgntgP211UhwQtbUZYNIluZ/77hsHickzOaT+O0fwHZ6yso14YyOYFszm3qN7REM
am+R4urc0b+V/jnEZOdYVXsAzHrA0ZJ/s1zlTnBHoVWVaN50CTEBo5mlfYQBzK1P
fW13bOHqBdAr6iRiy07s9dS6tACHWmOMSiiTiu6SCthg8IIvlcXw1ayqkzRrN1yo
dJEjdmq6baCXjXl3EyJor5TNwuInqAa7qRQ64WbC38rL4EiI6zN48G+iYI/QyYHS
jh2iGa5Fb7WO5BKJjxwfWCBZufnheTQJrHGqksJDHzt19chxwfXfDaRKTRXk4WmM
R/Y7vDW63WaGojB66vdb6EDlRb2ui3KqM32DrhQozuCwKNTbzh5ZGsnC7Ypymp4P
N1P03gZwsZeKLM2rYTMpNqEnH1DLAmpGAR84XlFCfJbg8MocU8pBOHxCT42EvE+y
Dj+WBIVrn9iwN2D3C/sN9ag4MoGDdfCEZoWGysHu90YzFl9uCZrvP8Cx+w/drdTz
k0ukB0jkiKQnTNIMCYoV7PQ7Cl2RMr+U8jP1mRtCNvBn2pwFQaQwwi8oJz+DqIX/
I8M3Cw2bZECq2WZYaMaudD1lB9nO7Gq2KfWOM8UmnrdsAScAE7t1Xd8rijpCMvjU
kf8eiakWmDhszS3WGRp1NHOxMX8LStfUnx8Nka5KmDGRjDXV2XE4W2J/SGP9h+Tl
wjEeBaUfQw2fOo8eweI/nqNtyHojaqbNElY/nR5hsgZm7RCbmseEpsPFyFWn/lKv
/WH3WPqNGy+fqeQ+18FrWeHhAIBR/azMBcFvwkbSGCxtd0Y/IGU2JxzzTCKUY1l3
S31jL8uWu3Nbfd5fQYBslityoTsIQFdMo67NtLjJHbcERH5LM6TJ1SUr2YmDQNNf
jkSkYofM9cMAiOnKbW6SVT/Tmrw/uctbKd3+6g9LA4p7MUZx3DLnMLLozQjSDyoL
8shCX5n4lqvWHXoSGC1Uf7d5lGNntA55axPWwAj8sL7sCRlSqts7W5wQOocFSgsR
MgNHg5d4z5lpZzKLwtIEUASTMmx73DYXIYruNlOm5OJ4wVh8V5iHnGJ0au6Eitro
kR/HAwWZmvW6XviN+rXU8Wh02QCNFR564vzbn2EwTB2ATY5mjlBj51FrsJnv3l+p
inxr2zK0rvXRSaSkt1yuOULhfB7acGzaBHjy4iwjBx7akdI5k6m559reeuFlPNrV
m0BoQ8M642/1YXbZ3Y4+RBD1VeGKhVjarXVNQTngbar+b9ndx3wQt5yShhfagDrc
7MvRhYLBgrQDRwQzxipg6O7+CpRWVTalrgQGyKbC3Yxbq86x62ZGFgJsLmxSViXb
av87FzKbOlRafaSz4QdGz+7DeYdrPJ5EQltvyRMhvjbpJSRnyBB3tdgdYT9r+agH
XZNY8uzoG4J8qEJxeAUALWKWASUyLNUL+ikqrmyoxs8FCq/NNZ4pLbAoPLWW6dWV
mjDW6SB1zW0wkk8s1gjjCGS+DffUY/qXzdp7JsVrMDmteYUIwIRxueODAGMOn4BF
mZn55vyT/12Dq+9l9MJ/RWGo/yyXTLOAdNDb8/+4KsmVit3XRB9WCXiwLS6UhCwo
oCCQxiaZX6sn//jpk5KkZSW2Ukn5YfeYpDJKTP9PThrS2S25SJ0Lc+Hb7dGGxjqO
iMmYmFLDu6l8lVi8+u9pgi422Td7inCrIx6AFdiya5jpyCjOGK6OyLl7BIz2dx7g
ZKG4uXw0Il5Sdk/uGYuzE1AkDheHcKc0Qm0vjIL9bJTRbAzZzniPdc4BPfopqFRp
/H7DVqKAC1VPqu5HQVOsa77p+C12QzDCiqipToEI88NlJVaCxC4YP9YTff1t5n+g
UkMYyx31DKVF8RevvC1ngo4ZwoxnwW16TSyjRFO1ksqyQXciPmbk+vWPN6xZMCRE
74vo87wbb3UQ4V5UkPzePShVXxNiwedqh/KlT1SMqCVcc/GKAX5jPuFsnTfXuziG
BHboZ9hv7RWPRefSo+F0Hbmma16hAlAMlRAbm6nweneexOVmWiIcHZi0OvV+rrlH
wT9RbhRfto3bwASFKNbdOJOJhZSzMDzZBZsNPZupGEJe1NPakNksrhHzog7M3oZ0
wLzCT6sxwMBmysofWt9B96YWfrdY6g6y6OgxuYH4RcuhMHtRgby/LSmeEfSvLTH7
ccdX0XJkXIfKlxr2bXyAy6nOtIU7cZEhGQVBYiSUGyB+NsUCTVnK8Ob6N75l2k6h
Vrz0JAtSWPzGnp4aHpeXLV2J0uTAEI/Kz4mVIH7kIqQ9gNIEnzZMgSRVkXX8GjJQ
RXiJKB2jU/P1a7o3VfKr5InW/QR2HeyvJOjoC4zlEL9WKy6N4GwoMf2QjZlnc5+i
vzs9iXcn46GGem1BbID7E7JoypIQStXhBVq6j8gTbDOQyuCSoo9QijuHQyXD1J1Q
Q+BmSinwB1wH/DdyXpATKydnHjbeWY+s15wpSrRcT2sVuIF17EpXnfeaQmzGAiUt
eMPzRhkcPvjpeu+RwPpUJgyoYEJ+d/Uj4E/MQknpp16NcjIbC33++ollyv2XhMVB
y3S1GQhd/mF4lpEq5JAt8SvMd1ar3y59+gOR6vX9kCImN7BKmGL4at9GaoZanUrC
jcvY+O3ZjduxWn07CY7+hIE1b0gRqZusRxmw+tLsXXyMQJEARxtryevhydUUhnwN
2eKfXb7vSMiQ5QnePhVBoFs8jsIJrjzNYXQ0B+LFYQtnSjYCnwxR2d4/Mk5F/vf3
rhDrPW+LNY7vSArKlQa4QytXe413nNDeMrld7USNNoHBDYp7uTST0JkOw9v5vO6c
bF9PZiKI4vB5ZZmW+XZrvTqu9JXJPehswufgo5KuRr32brSQS/UmzpNtcDWGE1FE
MV21OQdiXXdnx3ENnBsb21DZ2p9U1l8adlbebfdAbSiMVByV5NKvvion6siPaZu0
Qnlchviz1Bp4Napif3WgOMAUeJaQwPEBEBnsLd+PDFsHdhAmHuHTgpAQ7n8i3zRQ
OMuVQI4QmeGQhK9kFaqEcVpRN2epW85nRLDfm2/39I9nT686GxOhcPHKm9oap1Wx
S+qQQsA/RLm/nYn9jbnpkcV1UDt6mpUZx+S2iLY5EuYokgnrypv3c/29hxQgmGEv
smQULBVlVc747HZkn4w14CpJmx/v8UWdXLKDb2TZTFL0o3UBH/+B0bdxY7AQemdS
nETluJ0ZGdWgaYS2DADQLOKkGgXHfachZM5k91RbvxXur0iiv0Dj0thr2LYRGcOs
PSt+i60JLUShOV2Z87QsBlncou2bvsDh3pZlOYJne0WAOtgQZfi9wS/+RFnjkvr4
pVoQ7OgbfKHTgxFU3zBN1WFLFQipK9g1g3J5xkkPHe34t1htwtLanFUQVNIfDL83
gIprovTmtjAanHmSM+laLHOwCz3efSpuCrSomSI14CCqFEIjCn3EjOOXDksacmqe
iAaSr0Aet9x3v5HvPNTcPsUqyK38QbXjDfULxdj24X6EhneU87ydUAGF/ylHsB7y
aHLYPMbGc9tBgi5fzYLZaeI6+ksoyKZou3zZvDtjSS1FfHwh6db59vQF6lbWhkor
y1Z1VrtAW56fxoA57NqpYLF5RYDGJMpUO6b7U6MWHTnu7TcsGu9L6N7KR5/ikvs/
zdcn6huZAqQVB4qJx4GdjsPirZbvbTUHRPB6S+BZF0EkG+tLZoUCL4I9Bv6bWR+J
KaqaShmBVI+7ZV3Kex7bvDDU4y1G8TO+zSTEzUZK0+XBLnFdDwsyjpV+vliv87U7
vAYniRc1xLjwTobuUwYqtcDAW/lNi9GBCVFwzlE49dq4Q4iRi2J6/jJQgHiMlWJf
q1L86fw85FNNoxYIRnve+bNSiL/PfbNh4xjSzidj3CoG2qrjjXRgaWgGOoK61Pm9
P/xbignDcAUHyWe+qrtFH35tRCPvQnadyQGanb75HSaGFpUWsjImdPJ/j1gz8uXL
DKj/yEBTOZ+9T2xhNxVbActSmuzhEtp3MbiFhPIMl66330/3SjepgwHHlcrKNlZe
GqP6B6gHyIFgVlFhckEECXxTSTcn69rAfMilp8fkmL7xHU9Zi/SuUovM2ueePR3i
kiWpJDjJ7m7cnZNsJ4prMWt6AQYZKLwlKWaTpjUjulDKhDrPlE5iho3CkjiWbyFd
1O0dolttLR3GFFGhmEWtr1E2VNvgfPly8O/V0ayrbmlgqkAMwolSQ5ktikTtytxO
Q00vsMLhlgqvX3JIOISCwREqo4vUKZ/NI7HJLtT7Ghinl3ifeuMp9v7Cb5p0eiLh
tIyo1tuMDhwnGvVGlRrbB7KDMEythlNEHazIc5K1o3DK9PpL/2fc3JHJoeXXX6lZ
8bsNkj6wjZNRRLC6O8xfzIEKX+KOv66fLQM/GqD785/0TrodpUhGARPLV2+zUwB2
vT1T1fpXMgdOZL4+KXAxRFkd70ZA1K2+YPbRy9SZR1dXWJ7w4doyHGKnFmTyEmJ1
RhOhe4j4eCgjHrO/PTcA+uBHNZWAYi0gn8gZHM9KlTGMWtR9DaBGZlW18dRTe4UF
aO+P21ugoXResF5dWNONhodytYyjxvDGtR4ivk2iGZBbFlh9LXAtGm5DX2cawzZy
3ISCLcvNLEfrdiGvaguLWYnUMUy+rLuQd3Q05jzHC5yFhqdzsx6JIVhZm5McauWI
gMOyKm7L4zOfAdbYwSJ3HGO7rttCgWmGYstVfGsIdeNIKewTmxIRqLd8lZWHOh4D
ZqjuQKn6hlv2RGEzZ5Q0Ki3qpeV1AQ7rpOnPaAxl2/Eiqr9gkHJtwr1c03CYyfnP
srdVsqBOlvqeQwEmwKS0a1k20e4ixVWRZoQlwje4AwnV9z8erEh/gdlhFxk3va01
a674wUyzlIOv+0VEw4kU3xkvmT4Gojr3kMHJFvoivBLgSGJgp/+C5ZenBD9+3zVk
m8m5KhXUKxGr4etJktVLBfovJ1PbCwkzGslgjyS3SrBYe0Uru0YXLrQlem7WlXlk
lc2JGcX8PhdU74Mw63TtCjVFAxEpp2m+Cc5Zm76F1ddp6x3nC4iOWcY/Rrv4s3jD
Dr0jHPz/T5XLSXjGpv9fC3YgM3M09VpH1Lo5S+YiGZdB/1dxhWRnGNi7nME4tUAw
By0QLEO9Gs6xVLgXFAll6T9nhpBI1bjAm4ahoIE+ps/0WmnSCGS2uakjVQBdHTSi
1TZ6GinELC2cngKAQT0mXWZSfIc6d6+LNeNw5v5WjIGpd06iy+yeCDMuNacawh1w
A13aFlkwvoys5LP6tSkA1L2dCJAOkM3csND4/xkrnhOU0bH1UPvpMXFDE3lzj92J
N4vVGlpCsyQt6Y5ycxoAOXCO7UziwZCexhN51t5iFNFhgHEFQxwKBeyG+8EbIt2v
KwQHLWzztChzeoL4Co9Kmoc4y7lok5l+U1xsNFYvQklbygP9BfOy9FDHknVJ1unr
vaCU+Ueo63LdeVZvU5BFzeuy4+kbBh7lsXP+hSRhGTdPrKxbNgkMLAZtl3vUmKcy
oUUgRReqAIrfiQrynBZF5f/I59KsDBHvEVEH7u5qHU6ghVnbhtmpdIwwexfa0Hq6
Ah8wZQGo0e9IjcPbR/WV7s0ohKQwQjkk8HPAN6xJrMxxFzeHwLWrHwdyrgG0GlQZ
38yKGjAO1gXnhfVkuzKliihUWky4pZu6oKUjvbnJ5PDyfOCFLGz3YhDSKM23xErz
eJdSkwDHJtoTc13XUZmG5jwhXm6e1wNCxzf+FhzZDFD2qnq7OclP/CHivH3Ft6YP
jg6Ss04b8GlIASDgYMlCYeFXgZraZ62PO1A3CaUUertiDd+pSvY/xZYtGG0CoA1+
5iCIh1bC/rYfAibBazuhd/hFWr2q9dLq0xPKVYpoGtu1CGeulQGC4NPDomvxjkP4
uLJHwABsCKH0EE1B0irJwPbIthAhR4otx3v9gt2wOQryfuZ3Xv8NBYfem60pZ8Z/
xMVJkvGmi2mZCYkEqSr9USP0xJFDT24hKYjWytgakw3CKoWL5xv2BJOMnGnZcmny
hHsm12S4nxIycg+q9X/EVb6v4PDQZ6YAJvIsBPni/ox614k1+x5DJbdGwxl9OWlu
FHa4JHFeSonTOQZjGkuISRkZ5tZSfTB5rAfknIKstozZG8JP+bFrrykrVM/RRQhj
ONYPsNG2y6fuASaI8TsGTV91VDm9WETVClB2YeLrGUkjcw+ZaRRzW2zZUn4Mu1hF
jmqSpLKmJQwlL+Z0lOut6ezN5Jja5GIkKIruB59Lm+8iYQwllciVPsjM5AFeiUC8
DOFxQFvbbMrSuZKzSpn1iyInG3rnUlS8BmH4rIhtmhT4y2c1HS1a7kOssz9IDbQ9
MUIcdMnBha+FVQM1oepgRfUAf2osLxrlumQCEhDg/+919nqGphn6HQFs+lq2nAzK
CqJBzjI/lUTELq7q6faAxz1jAP4xXZOFFg6+fXC5Ip66+vcwNLhJ82+ENYtL9RON
omdFPLmEyJ7rUrlMbcCdHl80hbjlpTurJd8MozBoT+AD+OGSNugguNFJS1wNhgvH
RXDMCXUK1stpvOLxJamF7DWO1BqCSEEz8TfTv0MkrYt0Xtl7rQfMco9Oet8QkXDj
4qK9KYE9ZKpRdcHoC2sK0Tgj2MF7Wuz4uspZDTKx2oTgeeNcXtVAwToulE0UtNNc
KsZJ+wI02xUw4Ufis6idHUDJZMfNHtIkzu0/w13tpLhEio+XjMF8SmF9UsBHIpHM
zZsLdTtD6C6tuZHfqAyS9lkaAU4YQo7hhTntC2WVSpwN4PsnDU5+5DopZCtuX/+S
sBdfLKetxZGq/EmcPJFOx+qY1p3V75ZnI4cJkOkFwGKp5HqITvvXXCg9OQyeOKyC
fmOerQWMP1wm3Xu4wAsrS80n1BCh2gwQMbjFh+P4oBAyUqY2UdP0EYXRpjk1OwiC
RiG5nAMWQp2vWJoOn81mUWgQw7wIOgTwdTVBmWDF7rDFIXmCEgVvGeB78ApsaNs8
ek8GgCpVBa2Iy17wa7mpNXBy9AIryP/N25is59uZyUHtVGuprh0iOO6rRTmgC398
+OhPoWiilR2GpnraGtaQ8iLI/7ciSKaDvhbMrAgplcSFOm4xEhMdHuVuGGyyS0P6
TQktRgj/1Ph+nHgmqjxAz3shskucMbGFbB1WEB4MpDADSnjGBDYVRmqiBgYO8Vm6
tbu+7qQDYqsaFZIvcrkIDjSS+rNHF1pLJqdjA4Fn3rnZtE3JukdDZIFd/LCy5OSK
PYZ7VkhrnIjXZFt9fzAiAiRXQUkoGZ7lR3CRPRpWy/tAhKi9WdNVWbaXIM3ATJSu
DZiRL6DBhfzUwOD07RCdK4z6cyh0AtSIgBeVpF7h00NVxB+cCkWB2yhG8HcI3ol9
73wVI6MUei2guDw+8X/1UVEAUcAZuTGfdPdTKQt1V5bdwZXCK/D4kBk9DCgnanBZ
SlkF4jaSJ+4pXEarfmoIWDzhUockM8z7pXh/gvouey1TXFVms4DCuwUYWlBkITGG
52FDkk58v4Apy3acbgd0bPKbDGjFVWWiS4GOXTNZ7MVZqWD4ASfjFAMLGU1tzkBs
Zn5MqZCjpOflRyM7l8KbCqLzGYpH2lffySxezJZ+olvduWdBpsCy/HS38A0M/rl2
GdUOkc6g/2BnQxDWxrbik2ZXvUm2PdAFT2knaxj74faAnX+Z5qRWaYa4cAsqZ+i8
edwO7zdulyx01vPj1xLKAsi8EOSH7z1n4I3RZyEp2CR2Mm/wJ6Xu67fewkvpvuk8
r30anYW6XTt84097mdVm3Ssv+u0Oq2cCkfVW1c4w3/s1Tbh7ybBudOdfKuEikiYD
cF6ZycxXcfc/6GGOdQL+dfAwfpQreb36ZRS3f3UKdGPYxes9QaUzGF3zOGyzhUi5
ZsPS4yjQRqUO30oismEweZHO5bHtsHBYxVjwVyEL55ja/i66/sRREM31EjuCGwDK
QqDwzH3LMIHdlWg2HDLwOZSZqBLb+jPN3/CNHEnvm9OvnU2R1XuYkx+giaAWw5pH
CVkkgBRmxjLEwPHI8JdTDm9rnTQgrwcaVn3qmNCWN8nsEdgB6B8jMG53xM/D2vAT
hogRls/ph2pVACgvNEzFujuGr01SZXeR1u6lHW6ecxeZdrfCetIaD9djL7EHZjtz
WZG58qw8qGarFKp7MfhcNL5gifvC3siIx4G3MoFZv3go6c1VvwjME3Dp1D7dYD6T
o3JFGo0AudjRU9fIw6p+aKvYVYjCv/drpgKPtypPYo0LfPa6WkWJNPRi2ymNNl3s
X5QKkGjRMqVxuVVT/T7M0vWXOEFdGdNn3VTr8J+rmVjMk9L4n+EdbXaX0o7cHQqK
86XWNjDznDYLuNmOOGE5sHF6p4AvnqjCMwKqSLYYLo8JMDdocOK7yeYGRmrTBxbL
iw4lLSZQxr/f0WRVTHh+NkaiEhM/SsGWLNrv9clMrAhToUXFbGkyhtGkW251WogH
sVoTfP/Lx7DPj3OW27sl9yQfVz7FDDkLjOj0kNSSopfE3aKpF5hat2G2ssGGMo4x
rnT8Nm9UXjdNsyVJyy3o1+eKh0NQOzAhRWEJbmiqfDxFsw0PX8iqOxp6ZXzMfQjv
vMYkZypT68gdmMuhaI/u5cR7V6IZB2DlOcZg3q3dTDVu0E3e+7pG4ctbxUSMjygN
+phE4UvjYHmOYlRHSMheiREI/xlOynr9OwbBaGEsN6PcaNjFCuFvH4i3a6cvXJxE
oIJeICOHD2gJjaHkZLg1qJz/PSzv9wQO4jV7TlsntlP3sSptpqv/FQA05FmvX3F9
jg2JtuA3GjDqk4hGaeT4SjcddzwftLGmc988+W/kcTg3Wps2KZgeo7VNar4ea1GK
ILTNAecAgd6YxLdFHqDoZhMjaynUEDancQRG0V1PpckAL7Pr8mAKbDWer7uEt9u2
tca9hq8M35iBXaboB0RzD0coGt6nEuHGe/Bk/5u1etiD0qIoX95fn9OJGyUMFQt0
qEvwVlqKCvBxYJYI3amUL24+ebQqS+r56mbHibzJOqiou924OlXMOhnM7k3iyqCB
nJYQPdolp84yYbX9DoWEAjwhQ19jCCHFPdK7gfsZow7E+syxwrv+gozH2z80kh1r
K0U9dS84HRjBVBKqNZXRo+QveyTe/Yw8IXTGW364ZeBOvUFPjjJK0bJRSmP8vFj4
mbNj7yHxTzJXEU5kgE8DbVVWqrPfbzFRdvvD3smhpz1KJGL9TzI25QNcDkUjgB7D
OhLT2JTHYSEz2Hn5/jtQrfBPHmKOOZvnDTsbJQaWsQ/creg+aFQ+AlaokfvdISw3
IwV0pm/LdGvejOoORkF9bEoAQ63KZrZvJF0GXnhc8GL7IcZdjkILu0/0VyW4qu+R
QWqbo97twoY4gmXv00wf+l7p/DuWpYiggV4RPj9Zf7kM7B9w0a+5fHa1PI22cTH/
DQ4KVJ8fYnZIgILJaT+PGjwnDOE7mnLOCdEfkLI5cMX2hFVdc169WdGjtoFcIKSX
22mvg8nbppVjDw6mjklsXT+BN5yR/0WoRmqmNZBdZyGCyHb4sMEZBrp/+rT5OHei
1N6/Oad624wQ7kBuWs3N35XSYw2AQv+UJ3DEwGe7Kx/6PLv/pYYR/Mdwa39vhN6R
sY4JnI110I6QyOJPfp5yyd2XTLC2MWo6lzOpT3Ktgd8x3nCCFKITxIFlbm2I5LRW
haK1inqRXQkMIoZ3iPjPwwvyiaZfHbPlmcqUx0s6jgHcSocC0wk0epGMhrN6oSSC
IaQOhUaJOJVvIBwAEBk3r/cz6KXRJVI/vNMy3IeSzEJktwjarJnd54KiCN4Wrd9U
GGLpSs+EWr/d+mcLUFs+bUeL2fUQ7vHC6rrvz0eCszHUOI00g0FbeQBkJ0QXjSG4
TeeF/XhR1CZnv+4VK0EV9a/ly2AweNNEYOCcCRMHwj/4bHo7WxBS/hoi0jxx/2FT
Fy7oReJrYOsBjCU6T73yvA2Qn0ta0O9FdiUAneAAVTXgyK2hdMqDSG5m99UHUUiB
AhyFUAQK0+aSGzJ1HydSRSGFq4uIDe7V1GFeb/odphhVfOLxRjOQXWDD+5dmEDlU
h2vng9X/yn9mwcov+NiW3a3GIOC2ayAsBtLDmcvUIIAgNY8gSTpTDLHtGn46XzDo
Ap9PflqZ7ovGeqzrF7KQAGH4AzanIb/WnOLJYDmPwmTJdJUUOjWQBzZMnxFfTsOO
OUTcuncxt7XUQxNQz+Rcy9UaOlC8rio6Hw5euZbI93SCI1rs+X2Wn8SeOZ1cYhSC
0sf7sBQa5ZqmLLfhofZqbBjTLxjZsC4W3hQyPrvoqAoWN4gvIjjLmhKHL97wl3cZ
pmV1QIhPKKa7ntGLJotUszpHtkvZJX7BlSFXog+KptjxwGV0zEvKyQZ+983rAJBw
d1yfjU8UqdsxlYki2dch53OFLHGlvBW82s4KiG8fEtNYQDyrTTo/jdbY11RGzS8y
W3DFL4rsXV95bdPhwnLPHZuEyre0qdN1NIyrdVU5RSYk8rsJNHbilmhKHnPzKvi3
nmEpb/UjJJLEbP7u4UfdtqFttRtwJyKBpDaXjdkp7GFstHvRtdwM9nW04xkiuxtp
GODJSlqC8NqnKz/HRpzpr8M40i7fZ6OBD202hO8ZQaWnwSy5W9zXcnatjYTDS6SY
ZylCV6g3Qa3FMJi4QmwFmIHTkMP1Gg/BhQk2hGSTlAXMTZCWqAymqbO4ezbAcGz7
VKsuwoHvBSNvmljntUQwS+U3PvusOtoxSS5la1/qRvbp3rg8cHnhB2NPBLGMZmH7
2lQ2pR6EeN05bwPBV/V3S6CkAQ4STBY/C1oomXnAwMYxPJSz9rIdd25CYzWCrApj
mKgpyWTFkR13qmyiWU0Akqa1mGVWDZrXN0XmVUE/IpUGee0CAzUMo1H8EkIRSSFl
xnAj3sqImC4YvUX4w2FamegD7XR3ZIFvyyh8jI2jp3oMUYk+gt7/wcgSrzV7kRLE
5WmENgMkTIETWuaZWm87UT0czoF0CHY2TemTbCx0D5ToDO3y6XQqJbBux71UlXb1
J06xjRTeRZhSTmsvQOwwomxP8y/vtJjsnQfZiNy+IqfzwMjmKnJGDTLzCMMywmys
uZnkMzn3KUWOEgkNSMRWVcDEldSm3jxhdTgrNYYww9TuDz/rChqv9vBSLw5AJ9uT
T1S28N+y7YU5e8iL1iLvMemSUA0Uyg5efI1QKEl7yuPi0FeplJNMvfGzko2OrGC6
TrqMwM+TU4r06rWpGPBa8RziT//s4jlOPPrtPlO8i/2VAj3fcC56x4EvnN31YQpU
g456/o7KTCXXOpaSRtNvFA8aU5oZh8dJC6ANTvrxLyWakqS5oTRJ4tpcgOzUze6r
qyhiZ7mzWNUtr3HR85ELYQW0XwLTBkBb1wbU6mVW5kFYE2SrenV+wgLd+uVsT4lU
ekqQnawMc5du8yFeMLtFOu5o5caThDO5skOyHU5XE1L7uPNAgNQRSoNxly6JoGVl
aTjrd7tkY1jbkahrT+78Lb6U3PBx9bC2fdNSUgaGIM50W2b/XG236/R7jIwnr/YL
lt9T4IDHGs111rb4ywFrngYQoizwfcVtlmeP4/L84sw4qNc3apTP6RfzSNhbKSaW
dscedyGqC3FYIDWigfhzIRtzTWqHfB8tGFYSbB3n+HRkEXhsANB4Ux+ksNLbAw9i
NGVnPybE0yjSBDd0DYxdwkKkJWEV5VtXsXblIwS9Zr8O1rwAPAs/XKnAdxuUNi2x
Q9j+Mt2A69NK6fl2c7p0qdSZtwf9Cv/sHsWGLRwAvFr+AsxuFOR6l7j/4P+bCIJu
D/kcsyz4dxuOcAazmg9GltUtj0+EY67CjXbF0bRMxYogqwHZ62B833OyWzA5vRRv
NGZ7nPPIem/h9RR/pLwPGhkv1OVMKS4YOlLZwJzkNF9kRNxMSDCS068jdmfPA8LY
WEvKL3JUVonuQ12JInt5brmCFVkisNIoLNRYdqOEFt/az8p4q21UYis844AFrYyD
TUIGsAtfqFAHigHnx58oaNdtNfNAeTnJWIQn19ETFjVgz5jtDazcxT2gwKaSUNm0
NITzErqyd0wI6qAjvtiWMOWHjUP8pHH1g2whCVtkeE2lJNUlvl3nZwwm39dbJeaJ
3tRJD+Rj/xbaSQi27dQ2NOnqLz8sjLBlPeC3XYEAXDIkDorgCe2xQIF53V5DWMDG
0FQI3ms8RV67PHdlSOCvBT1f3wYjKZr9L2reBG9l5dagcUcrmS+Uq3fOtOl8dzi+
cfVuMJrWYE5zrhfvL1T8S17W2ci5DIrAfZsbVNsDgLYhxJutLfvS9hQVDJciLx19
V33/wfX8fs76SE4edEQRSEoULGvJEKnZ1V5l20VoJiHuYOCx0ImMDUNNdcZrXHFE
kc3eyEhs3RZgnpesJxtgP5EKk/jitKMXYKORTeM5SPIdLF84jtAhxhI8jcA6FX0i
od7MyYQ/0nFAkhBSH1GbC4DfN2qEP5ts6DVLFjBSVzosdxS6uWcprxvGphSn2Iqu
yZcWx1C1hJPS/7J9afFz27EwP1ntRvg2RdQIip0K9zVaTI0+Cnp0KRzWb+auh+EL
0PMvByV4PT63GoQ0EcRODnhPMnd6y+ZmtuGb5ENkSlIX7JqusG+vXjucqtE3V3aG
TjCK2soBb6aKOCQ6zyv1UBMlr2S5giIm70VUpXTuCz0RG8mGYVQLd7zSnWFNo6XW
Ac6VPC/s888uaywwAgMk5jjKIceYOZm+xz4iovaBjGCD94Xm+NMCAYLrttD5BrqB
MdpeBkHC5QDhg8yc6GiIfYP0cLNtsZqvGd3Z9foVHJvZrtpOUwmGBUgw4nv+4JPE
MgwoIiX8ERlWwI5YaAvbS4rRpEPeBNNxs8TjrxC6bFSmYmgAP090vzxr5dr9+ot/
j310I6iiE8gqE2MTcD+AiI/e+oVO/hqFy+zuU/UNWswGnzlNNYDOtxq+iGAJu1OC
KRsKag7+wmRFnv07rUJJkvB77+BELoU7SDpY79OY3tbjekguJeW38GbQ6kGB3mPi
NzBXyedP3n0CZwp0l4nTqau5pcG1FTYRTIc0WCgFFLJLDydKxObDDYU4c/HhE7wD
nkaXTq2AkpYj9vOwHrosLLnbFjAQevvuSS0m09Gxid1rzDiDB6FKk7mBaBfvDe8m
+/2nMw1gJkucmloER02+CdMwcItO8eD80A8PU+XeNnivBlbdw+0AwGExJMMgl/Tg
1C91xGDdLcfuOt9xqME0CNLQLIj/g7q+JR99KLq9KZUzZBVeSLoyXJE6aGjPL1dZ
IKiBC6UcCOkeTE37Pr4X/Za2S5dUyTi1UVKc1jrkUMqd73iGJlFYpo6Uew0zrNV2
skrFHhJcv84NJVsP9cI7Z0vb1LO/CO/z8IVU5VHQE8BeP348mxrjsZK7f63sygsZ
WSezetcPAGKb5QjT0WevSdsY4gJwYzFDKAtaJwDDhcROwAwFki1I5/xNDAPsPtiX
gaRzetEVRR5tpwcKNS9X6pa03nYUlpDaC9mCMz9izOMfG5TYW/iA9DyUgAnfnCkU
C/QIoFraanuBIPxxTi/w09+fkE8ZlwqQ8oaLSXBBg6rKs7erEsnVnp7v89yqBY+n
29fRiqVwBPkWX8BI2J/Q9siYupPzYFMn43s6n+a0pgPSa4QQoj0RnyDyMfkVxJ0w
wobQk7mQ44t10RN7K04l/vzvaiR7+FK1qsqtbxGkDNqrBZL6cpZrnCvMi6cE9MYp
E5CLiTEdIypafFBKVZ1SsrHDOv6/BCASQmbXyleIUS3xo9e/+f6hVr+uKEW7yL8M
rIURaB31oLIdab5bYFDpr1MusupwNkiwfxNMm37Z2HREbtWFSPmkY7L6Tlk6eQIT
nedHmKBAtSsrKlaNiu+20CHG0f84UqWoT21TCJPnp30XEh40rwxbfyJnmQiNQswb
DPrusFzD8wca3ln2YSkbzSJzjCjs5Ta/+i75/kHD2/Vz/7aswAJlkhTHwIZi1E/K
sl4GB/rgD+xfTKsQkmmTz3/T2ls01C5p0b9CE5Dxj0m6l69mTfXg9cefuCWaDrth
cTDVaYnHZWsMWDq/b4Seu5zB7bGkAqeB12Qhgvyuv2DH4NRs0XacQS4t1xHIFNYe
QPAviW+T3bX8TEm9kgQ+lTK2RnE1/Na8sf4A7Izb6lmewGNT4fFoE9doy/tk/VFO
LkNjtt60CIGqba/oLwWGtXxtXTLf/6Z7AMECa761XVrBUlupXmAMHMzCPo9Y13mD
leVUnUK5jiOWharvbTPxJKTVcII7LxHCZS2ZtG5JO96XtEOVALjh7cCH2hLHX0ZM
v8f4sMG4m7D+P4u9bc9rljBsPBhY7xEfVXbF3uwB11mRDN2236jSFTOaZRx7J+Zy
2bH5XjwHTGVNRfJ/ckzFcAJBqJjyHKTvNjZusfCQuWeCn2YzIzbmlUb1kcyAlbkJ
DwaPsdz+uDgv5BKgk4hhzZqHOrFu6kfzY8mbAYVve5cyPdss4Z8e7J5Fxd4vlcLV
jmaIMfbwwNHJQX+l88tBZtnVTQZaFZMalXi2NaXIyltXIVpM7rlKNurLmfS/368r
U6g4VgcbenG7SZc+R+R70/kPiogoeFdEnL626bzo4FpvtP65Ac4wsPUDy9/fPpcl
qAdUuVtaliggv9RVkvGiWKT/RiYsOQ4nAjkh6P0aGpHltrLvFtnD3E0976xA+PDB
MsFT/KelDR9I0LSW/yH0Mb6/JvaIOeqpcvBbBgZKrRFzdcpU/s2yOHBpZo4BC/cE
Yqp+rKLP5ctKXEJRyIYbDjfOO8Odxb3ZRIjGV0mQA+uQ2BTP3pK2NHW2vjAwhDdM
2s9EjiHS4MEbovi1ZEGlV1g05mHVxo9qEuDSz7TfGsI/ALETzwgOIjo1ZOIedFvc
naTw7oMYTQ9eMBAH/HC4MWXebktUaMwBTCD7qFphdXP5OrMoW0yq4S7EmU3Hr8dR
5tGYJwGzv7PEbX5e66pgGkWbwxDg96qlZqF0Umizw0O27FpuVypMq4wFYDEcpc+3
yRMMIraUbWe4BZxwy0smebBgRN0nLJk7yaqbImw132MKvyBcYM4SXKzeMi6Qoi2U
eFJ7YblTE9b73P9qqy+hEreeRNNknQnSBzjEhKXN9Rcygo3ZCgGrtPj8s/xUqbK0
EtDRZuWfMy3ZT984JUoOM5pvbxxo5A15tkY7I+fGKqp3wRi9wevbAmPEYAX/F1kS
WE5zX2xCDRwu6gywc6WjcNJLsf3uZzmcjdrDraKdIitANVegWCJDshAa1y3petpn
f3i5trMKX3EfsfSvvL6AFQ/hC5sO4LZMWYXQrEQfzt5eUTwz2Ex+xnZBe+MovsYK
ZgroKgTcQLv+wIFRrUeGrf2z6zVAorYHCDMMdYVIvuoTpDAWGDFTMQQ2cWbmLJ04
GWvnCci9eOG/OxxvZ6+Hc0iFz54RvC7ERUWeT9xPhmW3cduUjpV/tTmJDdiJUXDl
sBt6RyYQ8Cw09ZdwIPgOFjeWl44CPvObRl7GC5gH0MAtUHnUtMVkoX8lHBEfSDI4
UFy2/Y2HTzCntVjOFFcD6ISl2nIVSH7+eeCYQGa3H4aPZ+hhTmvqCK+s7aqzqbCs
Sj03+8nljjRcTPQhadu5qKWHCJOinAJD6RFQtoWlej6jAsuo5Xh7iUzIIm92emFQ
DrBKVr2CBNfWIGrbCEtFZyZc4ni27/8oCZVEaXzaH3Y1TowP3TAaBw2Ue5iVWDH/
/EhLt/1e/EYNCAqKgIiu36DnArvF3OmMgaVTdwwXT1neQfNRdeJhZTIFNvMegWpy
pAc1PK1z08lY7C/BkawuEAXF3DBh3v+ejU+lxKNDYzj2HfwcrdFM/xA0rDyVht7O
jbTcGGQwQyOYyZ/BYxRqDoG8AyAbfchCf1qEI4sxj90eol6gXYUhe9/mmu1BuX+W
iSi9I6pQUqTP6IdNnQQp2+F0A75cqau8+XNQAlZF9tzQ3w0l3Io/I7oeLKAhdTUJ
rXi1spf7I1iSsOvL3egzlC7xbyOJUz3CVv3Wlfw53+pTQGg4m57idOZtJb79t9fG
z/0IrA6NVD+lWgp1OdqTnRCMeDMw5VP8p2pDq79f54J9G+0PJp3r0Xa83pOYuGOl
yKMJt5ZI7Jqd5MxHhFwOnxvxMPpsc0MJASBPZ5uV2T5zcJ0A787Rt8OY6Q4OVbcN
Q+uDg8khhDtC4diI8fmVjx+LPKVawORDbWVa8YY3/BV5c0BjzYwdYmOO3shseJsM
T42X0EWs9CvYs9HM7AwSwSJSlhgEtH+cx0G/aqIt4dP0mMFEgr24gm4pzgGkO9yN
u+Env6bzRwPrlJ6vO37zEkY7CumSgt1N0czArucdFs83a77EuSOJpxMffyz0FkIw
QGCF4LRs419E73hkO141IBhe3hETiwmG81WmNDw36fcAyWfPwGqsi/IKKdEHYMMp
QmKalywSH3g9P3QaFod5Q60uFyaZmK1XE1bc9J4JXZn0VADoIcO3O89TFi+p+GgO
kiXTCITk+7BkVPxjVw5v2FU9EdkATCprBHEeBnHKwuKNf/G7y1OFZuAOvBZdY4zJ
pfIIQQRo557YAaiYhXbxwpjzDzZnQyYybRNdqvesk52lLe8Ka1SmDeW+mJOUHvyb
8gFhpfaThYDPdfnf5olb+v5RL66hGEbftZUdjAx28zbsqnS8BKS1QuLktGT6Ou1J
feO5gxxGL6vHxjyT3hj2brrPPsf1vlf7tYICDVUdWhInC1dbb8upld7ejinZ/Ro0
/5qNIWFusPiPPv/sERIjDKsd8VeMA0zG0ify2shjjeQhYiyGTZStOlqyfB1HU6hu
O5Gnlu3V0StTh0KC1wUITcxy/74aZ3fxlXydB7kwWnhiwUWV4Jc2e11LSt5FWaWK
NSIoOjsx/QS5AoVCqiNYUPo1ABuK+h+PyzzGhN70H/MmYmxajA/RrfA44yQPbO15
p0aZFGe8VgNBD9weA2ZBaeVzcanj/HuTZ5iXI0pkqJhTedoXYb6qbqECcKp5cmBg
32cEOM3331J200f/L/rwwB2Ejh41l2n7Mg83syWvs+2jeLzibyTMDwAmqWwuSqhm
O/0P9jKcze4xteXGkwdeH7QjhBTVPG8EHzsTPiWpH6wcfD+Hk41jUJFebnMIlEoh
OV/eq4jQOQ/tIiQxokXRtrnwytpnVPJ7Xe5kqLHYZswoWRTdJtHMdpn3/XTNc8m7
ROH9+5gRae61vK9c3MQZl1YYwDlJsj8fVig21cmxtYS4FGk11JtYM+n9GNOQNvSN
G0KVf3VlcJ2gSMtpc/1RVuAgxZE2cdr8TQE0aQ7/DF/TAnnRbdsU4uymOFIW/j3P
C3ypuSSZpEoeKjYMmelIvdBRW7VLcD62glLSMiUOn4jznJgcoi21ZK8k68pjBcfU
0z7HwlYtpWBPFd2YMJTwkCPRHRXPIuChwKH+Uhbp+E8+Zewwlo1O758Riq7uA7nb
n5uUZBgZMk3oTc4N4XU5FRNk1MdyRAVZziA5BPos817eDZvCDZkX50wj2XGO2Now
dgryjh8Dmi4Rky9+XQQYbmzrzdGkaRqdtWI+03jD4AP8gSHAht659EHlAkXkS5dE
Gz/8kH0vsXH7iZEDY6iJxEiIm8UDYjHkahBsJfen3j7Wxd1HwpF0DgIb3V91lgV7
Af8AqYfobweRX453d6SLuXxHybUuc5lD+O+RBD8ITTVxhVopYTn2H5iBY7iFrD1T
q9I9tSzq9ZvOJzwWHXeGkmZL0zRROx6F3wT0XWvlANDloVi+ftmfQJ3hpJ+ivx+9
Ic29ALhCAqUsx4utowS0e7TEUwPRY6d68pKqbmn1mgSmU0QGJqIloubzxetaPz53
N0P6Nndq/CxHdS5cK2CZUM/oidMwp8SCbJAVyNqwC9G8/XYD0iOLKnKQhuQY8zXX
Tx8QJ6Tvg1mpy2zyAi1p9GUa97zT8v5IB74V/sg+952DlTRGUY8tgxFJ+ddb2SXH
P/IDrhBl2NC8N9IhaWrbS9yQX0kxyqAAhi5uIteB9hzl/LYzKyeDToCQVk746Ujs
HJ1Jwv5lLuhsYixW/uDmmoKDEfvg0gErWVMz+pY9Z6UfVogVyUS/xveR3943GZ4D
P4TP67WEAOR3zkarj6jCDrEqa5a6ISzypDbjg9GX9K/69ZGX5Moqb+UU5HHscbkC
EvuhH/ZLk//XhmDiQsDRghXpTmv1mpSgMx+I+3DGcRz81u3HcrIk6jBcLhMWBxHO
McBrRwq8fFEnmanBJor98tRiz+YZEZ1KS2o646ITlJD8lmmU063+sVq3UrB9OEB9
jmdFceHop6UFT9JMBvacSP43IoTpmE/yKaa4qcRwSOIJvb5qRMz+hV5J1CfddDWg
QNXELdu1k7TjDCf86e19rIkYyYpuMEvalTXjJXm8j4aqpMcmgQ18WSb4cXLFZu13
VK0HERXvNE0aWi5QDFk2TsB6KGel9gSbaUhZcSanXgKt9Sv6jeojAH+71HvQFgAf
aBeYcjoAYo+qLHSvysiq/Ayj+wSkRuTcAkX1rpki/OAWiJUhmfUswFJDk4f95srx
XIMVLSu5Q9D92y44ZnFlNJumZ5zn5oYFF00ZDKnK62UAhKW0qPiAQO3G6DHXD1bI
0NBnUkUag/BIfUdo4gBTaKTKzX7JQIh5FSUtjYQzwOpp2WDHFD8KYKbFErXBiK3a
+qepeIZvYAc4g6z58bSfXSWVEqY7ja9W/wxrkmg49I96hF4RLzS5VHmhCDtnRfY9
yhMY4S7OOB9xlD5/Nqx905rJtlYMpgJyIIukRHXgsFFspHNLpAeIn7HVGDMtNCFY
S490Z5NK83mS+bvdBk5grD6LdxTiOc548iMoy/L/WKg0ivTgFcNLiPd9iQzhWdVX
KbDesxzQ3eKcn3Hzfx12lB4pbXJ63v/0EGa/h1OmEN8W4OpiToeJALhBrJDx3Y3M
pyHGt+uXOMzE7+bCaVKV+7qWCDLUGxCF5mQH7z/AuVcqoumuVH4dUyPlmXaJQIh6
iZXPi/eYCAf0M68jlg1m/G9UZD6XtwSTb8eWxWAfZwB+N2NqIaWN3RARaO+55LUb
HcnSewNuUFjOGFjQfljXH0XYkkwoU6yWX2+rHfGpdBxpQdSsQJk3zQTS9g3N1wJC
q674Aj9fFMLPpGVCwWl15oZMi4gNWYaI+f/fGcKXPkOGTRAuu+yvuWSOKWHutxHK
OEmeaUgyMYxsCTT5HgZnxavq3GyA5CQ8Ikpk98lSHswADjWKJ7V224sVi6pIGYK3
FlXUeq0vyWZhZ2Jn7CQ7qwCjmJsChGONAhY2KsP8sZl2pG3zKRFKplj6iYVMoUAs
w6tGKvKY2SmZA9Z448blVLCqZgCjk84gg3UcT23m5pS53GKn/oFGPGTldoiQAZTH
ZkguXMm0jFDSrb3mFph+7Xb3AWkPOj5JeYYPZXVYik53nWKVaileYiCNeRG4NYkZ
tEEzIb60A8zN8BYfd4wtN6wn5FbBQRymmkNLtZYdska+Vp3wp2N/qmK/d/vlQ43S
zG9P4UdRAnLQFW6RrXG9HJpDx/rsK0hssH2ZPiPlvombxB4Ayw2k+RbVQkjr8d02
QXe2OHrPo1vN7TkSv358yk9i7plK4yhC26ur4g/uqdbXtGiHC9j8UtUihwlYFzUR
A6nr7WmT2PqJg2TWUwbzNWrtb0FRDdNWOEvRqNp/h3o9eq1IEjdTET7zHBmRu3zp
+CHKw5cZLLvw0b/Et/U5kOsjbKAo7N+U6YD1Mp8He5K6q2VmHFRRAnMXE+dizmFT
2nrWAzWEXAa90BfcxqUWrlhwv3HQJLfzvVmHB5XULmeOTOS3r5EHPz2DCONoZUZY
I3TxTHegtKC5ynrHQKx1NIw3+Ph6Ib/i4CxEhL3+nDNJPbhCuyFwap+O35qNALY+
jGWc9JAayGSBOSjnYVn80lhcO2p+uegao1sgpb/WMCWvi8DDg08iQuJijDIdNCYO
THZSBDlO4Xm73UYDSExuMFI3jnJixpOywkRy6wLAOrbp9RIQl+hQ69cn+wyfhBzg
Tb3EEK2n4tRkX2yhZLmZV01xG+zI4+OTyxc7HYBNkq2P3a8ncx4+trarYBElxVaF
7YoG8FE9jRa6Q3nvnLtBITZ7KfHq/fYoespCvQ4u1EVnjBBQmVDUbAiP7qy2DzKa
tqgjv4eRmXBH939+yeqlbfOEbzT81psYl5zQy07aKRhhuxkhoxJjPpV5HcpvsS3/
goIw1xKYGDAfmeA3xdKbqmZGEtpwUCuGVS/ZADqCVO45iPl0247gHIG95c/pUnsk
0IrP8FPAAb0ljdSLQZznvyvcT5GMd6Wg0UAQubggu5XcCg+y3njyusEsmj9rOy+F
ws+RC8NEtB3Ri2dwl5AsrRh1sMnrrJJyFHo8ltm+UmN19Sb4ELeEF5vt/wAwaFuc
lCWv8kTwXPTJByRxJ+QtliipZpWfIg/N982hsyuN8HX7gUk8D1FYlpkXwDCfznKt
Gr4W/Ax1bKopybLVgLOoU+lCqeLeiHhCD1Ej+X3i7kocpRqY+5VyrX2Lv03ntKNX
EPyTb6x5qZCkYGffxihymARIbZW72GS6AwKrNI3oo/IqPwUQ1XTw0Gef4rsKu269
V6wdsPFylryIDYtaInvS1M+QTjcFxvrUoLFQ3mE6WQG600RnaDTtgf6TmcxAfIS3
txJusViqtxHyfNoDh/SxIgRuGYJjnKfkJTkv9rqGljcawvFw/7yLWjwkpaDOSYAf
R30DBolm9/5bvXI/kW2ehMhRsUfiEwfnUTjgF1ZyEZI+Hk7+YgB5Jt/FPbv+CIL4
t+2LOU573fcCLG23gpB0NdUecrKT/GOYxG0BWaMvm7tYmuYerq1g8npPizX/cZGO
kD/a50cGnvjn4MyYxNH4o4NKN8G32mwEymlmVKU5PMHrWawjYaEPSvb/DGBrby/c
QP80tk+wHcPLQ1EzpngoWVJJQKSUQ1Mj6dFuY4CslziZFHbg4tBOXzuKEvaPfh4E
9sKINtI0owL8+aAjqNUWPP32Qe0Rmz2B/Pj/3Uma/Zf2NWBU4QVmLfy5e7SqWpSd
DqnvyuVd5hAeNREvHrX7CzSW3jCkCvq+RkrJAFtTwpwDOoaCbMAAIHGlIXC+AesF
9oOAkX43UT+XXkyu7mLXjMKWw0JBtL0g7SL5ieO2nsc339eQszCfB8bocwZKyjo3
9dtpYMHyQFtu3dDjdeuqOeF/GtNuNcrizkVqlTY/qncdfBdsvYMHMIHkS89ojcUk
S1dNvS3JIdPJKBh7jucFOySybdmDFeWsEqF6sEdHxs9l49guUVph4C7C+I4Jd/YQ
7Y07Vid+yw33vpqN3wYHgMfr8hGLIKz5NYBnlKqmsh7qPIv/O9eZbZt4gNqEyVb8
IiYdnZQo6M7CAXTeklBHMHAWGVxxkmCvtRkho7uTy+SgruTLkHsbgqAiFCZ+aqUw
NzkwaeU9AMrOiggfdQPSEgFM6DQll9VKcGXjUGUUwOPQ5w8EYE1vOggss3Nl+CZF
a/6oFRwocUbM5k/ekTWRL93PwdQquYu7veF9kn29PWixLsFaKexQTtzQmRAbqE6s
j8Y+BYiKg+Q9Zv6TiCh/d/skWghwuK4iMkE2KkPBNRQg72GYTIE51JhCXjX0xs74
xi1XYA52Yn0shjICJZyEmhEGNLoXHfswRlQqRHNZgSVr/r/0MwrkqRLQZRkv9smp
QHPme4za7iRgkkqNOp7GdfFHrS5Tay7A2NtdkMRzMypswPOtFtWK6Fvb3MuWukLy
c14wiNwtGZEU5OKiaREmXpjaN/+NyZPLgUvyKULkqI9kPG+oE7E3RrqtQsIfux2M
8/kXeoB6MRSHGhVtLafMX8Hs+8KpZaPmFoAp/Km9stSOnSQ+vsC+p5xwI0K0M99G
vxudA/zgho+eSHSy/38L+E44LJA5Tf3C7Ws/4TO/sKZ5avQMQCvxlUI0JZQUpXDk
VcyoPPOkknpaoMNtdHs8RmYB3agT+CEVa2kaYDPgPZFWYRb7zA+dR2V1eW1gvyfw
r8W7dEivOZWVECnc5j4nI/FuPt13czsJiFPfhgrXjeoxYOyYpcDGS7mhFb0Iatb6
7Exb0cmUWX7ISauYYyrCscrJOhAJnK5rdUSTCnqUWKLRMh2jlmJ/sQ7/9aR9uXaP
+r97yBfzYSOt1PEM/XI8ylFsvQVGFEML05v9gNU/shJ4ojSCB5E/k7Bx67T3YMwN
VPAa69X1f3IQfi3nmIBAY4mZS2wnm603qpFE24/XoW39kmKAabWe5mnPFJkMAix2
cVxddTJ1GargBqDmBff9HMnS6U4+EXO87qmDA0TKE0R0flYJcC2m0RGNJfPJRf+a
/WH2qRDTMVjI4xeSX1QbWjFd9eZeE1hv8cJU1kdDkpzuVIMfsBJYd3G9y4n+Dzl4
LEH6ysuvAyT0Y0CvL+s+4xem+QZ+cF16uHQq+Me+uW6bRKTHLXo1cHiT8i2eZ9ve
eyEUdgFdrb0uHLpQ/URXpWK69tToJDt1Mdt9O/FatVb12DjL6xB7BJjks+Lb+kKW
/GpqISIz5rG6zZDEF0pXWqoN4QU+TgzpQ5UWkohSiv2C3dOJD2yJC7gD6BwEVKKl
RlDJW3r+gQ0CIyWxtEJ6SQPgLQw40sUwLpiB4mFDrv9iDzCYrgxDsREyZ8QlLiPe
ALo3xAVUXy3I8LXRaaxpkxBUjj7kfbAoP8V/c1BZfG5O+DvMR8RBL21QVrpBkuml
E0jCMvZv1mLDw1Ww49zxJM3WYQmR+Odxz0iMMCFDYgX7gE7aPEakGBOo5uEkrAuc
byy8k1knXiNxp86GLKmsPDr7P+jWIUioh02SASx9qTZjn/zBA8zFe3WDJL207p/O
G2B2MEFEpwto01SuU9HmQyOCx+tHJuVFrEgBQhRLApDd/5ZBMmev3uPx1iF9s4hM
WHpo3GTDdaeHXtCCcKnCASfy72URFsj422mliLoprgFlOPkVh9h+gQP4zYAoorSS
1Dp5cJK1YQgfDSwrOOD78hyZVvUe2AQypON+zW7GPkUAAHbbDrxxtqR7hXhP/ody
mIss4/NtkCyWEMdxiDP+fMm2lf+Ou0XblDa3J2LEM2NHg5a6ozy+Yz4bfzJCtJrO
GASRGeNcqwDs+hmWdr40610N8QHOkFUAGXVo1d4LIKXC9h2dReZqR25NetJFrSR7
aq3iAEUnWzwcslzFqiQAlr94NHxLSpnhyKHI2oyv2hm7Bsh7wd3fZMVzBNl240ML
a3LPEhApRY2h5SSMIuQQg3q92wUHevTSRDW04QCrUFyURp6v/4zM600EifskBzaY
bWlvrknAdM64q5t9oNZm1IXlykcHw3o0cQhYaGEqZ+Nr6xSQL05w7TZUOGo7TpUl
YYJtZBc5Zq0xxyO3HWRBkiNQ1pewREH81WJlApwmfZdKWApU9ZJGh2tSFPkL5MYo
pPMA0UpMt6FvE8uPZZUkEOO3bnfTAilL7Vhv8qFlAYOpLgqvfEv4Npj4yYwk+nzY
EoiblYPsh4c26Ui2nBVsWYWLjt6TY50A4y2qZEairdZBm3TXWStQTUkthlQtaXhi
klip/79YVy/s+Gq5r/w3p8sCEEnTuIB8w28EbU78TCL32LlydVdmg8+VOrWYsk9U
1oSmrLD31+/0QfsrapJgo0Q0NDBjXmTWHjisYsYgZuDX8FyUuVitrt9jkbAoFRGe
f+YJ8bikdQa37u44qweXVkHrmXqzA0KFpLO9gug9/FAOMeZV3oEVg5VJXQomBZrx
6Wf84YwqA9rH/jF7QcTJZhPXl5FEA9nvQlqxxCPjiF1OZ/Hiea1/oD3r5XkuvDEF
64QmBPfD+GJj1yiBICmDmpWFaLdTLllSIhBk65AJkpPN+OBV6X3a2oNQlwhPpfrB
ntSKgzgY34MSbq09IXb7yJRn0ruJCtjaa901M8CJ5yVefJVJveCFwMexglAasmI8
eEZGNed8d7oj/UwcBMPh387r0CfWRVy0GTibkQkfgVERC/Vsw1kWVAq49CLa1HdH
e+rNJWEfuxN5VDWdxhdo0qBnoH+r4mnG4Ji+K4b+/z/+Ck/A53wt/+jlquVPyETu
1ShX+nIYMvZ1iBRpUbBO4i616U+1t1CiixIdLuJVl5jwJPRKMX+nMBvRJ6keYTxW
naV3uBsy8x668G8eCMeO+TYO9FiG7jgwo/x6egnSTnSjw60+EFx5wRSI8cVQUrvB
m8eBJNuGN2Fns+OAoutN5ZpYRal+M01FzM7ujiw9p0KdGCi0N5NurHbX+rXFUkY6
dKxsQwW03jgLqxkgKPBrgU1pTuHHFZMMMjKDkCxxsuOyoFuL5g/F+IHJM77QSfoC
gcpB3BWcwNwj5bK1eYrTfowJgRRS/fTJlG7pToA57NWinU83mvx0VeEMe3VtpVuh
9YjKFDmlF8zXj7sPQzE3A8TnUmOJ1qtOvJ1AAm3eQSXjs5B76yOffKbwfnTRXiu8
1bOhrGCezR/W/Tnf/Sl4SHYTsRNPScx6Gk8qZoRRCpC0mAXCpjRkLxX5EyDxaJVn
wrKZ7Rm11kIqzMhXFgHc4fsJzRrut+P+mIMTQsrQT/XagfAmJ5M2rm1Q4ggbAlh6
KMW1ngKc9/FPyVC68FyZ3JjIXlZsqvBnOF8KMuLPcZFkzGrfE9no9AI1jdmgpoA0
m+9jn3VTajSM4NtqwlAQVgD2XcnbQO/UA5go4QYmj3+F+umbi0qvP1MFykuLxqSC
CbuzJP7XIOAGXp9xalikC7d8ECgRMSWzNMXhcav2LudeHBWhrq1F5xBLeS3sIQAL
wYvJN03NzPHQ+Wo+7JArpuNDxCwpn423MnE79caPFwIuNdF3IjQLcwpZQqYmRAt9
sNdkNWU9rgJnGLMIP30iyy0Reppw5kTlRZo6OmgyhRUfwuBVedAL84y3yWc1bDVJ
FTQgKvMSO9zb9uklN2fPoTtbfSY2PwVY1CBOF4bK/YU2mmBdsNldf439wwSTfqXY
lWwXfYAYDjBNRudXDoI4KpCYpMi1mOB+bHd8/qAs2C6kMv5XUu3RzeIHqR+BQAtE
mYc6RWdaKGs8YOFCKIgb2oT+bpqPgas104sb8EPkhbdzyJijKAxkqTykLwOYz11N
wN/OKxNXx4ipeaXpxjsbRGyeyMtyeLFHybOMJwDWBbjbmLHQBiw08JPLBLQIB58o
DDmjIf5BhQzi9JyGQ5rz3WEGmsqQ7IhtKw0me4by1EufKgMpKiZPbP1uJUdmS2oN
y+2cFFTOBlb2Qlbissj10Ry5+29tkvTo8wSC7nQteA2/2K2oIyoymAbd8v5RPWCq
lUagvg+kYl8oZnHI8kF972NDrgRG+obI1tYVCWWxT/pI0mWw/CglH0hBhc4jMUqw
D9yWC2TRVv5PsiwqgEZo2Ffw1qjxWqAt9ZitAlPDc/0/JS+VcbNinXWDLr1OLQp8
+JD0mEiexC7VrghGB3m55pbyRNm7Id5sng/58pINv2k7zhjHaCBF1GyinpvA3ZjV
BEwNSQy7V/yGe/ENeK8XLUFj6mXf6gzCvZFGO6okQHflwje64rj6kXUJTR/J33I2
O3HbyZS2cctjRZJziijLarijX3jpFOkISNcJykO3Nku579v0PRVIPgiZwHy84Eyd
NqzL8JYb2N28/MxTy8mrDXcnMoz5+eWhClR7xhiKfgq4V0A5h6Qj8ure0mGGTmN9
X0ZIPo5XxngZMwvutNsAD+sjT6d53CE3FgMmPYrztVEi6JbF7QEakWqDhy0kSDJ2
bmRsq8k0L4fQYYd+M4+wne9QOAmhyvhrrRzM6lI91YA+F/6f+zQHxx5f8cuQLiVr
Cx0kSCUbo8hvPu2D57wTwe3MCkuiLZOwxa88bO+TJzn6GsHptVNqInBwmDkbP3iR
4YQ7bcUNNuc/ix2tJwUNQ6JTY+YSfHTju4wrwreD6vgvm8/QGIEiJEGwGkI/hMI2
XlFFpjI6y3HBEIdAjWqDSgAq0fguerFMIih2Per5lkiQ98/G8dHF4kF3YZl+8l1V
OrEtEEga1kd3Pj4T6OTdzYA6d7+OFUMZPtcW+ICmEoSeN0xUaspP/91s+SZkuZH0
xV/aiQ1MoZD4cqGBGMB0NhBU3aBf4lem7YNGxjTSbrgEnOSZORVFsPc5t879+aIa
O8cQMJC9q+J22QEFww19viDbZDRDhX0+QJopkHviIaH/MRUjryeCgqOLO8cNCWVs
kRdH8eVTbJXStDqMJ/l/AAmuY90czdsRduZYf2Hlgj+N7Lr7i1kOw8+x/hhktVmw
xAf+HcaeBub9lHh1emsHmDkDHx93aORXSBcIK7/eM3kos61/JaU9CqONj01PL+U1
3axVDnXS4UAaqJGwSC5E76yU6LrPOm+e3zCaoWXm8jBnuPNh9vjVgRDnXSCgZSvf
2ZqblXIrQznYftyowB4qvP0pqcgBcGRNhTas88jUdHNNqiOrjuXoTnbzveZX6oVB
NGpv6pVYD5TrBg1xJ/8hHRaC0kdRt7eAQcCK7J3O6QKYjllJxZ2p8ZAuuP+V0HbU
k/uBmVEIrHAnrkFc78Bfk66ZrF98GYG/eMZsxBAYS+9/IAyZIP5wjmglmfsmTo5z
mTxVM8VPNvftah7wgAxwpxSYlPxOVimG5cTD9JPtUNhmsiCDCB0/GwDwiXieFzJE
B/mBn1rV4iPHEo1EfYQA+FQAOxNPkjqA0PsFKmLVxb3hYCq38c4ghD0ivJ5Hdju0
Xoj8bmqxUKsG41ArzEKQ1aANXx71r/pmpzwiKImGCd8FkrOIGPflyiS0e+mzbfb4
fIbphg1800xUwCHQXkVsRSVy82AYtChLQKucCIlaZeFGSKfqjpoDzJ4Q7In7Ch8U
FE1QMtkhCuV/ksl3Apt8h05fjJF87LDZ9kj+9De5kSRr2qn4yiKiIAn2d9MxatOf
PDDbr7ZpmyGpa+lX6tjPeEnTCZDc5W/CyzkCpBV8fp6T1DEpd27M3XP+UtZrSNMg
a5kuw7qsh0VOTBtZzojaQKMvjl3zXhoQSVbsy7F7UhfxRKg3F7mYh+Xj7seOIqkR
oEDi5pX4CG/WaOMB73mJF3omSDICen3op4/qqGK5d/hebCSflgx+S2HHC3F1iEPc
6ELkEtXydZwrTEKH+BPh03LBRREGeZ75f4DpzNDNgTivTeKPLZtSruXLXXocHJON
5QlxYEzxuc9jHKpA3OMMT0tJT8dF9XllseuCKk+qKPB5WUkAX5ZBQsE0q7fwSNVB
qsnUkYy32EVz7DQ7WgXOnxINP8cvxjpss8b0MRv39toCiWV4WKGR/36nt/mK/06S
hJkE5+QuIB5IDq8pvkKj/LIcrihykJ2dn6Frtrje+wKgW0J7xf0KNhfmKdZT0uF+
YKekLlPm5aLa+87xNvNGD38UCUlDcORJ6qX+Ymh7Jtio+ZMF5YOzUHiCl0SKE6F1
caQ5YvwWU0hGuf5mP+VT9AQbo8fJ2O2zzL1BrzHIhQsJg8z2q/+FnNAtU974Z+Ve
byxashQoHR5r9xXRApH7GnTAaE5Xdc4JyWcWKKLi+CCsyFbGdWT10CMQhdVGfh3O
wra52sSf7bzj4HqQO3K7BNRKvnUSBcS8DbQ2FcsVPgKC9qxONjTo4PQpi3tQTKIP
clJ8YwH6AJ56GLpHT5enEfCc0ZJDjdgezzIBKRSowFMpaBAXaYI2UV0GSlmSm1Q8
zjz00VZgtVV7ORWzjniLl5dKpcVYqExQwlCwiojKDFzRh4q6bF1BRvdj19g6UOMn
tSgHpktHGac58/6PVtpvMA6TLQDYhnr5/+ZllIMXdS6VZPBkfdezs7LEUoX3rnmV
gUjDhwFoJUoEJAnLBeo8NM1WCQ4i3b78uYKztMDdUk8xL3S/qzfcliFVPvqMy8HZ
ACx5ic5OTWbFgjQlAvJQnjYfmsTa5s3zQwJbOlado91o/iHx4CguVQe5i6pdoOVb
xQZK+mYlesH2ujI90smi+jmMsWNqyU2+amHDLNNqeB3EdLxdyeMly2nVwNn2fSBf
fr9dvXOwZoO9FgaGv3DFQqAnvJkjYpD9AxSqO+dopfDUYuuP+LN8379XgkWIIvU4
YJOa037JGsOBFTxvNK+4/zT/e/4/NN5hbHeQuy8GPETO8O+317JtNxsRgI1awjV8
pCA7IQtHTnL42gSgrevb+49zSBqaOkwZYka5TSLUeAbxBdJrWjIFny6fInXR8hs0
3y5pkwPH2x1DOEt8cADDuYRylW5lkf8qbu6p1cwhA5DWMco/Dqdzwcj1RHxStzZv
u1dcxo063qiCsqjvuk50mLioTmM+ZqP6IVe1P3o+LaYEYn8B37bEvts5GPIZUD46
wHBLquPx9KaxWX60HmfPS1/KSNskCA586Gwbre2TizdlhWAssXjM828sjFnrXUcm
OW5xSDksqm99HoQtXVX7sf82FzXKcVbH7wF16oFzcNwT2Dj6VUxVFfqhJVL5qsfm
LiAauGFv302V8gavbgueNrgQGdv19ewzaak0Pt9TCo9BEhlGuU+3BY4I9d6qptgZ
wgAkw+1sG5jfxXxfa59LebDkorQjajadYtf6m1zPJbTeVtrm5QQt4fi+qbqsZcEC
I+zHAsbytIx84/l5P4s6K39EwIxFnVR4wW3GC0bTRG3FNULvHteS9uwb0ZCbNa0F
B7pRul7vaPgAFGFtZv8ozKVFALBSyau4VzrF1Y0qnuie4ryTvdeTjrqR29LqSsxT
Lquvy1aWnlQZqf2dzBJkRMHwRDZDAcCudFc0qAhsbenQKGO4kR1dEeAbXDg5GyC2
RwFUR+LH/6rXjmtAIC+ZteFE9WgBlnokwBhXzJ8cM6m87hT+d9Fe+6k/60smjElo
AV32IsCgcJiZE65htaNEFYxSYTZ7kqnYV3V0N6U6WxczZcHtvuQuCFW54tujK4qP
R/dy4sthEmEhN/6hQaEvQJnYsHUy06m3c6iB2uw+bX4VhbK9AUPVVScpLRp8ozZK
L5m6ct+OJZYfwP+6tBL0p/wDiKofmr3Q5KGs36+rlK3bRH5TxsRlSNavTl8bIHAo
p4wS9bzsM6dF1HlsggDxlRtBO2gcR2tfAUUoj5YPYjY4nO/iVOgD63MecYYQY86U
i3Oc5M2KXBc8FBr8iAd0jbjz4iPuhkIgcyu/IUrgEmKR+8CGfSkcdOcMJ50FgvxT
rgtBB5Kjqw7R7f2lhkw4kh3+AcaiLFgzatNjwl+5BNEtoUlEAGv1VprhKSeW+jqU
CO+ZK2AQi1ghWwRFtVxOuWk33IXfgZ2CmWGwnPwr77zwPNM9VT7YURFXPAyXTDwT
/4zze3ea4ndCq1GCMSs6Dg1v6yn3DwdcfLBGlY8Jy/JlyCGAU832X4eW3bd5lTVr
XRkEjBKSBYKBJ7bTAtd8xU/58zlXCyTk3a89VTfykAY4DXO89M4QfrzqgbmMKWY8
/19efaeyo2nM9AJLTRtvQQqOgfo9UWNitHCIi+tEzlfao/WkADt42MQ797jHq89X
CvQbPrYvcI6dO0tcZ24d/rS9ljxRR+TwCWCvoDsCCfNFhA77U+7l2fy+ht2IlUiU
CxaAKKJZLic2u2oDS2M63opsN+Getj7jd2CyM+qGXbyZO9tWO9WB6q5zVsa5KfTU
STCHi4Vr0Z7GOVGRMvMXQMYL8x8iLpxFcoD91i6+GhR9aow5CwqJc8EM3z5eInX4
s0PPuTN+R+oJdKjmpaVv7CMalG/ARu+o5jqPBPGzEb1IUtrHVE/71+SURmrFgKjb
7Jj6eUyS0MUfb+vD2EM55AeQuDd34f0qWCd6rxErCuKP7rcNHVnjR5syoiLfkmJR
VUcnCRitfOMGZNSbzXdAfAUVjp3UCBcGzGvaLVeRBubioXTURXthNKqrF2KX9qGb
oNOcnS9GlPT9y9w/oAqMy43ctbB7g6Eycp9ZAzCyPqD7S2AgtT42TQYOCfHB7oJn
9+BU/LjtPkBqnEeEWMF6R44dBKju4aCOBdBqUoA32GqqEKS+75dZNYCPMzHI2Lwc
aubWBwVzbuy++OM8M3D6I34TW5mvqjpXMewWh0aXQ5hccAEXAZv1y8VJqa9V3uSs
3Ie196t8I9/X1yztsKxLBjExx9V0d1qlmvDK1IbnEApO/ArqbuegrW0UImOzxNVF
4g0R3+BNvKV2N4i4VbqJSt05U27X222fn2kFXo055+lJMpL8VwYXGZe5aXTmV2VP
eieN3WQAM4BGZchXjoQOIcOW4aOYxg4g/sx7pExzylb7++6yN2f2bqjNC6d8ENSL
AjBdPLBqIR1EX8qQCRP0t/Ruwmd9W8YPOahFzV0aJ7qhpGUXR4W3I07wjuFwdE/O
SvXbZyNdJ3PFmBb5Qj36GnYCq7X6kxh5Rsaa2lnzLAcW3R/wHar/3VTKKIrg90Du
Nx6TNHVeklOQl220FWo0ERiRaW1WC/YkJ7NcSrB+FzfoQfDMwieAbWVwNjvxBy+x
b2jhqhZFcZGfln9GnV+a/xcFkVhv246saQg8MktfXXoMNoJBhEhM1joF5AfNMBp1
JExrAgML9JS2WdDi9rLcn8x4jsNkacgoxK0GnCegRWPp/+ysPcFUVv+GU5E0WC/q
V/sJxW7pqWdCg2SYdzqvF9ajg11AcBCWY5qlyImVuMMn6R8bPdui4DvOcrkejzwU
xlM6CaRQkoWWEsQ2HLlElBL4IJKzxX7hSHGKyyimVjEIyqUFeIj4e0uazQ1/VdQ4
Thhf+tBbGAxQ3W80xmqM/pdzgOYzwAvW/a19n7rsiVTdvsF+lrc8TVvdNXuF5DOW
kP2sdHc/xsxMyhiaW3SI+X9xp1Hn+3z5m2mJuM955k5NpFxaozLsookGaTSOn8E1
1alEN0rXktSe4GQZ3NLNJxskQzeANkvb+386ZIfmGhGeU6SyyPjhh5iKoXlwmMnv
hhnjueuNW16uDYj0Fyqrh9pkpr3Fo9bNzXcm1eX6ZY8ssChoAeSmuM5nNQ3/0Dw+
MknibDOlKvVCgbtxcrxnSdXPay7ZWmOs0kgnaF8BN6xl4o7nXCjVGbFz9kF7aOxa
q2MJYk6cl716cQoKzgq3NFmyW7GVNIwBDqwFPwO6jW0iTvKcg3IU6IAR4r94Yyb8
+58+cMqFnfAXK2oMuzqXnooMeP5BGY5FjrhujERPOKBvkrYWaIkmjwwwsryNiTXG
iFjkRywItqfwgVDA++H8tCTMSrPc4TOueXWzMd8S6dF0b6zztpGuUwoPv6iSzM2h
YD6WAMJuMOjxRSXIRlIktPe2JpK+uRVTZeueMJHmOvYBL+O3LeArc/DPdz4bReVk
io6//4ri5U6zfi+bdzfbY8TqmfNI+wCviPD91Ik90FLAjL25Ib6oseauIYtGFmky
y9aRqxpdF2OkU+GvKzix0wFFHHhksJ/rSSbQ0sTR1ddVfWzkw0WMoNIkSvZ/MTZp
AcGa86a7GTXxw/ssw3Mds4aF+y5qt2cVlnTwk1oq7W5k7/WuO5GmS8XG8Grw/gtu
7elrhT6yX7nYNlu8vK8hKYmv6MMByV7D/Bu9+6kJFXcuOsW+ApwyXuoyEs9m2ke0
56DZ4uQmorbEIlrpzV5frG8rkRafXbrKRJYMbA9fsat6x07y2HRFBQlM1X702krF
k9hpsE9ZnVkpFti6tGggBt+vs634dgtOImPKeDfySrTx78l9TkXy4qmyC1slF9TB
2FUyAj5QFaDYMt8FeNUcsRB6VCEa9Fv7FLuzOahxqpnzRiNXC8vhD68scpxQ+knI
VhqCxbOF1r958npASGtNEZzn4JynQGzDb0DhElEvkOa5cDtizl1K9zoi8Wz4UHdE
/LXyKqPgqvaT6diHuacMBO4WdbxYPaHon0kP+E+l6uZySHj8pPhin36Q25d7TDZo
hiHMr0cj7ErzRbMk0JvYSARJJ7xXhRy+IhWypL1uX9UTrAHCl31mJEygzGK7BqrF
5aEjqecde/hb2WkIZS560fAyQhPO+oyfsT8CWSFzMZlkm4BaUQgK+MPIfnsVzyxZ
LeFGf46LhbyqD7J0C79xgUcvL+Tr456wVFW6MQDw2Z5iGRp3qKysvTsJmUeGpMQM
CWy1SVLm1I1zjnIRo+TcojGJUw+xhQf1B4jTVcdcKZ7TD6e4kv5iTuU9/m6nuowb
Jb8cXtPsI8fRcDdYGDk5U1xHxZux9KqSLbUHGBfbgqz0Z2rvqEkrpxm40fYwKQLj
Xx1XbWbXyz1rnN26tYTSisXF97iPbDelmr+6IQGe7J07xqK9fvZ+t0qFynKmjbBN
vFlRBl/xyMOLudHrs8NnNiCbhytlneMisKJPAJ9fVQJI1u+dydV5HfxwQ8lwUfgF
OpvipJoMaZFnRlKk24PYvL6qd8sXhm8xk78DVaYRaMNu7ExjT1g+5BlCQ/F/wyie
8vi4I1zHOFwRT/RJHNN6tOangRwaAFKzkmveC20TaAtIiPv0vrlQri6M9I9YJcwI
RTdEy5y9Gw81RU54gYEtIi/2YiJj7r5pXhFL0R6leyeZT75WAU9g1PZudFWUQEdd
lbHzvIWRrDjMn6UgahpHuPmHYbasG/ZgZlebK9ClIgatStlwAGykuUhHhTWMwdZB
Z4RgMZzvGDG2W3mOoYoKyLe2gG+18rf/XGHd10JaycgmVGts1rcJEAQaMe3fwQAt
jfLQ7wLmclPBwJchAAaSrCC4NHIb1s8z3YcQIMxzBnQ+gzoOy8LjkL1PZW5v1Wy/
Ivu5uExjz47WSvJdFLBjNh6ENFZSgEqIe5LSZ4I2yVy+KsO40vjJB1mPT+GG4RSD
6BHBtMNs9t8r/YNaUm5XLlGv9oFz2I1qbCUnk8oXU9Cjgp/erXBvtLdIvrpPJ9fK
l1wVrKS/UNy7K4jxze/4ktl7tpIaW/GhBIqEOqNpQO8mN1HPCNLCm18Z5ti3jf5N
RCsXd2Er98kz7w1QSDYd9rjIbRjJ2PJHPND6fet50oUlXCs072NER2FWh7cY0c05
Vu1v7AmeDC+zGVNWcoTIlv/O4uaErZFSt0Ug6u9oKOkw/xRriPO7j93y321j5psn
NpIALI2RJofYiiW+YZMOfGrwsx1EuLjUty4eKJjwiW5DGmyk117s6knM5b83ErEE
7tV+UkBaMVJYZa/g0/fRV5KGWiwQOPqCa3La1abLVKVcDe58bkUO6iuov+bgOuFt
sABagSBvWrBW5XrtSdz50dKSkeydBeMH/olPKc0arZOYiGN+gANmTsMAQ307mKL1
/ddpP4yV00cFlAv7vf2O8/sg2dm1xsLt9ARFP5RO4b9bU3VODcvfMtALXM3do+G9
GgEQUPJd6sxIa/vAa38SQAZ4vrNtlSs+skQCllcw7dPwhh5s/BELLz/K1JO+6dNE
On/jI3ZjCbDrZDW7CRMdaf9TcaV2lQJGuqEpa1iONW0uuP09I6RxKgFBy3uAA7g/
zqxpSovjlIZUDTZqdh7wrAaKhNa3uYow73eZqGRWhzDw98m+BdEULMoMgvXq7g8f
gJawb77s4HOWoJve4zLJvYqnu6r+FQxbo2wanAkWt5lfv7JEj23KWNO1BvC0ahm4
V9Qr1HMyfxCcgVc1+1jJwn92YyL6RWnwf7K1upQK1WdaV76dvJgjoWdddkWt6fsO
VYqrFbxtR68hCMy+5Pwy7yKoIE0R/2T4zrZZ+Dxv9BaKxUx8Y81u373TsdpYryl2
EIem3IEYjxf3EB6yiRfcWl99sksSDjgNCASgwdg727SgiXfVnSyiW5Gzop3Qdh8x
NrMutokWUfEtmXHFenTXe/6CZL5IaeavdwA5Ll0vdGhInie/RLvJTUKqcdaagUaE
ztX1WdTlUAU8TaSPMRi3ItrUInwWaaIGQsugdRtKxYXo5nuNd+JpNu3Hjg60QzT3
ReOFPyxZt4fLJOpPdjzbdi/aWoFnf9Lvp8Dy5x84UjAzASabUIlQVsFDSo3rodlI
2Y3E2MLVkzW/SIqVjAtCGSy5M6wuGS45PGw2oSjW+fMziU8yab+uQAR0oISSDlKw
oUYJfZ2fYvTYAJ5iOT/vzUFV1LWOY0JEpU6JKAt/1xw5u/LLMw4MhiMaInc4ICZl
/uHxofbwCTXSb2srQQ2YRpM+BPYhDbR2I9QifotVFsk3MLb6JJE65VZx4j0pWtF+
jEzx1MmqdbkCog9xfsO4pilGhltssnuHGf8+mAeECutrdEjn819MYzTdyb3y+laQ
kYYo6EDsrf5pS4NOkc2OBWvkbW5diiL9xaxURYgJokig+D6D3D+ngqbl0Kxw7M2L
nNZ7MGM+rXU2nrC6z3H9H3BL9CtZ+dtfAUBuncv0tfxVqHLDsFNfxb6yOFUtbGvl
HhmwiKpVdfpGpNYVSgoecgvkAtrZwuZPirbRD4IogGVdOlUFUEZryqmN20xs2M7h
+xamjdTHVzEUdrB6FjUWA2Tf2wxG9ccFwnlWSRxPLVY2k4wlvjF5AhYHqwkfFbAc
fS8jNtY1T/OgzxpfkATJsiPuxpA0czK+NU1f+5rmcCtnBesBkVr3LU8ioBTX4eGD
1+BrWsn9MPx3uyw+IT+So9ugh0Bla8GzY+p09RVhg+l49UX8395wSN/kLuy1qtFc
zdT7L6yxqEL7ruqfW1X4/s9sBHgOc2D7wJY1RVFBZtAPOCJsJUvg868ngi0a7sH3
lpLb/8CbmiM0+fKruz3gg6Lz16I+GSyQwagRqGH+JOrAW5Ww65ELsTP8/7u5Ej4D
eVMd5R3st7q5h8ZOlOFf5tmNSLpnZFm6hQ3SKfFCyMaRKxVqIKYY/g4bYgXc8C0/
Nc2EWw2B4ZR3KbjGGRf/4X2sCNZOZlQzrjzoWV3uOSrXQd2eslFUPbGNnjLlvAGl
dZb1501UDARW2Wfhid2OwEKUxPO4AXNvqhM99U5+2tJkIdPA+CHU1O7TpehUM5nA
qnHACvYZwQJ1CINhNUhNblObsCzRLZx6O+P0pR9fqqVlQy2wVywYM5ODGYuM8skL
V2/8UnhtohhccTK+Ue7CE+3vSaRg1//15YwDoqJvlnFNRv6WxhPaHZmeY1S9xLwG
RaxBlBlQp2y/eWRGdjoDEbKICn1WkQDBnR3WnZryMcU6B0EMGgUmeAttZbsiwLfz
ySNMhQFHpLO0r4ZLDABv0kuKja4/teTMmxEtbw5h4S2dWgivZBRgH0CkJliUrRLB
Qxi8hlLC5iUvHEb03kkF8E/miFbe9myzqbyDiK2ERJqz02iPHqxaSZtyYAfr2zx2
/M9UXizLO5TxNwSfcMOtCqnqfaCzmGR0G3h/ZRLcv+Nf8gacCU1OKrqj9q8SJ1du
ruomS3LUE94THTYQkRTTwULEHAa+OYIMk4GdW+gkq87HBg4dBUNWBosef9VScv2M
iVFfRsgOaMeCWG6uWTcreNiGu9wAxJz/9kjNZd+zQuah2eyDNuobICmVYDX77uI+
0hU8E+U6yuW7SQWiztjwrxy3tejaQm0EwvC6OhbgCi5wDA8NGy5Ldhj8hN/sLkMR
FUj1KspAwBKWlgSd00Grckwfxntm15oZReUvDaapP29zB84DYFfrBZgN6ac2vxoH
8MfhNONmCQhlbqbVlhdGmyuTvHdhNA7mAz9g2ZUcFizGkP0UP6E22U2hHcOFAqyH
yjyaaH+cAHL8WsNv+bMtu2rXzDzfdWzuyud2NWka/LIVvZgIfU3MF16feiNHZHhJ
aBJzLdSyIKo2tkN6k/peP1qgDlgq22PnFlQ9Zcn8KNMtmGA9INDpxYElYZF+09U3
71l1V8qx3bp9b+AoW4iZaeDpeluh2zqL1ChW20hoTUy9M4IuuBKrtZRLAjrrn9u7
fEDgy1okfW5GSoe1gx8qxdlATKJ/OGTDZLV0sfZIM7niiBg8jS1md7362dvNkwGD
G7tfcdvA2Vytq6Kh8sQX00eBTjVSAr8Y1U+KYfJNj+KYhepPt+KitOY71Cj+T8p8
MQRC/vPoQod2p+mcCKskVrc0dx7qkhZZBZshY6OwEjRzx91aQMqdWD9AnZ582n8K
2MkT1R0WDVc8eCDLTsnzbwRZc06s1BybFqR7fiwV5IXwJRL7RZSXJ6BlImmE2w2D
FqHYxQwP7Zx+zuBSADzTHWSuyryGew7rRLwymKIkhI9ZO1j7MHMBG46Qu3A3ImR3
auIQDeu45yJ7Kx6GEY9OBPdpDoYoNv89d8IJqFmarUWq312hbAvoEsi9XB7wix8W
2ASUbm7o7kU4On9ANuwsLUiASMvwwMdEWVWCGxz4oN/tn1ART11GL3jaSmXpdqjC
hKV/7WCEvssRVM0W2YsigtYYXm0ooSOeXW7d4c/xuBm71SC+fAMoxcF+DYNImkdv
bD+Bb4/ZY68jbsTTBFAQxyvVWvKvORO2+fag9spRNn2nIKYAOnr/dpAOSD6Y22Rz
Zagz9onEjYTIIvo16QS8yDOi2kRvtNh2tLayno17xIANwSX0IPt3zMajLKmEkYdr
zWOAdhMclyDDoANHHJTp9V7sZz3Eo+rlO6OmDb8g1m6rqrXLELrcDmmUDtn6Ekm0
RIHDg+3r2C3mN4anLTt7WueQm6G6NRFRTGdaMX7bBTF59xZQXVJgc3cEsoBfQ8jh
iba3K8WcSW4wRrfBj1zr6wBJdU4Mk9D6hj5XSRcMpjzm22t1LHwXhcTIEHRX0Yfy
tqGrE2vj9KSWej5N4N09zSO3RXTYj+nvOdfptvvjoRDldouT0AakBZnouaEMiA0t
lmwVlizphLiE2SyFUGZFwCfGD26iS8EAoBmXVXbl7Kj6UZA/0+sg4Vw+v6KnAaCi
Ix5AZo+P1Pi5qQVMoT8a1lJN1NQ8DCtJ254MZ7O0/NX2AK2qAqN1WLl/BNxgY2kT
NgLR8kHMMZtZKyPcs0Z0JyY6Wyl0UZRq36bNCiyI49nf2X3yca/p+jQQT1DppYpf
PA/HzooErqQMtVAeUbmAqB3fJ9w/Ug+0jDO62ckJXI+ANuJhgVpztn7r1A1EEV/s
Q9LSrJ+TbqPVvWPYvMwaIxXdeVOiz8NTa3dKnFf43VRMDF21QsDcArQiVVtqZmiv
Ut0RZgTUtfXxy6RY7SxmQZ12wXl4eeC/epy5bTDKdmLBdKHhDUPT2kQadS8+1iRr
mbIwKmuV5ab8PzCx+VL0pCEGgrmIr/Psv22FSYEdgaxP2GGbfdiyHf2tlGzcZCFL
6Of02YnkIw+WQpyXTDixrzxDNHiZGmN3i5KrX4F2QPAFeDoXv/AmsIoG9wdBWBBv
Rsaew2sGZDyN/sB+bz+OSjNFrcH8Oh5UH1ca9oVh1a/Ei6+oAk18pNQIuiNQ/6vK
LVUfQCAGlgkvYDuA12uxZ/77Xj6h5b9o/mJCuemKZfS/XHyZfK+KeTIhJPcicM3S
3zM2hVXdsMJ/MMwG0D58P2QMmngOj4+s8SuOEABvA1ocIb/rK7lApElPASqfHYkU
t+1S9MaRkBp/bV3u9BXzMYIKgV9x/WJPED22JYLiVt9knWDeBV6llNy5pmE1euMy
7/jZq5HbRZyJZ0jlvpBXF1JZadgo9LgC3CWGcyYmRPEMNvpsb1O1XV0PiqCR3kbU
wNC/6cl6Rfx/HsWjI6J3Ne1/XgKAEwtZkVI14UPCWlY0W/QAdcfLlh3+i8I6KHGn
ua3kmvHN4jHE1CLNBrRDo5IRpIrddYRHYkgbsvwuqGm6BucBTTTgcumegSg2nnGl
pA6ktbd254T8pQ1fU2sAdAegTABfY3BH0JmSI9cTwntnmuCrpIS5R3wr9VoFVWH1
3p7u5QquB/SvfdI+/Z2YOAYF6kPaTclh784v574P85wsHG1hXlFy51g/jZHPV+nk
40KHTLTKmwAq5Z2tMcFABqIWOFWayCa+KoD+yRyqfDzhxk8LlXu6Tp1f5yh/Iu2Z
3XhDKI6KVIkxqLbiAehBKk8GEx2wCUp3RZE/V4wLbt7TyTAoAXK8tnO6574bNyBj
p2Zv17Odm3ZX0aIJYdtGQ6CiFFcCXtZH5EGps59SRt5x4LTkKwmmLYSeAHLyV474
GE5Wy4jXI+D11/Xt2m13Mt2ZiqhCXCT89iaE2sy7CnXRTq4ZhBj8ok5UxQL4MwuL
k8DdxAHBqvkRmsN1LoveVVqD+uUUgosMbcY4Qowkh9SmZcORedqYqjBvg5smsmvD
YMRU439m1yjTWGILYgH8G3x3eQ9u/JgaEkbLc88ka2wgtHLn1KtEWWTKTzgptAgE
qJnVE2BeN0rPXLabxk1OK41ea3doRC8bgPgclguQTjiViDYoJOxQy4BPb91YgRDL
wz8HlR7xUv3oWRU0jtcPZvl9XFC4fmNiWcuMtmoeQEsM0J0u9jKT5lkeKX8O9uP/
gnvNH9p5+EULsbgJXTyf98nzqI68LEGqIyiTmjbL90JGpyg0ADiu17Onn5nqwP9a
Tojtk2T1GCOlrThQB62mMUYnuXBldjGvP2wKdbQd3PrXdsirYjf3k3A+tfAmwTh4
okBoWx/aNmX7kzOcqjv6EeNUr9bkIQZg1FmYkBhcSzs/aKmFNZpCjogCi1yZ9FSY
eRJkWWaf1PTHuyegKlZWN6WISfrKUm/NWJwp4Yfz0cwH6UWMNphoTJ56Hkd4IFeJ
UGLhxW4j8YmChMKRsGvEQGOzNeCNciHPAMRwgiVOeg4m4GAXJ8umvd8oJDEgp2V0
sp2lFF3UqrQIV+iLQXnMF4QVg/dp1lkQ323UpF/GQPgILPekuD4LRVfx170rLKhq
PfNHZyUCqMbAqEip4j1xDffhrNYCIM7ZiLUNTZTWYNbpTH2YWC5cGSXC6ao3sbVa
7L6jXOWfykwuQOJdH9iAZqSToShFpsXS9iwvCyEjygto0zoBPKhH4esrTcrEwZkk
gcZyjAu20T+KbQgYC0DxU3v1FmekkhhLdnb8JFUXSA1tZL9kM6PhBUvykVVXUSkR
tPAmI/JDeABBSnTWd4GrHzWeUkSKzKOSb/crLoj7g5LeAtklFbEtf+1VXEwGL1lf
kXjtHQVQJa6zI8s1cC/O3KUBcUg6OlbbFzExScIzf3CjUtuhPgZK3+TpJWF9/A6h
WbLe5cF60UOXzSG5wrKjlSp+YSeYKvql4MyahaKzzXx1O9TiqOuZXqYYgqnb7CRO
suvmYDLOeDS56w+arSpTvbOH9WMz1V8el2MQFL8lRiCaRgRK/egbeyNxSyBL+uGX
ISYQVrIFWRrwbiyDPvnn8FUbSzNavjfEnBWlXqvJIg4I+0N75OJa55yNZgpHLzX3
jMcQsp24klGmwZvcVj+IWFYDGLhoNEtIXB53BOi8rcaJf6BtBd/0Jo2DeI4IOG/s
304wcKHz3mlLgkat0t31dkDNULN0WwcbyI6DjjJO5l8y4vvMME4CSXVGk4Ww5U5R
9tTM7X1H+TaTIPzqrYNIMKBEF9GfNGzt6RaQa8XmYUk53zWF6TKRDZMXD8cmdt5V
vZlCfRCB9ulrDfp04a3wxAAC7q9nnGnaw9IJ+W7QQI/Kvu+x1MbEAgeuLLNYpbu2
wQCtWA6zR0b1gop6puXBmLPQaJ/ad7bCAXVBcRD9CtbeYazujBlJ3vbAVI28t1dQ
ZyUwfgPx8V1j7zyKW93nXUOPErv7KP0c9tdw4M5op8Jldg7yvubB6qiekBuMG9Oa
yXmRk/2NxRL4rg/WXbkFIN2WgqdczA/ShcJbUF5FMCpsDtkqUtrDoYSOfCiKfw/I
BKUD1s7Db0QxIog3Iay0H3wSBg5I9eITHEawrNTsMhZiszab7k0yoE+DrCol1Qcd
G30KKbtZYZvvlRgV4NEvMWwmP2Nui/XFx+N+5mB1f+fyh3RcZT6B8Q619bc7Zn58
WdeO9qZK+6B0OgbDsOpUYnGU2MyZH/7JBpGqhG8yTtQupGBwLwQhn9JBQ+70NVlq
k+cdRof60qW0h0VNkqiuBYMFV6G3KVezgN3dVsWtefRRvdQbkRXM/7eheBpceZj5
+KUM5nNGBDkH//ve/OLpQfSRRflVALMjiYMiI/1P6ujWPHioFMC1f44dfEiZ+eEk
/EGHLyuM1g4DSREB+MQdgf2rwmnAGcj0LcGbg3/I48x/smbuVZ2V7JhzVYk2HD9X
FiwhqfcNwqjcTwr85iaUQHbsY03/qFqhVC+9Ta6BSKhTThpUMhS9yGQI4VMnalO4
ThnVQCNs8faAFlF3cT+EhsMFQVwfGatI3DpucoCQrCa/q6cM1qmwB+AzDWKrBazs
bpi4W0NkvTd7q7UrTBV1jN/Ztl+fCTaWwOGnhlKen4BYg2rwfF7ey1/6G0i5BuTF
INkF1vjv2hb7EpxRfu0MkYDAFtPO7TN+8F/erCfIJTydiGrxJciqqCKEyJjRI9WW
K85vk0FUmalYcOKOAL7VlOozV6OuYJ52ODSRcGjWXtejxw3ih1wzphaOQ3DeAhuU
tOYyjKu+B1ysgKYYTZSDCUFbdcZLeJxUmRa9qjZkxzL91rdy+oIa5Kgd46MPtp7V
+YGv3fO/b85JVHxYBrN1OnLee8/OgMSYjLdloveMHPev6xZxKR2XEXOhdWGNlZNg
icGUfsLsLiUnrwn6nPp4hr87EQWUkuZGQXJv9E4W4mgMahPxdZtfpUAaQJn3pPCb
/ixXKqyMTAWAnVqtozr9jb4OUOCMCWhp66bVBjImKz3fYRiw7qNuUeiBqpYXmc4N
Iine5dTSVQkqvIwSE+w69H6l9/mGs0sKg81tDpupEWBodDG3kQVUu/uaFoaja4Tf
wzL4fygngBfZoo6D0uRgOQSmUBZzAznZ1IOF+fqLn4/TUTc20UnIE+10s57LhYlb
r3Nm4SEX+8eJ5NhdT39C7jI7eRg22jQKPmfJAXyHASMQfvT/ZJwq0ED13G+zPTiy
Of945B23DqN87yw1P4YQ0ZdlLW+rAnUKPOMlRjKWL/JuNKweU/OnFxTGVTBn0ckX
DwmZcdrhaHQQm3rctMebyTzPInTf26f4/xRP4eWFoWlfXmI5M7CFYjQJwVyRT1iM
IyvNi1M9TJpFfDkc9i1sOD8QEwFi0WpqdtJ6SlpEz823Za1XBhl90NuqbcjtJp6I
71rIEiPKSa5ysUsltLE98cTDz7YHxMxGUKqAQ0Fi/yvqANJE3QdaS9tgnkSmXNNG
wXqR27gw+z0Bmvy7DUs6t7Cx2fn7elf8f0dxib6exTrpsNrkhnjm78WIy6eGq1ov
f/vVNFR34EGoWhppzgrrMfntJyw6wkGP3m8wGdo7WU4lKgHdgizl2cnQzH2h8Jy9
LBKK/PGKXiIh4PohboDP9ywWplQ40R7KrcK2ul8Y/irN99UW/pu/u5mcUitWp7Nm
bid13bPRRDfqsxlLz8QK6OHwLqfiw8qPMfEoUa+xPnIGKIy/hpEo25UJL7UBjS0Z
lqs8Ml7GZ4pV6gdmnX0JeW05ihUXiGmpU/jav/69RnutN0XS+EcSsnp2bpPeEDEd
5xxH7MKEKcLrD/S6Kp761l3nZq3hCzqkfGrAiqnyVctpRWDvGKcbw/YOeFxonSpD
lLwYY/W911gML3WvqOXMHCuSY24hARlNh2p0x6FQRo1tV3TevgL/sVCgwREUCdyP
/E5V3aCCAyG7UbjyT1Ohe6H8w6lfVSC6n5C008h6sRGkhWh47f8ygPsN9OTvBR3Y
QnSUZanu9ChjYML8dnioMYqdvSLedE7YYBIVLSD1y/VpfHnII3KAB+51h/Tf/ikD
a4vuzh/ilSowcGpn96aM0rLPeb3FJlvs5nNSVjYG+c+1dobn/Onr8hDZBKlnBf34
4Skg4L1oFhhsYwLJqBAeKKgKNLtH9sAY764CdqNKN+jE0nshKtaPmaGN5moqpp98
jorbiBbmxpM46Xxpdf3DViiy2CeqPFxophn8Eb6I+ngENGXoxx3MHagi+dsrw8n7
LemeaQubUKOsStYW9R+hVbXXee7amdtznVD9ZYHET6796GqVMY2y2ehIq2/CU2+D
2+at6fFEXQx1Ptsk08Qu6gB/gr6G2pMf4RuSCk4+aWXF1Zncf+hxVADEy+fGIYSB
Jtshtybg3ZCU9ab3zIB2XjTrXGa8PyTmhcOL4XssuVJ0DTF3B6z5Y+/cbz4+GReX
H2zbFoSL23R+vp2V7qb5RK3yQECJRZMqaDSZQ5idtmPjNSYztzzdnnbr5R5x1mdX
QFvRpG4zTtvtjQQyKXjUGxrneJOKTnHNWHXGbOVPyugdln336i7Eb63u580JBe8E
Go60xsvzs9Iorj864ZCxZ6gDyCFItHLZViOMZO6pN87aD6E2pTeYN/QHwPCrNSXB
Ud4tPf5Q6DUBJJqdSE2satwRzT5q9BzqHftXRnSsX5XA4V8MVv+5bIq2CAoikw0+
SWdlXLJNPUR7zp+3krApovmvkPJZ7LPxU8yJTBC9lute741ISAsepjMtiZfbYcR9
Y/Wu3Cga1WYMbT/DtTnTpTKGn5Z8QtusIKuDaa3oqzIwMhsa6ipHPNwbR78HTiPw
dZlHh8vLFidkFT2S5NWhY4nium5wckWnubQs6J5tfRahwxeFT29mkIO2xl7SzwZ0
zUtLoWb6I3qlhgAqk6UAYZ9zDNmTEvM15n8vDYY0uBt4S2FAEWVEnrOu8xuOA4OK
KI+CQz69RoUViJhnYW9MZkwtjD97x6WCQBS9nVxhcqhqDBnkuqxhl+lxzYp0ZGKc
db/syAUnaBnSBTMmvTZ+ytgoZzeylDNj0NMgWuN6EQGwp1udrdSLYougIUI6WNZv
jeMDSO3ByLgO0exBzjNPVJaUG7ml6lwrk9rn+hbTzHehR1xjGtH6xsPL1SJ7h/t7
fKuqOW8KVwXnhs88Cl9pfnLaTIlt5nE87zWlpo0RbCNM56Kv7QHxMCMSK7kojNav
BcYN/+uFLLloPQriree9oF1z5+OCBOI9YK3mT7/gKzLVpxb7SvfzMwnlmUwTQ0bK
9xM9RAqVXFL8dWZk7ot2dq9MUwGm4jLi1SNTtaI3rOFTZxtFP9rLD1YCs1ygbDhT
4PEmkU8odiHTc09is/GP+FgJyvOU6MgyRgEn4nxdeBRd7PEk6haEewOLPsl/oTq7
qpbV5K6AdG8HJAhZIjeybf3tNbE+ZuKt249iozu+XIL39tPIZSm11bg/Iep3YwrM
ce8h8vZ2dn51pQDutfWG2W3K2WlCInauQ11D1xKHe9qHIgqbEH4EdSggQ0cQKeLY
NmQ6UoYgtic6JCseStWfnDu7TWXmBnub6XNr2vcEVwH/iylAPuv07bSd2e1eY4On
fyboM84ei7OK1zE3eJeYMpblZoBzjEHnDcc7BiLHAZ6aZmRpQiXzHW/K4uipUZKk
Kd7sjHoLTfdXs4duSScHnX5sW2UEln5YimOfUFihKLhJjEv07eNMOYDL8VsInEbk
PE5xZ3EBhk+JasUeI4AyukLyPl+OdONOcOdimefN+W0eaA6IIqIZCR2ZWhgJ3gb1
/pBOAztEW3/jVhNcdUdf/D6LjB28ACC4FPLnGhO3pbQLpLsd3UX5s1O262Acth6N
VDlN3qXN0G8ygH+90NeTmXlaUH0wzTJjeY4oL+NOSx3XZhPTvfG4ANci54f+EmgQ
ZmemB9fdqMOJ8pelu/2h16LV03rGFFvchad8etwDtlYW1cB5mbFY3g5O2GQBD6fa
2Xaz3SlBfo4tY9vUNtS+erSQXjl9mw/GUeiOzPbnKME2WeWgRXQH//1WSwHZArcl
qOzJ57M6bRg6bUFWahKDokQbddOMEVqMwg9vaO+nbIl1xXCTKYm8TqIQv7Oy5FmY
AZS+fiw66APV/0DVls7hvg1u1NgfLJe/zwnFLGn3ETKTkEl1WeHqm/3yQt5IY5eT
oJbt1mFQXluNijIFm3FSVV3yPeYKrczWSSg3+rEEClP7GUsTTu28vDJg/PxqSDKq
keMysShM730i5Jzc03yIss26wBdwDqjECl7m8RBAD6M3FgOA1r5CyIVmThgq6AzZ
eJCvWHEUw/tT/M/bkU7nD/h8en1mfcavI7U/TEzjJQVRac0LlbmpR+v3Wxhya0Sr
ghtr5hr8rajr+qiY6EA62F0dEp6dYhAwCu7labihF/KY/geZQezAnrbMzoA+CinL
FR+movFcDif4SkGVTBP2+CfV85LeKIqa6rUiqxxacmc+Mg9bZlQ1bVvf/V3uyK+V
slXeqW5TkiqXH5g5z91dsZ1Y4mLwI1o4rQUQAK3CslgNO2CPZrecK6TFJxPpbstI
UXmdSouwUY1BZdzbj1Zw+q/ZVWnjRFbIbIsylJ45k0OYQxuWNG0+BQHVSMaVDJM+
3GsUjL7+CMzp+AKSM560jFBHkq69xo9uemjyOjkRD9R4YETnJS/j4+Hvt4oymdLJ
yEFzUDCoiBi9fCCwcddQ+JddwFwtaZdO1lmRGE4qNUltJVrBtqiw6jEWmH9skwqW
sajJnKcryuv03Okl7ira1Ws5SmDJnCo6ITM9LAPTizChFAWuSKeYbd+qBkir9pNc
f+6fbCMWKT0iKq9kdehWYzu2QLKogGk9o0y7VYGVtOyod8Tm3zsCXstZYK/VWp6E
5Wn7MHimopQQs/Yttna1HO12snctaT5aTOv2BZ3Xm80pA8l9dyq96SdoioM4B1Sy
nkwyE6jg5V3g1H+XQk7FdogxErWCStWEVX3Kly9NieT9+P5yrbI7122Apv1nY0U+
tI7Bj5c4MxhuB1Q9Gd4EwzwUs0/NqRljp01CBYhRIsLyuyPulbscvKWkXrZHFxqe
MMYAS11FUQMDrBzmScOZeas/XuEN1lGAUt2NY8kaArNVdj1BhobeUgX5MjnOaS02
LF6FLuLqEOkd0aC+oFGcsRpesdhxgm06I7/I/P7VgAKj51eeMdBZS3QGhRry3+0c
UAFFB4GInk/Q1bSdWOam704P4ZEM9UJUeCHE9pw7Ziwf8LdhI9kUh0Ob3aYu21kC
/8jLKK93zQPUJxg4tauk4IuA3bx5DxdIYxkRYnYKjWiDDxHrsOqDCJ1IZH9MWflf
C+fDOc/YfHkuwuZmE2Jrqtwm+x8JemRz2xJ4y2MHfGwUksleGaZjXYjLMzYOUzwL
DLFfkd0Y2btXhgRUkISjC0G4Ksoi0ptIvkjYOFbzYXqegDLSWcWQy0lGxsCcMesW
eYmzzrw2P+t5qbU+FdcRHG3P7qBgrfuuAnCk7dxXJtBgpeGQ6C/iFpY6X6LSjhju
Xp/CHCqJo/iol9qdpTn0QMmkAiSJrgqlFCllSNKeRrLDe5bEP78gVsLbWLxSxm3G
Aq7lESjDa/TPUs5BK4i/LWGXMgxgPEoZ7o4+d89jnY4PC+vVaHhvotY0D+DTykzz
qxG3tsWXJvBHZZqTUop0dlf8wS4NbpvLaFVhk7G+CwIByeuFN+qeN4Mhht933x0Z
/L9EMsgij4NIE+KAiIfdA2OmrVCzv7ZRc9q797yDmjcLqOPxZUnBAg5k6c/V43b/
q1hKSgx/4K+psOlr77UgQYnCilSbqrlleBrEgZ/bwMoPjMFI/u4Y1ccGa47a/drN
N+BblL4VjEgS8tZOmrQGpGVB7+V2tvsHRHIuoX2tLVcdyc61BmIRk9JZYy2+qqMj
ROltf0NjQ6eIrnqgngiOH4cQMIXGw8U+/xDgNs3uwBp7G50YdN8ABhm2CsT9mZgs
pXTU8IBS0K0mStgGdLFgRF+D21gYzeDGvULNC/xo6fTnSjI/5AxtIuiNgo8lDJqE
mhU9KOe+w7WwJQkc6cu0wWx51HhGqkrBS1vHIFjguye0bNBl3Cp58IvCIFKD5zN9
dZQ3elKc8SO3O6ZTgGM8Xsk4M9fpf328J3p4ew+s00Fybv/qi+/zBjwrLC9IDQSL
D1E96YvDF1Z6S1NdQkELeCfpj7ATBo90+/ay2Q4s9xX/x+msbSdJ0F500fuouAIn
kQNvaqImw/jzSTWfxV5wWCGDwkKreMgAff1iq+Onap4yLmGgF5OXaQ8WIFWIT8tr
/am62wkLRyqcAYgDWOLjoducwCQLHQL9Y570dB9YnHt00LPAlt7OVREOr/PA9mY9
sNK94vRP9ibyDGlm9ht7bSXzzJx/b7t+fW9Qd0YXlv4aFxsGR69FbDT6xdcTpedb
7Cn7dt7yR5Hs6euh2YvA9S8zCLU4KcMmrSup5QIwhACXi4JMl2gBq5YyT9MX8ruc
/VaFmu6pWEQRHeGDZ8nGzIbhu75pvufqJnjJycV+Z8UNPjfQz9tdbzxCWRpUuv3s
MQGCZYOg6pndX7hiVBroNsAPWrD+GH3GQBQS3J6h6ErXFpsSDCHvOc59JJt8QfJi
oZb4NI6W0P85qPMLKxX/4zlpQaUINadWCIlHLZS/57DhOTx0Lz4hADv19ZOHPElk
50KuSh23X6zIp+Xp7urTn0Fc7AL3u4B8R654hK7u41If+KK29iR1PJY2rKly1t6q
Q/5zOWRo6sO6TE2Yc7+tNIXbtmNua0Om73FDpJcPZEW1LoCPAHCF85GnpkpsJRCn
MJR+X4Ft1LGUtSAmwZH/aygnxIrnSzlJcjbkT9oud4MwIyLHun4thtXFIq1aj3za
qdeRGDfAYvKOPKA+k9iRopIxgZ3YDVoABECJ5LlYbpR2ueeoGv4Y2SSNGnIjo9ZN
shhkxYBF4b/aMDjp8qKERSJpK0pkPeXFDkI+sd2vizBdUl9BgfA+8j5UdOBWuaw/
9oA8mTHAfOG235qIXb81F+2MG186dtD2XyqK44liOs7ng+hiJ5Ajb5C6/bOlg863
a5rGfyIMC/e9/QyPh9qfs9AblTVO/vGkj/bZNZifVj7MOiTwIHKGF5Hl1iQ39Nvz
iKHbX6Zm3aQdP3nhHMBqS76aqIfJi/aP1CO44liqNS5J+9B+TviE9Rh9rpqLUyKv
yebTIWhENd6MRldwrkemp5MqCHdLE9UWqqcngIyF1J+4UFPChURDsE9aXchOi1XT
wmkH0wx8T9UjFzaxqpKd96RlhV9iZRLdt/jvLZS8mbZglWsD41PokzCsj/SBrjxe
Ix9mgGZyaPWO+20wP0h25eCmMebscfm+AUlCNfK9tPWVlmntm1u/eSiuhT2t4kbS
O469JcJsWDcHE6pBXja52QrBzquUY/nREvVAQPwiD2v+hl8nlloxyaBeVElzojv8
tM1ThqJDfq9bQGfzni+ISTQJdSKbW9GLwfq5SXfdA43S37yDPIzhGOVNqbdB7GVB
HhRq/KYIfY87TTgj2Zhabt0O6JjH8VWZxjVJUAWuJYzMSP2t47bmOyyd7yHjW6mk
75N05VytKKCwFRZS//iURmgz5RKSeMbCBEojsRzcIGyLt+kZSXvNMRuk2tpm9vx7
POyzGMrMDDZQxZwhQ2qw15fNnaYfvPs2vP4/na9y5fj6p7FSgegV2T69o3TW4bwt
sB0rRnxmj7hshxua8tcTVLo6ECvHVkEYu5YI5rcHBNZ49PV8OzHxPVPs5mDf9KhM
tXAoZ2McscR5YE9sIkeXwWz7Bme/aHVVO0OMaZYQpTyY/zy/ZN8fO+9AH11KfGd5
++yGSBHLz5nesGwN8qqreo74NKuuZ+g5EHfKtYqCOSShp+q0okwfx0OEmcNBo2zp
kDHyiMfMRQ5K3Z1RLjcvlXq40e15ChYoVic+1/+oiGsmVi9Jp+hvBOIER2I8RvhA
gEGkO7ptLtrl/WL9EMEH6nxS37CJ8LsryNGltq4VhNwrOcpyYrhbT6ZuwbuoJM2+
jNlXmhyFyBLeqF1I6GvB+KoPBhiHghb1IyGFnrMJSlkXzaxjPo1krRyXyPKyqEeX
/SzkymGx+e+6T3BouT69ohkPfNO9BqCk6aF2//rllIQgjmF8cET+vPND6JGEciTr
ga1fse+McC43HKZXHKhUES7HWFjBF63Mi52e/PN/mt9s4r7VnEvEmRTsmKzqfShE
B8U3NYfzfJ8sS2gBAS86IPOtDxMEIK5O0+s8sAJAlyxdWgqq06QKHBrLTrHrRvF7
WGKndpTssOk/T50jY07/NJiBAQMjyXU3TTlYs8Ww/jPjxohBsahPChmNi0xRhnaE
tggLjr+8GWq4K2mnSYXJOUwErzkfp5AwFTb9IR5ONMSj41VK38Pq1QEqC865f45u
Kdo45RsHcMprud7soneJbVUVMpzd9mB2b1V8ggMhM2D5vBDVjmjnkxis8+xiFzHQ
Beh4WVUzsRcNnjp6IUbwVq4n4Ai7d9/zMFI//WAvTp+FzynR2SbQ1awQ1Oye3YHv
8LzSwHITJVlIU4pNwHxjrflS3mlAeyIEG/V1ko4rDcMVLcrKxfI8vThcp0h3/eFO
NbLUA8cH59jNNv8GBNnlWeGHLE1XNewLJGN+aZDrVce1dc2gtvZCxdXmsmmp5T2Y
5t7EakXwIbD3i3EcS+rycdXslWlcsmmba0ZZu38rVz0xMrGeHRwg8/JE5AqFoKRE
UgWrnjkavKpyxT6dOTNKwL7jAOC50hZg9ZeX9Bb9emy3AOaIntYBrn8tOueWLGL8
tv43H83SMmoc84JuFnVeqGlHjSTyiW89LpxDsTJnkd0/gsFkFUQEoylpDPWfjKc/
dMbY5ycjbNl0ataIbvZpEZdnWPlHnWIOlG/vGA9DpB928g01Qmj87t0Uh4KaiGOM
DowxJ6beLQKiw7TQ+WfN/YBJpWTBGQQTcWG2CBaPFuk0ZFLwtVp1fzNVo99T0aAT
fzK5TV5LxiP8wEPJ5xNtwsFzKlGtQAs5BzcGyAB3CGf2vc6oxC+2R9vzjc2yO3oh
i5uqiUPT98U51u9EsLwNIEfnzDFwc0IlOqvGhgBfPxJYNzSN0leDTKsMKNATatJL
HjZRqf4tOaKHVp+WgOo74NihEnbbaNxXuk/LFsV4jOzriVMGodhd3Iz5M96J6jJM
j/x6o+/BwPat6UUXBtHuEgyPsIEQCJgzMaE0xxMEVExLZ/8zUuBMNIGXCjo5B/z6
JjqEIaCrmu7m2VMZiz0txl9UsC0lmYBWPzd3+0CnHa3z5QtiMk7yPXfd+QkUQDxS
Ysnu2bxK8xfGFiSHrkD/QWqioPXaP2qQyOy4QGjEG+n4sUkfsfCLc+Tg53fUJ2Ex
aQ9BOAXIyIyJL6fjWlWTtU6GBeDHQAgxQBbzDRzE00vyerkMlXIhnWCn+tuKmbri
QBrNRxivqpwVkcIgG8xiam0fXddnEHMN5eipD0jQb3MWYSE/8GJfsQCPwr5fPuXQ
JByl8jLpSR01F9VIa88ee4iG4HyJi7QeByRL+zW5+N00k+kFK/1f7oxJzjpoxgHG
nzp9whXShkbUihVXQdRvXXgMXcGrRECPqfz8Pe4XADlFTqulOUi2gtogT5tdSw0Z
tUkBUMGPbhH00Drd8g0lfCyiHS7tPhQKZMuBL1hMZLHqjgyqaPOv9oQ9G/L/023/
zQ7xA6ZR21OZqlMax9JOS1E8VMESb1b1bBOMrBZ09IAByvLwrmyjV0sKa5Fcfu4j
Mx2/ptCTu4WVR2g4qKjgHdJgAI0L5rblEIAK5AZUL+HvJfmJDFSmk6F8jQA7K/Ns
zJWa8NbiaSyaUxdk0Iibkq+A2hu6QJPLu9w4RkfASyc=
`pragma protect end_protected
