`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YspWv/IEzD3F5EyU1gMp+O5aHQOa75U6G8lMwI7E5X1pJjauO0VTcFLZIopE2mfs
c4w+ME9QjGnQ9kOlKt7hBnf0Xkyc4OqZ/Emf3LKXhMS0jAFXmVplB/KMABkYftOb
h/gcCGQgqKjpsqGnLmLizCHaI7YXrRnlMPzdObjmStY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9552)
2BBob0hd5/u8Dm1hxJgm98c1jQKsDUxJneUfMw/GsXBcsp79DUfm6pYaZATrl+/e
ZIlW2cc3N0Kh+MaVE+HiJ/4LR6cGhjN20Kaha9IUYfRmhGKWFFvC6/AzygdxCxUP
0CzpOYGfdV+SrarAa1+0UfDan2tKZWJIUp3p2pAMn0QEcIeQUFx/WyQrqZCoykmA
iYdSD1meereLtsCcNlpqsxE+EaY8XGo9lyqJajXU5bJSoHwJp3Jf95qEpw2XItki
A89hvSjfUMBLcnkaRsCCug1/3OfRhnHJ21x6twcuoDiNQd91RfBZvjBlapOv8LAd
+t8E/PIzSHDW6BVmQ6WvTtDzH+06W9FGVPK14h/FlAabOJTlODviDYnMthov35KV
JO0rlSxOCVPnNo4okrsh0xkxrNjaLIEVFJ5ua/pG1/XfSHDN7+z226PLsYTq5BJG
y2FbmhLuwwdXLlC/8DmJONZe22XjBQj9hmACHPTWYcC0ffmE7y4zTKnnuIK9Y96m
RzzjDMMl2jsJD+P/ePCYusAJ73kAz04xL6f/5MP95CqWVdTMYRvBC2esQC0F2MwG
hhxWhStoKBvdRlb+BpBDwTVUZlq06owIhVs1ClDgqsIEwaHgv7dMC9PHE5ufYwoc
LJL+7MWR08GAhPUftueBRFfaJo0GoVDtyiTvAHXa4/imHc/cFoXCnKKJCNp3OKiR
uVbhfok9pQG/7mX5P3WzgV3uUYSP16UDYtHErMzZcJAM0TkfriE8ImxDR8X7ahrJ
Z4GjDUOfNC5w4fD5Ke0NoT8hlOvC6IkyU6i6LZyM7f4NZpHm4tlrP4EvKNWlDJOC
roQFsEt2fmIasKfmIO8x/CnI9sRvmlmQOS6tBdqm3SwbdMjyTm9oM3ac/1lkEZri
GmKeZYgwfJQbff0wCe9tGCa8ceJI7A4BDkPLvRTnMSrO010uAM2nFlK1/a9f2UH6
APicvXK/XGjNNlNM12RLvhMfJW7DtrHjuhFpif/vylR+3d03BjmJRvePqnSr9iLM
N+juohCeAV+tNcdHbsW3RGsvsnOMmRnluhNU0iywFWBc5NjzctjQJv5YKaO1qQVv
T0WLtFeau6hIpTrVCvhoVQDaac0E2mJ6TjInNCeV4NnUJl6yc+BkFyKshf5FaKyD
/sxy2CfP8guzzTQeX5bQFw6yXjH01CeLWNkuXweLGEPx3i48TwiEtaoZ8+o811hL
xVvvk8poSYnFK76brpZmW3VU0lkyL4ZvGlWbG01u94CmCQOe7Y2U/dc5Ev/Ymz22
mB8lV9Gs0RRrGvS4CsJNquqVn95vTG+vkt146jPeYasR5qHzBgdgJZCLKsl9a98b
pRDxRilB4FD9aFAN1k+54bxcx9QdMzMF6zNecd+btT6CeuXn6helP4jTpxr52eMv
1wLjN6I9XLpyPR8gjdolvd6p4mlW7UikXatF7D3Oc55KXoHKX+R96YKqDpKvqYA0
KnAE+qq5NU7m7J/5pFllknGt+5hwR5EfQMH7ZdIK/uZMyHplGpBWDCsa+rQ5YaXp
dBQ2WSaSzUa7XVJtrfAZUd1A9YsWvNLroSQnPKH9DMOyBjdwgTelK7jiQhgxALRu
37G35sMk0TECG+vtrGzkwLjAQ2o8RC5LQH0SgAfR0NdyE0bTVceobO0znslKt/w+
Qm8OCOMlv+Yd7PtCVDyGcI4mnWYMs7fUEdHxw3K0utUPk3bced+yCJ1nLBhSvR+L
EqOorJRz+rdW0p9gp+Eu1uIu3pvWHJtnJrghau6GGJpuTCRdUPVk4m0jHZVHpYyT
XxbZ64naYmY5Ajd1caksQuODuj7Cx27a1aG888HvMCasC4yGij5Vcy92tUaYKSPa
lZOotDsEt11aTSVBiyoKdVD6wMJ76iWSfAXPiEuwsopm5e6u4Vy9nV906YfhxEw4
+FT8yGKwh9oOeGXnAg0CNB+m1fWAZuQxwehK2PtB4ga0Q7Weg61CfXSlxeq9YyHp
tHAgrTq3PxlNv+zfy3RI+2Iqq7YzP7wv1kO5Y03aGSjFA+orlnRxYC+d/jvBTkNa
sGQ67N3m1kdxjHaC9xHfIKp4lOKe7e6lsB4feywMpLvOceiv/ZZ42rwcU09L2yjH
no9Uq1uS9AF9HL+kZo1PQkON6nyyyFP8ey3Ydftr8SNnL39IJGqfSreLYveUf0Qg
zAhPYX0fH7O2MslEt1J4dvYw34sg9AA98MiXp38ZMY0/lurgBuqqB/Jnt7s3Su0M
FH8x5Xj94fhtUiqR138ls/mL0n9lUiJIAmo8HSlEFvnmCangC+PEfr6Snh5ui6ot
ov8zGWZBOKANagXSoLdPbHupUXE+YEjanAhBGNUZfN490Lzoj51ycaoxmIrYNSQS
AzgQwiaeFMPZf48taT5nEc3ZASHiR12Uu75JA5NrXV4KR45FS7Bvuo+qiZVv7RZ8
ynGUtfYM9yiwK1l8nRRhCXBbQ0+AEbaXUOb6b0qELPqLEQ+TP4KDsJCemTmYuYyc
JhsI3A/ccxvLkiv29LPG5rxqk2VBWfKdTK7wVrsdoXZFsravIBoXpzW7ushi4tGj
aQtN1GNjSbxuxoyDPkxLTxBO8tmmgOKYWlA45Qn5vMXKMbkJEru4nrTgGx+xE3FZ
yyqShXuK3N6bXv8/ZyxBe4GyyoAQjMiMfSU1ForotCS3k6rdqxpeaUm+bAktFt5i
N0M9rLVXma20y2gnbZnTwWdNzHsZO6hxqq8Huy6vRwYpra4KUfEXo9uibfwFGnYX
savaEhh804kwYojdaUSZei5XLtuXKzeTWvjeIdTwH0eI/2+kqdVlhiGI91ruVb/G
lzFtSEzAMAptZg5kvqsk5D47oa2AeYFfrwrSdV/awdXPOLI5Z3epun/ELJRqFP3G
zX4SSM5SnrMPQRacCabgh2GAmzmFWdg8rg8usgqnsSILPH6N4LMNfPS7U1vStOdG
yOAQd4iDlZLWNd5acYG15h3Ce/pbqwRvUQKlr86TiQNsI9i3gnsr55C/so5gEh9j
yfkGb61XhhJicXMZnYig7VbQz9mMa/5ScLZBP+uFK5cUTvGZevOdcQa/pHDNGtKY
/ZYoDqN+LKSeEZ3BJSsJjSQiw53TMKbdGiegjyxoAmhEY0ch8AEkH1Sxo4l7PQje
5jZXz5ZCtbmI/Da9JuSiVmEx2nxNvEWC3Vr28NM5ZA9quVVoeqgVQDj+pM9Zloj0
BTSY4BtUDZs/hYypgxSvj60uj2eWmozEFK3tasokkJj1Ut6zRKRmipa2mN+Blw6A
FXMlF2wXgLrgozGtsxZJs3LQZPAvx7VKSxTyENIwpPZEsz9cXFECFhDyMbA0j+XG
cq0Ic98RrPuGi8JKNxn5JDWF/4b6ydnn++LEn/HdeN+WtFoXRvS7gLsDXPpABKPt
ySqAxj2yQcsM+/SouXnb5mauTBsHdV6YrQRRIbUKpoL60eiNeMMUc3jRlf3Q2S0Y
PAflg+8wZkvW1IDSh8OFuUtFikFKAkit0XR6gmEhU3LNu56pl2t+t0bs0ifNX2fM
MKSGp+U0tdrTvscwQtwPWWc0jka0EaEEp3o2JrLewXKM2LY9Ov7TlJmhVFn3hDYR
/5a8CO+tIbMeiK6+c6ffIjLSRAemnIw4Z3hXJ4/ACUDpvusEBE84kM1kF2sE6o8H
2rbMtHHXB4LXrIKJL+0SGMitU3oLQ/Z6iRkWTF5j2ZF4q5in1IAshOxv0OPUxOY9
riTlzOQh0PzujowgBYS0fAA9Pcygxghwf+bSYKTa4TTOTm6Oitg250O7ClSEjp3e
W4RwA4FZZ0WKIcfTbxD1T4XvK4In8LwGH1EePuXIuUKyLjoCvsfzfLx9RWQLsFsm
zJEG/WkYbsDAdAHtop3pztmoR/RCBSKP1tpVzwwSwyWBT2oI6wgygVzGjaG1KLqD
AIt36nanYpZRiXNokGAQBzvtVJQ3ug6guyt5GhhlUo297wlyq80ok035EQRPPefP
63ZQufYbSu1zA/JKQ4lfEnvFoBhuQ/abmc2uFcCQ1vVA6VwSAWgrZvtxESxI07hy
zOgwlooIx7eALIvHWHOAPwElGqyEyva5dq7n4fXuIXMAs+6S1tyu+cefZTvcLNA3
S9s92dTM4EXXGtBlz4z0bqnFsGELj4VPkgHbzP18Qdr3HkM6iWZSth93dCIpJQmd
tJOUGGuVuPm17IW+jrWeytdOCYkAUE4+85WhLVcCMSou80dRizrughmzXlP2eMSB
fIIgm49sGxmVjK0Uva+1ZPltj2nL94KBk/P9sbRT0js6pxWeMIn+2ZJOH/9Xid3O
P556T0v6piRVYa2YGsqnnTVBqIRcI4cjt9lfMSDGdfC+wI7tCb+ykQAATF/SDOln
M3wvOmQ+3X+E6E0u0GoGM472iBTl751/OkWmoceIo0fLuqbvS1z0QKFixKqmVkby
erTSO7fid76O2rtGWHFSTa9ETHxGfDzJtCO1xGim81UEk7hgogyaZoRJBye9yuS6
5WrT1s6RtMhcx6Kd5x7+t/oSvc62/Evbr7xg4ar/eH3zzAjUfMIxfEVbvxcSWkUS
nI3+l338ZgW2pxj/VfHaQbBL65TML18rzwM6Stq/3O1AHjVVX65n6DQAMCBoXrzY
s5yQFV2wP153dJ96AhWzPpfzYRbaJG9NR6X7Cbxl2LKcORoXcJ0QYBgILz3RIwsH
w40r3EBJmkhn6sGyS+D/343jcQm9xmDiVY9YvM3f21oPPbsmoFHQkxU33/LhoUJQ
7X4W+rZcvdcElGe6Zwo5mOu1ISkOX3XQyZRulh7e0T1jQY//g5Avn2bqQ8wKtvQc
TQDCPESCvhrIaBGHjeaiOKVoFEwgGzwPyLLT9RBqmdjmPTb5rGKWEwktVwi8PIu+
7Mb7M5WHd6xVD9G9OL772BiPA6eHfagBZdrjetUnHG5PwpPzqfjk20JnTPl+g/AC
wW2tt6jjQZk3tMzFgnCmJO/+0KJ6lk+D5/hYSXNMiS8Xfo+06KRKnMIzkmijyGgA
auknIPIt2zrwEhBNe6FPWvDgXiFhjJ5MR9sS0LLwmWKqbv2chcyKkm/w7Un0bk0O
B/3an5phAPYGjav/HmiarJtMgkwhgB2u3JuFQ9w3MaUJIWwBOex0HFyJ8cBo38YO
rp8rnzbbZoGtKesZt8oq/TvUblgNxFcqIsydcbC0U8/05cFrFbFGb/74oxLAS9lD
ZYEBK+u+XKX3IVbAKekACOhS05uNI3vqKr3zICnhe55In9vbYV16M3S0f3sckstz
wfULcrwUlh7ggfUCS0GAHlQpZxs/90visq3AvcJAzH1xcaTxg2HVWQuYN28yMwks
NeH2hdy8ni5AphhZujGl8S+hDmHAiWCyEtQr/S1EmTP4UYMd+hbwQyi1FOgSvjqO
V96gNY49k8kOjveY1Ewb0DfaB3QnE/C/Rbv4yOF8LwgBUThRvzV8Xjm3ijZoNV4Y
h+Icb/sH9ohz6YfRGps3lK5zCMQ+0K+NGEU3P2OVXAge2B5HE+LV2YT2AWRRmAcA
f3n/4ZPlrTQiT1Lx+o3Y3BX3G6fK5hohvuG1ZjwDqcRuM4vLp1bfhC+TyrTaPp91
R9YSRydoXpOTvAx1HidgOQloByWk2YT3XqHxs6GS049nVhYD0FECrL0Eb1C/0f6M
7GnlGJTyar5DGgDyzRgImCfRdCYjYffalKwYVV69GJ/0Ek6vofj8FV6zWPxh7U/S
i9I0Re/+VdcjoWm8H0hSB6QLGNPlI2Xco/X36Ysg2bwihduz+PqJ5agT/mMDUdPy
yukogVw1KyHw+lOtXF6JiM119LyNBWS+RO6rrxQFYXloQb6bbavQGSefeFXRMc8C
8yFumKbEbtHpap0PslfKslvWygBKJU4jF3hj/YVUt30mCeWwUbOu+PbxLZobweXK
L26q0BiYK92aV0LF525dwdnBr8E/nI5A/lOMio4+qkTcv1f9YlP/FFAPMHXZ6G16
usjvIh19qjx/UJbGDkGW64fIBgIhlqJ5QPqlR+oiaQhkiV4xOfLG/49Iz0bOrB4V
LV1BsY7b8oij6wfkjljT1DsR2KLLdFVHgf/u5apu8prwxXE2c76BETLNozb2r0bs
tbbO6GE12nf0KWT/UZl4uRM4186Po6QLKTbu1KoEwxOeryyrWIBx87oI3PXBo5u9
2ffaXXTh1esjGFB4snohlvE5BoKQ/i9mAES5Qlyerjt9kbeqqiAFNfye4OUpek3W
WdNarnyyJzJFlLQF3cnpHt9RYAEeQ7zOpSo8KGeIyGgC5DGhTnmTjSnft4pDc+vD
cr615gqNuiq40DW7lPxMa07pTfvAbxBhoXT2Fda+rsrUSRVj5fmPcnBui4pdrNoY
DHLbsOqLj3S5jOWgCflqRXE9KIHe4q+MbjN2UAj2xT3vzJJLlv5So4t1ZeKxongZ
myWVjhJ7dEG4aKyH8U4vfbklUTuAWXIVr1/KrTNmZN9PKczWTdzK/uXeuOOEHr2m
2dkVGitz7n7TK8YlxUBAhv65/X6Ooz6ELSlabBCsVRx7TKoKcGW5htPgpEXfoxUL
wguJp+vYcRmB39Njqq/IOxIn+TnG8iSf+WK+kfqkvgV6l2geCO7TCDChntX2ml59
dPtTe+CuSaQqtB4RH21A7yiiQ/Q/p0flrbBsxwq+GYvKX+aBXy8iicNepDs4WHqV
Zqk1QtX2MV5l3dz0hLfHClBlwT12gdsBXu6haM9l3d0sIH4sXo1cH5V8I69gsTHq
r3W+fVQOVvvJfq7BW+egZ2v11yly8wE3+VwYwadwyrUFuCVs1RZKvX0/jYd1wE57
8/TYAOnPxQFcg/Bx7JXwfB9cOceN2ZXI2jsvTegQpMcKat0apuvQcBJnZW1pUdNM
FWrbp0c4O2V9xJIvjg+daKDca9IbTU/st9/UZxyCHrAoUS90aVxNtyVAkn4ZWnjF
6ENZtY2gJiIfTnTaVTMs40RqefCM5bpp99PsTWRVxzpy8iytM0ufbC8M4l8zaNcf
OUNnYOCrpE/Y/sKYFvaWjrKUcXUGSVLSjpvY8prCMcuNrUVpqT9ADNLDsJX2k9EN
6ZIHlW4KYO4JUjLnldOashOwU2itSGlnw54dyQ/u7Pz3142MXsmsm5UyEGnhLkn0
3HCbuoCCH6B3EeqJyUr+hBR9rTgdQ1+mwnocoRZyln/5DO6Kz0w3biu0RIUzK/rJ
6Ok9WqH+YO07+2i2EZoco8ARQjH9HRlDh0JKJ41c3Owfj1yR3mCIbIjIXa3fVMsD
5RxWazbMe/dxPK3H+Ijkksddu+lrwjgF5vTsikcFE4Kr0ocv8R9Jx1CpdtOwvKXC
W2QMbAwJ49yjVaO9YFRzteoQWSsUBWIsMQp9MI1ZzEyMddTjRcW+g2KsUdgUxstQ
FFgjs9NNTc8/d88XycsI/lGyT7M0gfNJ9DE6lRomAPwkpOFZhsjVZ6UtCHnERF9Q
ciFRU40WWVjkXayYFL1vVwm7AaMo5QfJkUSUIMO5Hh7j0PT6csB7MYcgGOK054gm
PTeVm7BNHizv0TUgV3U+STpH8pgqTpjnMAs9OwbP1QEVWj4lsKFGsUPOol0wrYYH
E44CHy/PHkPYm9Mn2LYfO+6AWEFbfcbXwrqtJT+MZH5Hwhk0U1X0xniBM0hyc8r4
/3SXvOOT3LIfH4bCi19cSGPMdBbpg8FFPLQtV0NfTtBRqVdurVVLuib2u8fFKqSt
j9Xj3fkFWoKK3/uXpL/iXTwX14Bew9GwmMjqW7R8zKCxG8E9t85zAioU3m8d41OJ
+PckymQFLiINoHpAT6+Qf1sJ5x1CI34wJzStslCvao+quqI+9/7TVHuSpIlY0Jk4
w2y9OaREdZkWsMa6F35iQ2MTF1BDc+Dftug+tgEoB7AHCbarK40qwBqTF+fhp8D8
QChZmMg8H6rKv6TLHBytPT5twTguzjwFPUi+gW6HcmLeYbzA3LPgmfIJi84z2/ht
Sbskxc/rDoxeekQ1c5k5Qevqirr6a4Aqx/QmDFvhjtnauEBGia2rHOWo9p/74g7R
9JT9+Jb9YAoPPXKqX1X7zUz+FGCiAG7KNQLvdN2F+7i0ztNhjfaNFBIUDUB9cteT
ZLI28jMax78O3OgZw3UXP7YH3GWL+B19Il+3GA/mLCsjLX2se8mXQJ3fu84eICkz
cMi3ggYbitW532gIwRWavAetFpYw19KR1Xug7iXPAY6l5B1EXPUxmnJ6baCGUgWI
vn1vCw8A3iaCyjmeqtnfl1sbSJgobe+AsSvFbdpj7CctnjqxRrK6QoCw3IaVoo4Y
UcOLIsYn56zNBn9HjoBMHWtz9IPssmVun5/iebxuTpZzWugBNZ5SB9P16ABMDfzf
N0KNW0Eu2PK2Vv6ZGbrpKBk66/vLqdIE+g86NLqQnxCWGIB5tEh4ABCVkvk0eHfi
mVvLgqT5KaG+8mjQMZysdKJFbhE9KtWzTJ2bJyzBXL0Hrhnc8P2JbxCnM5L++LO8
IJlwvzTXDOw/InLraJ5UsQPh4QJ4VC6ZyLw23oBA7IxHOPR+DCkhB3cK51M0egGg
0bWxcKkAD9/KNKk3QntDmiMjVMPPBkMvWjkyQz+lohWLhVyalbuGOe36TWisJN1I
6uLwDMuo6IFbXvW5kR8ETMLmFw7SHev9LgklDCA5xfALT+zBADQMSize/W+Uik80
NM0cOSCdH7rgVt7oJGOOpzPib3TlWPPRAe87ZgCXBUgiuLoTzfYbya/CLadSgaSF
cRjnG5DkZ7d0dTJnzDSCaPnHqmPJ0ICRCM5NAd7pxCO35hAkeB/sghaELnn+uikZ
REF0wPbO6ZmCZ3Qdu6HiWiUqE78J17C2mLHMMxSdmzdj00OqIxGcvFcWx7kcJ/vC
CZAMamokkgk2xDAZPIxCweakCCZ/u7NNgAcHjXmqVK96t6dNYTAz6q/J9QXb9SgY
1cuUWjpMRlXV9ELqvWSr6IrfJAWmgx+YSxC7hX4zgFfYUv1uUTIeSAwemlMHwPDK
SYOdWKRud6B7DkF57mMV0ixr6vfcrHrAQHQN1wmub/bCLM3d9ws8A5OmX2x7PrW7
p2HjDfoQKKY/rd5qbH9Yl+YEZAuR9MqxFkO+Q12GGOWKCY6TAD0IFFfIdy7XiNF6
+BUzw0AAh4NA/js+0Md/lJiRSb1OJUdb9O5o9sXb4ZnTNcC/Ya7SawjgouHIFKra
+S3LQscpRkdy4NUkXWnCltXaDYBMiEqAwcNVxp65Ly4/0wVzfxtYpd3BHcb95lgj
cbHKlk+lCKZUJnSIMXMmcwjSfNX1t9MD2cJpBmwfV+oaVjP3gh3o5WKSbyHvCiSd
25vVka5Qf5LaBrtz1Ki8xpuznVokjXkdgI3fDAF9Q5jJ+AajRtbCJsFdJZH/LIwR
szM47Zyf8HS/PUXrHDZEufXDh6o3HLMFQQwrNjx16+1u9+s2srwjFfKWYHVY2QsC
cBtV5dhUYbUC82/U5qloNVAoPPi82kFBJPhqN2xaF/w/w/lf/5uA8mW3F32RzgPF
dRTEeV9g4O83b5yGo7TClroWmmlvOelnzygvzIZBNTAlxPnXDT+wXrh6xEat1R3X
ABCMe4w9FISdXC4h3eWP2wnHSJZp9GMKO4mlduqFoJEBXIJIoRxBBG/ld498eGxu
f4VHzrB2fAlqnibdA+idBgfWN2crqqQrVQQ60O37osRdjYSjLZlT+6E4gZdNum4f
H3jk3/Czl6pJe88b0yfGToqIhqP9YjS01bBlO7T7+sR1SZ+bmjEWlygxiaBu4mdP
klOCa1uLn3PkhfqulzY+uqn0QbXeicrds0yOq56rRIwf9CjSs2C/i6kv7JJ7FVig
EF9qdsR/opgplD++3ATWfmJp59R6YUQ6COic5ZJN3rpGwvDi/f7dabPJKrr5Gdl0
qKeFBLNQdAyZjrv10D8MPJ/Vakhzc2oUBOu2B0E1jKHzltY0K/vL/ZC4E2bcbDTz
K193uQ6/TkgKyA0wrcIxKltmrW3jYre/dWDXPMub4T1mV9TKugtEuYNex6mmtGV/
oeW9roGnC66eaT5JZbSFV6yOfpX7ZzQIzKL504aelwgyjnjvxVtawXC1TqP7sdjQ
5nROxiB8f3xNyCi8drQolaG2hrimMp79RMfQGE7r9KdvWPxdDcVlvRViTanZQfHl
O1immMccDQqTEG8a/7KsSjXh61wSjV4sBErivF5QebAkthUYPYO9fvEjzOwr3I+L
1qfMDU4Pq/QwlQAiA6mhvPJGVR2NoeZyjqRNTjBUIWWhTyx8SzQrXbhYoSLCAmv6
AiR9lbTjkxBPlQHQ0MMvnNlvvipd8Qhml4Rkd9H5PdTecUDDKLrg5IYp+eSKbbM4
Gf4H+XoSy0YGpDXtQxdnwGMnvht5y4YfVpjg6znUVHjrCcjyHi0al39XO6Y57xLd
pmoPi3aC4HxJ0qOhmsG9J0HedjkrTa8UqkQzRXRfu5nXlRJQKTZhWnlNpNkurW8G
KU+0dUcBPqy6zSRs6h3mNFyr+DUudjFLpw8Qmzf69XpWkCLSEwTm1n1qWWRJVLkC
NC1sgKRJWT+DL0WUrY860mL8ViYwjJ2tVXPLaMEenOXIImHzF6kAkh+i4ZA64DTX
3Bd+YOYZmhXdEluzrNHYsMBPxGUwghzuqoRg+nVcfyGNTLZqpsOnZjeyeEKD0kP/
36wZnYi5WLPhDpQtmZAcWkC0M17mOkWVzNDy6PqcHonMMdhlpePBY6/Wza91SxLE
D7XKVPonJ0aJv+wVf6sMB3wbExU4GoP/Kf1tKNTiLbx2LcEXO1p9pzYJsB/8gslJ
+mntensmkR83iwmqKlSBhArY8OxwI7BH1uO6Xez1n9RR3H0kMLD6L1NivRZFx89K
Eu73yWQ0iCXgKbKMegglA37lMNJj+7pyX3rr9G8V9u1u7JEJFx9KZdL3p7Z/jslF
48lRYMHdBIV8vQzojYcm3o/5t57nQQag5dBaPz1HKQN+hynGMWc6Q53KIRt3VC9t
z6XM0mk6mL8DGeqTxcpGeNEwq6SIHkMtWOHH/J20ZsrxOZ7LZhfi2Ja4r3aB1oMf
PBtQMqONZabGYaKkEnxtEOeFuOKvShQ+Lj1eWz6IGmp2zCtJGtf3zyQvXIDeZzIV
aahpGWpF7EoFxN+8SwVPrVpuLsb0svK3nqLYttfMf43pdSeM1GgscoM6Bz2pe6q/
xe/Br/I/Qxtxe/9fcIl/uW/WSHx8FcuKzeQfxAGlTx5U/9m50+2m0AB/C2/WGalx
aF27XOh8pJzYMe+RfqVBh7LXXzX+WToAdk8GeOTzceu0QEqIvZyOFjRJcf6JeD0/
wY3ky5rgFXp0Y1EIhvVtw8DyWABGn4ZvrXTZvmcLvkrsaZx2j4M1FvSHG35GGX/Z
KZJFht5sG4dJmYSTBjctm4LchzQTAdS1FP6xF185f5+EEJERN6escRtkCk0KI/Xf
CFKnxE8OOThB1ED9eHAjFV+RisYTrMgZkf2fg/OftfDSZxwq0FunfaYEq2ZXggKE
eoK0rehChvEgIyyUY36cdF1Q8qnE8p3AG7j3gNeiJ7QAhzZDKf2Recjl7E1pfJOC
QitG+Rha2Q2/56MmHxNda2nMPW2dbtoOguiYx5YkXvKhEye5WrNfDOHSFsNM92f7
xtt+Y0pkMlksK1dk+So56if3UmihUxLNXtHIms1rrpyCvdFd+Mz4SgqHv+7MB8+N
d7tkbbj4Ec7f1OyQaddgKKe/Gu6w3PD6ysL4D7OF1Yz52mcqRdLWNpWmM2dgQFu5
j4RfIwRUEJ2nGCfWzX/sBqGsJ+E68W8Q9XQBY6FEyThLLYxMNGeDQVScpjkeRkiG
Ih687obdcX9oDv8MlM/3sYEJufNF3RUtMGuBUAo4XQcmYN3WrsZUi7m02Tm0flyb
nFqb84+mtHix049mLYawUyLwTi7dqMiFH46nKadQs6zEHsUPyi9TNzXzVqIlJFGS
K8R0HgKc3HAWEmIoHbAmIqEAOgYEG9o9T3j83U5W6pnyqxT+7RgPnXAdhI+NQE8E
LUJz8vnyTsnemK9+VUW9KPxWHHsbWsnUQv6wg4c3DPXeSiJlF+1zUb7HWd8E/omw
YkG+A4N0oaq7PWqs4L6TneMF+AXL83Urrk4OczxOfw7V5EtmuKsrVgH00khsSDXC
vf9w69RmuBVD7j650gfilOudomn9kvBgWs5c2lTF6MCtSlHZTN25QxGaAiyZITWl
ZBMBCWDF0+Oim/zSUghFSV9h1l3XJd8GZZN1JRLPLT8XE2PuQ/N79uv7ni1YxMR7
Ipjb086Vhk5jGHPAqVltVQBDjpCyI98G+XCBq3V40jm5dTcvfwyXVp/NfwzL2VF8
FCf35T0I38fZRpVnLs46zQlIUv2oUOp9P4iyYQPULFLtBWm9lWLPrbY4nTv14/IK
1aG/+bUh2eIHusHmxUYaqoigrGqDjAnerJi7pBxQB3HTqh41/lE/p/x4SnXz2BLt
5+eObFJILz9LooXyeiy03cU5LXFFxGsReBL7oOShXjkhI82dPTWBhcW0C6/w/NaL
p2hBvoKLdqq7/a8uQ9ZEEdtZyFx4ND7goNzp2PSOj0XioE/NH4drHiXLR1GK6oKU
ayznZN+cA3iLp3vTdInzSovGQFFpPcGwXAZBZUHp2NvoyvNFN5iLun/qey1Ucur4
Q1L3tEoY2403jswhNvyVLbPXqrs4MwHMuYS/bqiUYfk5tXtU0+rvMPU2U/ygt7ru
w4MajfP6+VGU92kvgF3kaKUe/ZiRJYmaD8fpumf0A01XdkP/Bx43WfqTp3Fa9k8A
`pragma protect end_protected
