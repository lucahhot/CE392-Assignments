`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jtDhL+WOyAtTYaVG2Iz/q9WJYymRjXahga73IZdeKbhOYHPgwyHXPqaGwd+Gm8BR
7U4usu+jhujHrMJcXQXpHQ92dXnSNqBRfNcQcI0zkBwm+ZWU3YIN1FG26jN6u5cJ
ogqDrJrMLGR6QsSjp3SE/NEGB6Cm8AyFCAC9Pi7YHzE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 54112)
VeOyZe5U42MjGnxLNMphshH0bPw8/q5FfaLqRZmPNQYyLX5E3OZD+YKyIW4AUIvY
SKyEtf7NkdIWvWPp7xPcsa5BcZGxT72d5TETCqeEaKVZZbnddUNRMKwtXepZ0U6r
c6nTsHLljHtVsDjaJM7bmr34r2+IeexOp8iLlvx66J9V0Lz8vMTDbUcHo0nLZQto
wAGx6hN49OXxlFM6TGoFh3PuyM3Ji0CSeFNc9VO4bL6EKF+etxaQ1IN24OQk8PEL
mA0/EyxfL/I+/v37/ajCDBNItfa8repf96Wki9gTUhvuYzqYO2WkGy318GWKwSYz
kKfxo9OgiSXVsiZIAFEwhtkbaWY1R4Jf3pujNKmXe7kBp+THkznYUoE1Mr9dbNqX
nXRFjhxJpQ58bkRavk7jyeYfA5C9QszzCRNEuD38SPB/tX+EhhcTfKPYKgn9O8pM
QUMltaF1eXOGkYCncJ2YKcFGiRTJzpsAmlBP0IWP8HC/ekZ+mcPlVFc8gtuMH3Wm
FomXGUt1UUo2sjvhLoBTIc2Oz5m+N9hfI+7ec5thMzpGka9Y8NWPAfOprphYtKGi
DAKO1gNiaXNPtnUXBWaDM2CpBunKvKF2BIxpGatTHa8UGBgzquqjq+vOv/PzyLON
7pj5fbd/VMxqtAhB/m3cQKFKFZ5pJUwRppcyw1tDBBS5RLd1crQ71q/L2xGta2BA
HWZEtlO/2nTsWGFeDT+QSlNzK0ZJ8vEQWgiPNlJwQ6KwL89XN6cMaKJtJhwA71tw
Dq2KRW/mcfi6U8U5WbX9Ka8SkqhoAwG/U1aKLODmJOt13/ymgVhHFuZApS4eFQde
MsghdEhN1i7r9rLoW3DYxk3cDUMxQH3XGhM5jRn/H20bEPGePKCSnFMVOmtPePLj
OY8wn5K4FcZU/IJnhQlbEFRSoVJCDBdwNotWbkkhlI7P4/Gyg/fr09zBYOS8A2RL
EUhRLL0ytBnHM281y1yN0RFd0MoPQW9Z6Feh27NCmKNtRASB4JJ1jUj1n88SBDVE
yZRi1rASZ66Z9hsQkd759feC5AEDk04JBr+49dQdseFBEtuJ7jKjh0dDwOJrVCNy
JN/2B2T0xnNcqeuPySYF25gm4CqOo5t7xm7Mja5R1Cbt/eA23Ij//GaCNSofwm2h
IekIfdVDspQQXKpmIcvmxFjCpQvoVchhiO6+k+WB44NZx0uYf3ZDUpjbHMPfb7LD
V6+NHbf5FtO0nWuh3kq8/jk7Bw4S1U+XtxmuWFvqmhCTEreBAH63bsT4gXB+K2LC
ofUUQBJnvHezLDvvU1cFkhtrxWuHWtksbZvGqftLik72VubIXBACNXrvtENmzUZj
srboUyltZLLha9Ef8cq7DuhWl0JJtcxmfP8RZdDM9tM+qiiYpziMY5vSiUK7vfKm
jM7p2jf1L7IWSDewgHgBTkOipEbgVv7C1K5voJeRM9ahmgyLzqbJRqfz/x+bpvGT
AlkUO3+fBoLXUyCRtJpzwNC9RFmociWtqG11av2idiQqBvEYvOlTPrHaxGrQwqFw
ElsAnCbtYPdlRQLtMSprJuWlHQ7TN/AXXxx3PzuW8R32ieIWLmLpJsGdGQlWTjmK
wSe5ACcfYw1HxTMe/hYIm33Sf97ILHsI8zEexqFjrO6p98cxhq3Krd+FHJPw7Std
fdj2C96kSkW3ErsjAaGrRyh/15fBN1cRS7fELYkjKpolrJ0/zLq1687VrLYAouOZ
SNwqtQ20JHFH0QQdiLFQ/+N+wvM6zkPGT/gJ3NboPJjOrsENwlViCf0S76G4GuQB
A3l0aheKDfNsiQqqmOOCtbrPQqeqfY82IOhQ6f+Xyl/qIVnfhgKKi7ez9p46Lb09
YLDaUm09Bvsxo4Jy+1WozeEx0XwcQ1pFl8ds/49UYZ80nU1G5/QFxm/nL0hWexMU
AncdSPmeVd0ydUCGYcXFLmsTk4nNOUCPlQXu1Aak1O+6Sd8skGnOLHWo2QIQ4jjA
XF5FpHyW/hK73n8FWhoTIzP5IerNlSqdp9qkpOFdW1YEMEBVJIeubUP6EIb+EOgt
yJAtA5/kCzpMwXgl5eRm35nRRspF8I8wl450dAZbEXiyUZjfEBuwwAtqftZb3UKJ
snHLBEKO5k/vEir8KTrEWeA2oNoUcIwZflG5DyakmsJc1CNKfwBGuJnybp+Lttnm
ZOu3WE7wVg3kgQvcIweLeiaaCB3jSq/s/yiagEIbsLJ0+FoTz6CiruPw+JL78Lg9
jBiOcJEdqhGs4nC3LU0h0WZKd1koC9yMlHa6HOKXx8APhagYYFsd8Hw15UcfjqiH
JV7vquewsi8K+en+7eQmiHd8TROGCGwebD0UXNQEzWNL2IzJQ2qDBxGViOlIWZMo
l3j9i/E32Y1hqVbAbAOlLCcUepAgFxcDK0E+h8MWyXE8rR8ONVKuluPeRPK2pclV
2kJdeihMyUuCiUKpVLJfjx5VetwR06YhUAkFee5ZNZ4LaTX7+ju/Kvh7LfzI7dL8
dV51iFpdYP6rnUI78uYcXF5DdKE5z617zyCERPlNAtZsmDLs+CVYvOHIcEyMJ6lG
i6JtYoG6Vz7JEEGza7wz/VAF1ip3/8ssIzKg1QFv8xG/dL1otsJ5mDG7wgx1y5rO
gqiamR9QETbkZgcCABl06l2SbYirU32BkX/jsxP2+cjbdftqTp234rbAkSK3+MU5
kV0OsztNQvU7wU1DpKT5kQ01fPrz9Lx5M44MgFAlE2rtKykAscyX06g00psXc4Ga
TPTk504/pCn0zsbnNkkaDOQPEfU4HKRZWnNruGxFgKNNgL2TOLrdR64ez1htLchL
qyfB8CH3WzXbiGX08zmQclqwMvm9p1sDbgu7QilRHTim9BgKWHR8TlRF77NQSObO
I7RwDv73nkN0ZhP9k+P34twDHNL1VTGtg4JhkzllWCPcXFsrfwzJtIPZji7MMD46
xZItD7TUecBKotj9Ix3x3WpPHtjoGm8vA38l16P2Rxd4kx1bN9JoohQtFu9+myC4
etm/O6BTXUJgiq5uukJBONfoD3avbGjmwyPCSX3WkiDp87SotLi/GhGK6hPp3nbT
P+SCsuaW4ZPx9BbW4DfL9eoa7qzbdqg6xEkZQATq5L1JA1eDuWV84EO96quTKZDZ
Cqhitkw/y8MvQYOsdFM7z2Z4RRst/CC5X63gfCQA7Ewus+k+4lJdm0loNbPYbpTk
2B+nyMjIbjRNUkezzDVa0xVLLH7y8YLA1a6wQ594aOSfhQV8pn/xqkA7G9MUGgOK
fNF/C/RJ7CsBjQSc7t48cA7m8uzbqfH+lBf2lB8As0zGG9eZqsnLfrrJp2LbHZ5a
eNNBW89WSmnOO+NYh7sfGEJIOuJifzMUkNmvxSpkXPrRYk176igXL0H5RMamQQvK
knfhf/jVZuwzHmSvtqHPqnjuQEKfds3J5J7CmMTi377Nq9bcNAM8QUPIxv1mjIne
TsUBkS2zZ+gAQBOB/c3f4qUUuTlbrWNrO4NP27wP/Cl3Pa0UXEhkx46/BQ/oo+FJ
C0Uni14s/KqVz+0slCga9QyQsvBq5QATpkg+H4ODUzcbqYh+S9Vprwgjx0ZWmiHm
Qau1N+j04mSXU6eM++nEaET/ozQtwo0wwhntaQYd/R+JDGq08Uwl2YFvfkGROwg4
g/U2FzWx5gsqyx6/50MOwL2xpEL8AaSA16Ufdiu8fJlGbuotn7ey6ihFFg57Y6rt
TP/I4U1VicdxZUjnqlu6Ucd41rEVyT6ClrEJ2NYhesoWQpkklVPnktTGMibutbVu
ieiSaNB42W2M/ECGanbzJNtMI0li+HdOysBd0Bh6sD1qhdXHyxWbgAXgG4jRU9eD
nfphrwG9IeVRZSo6tTtdLkKpoofogH8Ky571AKgluYqR0lXz0j/BFN+2tqfbAKTa
q7e7VKEt9tJJl88CrPpvhecDLKTo6l/psOS4aqT72e+fuP8FGPTBW2M2LPLwjORF
iUt+UEbnUu1cqWOrJ//yyc6a3cCLVdc1GlDpkW/d4vWmc6hKeDFxnPApAYuqbLWQ
fR6lI+k5tFm6ziHAa7wvlREBbr2xBu++j5jbVBnBf0IVXucZZEID02p6g1mpbxzJ
D8rFx+YGXHGWnsh9SRWfEHwY5H2QEimBXvRJPtm7jq8iSLizZiz5CwId2zyMIXte
24KQP489+FK83M7dIHt2mITiXi2ahiFYqEmkEGIyXZJkzXONhVaktwcTgCpBPb+k
oMsQuR5gCD1bJGjbvDN0bISbrwc4TjPrqjjkb4RjkUREUT0+hmmjUtdgmarygCnP
C6frDnAjqPKunCY3x6H2lCHapF83EOxZ8xtgvriqQst8zfUuwDJhXnYs8D+xamVx
WoKELcpSxGfqMhMKXJfNw4c8mGG7gJz+atFuNoqWzRqn5hV4+sNvE5Q5ZjcllKrx
uh1fhRAaH1gC5sTFP6aK41XP35Zm06pZ58eLwVXN8HIKct0G3Faxa0zFjHHwgc0m
rauqXBMmHYPsl3FgMVlRnb18Mnzeo4sVTvUNzDcdBAPldSljux5cvmC4EpuDHex6
5lWV2hJEblnWEvuWI3D+RrwDpVvRtMP6EIkCzah1uMY4kIHlG/00fcDdgBXSufpO
RCGicyv/7xOejn8Tnu2XWwfcLtULfHRmlx1J/x0zhoFyLM2baOLRlOEJXWEkWlbc
qqg+NS5V4PWAA+3aKzFTKstVrgU0V/dmXAna3zEoMlvfIifWqPb9UYc0b3rGkrXJ
694WxAXR+qE8bmeNhm+dSps8Bokdpm7fgeq4/DROX6q/WnjSatuxJhHCxc/jy2Rl
OiJt1/UX2Uqc7c3HtMRmbBnISKvlyTplc+ZVADu0QAFHhSoR3lq761r7QVyxIcMd
fk40KNR55RVF9H686gRWHn7rsS2U9OhOWJrJrMM/lgNF8qh88k/JpIttHiOmBrVs
ezMDv6fKjMvJB1o4lYeGSa7Q4m49GUKMnh5+Nb1j/2hPf8LEd3ATw60/GiRztzOE
HBz9E1+wvms8QeSbapf9WYkcMUmti02aVhCyKuousyoce5vPeEUtrJlpfsHh2Bzt
adIIpKaBE1Kdg/H/J5jul4gflD43SKI7/6UqrvH4t4BGjFuaoH0CzrjuQpAKSIzF
Kl5SxrGIbIXPQ1fMR4fn6LXj5ng5v/YpH9zTmPbrBQ1CtGgDgZ0UQcyMvyEebObg
w2i+TdUMYiMYrhni+Xr3cKclEYUrsffQxI+S2W7d6U94TwfTC1W8YERpn2OEIptK
x+Lo7/MQuPyY0NGdFxxRHinZZF4rrKbvZVL3jeCO3Z4pG4PMou7/42xo0B0FM4T9
jmXySn6Aj6FbiQYLC9zYFhTqgnBAwe+Wy6N2Qr4MzQLnpxGgv5n5JLGVnbQRkoh/
t4najUSDRX7OA4EEV2ugMi+jUpcJl0MYTCXF6nSkfcKTzHq8PdVgFffz7IPo29wZ
341beyInpIbexK8dCuHZEvzfE7WlQjB66/X/X4tGwljsjcKgmRb3g0Rzf3+/Hm1g
TWf471ucaPE5nPrT77uVsOaYL0BrWdec6ndoylaPOUkWoG8Wsoh7wJwlCYTgxZD+
WGCeY05iT92dLoIL6cM7IBcv7D3XKvI98vBHxp4hm+pgfMHYBJcmIqqwA4aNpIUv
Z6kY1GaoeFHqbWJwkEAfrWQKHbHNS4ztu0OgdTKR1OZuz7V5gAScuVQlrs2KqmNy
HoXc7TjPJSHLZsmO1Z3iWE3aMUWeqtWhN3WlIviuhbGy9vafCMfu3wHOL3jpQv8z
rnEvb2ZQ021vLymHLeelId5HB6WPVGCGIbMoryzg3Qk/brnpjpkNsO1iea0cBPc7
dcehr7qvioFJcP4yyI0i/cz/2tdFZZfgh0y/zFOcs+UoAAEItk3vkQPXJZ0JHZuQ
+GfiEoe2dAUum6AMMHgunFrbYRjTCdbT9TKEAeT/l0pp2PNqu6GpiO0D2vFcyXzh
0I5q5HQXbD5Emyd9VD2IibDZIg+jMA+7ouVij6ENzba+METTaYvjxXYxQX8j+WHt
dLTilSRCCdQAY8mueu/QCBmOML7zxgmNXSpFo/8BCMvdmBtKAX9yPkIbgrrTYag2
UXS3Idko+6PcwgUqu8h0kLVONvvmKu/0RyAL8OW2V/dzpToXO8x9FP9Bo65i8Djr
yj9v2UyGQXPhxI5IMDnUWg6D4rMJ8jG3sEukqjJaWWtPf+mokp+mKDrQeq8Fw1tB
BWP7akeqeUYcYKzJkVZLNPZI1aDITDwveOVX4h5PUGlo+iY5e6cmoXPEjiRnZ/tG
seWpR2cdyUu0v1tIRuG1nIBg1vVQC9T4iN92tqvsbg+5gV/B0zuGOAVgiaO44Yyn
Ug4b/hcZsYlGcwRExJ2sSFdJa/jXWsuiWgXiWean9+37e7FkV58bsVgPkaULJL0A
O0konvX55mpVcWGjcMDSiJ8lnAOCb/q3ZqnPvcKM8JFMoDzY29m764czQwkyhOJr
4H4Ols2BswMcczAPF/77429f/yZOOEt5Rt02bW75b7mazx83YnYSSaKm2rbfJcqM
KpZIm4bnBq5DEj1U9ih0b8C1uMD2zTub7rUKNAc9fSFb0wu3LYBEZusazKYaeXUP
LLkoGjib10CXr+61MQP28jglC6zv14e5McdKKEeV3yRtVZ8ErgroDUPwdPfYdgS1
q6wA8hC84aPTdoaw4pP0JPY0wzBhjgwKs92eSUX9s5cZnMGjLHm7Jrt1+4rPot9H
NLWvEVWdYA5arfYBzc5djmpcfQ6OpCE5HhgzMd+lX3wPcrZLeBQGkr7BPPU0xHWE
/ownX6Z0k5KQW/LDgGeSkgeYKmjgc550FpVsm5yCVNH1xhfg6EJ89GABsgYYA1BF
2n/ZFeOBiP09QQtu6viTgIVEjd+QXAqtj6veVCc4UmVPh5DzKxMOKZoE4y0vrDaV
//R7yhkueNubeGer73Gg+ALIA/C9FLhKHKJp4tsD0z9qUJyxKSGjd+bVqXTRVDrt
8eEnFVRfj+FeL3L78vqai+7hP7sWrzw/HV7oIUvNhn1ro9m+EGc/O0tGQy0ICcFI
SqLnm1bYID3YSSEbo3zWQIcdgoCdZYu0n2uAJGRHISrRwsPCp2M9N0Va5K1zivCg
my27tSuv2m5xKkhUMcsAGL+f96QYU75ClVaE7MBqmrQ1nthi5ldEbUI2YmaEWgeO
U6FGISzYgwItv3Pjd5In1NsVrMz3U+hhwTp4a+bgfCwsmHkwomMX/frxgOy6Ahjk
m3VOYFxy1Ays0HvnaD5jlth75eLRJeJjGX1x8OxD16AgCTrtPmHMOFZDCR+v77VQ
ktR4YOcc0tBOtyTu5UwA3E6mC34PC1i0Fe2rjUhvNOxUrkmHAp/hrxZEbxPZcuFo
rHTtaqNsj90LTCI12C1D5I9u4T/xYrHY9SfqTt/CPYAEY/zGLnHd9tx8uuIB5wiO
JheJecM+HFDIM5iTWMg50y86Z7QyBh/yGvvXEC7/kJ0GoFK1sWY0FmPbnUjFcQ/I
V3N8ddncSaVRupsesCoEd5gr5SN7Yd8fLHi/UkU/fMhbQM62r7WfA0XSMnu7tUZJ
fX+EGQmmD6uuPUi+wAhzlj7oIfnY055coLk5j4END7IABzOFbYMZUwEqgX8u2VL9
0Ool1QwtvePCA08V9VNenyPFBi3bn4QisgVRoXP1eVSuuYgXqSu6CPysKdZiGUpT
i02Ddgnj/P4PuJHMKHnQVLeKA3VFuS3V2CDUBlPNY5TBHeCZF0i+N1BVHTJ05vhk
FtIvWgTRVyMVvWtn+ybE/907sXzD6v3gEWluTjDT1pgESGfN4rsf0f0mbn/9+JpC
s/nso2NncBgPPijsE2XD+HNeXVkhGfOaJyFDq+m8VQZwyYpKULsTQfG25pzyr6fb
1ZQBkeDT8UJuGssaTXsGqwshL1y20b7RgbdWxE+75jG4HVg8Lw6jzJD5LdRZpEXc
9aY3d+NTZP9uviK9dHYgoQUFXKQHdpgvQ+CECBfLVvCgvlVVCsgn8GxLgzHSNeCt
TvL4lFct8JWu+Kk0F4xJIIzs0jNeGiipxOU6SwvbNBhGTTN6fjnP8Ih/zKEKpbUr
wdJzhpiTf0J3ndYfQublbvEEZJ2sMJRKO+NlAJ1VOULfFbSzHp0IiYKBi+YcvAVu
lgavNxr25R5NNdnyHD3HyWyHCwBkcSjw/RaAVRO/hosWOInmwT/bKLj4hBb+qdlK
0LAZratD+EFAmrbkqZW6aDtVu5xY+TZU53YIgHApJuRJEM5FfUWwejRL+2ecuTh4
xxJcG4Z5TH5IoCcbjM1CNqFFiU3Oy8bnymtTxKO7iMNYKOQY2LEgvDx7wcSxR2Ca
zgelIDD8MSlObt9wkSVocxP/abBoP4V8O0zGbiawQA0IkDc7vU8cS0RiS40g0CkJ
CmoGaaW4zoPsde/Nd42ImFkBCTpy5y7S0IDN/pciBxwfBllGWvy6bUCxP0LJMHIO
LWYUUi+/VoPFzFPbG3BBgcgmUJ+7Nl3k1GF277WpQNii+MTj0Q8nJXZjRUhXvABs
hVvSbH2nO7FftoUgq5fW0T/uveOEFkNKbDCLzh6En3A0El6aRmuXxwTIhzWgTipr
p5e0YF/YBaORU2tUNrh1DfSOYH1y6OJjlcTQS6szm8raudlv5HuMWLHcFiNUh8AZ
HJ8IyUENM/5+D51Y9CEv41WJj75iV8JRqmseJ0hkwnJa6YHBmYqUuZ8V2TZ1D1FD
a9JSMyXg+TOZH55iJTewW3bhvdhNKfnYVUGfs/RidTygPqYyf6sSZt13H5sOMPuX
U1tpA8LMaWjPGXInzPd2dLShdlJkzuX12c3BISjbngw+eoZqmk+KknRCBYgrv5we
8K6PkKjzAhBJ+V5BlJLhGAyqePmXVY1zFCwurarq67B1Wj1s+93nKOWNyCi35kgm
FfWDETmsxpFerHugj5t8NABegwSrxWfXQTageSc7K9JH0REehQtBl2Bzp0YXFK4f
EX6w00Gabjy6EBqAA8V4bwHJ99TjPrZ2Ev9hlo5Kxvsh8j04tAHeu3hexwctx6Wz
+nv9GmK3SNAwtzMgMKKmgQ40ofxvFCXl02FcaGavhQac4/j2dAszU+3mlyArODxx
nb4a2MzxbWdvWhOhjjP3gAIAfVTge6dKPOdku5kWMqpWmGrxo//Qb2KvWMyrrRKu
iJk1sHvveA/OAa4u8ihgKNbb1Y4/pxRFCnN0Fm+jkMCMUfCpWP33dNnt0XTaBC1+
n5IkmmNfNo/swm6+9dh65aJIUg7BLb6ugxJKL1bIQECI2oXNlEt3oq4zTCG0GDl3
zRTHGzQi5ZhnbwRLYLgGIzzVr44TGcHqNUDpd7oKTsTMt1yapc7IY5YeB51jxLYX
MVqg6xzGF5CtkDP0K49VxJRLNVAv7JY/PDr4Hz+qU7KS3stGDm0/MV/Soqk7m9pv
BvmEdHnQ8SvYEkMgUxUjVBQRMZ8ivAPeVWM1uUJu3fZZ/WF+lTKNlVYClzTNj3DE
py63s/A8E3oUNcjD3KWblzdfIFabjVO4Rzw6YEkeUO8KHKzzygF/JVdHpio9y6tO
fapu0lJFvJ4FEieIAHka7NnZVRNerDsu0tbXYZ7/9abRPRALBu318Qwkeu0eLj/j
kQOK1gool66eM9206MTBWzBXoIshvSEkgYMRtTwKrQMnLj+aP4BhAWZtd7Ln2BsY
aV9oPgvWy5+pepUvd5dj59kctmRB8/WAq+O/ar+Hq7xNTidf+IfCOdQbWM0/UC79
1NG4vyfUYP06v43bGF/l3eTugUXxirYvohb0XFUm47wmT4j2ucVNvxlooCsMtRLb
xPuHIuwcXq1lSyvnzw8n9IQeP9ibLHZpDXhYs3HlbVairxDEihorVI2z+wzYlu9E
MjYhT4T0YoKLgn7K4/IZegLhUcHG/y3aox3mNLJjtZjI7br1SSaG+15KcNMSktgg
W2omjdfgUVctKN2c8Up7iDY1g6ZX1wnRUFi0NdMXxHtFd7piFnqJXUJ4ysqyx0Tu
iidwI6lin9FOsdztSjXp0i7HKA+RashO0jICdeAjkxHd5Ny38aNwDUiRo/Vc7h8X
nGVUp95++Za+fet70ckEyYkBZBkDRaGMCp1sAzIzUl6hCnyuZyGfziBhqDHUM+Ho
ApvvMSJO2K9ntmfsm8sUEf4p6c7wjvmWWNgzAnnn7UkkNWOq8pamiYooBbc1iFQX
RjWzHsv9iJvpp0vpJtMYe1w5Q4ifE8+L7RH8gzsnHE2mMFwX78WG9PNe/Btk2a0F
UTJGgj41ZLpA9bTMEW+K0IyHKhXmht5XhsqQOz56cE3nBqa+GaQFaEwWZ7hHzQJB
xCYdefK7/TJd8ADx8IVOS/+vfEzLBOiZB6ELQJnatuMVpQUGjiQeWgSh7531m99O
GUqimDUNpmQrR5l4MqUU3kXFo5U3FT8h/MXos2fJmcwkJ7shtAmJoSCt5d9bzzBu
dKBTiwTiE0MmqJJEkwXLTga2YzGUYN5yIDwQ3h7KvZC6VhETLm/dE/1DVAs/FKwB
9aDKqlw45LvBtom91fppo3F07S+txmkKOeAUFBer0460nU/aYJDoSb2ZmZSz0dXC
+E529LTEAjjCMUsJ+ntDU4mC7Mm/A/3xBmP9BU425Gbhr35DXDpBjTSmokz3eBWx
8sz5kzMeT+C2uWvzPtDBtPnb141ycsmW1E17S33JEat/QdYbPpwCyVpwGKxPdxbA
s4og5hXL4k23GamMDhyKlF0qYvi+2Xvb+7v05u1N1GCbrLtSnfACieV9YPi8N/g9
xqOc2pUxHnUm+QTPcK3efx+33+4neQ24UY9O9TKDhSNxDr+9n50AiXLYOn/axicH
A0Z4vhjca+aktAnlTw0OnJD73IIatxpJ3xpwnuQrtEQkNH9yHQPXxFnUDxQf0Uub
xxEVkvQwZdaqUsvNFXH84lss8z1X20jFObvLrZl93SGilN1RvasfpY9vTpLSH/ya
eDLjm/Hm8XgqAZpQD9VnY/zwmmfLAG7577uILegjEoIz0HyKo5RHjDxN2o4Wpk67
JhIhoerF2tI+lKrd7cZYxZLEY1YRnMJgYy+ssG2Bnmm3ZaZoS5KXxApdNTXw0DyD
30OH76Zhu6KYfzPyFXSSwIa5t0dBaSazX2+EMh7JZX1t4/g/xDWjBarRBasdomqh
vbw5RQh6HiUUhLP48kJ4VWWQx3Q1Rjr+3siRhjasytpib2Jq4RWKiU4PHE6dbTax
cu8h6XiLBzGcR/0VGPLiFOlT9yhvaS2U3cRkFGGkQYmLFvkBf8ySzs8dPhuZ+Tkj
yosYfIuW8E//IGuW3iDdwCFvfO+wiekMDUgajoFK+7Wp7i8CR40rl420uXpD3TST
7E8e/QHvL+hNIeePBqT1uco7NrX2mYmAE4QkhzQ14KCBAwI3qHL/B2ARqYBkxwfS
Kbg3xIHnTyRY7KRzoXwYECfmxyphpH2YwXwpvihgElujWlsKelR3NSc2UkLfR/ea
ZOpOHAbEPNGGia1oUKHTnwYUvnlo7hpUdY3blS8LdmLIlkgruSUenrZZ/0tGUBMT
h5A6rpd1qLN5cefEC/Uyn1JwAG6/0qZ36rrVUC0Kk5xK+dMHqBheNH+M0b4ZbSLY
HmOFvN0IDq0sBI2JvjCShHR1nJ/7io/TYSZAiK0K3UbSrm9XqiZhfQVraAFf/y6K
fHFJlUPfj/fi4GRStt60FIcTrj82yniJJGhUTb9IP51YLbvx4t4uU8z9K9p8Qrnr
APid+ACZ6sek4LO1kiuKhkhAJp8y0+TJnrdwRHQjeXBY6EycS90VMGXgQd66n8ax
a0Zh3EMSnnDvJqr0/7ZBrf0+teApxxhwq/duddFEaHaJc/dLXAbTYUE2ospZDDIg
KjMJEkSiJvndow6a+b52n36ZRSOU4wuw86XAG93xYEJOfvs83yU7ulqj1PvrU8tY
sOyl87VZUpf2fhpoWq4uKoL4RWeoZQxK7189EYkiR8/0Y6nbpMo7KYCv96g3QXm3
VI/3JJTAU1Dr1yvfmNtAKalMrNnKMxltTTMEk1wohKDXUr44x2KNwI3DqtVwMnJT
xcJa4yO5d+DrElziSIJcQnpFM9x/Docj8W7G5qPeD7ELXnzNmQxxb0XpJ1IW88Zp
6n8hRWZxPr0X4h0rh68YvxwFC9J2dnJPKwzYzJCQehF4aDAd1B1+yGBjmUz2cOEq
3C8pM+CuXOfZwIsc/Gs9O1yajxcNQ3n2xiADRUYnq4td0/X9nR/cC1yB7CK6QU1J
iaZUe7UbH6wM7YPtU/QqBC1OzEQa5pHBgSrelM4+Of1PY/3pA4kH6AJazSNTlCuf
BgJbds0iNHuMBAK+IBRdGuHaT5AMVaDLwTFyfZmjwJjUyGKU6d0KH01lpHslKLKp
KsZRZ6RctoGq+RFBQVHwcEAPPkrWRNygctdzhpM5s5PHALPHO8f9QAHZa4Bt1kgL
Nw5/Lo1tRmojUQaIow3oj2HaBBX+X+cDYMecEInoltRKDdWI36etjSwBisM7Nm88
OXrPD8pB1hW5zuQibND1TxdeR8G892NEw1WcHJOJ6Y4pkL/nba+vZbAFm/83lS6b
ThJ4oE2w90xT29+Ydk7qFhisrCeR3hqS+P4aO2KJvGXJWVjRWSyEXO0YnfnwfjIl
ln3Om51MqK/5UmLXwWfXs8t5Nf+jC+EMMUFK2oLAH2uo1d1lp40CzEVOJbA1KF7/
JkXp3HcOTl97nS/sa+zQ+AznNyTOENrJJHvBW9v0utmP0WTMmfiKxRkrakKFJw42
tyQsd9UHqH7W4Aj0NWLUW2yB2un2f5c+I5Eb6uxU8C7B2m3T5T13Tpb+0nB2Er6l
9WGd6FB8PncB5cvSd6wL1ehV2j4XtN0jy1qwwEV/dMn72NerzwyxI9Y06EGagkAI
9nMtLmYePQa421fHP/41/iMWxUtGZ4/0IM1RlIYiZdOTLTvrZAEJAw1LKtU60RU+
omq5TfEjRfzzIhSEZ4mqB8F5NqCUhlRLUYy5ORMgWNarVqL9VHk0URnsJR1RhiSI
9enxT6c2NCUm3WtBj00MJ9O1N6FNYZYWKGxXWwShzmckOgg8s8j8g3OIVvQXMLfP
P4a5+h8lnnp9689F95IxKI9uFRXv/UuhLeUaj4i7bYVVfzxTopjRrhW8QgsArQMw
k+HEWA6qPCshEgEpcS+dz2uDcIEkTMmTV7FZ/jbJkI3qmWfWTd8kmUo5UZC0nDGX
7ZWUPSskJOo8qIKDjD3pk6LWV2vQJoYLMBe0j5wEXSFeotU/l8n6XVJ9crOhpSMy
k/HG1kwvu0Hs/QIhTdhU7k4l65yuBqyz1F8pSLK8i8t7g8jbyJkdLmm1HsEuMb4Z
L+54/GDK1+3EHXROZwFwzk0KZ0Q9wc59Uun1FCr47NbGmDJJvRVfXe17G4B9ioZE
5vk310cszz+ulA/H5A1srwDpIBfRPARqizneIDisH49RuXdzDp/YuWTd2tPyo+5i
YZEaNM5JJ9pEYKWLL/H+CDOlwxpON2PYFk4ELj4o5EbjpR3a+FHNDmjhjGa2riMH
sANuXS0pqctLMXIQpMqZsOVxN/MFqrlC044jNoJ6bUDhWtLWa8xPHZgWpNLOEA3Y
XAVxT+cdEKVpXnem9y0Iaqt0uB8U7QGB7Bd1d/KXAmxgtsE16eI6smem2387P0Ek
JdXcw5H6E3mlfIk1GZB3MIsGys5dDTV5J4Fd4Cytlyx2UzthPFwm1PqpruKokdFC
SfkCWAuKKlB1qFSFxXIZNjpwr0GUAQ3QmMTkiX7fwc3BVcYgwk/dn1ofyn/0ZqoD
/b7JwWC3M6h3nouOAF0GJoxsQ1DcXltMf5zwBRy5ANbPIZECioRv1RHkowaTPOIe
RveFe0fzYYCnEIdSbQ/GbcenTEcQ83cDTXrZSxhQhfGa3x3JIAahBDLx+6X/RAhk
7E3Wzr9MmTWjmcqYjyIlSZDVM8d+vpYJ79iaDKK21QrZngiNcjeK7mvvSNzBYlI6
Vu4VRRPj/1WtziNIpa3CenXbG8SIKnrqCgADxtXJM0PA56jvb4AnelRYEcPQYH9N
bJHzBvz19aGQyYdS69zRvPNNYvSMXTdOzHtkPULvIv8dw4G0jVq0rnNhpmZjkZvq
l8XBcFovUmMNTj/0ICb1AA8g8Wg069URafQc93I4vzxMPURaBl6bJx2GnQFO3s6+
Zkk5Q1FNRF2A0XwK9EKVMHa63HGMtdnGgSuesGZAVzUsKnNjjAPLwd9h9O1VjnMf
aJl6cLN28Wzy6odNHAQJj1THE0uYMpmXRNzGMuPBya4v+V1gz4k6ecPFBrGTsBBc
OwwggS+PhXz5+Ipf7Bn5jFpqDqSXt/yia0Tluvi4SnWTGHVJRQ8vJRBckKXTMdvq
wE2WrDQcin+/O4gWIlbrLZXqTaxFG2uBwJfKkNJau6auW4mnI16yA1w3qSrqwzvD
5wnmCXKeA64iXEgTe0o4RALIDZTo2v/On265x2Zs0QoNqTfIKvfzGTMhfRdNhK5j
4+5s+BJpz9QLY5GfBFseFaPSxfGquUt63t+3YozBAWt/gqLlTkhh4UlFrFx4YMCe
3zi1Jx7uh1AUfh1xkRH1wWi5zLKwvHCjSF8ZHWeTCR8lEosHugS659MPaoVlaPWd
UAgYctcN8pnvQCIg1gv60oV8Y6JgdEj9A0mHQro2i+WhkWVMFjrI+apgAHNU4/yd
Nd+6TOft3vpHDQZ4GfxCvxre87Ds8m/M7aPCmhirxYcw7X042OmO2VHro3D4UL0F
geoeB4pjfRI9OW5SflaCx2lN5QzmhVsP/h+We/LWHqR7GAnNn3BjHa8SmE6YyqA9
7283pClFzooQbBCnQ5Ypz4p3xaPwP/N9dQUCCZCoOPHIhRrg6rAJMdhSnAMZ9nHt
gR1Hirxcd+7Det28V8sI0e1tsHs61NeAmFQuCrt1jfq8fESfkoMRU/0UauLzZeMY
ffDUqxl7S4nsLwOM/4UwraBJe2hGjpJkLBdHWZPhVmjWdRh6wDZWQA121OGZFTZf
N352o36f52b9za7Q8muqU2QlAQsKKMhU9OSfL5bVcfL/Zo/XDFX1wTvPIuXLHC65
eKfCwZ7EeVfhDN72NDFnrFnN67Kb36RA+RgvN4hXTuSCOW1irkMTmJQq/JJe/XaV
hiR6iKyX7Qmih2XqxRbr6pRXLwGi2XYb2K/VWLsqf4F50Oi6FZYNqFiWXJmq81Fd
1TcHJupuzBI/0RafLjSj7wskkmcDPuIeaJZSIJ7pXICpens+cIhI6fOhJ8Vlm+23
/3/DONQ8SPNYrPoMlDvHrQAD1I9PB0JKD6ophwYgJ9SlOyM3RDbwI4l3Gvxvqdrw
YbxlKnwqhiwPSN35TWOciF2v/S7fVYf4r6sHnuGEqLgKytXzW7K5kOyHrvhDiuQg
DUAx7x4pJ6GEBj404CQw9EOgXxlmgUdWEleGWc7o8RjiX18gKerTK5PtqO6eyo5Q
us4vxGuVt6Fq0SrWxZQx/9H+6ol5VgrLEzaQM6k8xMT+ye9xotmLrOlcEjhJE3Qk
Q0zGHPtC4Vex4Vb5m1s11/WK384WMolqa0+HY/yTf8lGrpzs8Z3HVTS3f/JVSJ4M
yBmpISvao+T+3aZIzPEEmL8shS7EJCk4ai3PiBwFEcP5pw0bKdVtBXLA5dSJ/lqI
P3tMBR+P1sTRnPu6lORVt5QOKVUeGKhwSwTpsgshQc2tLqtOA6+u1ZjgEnBw4Ybu
mc6VoDFDAHT2+XsxtUnFK+YjZZoDE86k73P/w/Vdf/j4UIP8usvdFtWhjEl9Zeyo
p0Bj+WTQoaPi1zscskQWSIxN0KPkSagygJD9LUC2m+PLb5SBXkhvZmGpnStjdJXN
WZVRJnGkU+fJdKdvni05nMNM7hyTAMjnc+LYh7V/WTkgR6/5xlghFGIoVYts4Moi
iXhyoyXvrPQnW4Va1fA6TcbwKIrfrBEOd9K9S34naZ9giDPEl6nJ8dJ8cQllRdhd
00LOQTsVSWiO/77uWOEIaZB3OrVSE/QD6bOLB7+3yoFtd7W3Az96zIK9sYiojA8J
wv+3/VuGJVBPCFwPnM3VwatTWRKG/1Eg1m6R7Rcr/kogSzRSSM73oNaZXA4PSmMO
JIBQC8hJU3Q2ufhwnhMQSfXM14lZbvptTJjVro0RQpQZ+4+soCafiX4JoQW4ZWR3
ypbDWmw9Em0suqV8wBBKzYXXzWB/dbwcj0qjhFwl+GwUHC7j/jCXRhlLqAQH8mTs
7OfcoeresRRG0bm56Qbiwn/WGShkQT+kZgBQu4fRiKRuq06h6DERtKLH1fjUt3ED
/e++Jn9Gtu8NozAewj0Me8ngHZE3lsd7QhI1vf3lRU8Km4sMm6FTF/OQof4F84t5
4dR3xm2uZ+EvN6PJQyNgqS+doWj8taiq4ysQeFY2DyeM+Ctc4pRj1QrcE2GNtV7O
rXOhTlvWIWZRQl/QIT50TlqRagcyu+HC80MaSILRlwfCPghy7TjE0I2huCDjdviy
mo1I9Y1obCLepDfyLit2N4gUIQPuKtjHkn+vY1Mv6awOEkEuvdbaecM1Cjo/UD/r
ss/nORz+Zp//oy01bqUAsINvSmgL073Tu6pWBT8bJABF70Vifiv1iCExCBTHVr1g
Zeem72X88rjDpzmUj92jtXb4My3jApl59UZMMpr93uqj2Jn76bPVODqV1fJddwWn
j0r//A9bGfKV3nRNORjZ3Y1hHpxX+kW1YIquSiIZBhGDmmmsXk6AAX5DlA3nY7lt
vBneqokfSMBf2s1RJUCWimnQrKqqGq6pKOPxqYKnpBb4amO58sK/IEAfx0ykDHro
X0bODgp31qJOtK3D4bfkTDlSriILr5p5iCPT6w1oU+B74cPrcPCnQL6r45ERuYuj
KMWhuxDhINrPZr0DJZei7EkwghZZddCv9uAuQPVFGrQsXJrBHAfterIndW3cYVcu
S1CyKwJ2JE2u/53+371yrCNg5SYEFGcWaaZhWoNvVQCSCWH5lB1VVd5bq0GIDOsz
gSZERFfoCBUXA9A2LvNanAtPR3Q7/TxtHvwYVfb+SZn67yIOgORbvBi4wI5gt+j/
vEwSBHZHSWjQqlnFRiDIQGTk6mO7nyOqdHOP8z4tkCBfASiDdfkv7UrOQ9J5I8VB
rpSeYfAfIxhSQ+jbPs4Ms9fX8Y3Um9ZjPjDKpuyXYKwtySvrUFpqzWuL9gMKE6AS
BvZKzrjr6SNtyStnnv1OQNZsdTpRKKM8AIO48HC7QBqzYpRXuTuo7Hv3hx1WLbK5
qlgAJlR+fSSpvjjinw32+yOjWlC9VgquqWfGQx/DBZP9ta/BYMHMn4cxPlIp2TRN
EhNIRtXBLO4KpOGAQEVvzOA6gRud2hIhjhNRb8ihtbVCq9e7u/RVSvGQVoTutgk3
V6ya43iKSfBlinl7X1QtnuOR4JW4qOxAqEIhqpYjjxWy6Fdi23SnRH0tvqWrZfCu
C2+C6lRDgRJUTn+3I0hd9ha2OYsmDPLEP+0UCHF6/eayk3qqKVVjla+YG3wmNTTt
CLHONDzVBRrrQ+AzNfOPqfsN8kYA0duoE8rbXqd2L1rh4Ycs5SxGnSXqThs1idyr
JOx+cV+mmDng1Np/p9KafwLP0DzZh3Ep7A3ZEkroBQJGAex8bG7PmsRaWpkfuP4E
ZR34AzvmVcSBT+WwC/4Z+eR78uDocmCCvqaf7xmo13c9p53AG8zIIjr+iXZyFOU1
eW/yAMmdGKIf2Np3KNUK/BrXEcP953LLnXWKdnghtXCaIMScZVtAFq6hbBtAWviH
TCfzwphFL0GOdTcYEMHHFMoSolpP8rHDAva+C7ExbxjlsD2DaNN6qosPT4/afkuF
vODPFHFHyEyeSnV11fXQusg8dDjRLMSt4Oez/gtbH23Tplr1VpCFghnqrMFjR8Re
D2Umi22N4yfCQLzxgzZqtXX7lUH2+yVGtpohYa2ijo9eFX+qOJ9ScBGiVcmR3mWJ
8oWMHN41g+N1MDi9T/0bgx6i485kmxSeUGuwvdYeWlcoDqkOTBUTS3R7VT2IawRh
IozsSFVJJG1otOTZt+SCja74wwMxdMhKdf3v1+eJV5XkzYOCbnfsIEZJOqJbxrzZ
EQGJbnyzhjTG8j0uar9ysMSj7kekfQE3nJhXpXBllAlS3Qv28jV9bbr+cww7YTOd
sygicCeWOW5RjBzVJhh2n7fAq9ysjuyyZFuzETgVmjHuFyQqVgxznGUMpIYWH6o6
3VKqsrPmp8wXSVMIxOyiqVk7NkY7Q6CchMeSYSNd81TlRCISTTOl+yD6CxJV/Z4p
SCcYubKKrEBRDT28+ecci1FfpjRSnFcI+TZ+LJuWpxnflDsgs7IrL9aL18HaR2wI
zqtjzZSqnUaNuwvNGf7wT5NngnarU0hTmRWa6NoCeEWAak9X4abXgihopuOHHytA
FdwnbMJTArw/X3M9pMW/DRQa1OA7k/iTrYpU0YjEoCKzkVNz8SE1fs+0HaBSAs1g
V3chwC4DqU1/Ae9cjlebrHAUTcUk+Zy69w4vEGIs8jqg0i1QcxQMNrFit5tu9Ch4
1VNh/oH3f0UJovqrqpUJvDReq33B3Ib9pQenDymiVwPo1npq0S0uBIJDs7qP3BqR
sbLFqT3yk/v6rapVyOmrTFRRr0UabmsKy+1OHPk+dKBHb+RqSRaJbCUcjQKnHl9B
Bubr6PC4hcLwHJdMvaecCjLIv5AOLKb+5B3o4jneXzGqBw5nvxQVcQq5mCXrb8FL
sE6leN5PFzz9HOmDdGBPlrDqsZ0iNpDdshycZNr20jrRAsHEAiRvy+6Y+0x2qyjf
w2GQNA05jQNnSzmh6juBJQ2D3rHHpREmIbv69FgyBes33lYCa0WvQd6nn9dqduux
I+tpXxtt4j1jFdiKbcIPgzxRV8uJCUCO3yf1KcHBv3+UfA937supqDahXBZwUjaz
xV3g2fg7B2sWLN0NCtCLbm8xqlk2mOc0Bxc9Xs7B137WYoZ/OorMlllT3NJElplG
7opseffhP3NlW+CgFbL1UgOW7ftzJ4aGKpwAa5cZcoiyJcoNTesKaPafSpsgC3oJ
cEPwQ4Of0HEy9mzKqqkd+pIpBQec4kJd5+K2CvLjbAB6nsisUrJsEU5iNfxEppjN
+wO2o9YMvi/+hZIq9he0ONB73fk7nFMQkRNsWpX7o77Xf2BKHPOTZkWQjw5D8yh/
UmujAP2KCPqZ8nfTvGJojRxX2DvMW3bZC63jqyirM7uCTLQvKrJcwX28ImTOBk2X
RQYm4eK5BpGYUFNaezwR6AcggjxxIlLbJ3aM7OG+5mVxXVuZVA1B4SpRm58F8QdM
cZCqqHYMv+6eeN2UAXUciT+2mrfk3entiaDHKGBu6L/xKoEzmLeaAxSpu8LCerCS
jKVeLI9Fd/PUqphmdKRigemn012y20iEt20z54SIoPp0v7xcLQzM1V6LK7ORes7A
MvLvrQz2/8QMDnUKN0et3H0jHaZ5aUAPIFOD6wUxHyuaNMdml6L75/3cgHfaKiys
hSWV1ZucA7C+CUkySQ+99IcUYhtokcYn6uy5AtA36wYTpTwmbVDpGooQpILAzzjl
jTE7Pu609wTslKnIOwqqpNm5L+Jh54fMjerJf+p35jrxEtbjIXPY7+DxpApAWdvC
NizcqSX0OrEx8Q5AktUfc9g1euegJyehfuLrdmypkF212wgTTYOSjB/oiG7Ub8rO
IFdm4KRXY16xLkAhUP3IHVuVHQ0zsJKMRglSFb8pMOmyKwqw5/BfgbCUi6Ks3HK7
K4QnwHzbmUertQlUwEa5iX5/XRzbj5CIfAStzgQhDhbzmrQmtbgfkg9TCg7D93MN
cUVa3zl3ck1ZJHTECRYS5iaj8TMZl2ftgLnwYoRaH7Z4WiAamaCQcpGMjHoM/m6g
84epB1UzR/Jq143G+9R/iJ4ustDXmUDJgLS7NWPLPoKbnUUAlNsTWpHix+b4ETsk
62CF1DTORLjbKPOs8ZFDEC0ZNw6MkzFSwJjhYyMCX1cj3GskxDonXUudQnr8qMqs
7PUXlnO0sbDQLyPZD+tqZnBOKhurXITb6WKAwub2MgBIOH6uNWd7R9mLnpljWf/6
KhvJu5me7N8OYsMSImFHLJ7Y6IbxUl5DVwFHpHAUDNAkp2u5zhJRwdsedb6Go4Of
oY+CWMoEUOUqdD3l720UJuKdvaHusWRKVSKqDPbhKf8PUyVLNfWPYZ7P8EEJFm6y
aq0N8gYgzbilcYB8D9NvZtKZqUYxUhtWylEgcJrBPyP8tvlp3jrHIpbFygWAHVFZ
imwTy1UAG4sZfy4Zkp6xbZrsb888fOoAQDIDuj9UYiNhgFHOiVZgaSgiuv1eHHBR
60FrgSDYy2LRuv3cWfzzRePIKoJZUsJTwAPLgrNGbOvyrsDWHz6kgCPlMFEVTNiH
A+y6DqO6gb6WXZILwPBLbfhxyxs/SxlU6k4cT44Gu65szUpOS3tq6Y95TWfjv27v
ddofpU5pUBSD1My51P3XTCT3SzD7XXVWl5sLkOLUyX2UDQCFxJ27fJmTxLVqPIDD
2UdlTxM5luVnUZvdOkbAOpnUBOPclQhXmP6YiNNamy5MzewnpGcPjzYByYk85dcc
1pORFRv5sbFGnXJvoqCJhdotJkQt4gTm8haFEVR9AkzUqsYUNM+ywgv8PhQfn4U1
fFmmTInW/+OVFN+EW0tHO0UwLKrdJkFU47bO57LL2JDYfjFYBXHOOSyldRTvI1jV
S/UxVrT5LcvEUIhZUkS5Qmr1ORZheGkuL3qLfA7TBmR0xaY5rZUEo6L+3y96l7aT
WvbrplyQ/Z6LwzErupSVYExeV/afdWaCnyAIANqqQ2sixkN980Q9Ld4PnLC7BAqs
uLESIV9px1TxTQF/2yojabJ1r0/zCc3ZbYWVCZa1kJ86NcEdiuwNin/AE4HoQoke
1U5nb+F3rdhHycB6NBCH/3rL8q9TQnbwN75EstvORBmv8XVd+V9+xhJ+rjqKLd+5
dC3qNio/V5FqALK84j8xgVzzCexDcFoM4JyE1hNflgNaWdoQK8SksyRLX4JYoJ8P
OZg9mA5M2EkVtbTIp8F8Wkp6mc2xJan36aNKwgdjodBClgmacwIV3RoUAOKfRK6R
9xyAPh30sEtj2QuLHKjZJYdaBkWv8FCYnW3ktQyihBWWlCVHHdLZAHmBtfqeBMUO
qk+JxoQtGeuKHS0sIxCVNUyjOU6cc2A8fbNjHSh8UAzmjfdwMMTPENR4pAgw/oHg
9L7jYV+ZSGk1wT6JuN6NLPATMgbSH/DSSaJj0auKvtNaj4G7xoHEQDbkzBXD/kRO
DLNdSwe5NhtvmgyHK2oL/A13hqLj+8DYCyRlulxrjXd2qUeJDQMyx7LlnZsdY6Zr
/YFR+ZOwYbD3h4ynXYarZtYNr6/YNhcQvvP2KiLZl3Z7d9cD5kBH9Gpfz5MokU/f
PqRBudbZ3wTNADutG3g+WpFycPmBmQOgVrxvOSUU9Yb7TiWtanGeyB7ErXn1DQng
xC7GB0ZzXLRyLlNS3ndAiZWjRcM0DyKr0bAsF8ZO4XGyYrKmzj4xr4DsRYEhbr7A
ocy3ZFSnLWdIbJWll2FUxT5kuDHWkybYtbdQuWuAJ24ICaeoJAbCOvHGMG/Mw27z
pDTB2MHk9vNxC115Em+X33WW8SLDRMDiWX+aY0Q3MB0XKIqs5EKA2SKKXjejqKyh
oYt6YhPB696pLUTKhrHL25Cg9YRQ/3Hn/52vKbr6c5x1kHcPUSTTCFpLjRdxMZQ9
BrjxIxvnovT55hr//8FKGjB/f5/ApLEj3CxAcVITK1B21vGfz7OxokP+bntzC33c
e8G5Wodv29R7Mm6qImtJmaZRPzZ24UnpDjgpgWgYeeMBaVYKyfOjEHho7Ehyo9H/
EoWxvpl0SFAaY8+A1W0vRNpId/K927PPBB6iguMTlxsaZxSpI7EM+bwpM/Po4fqu
2x41PeHppqY9HvPlicMFuXnBWE7NxkE5iRW9HWQ/JRlIexryw9cmYQ9wcTNfXnp7
rgGrquY0j+aN9vxUngvBBDEN8uQKzkpi3smpFVGLd8xOxgCJbrAgV2gtPLWM7FZg
eJ1f0Lug6L6OH5rAY7jBtWKR/h7A7Ik7p9benSnTxlnrxRcJi/sYZilfiQvrFtC3
C+njiiK475qLW2mJfgMa3MpeX15BL7YoDVzky/DyH9yKB5uNqAaxg2mVvRSOrecF
ksH9vuq3fiscq9FAyDcdRe4F3Dz9NO0yRfMksD3Tf510zC6WJTe7LeVDRcRJuIhr
6Kk5vJ3coPF2+dqInPsMXEcQEuPlvX3KF4HrR3Hwy8jaNHToZy1+s4aXfsUq6k3R
PBTYwNoHrarfp++YkfZmrt6hQJXSEunsIfwUG8ljwWz5h8Bp14oAYDbdYkFmi96M
sDM48EH+cM5rQSyBrf/drjwUH6wDPcnSO1CqSkdFDOmB4BbJi8bNcD/jxvsKUlwn
pvieFxPiEH0bwSVYMtGeKKRWwjMVB2x5G2tScsk7Fwg11GSo9V1nLxV16bKtPJ6F
lBWNuzh1mi25Fp26Mtt6b233cI/svpqQBct2LBXan0zTR4HlrCuDfOVhv8NuwtLs
n9Xl2Fb4KHbr62cswYhcUGUgcYchY3Sqy5pYSg3SZl7YuwXqN1SrMvpNXZSZjd0R
+wZTfpg1VWAWyvotKp+zBXNLKD6jNQn20vkyPfhEaVOhjRs7lkFnvtEN4vlsZTrO
rOMH2lvKny6nHXe1bgEcasYOoJDKpSuHPm3S9aFjpc6PfC6Wv+O0pGxJa0kU6QPg
RRe8224X4qgK0ngYVYkKQR0L6OEj3sDLoPiexoFRtzy15xYC1uB26RTLE07Nkmvt
U40wZOgbNUCpr3cV5PzmwatauPtuyitGgOoz/4Ds9N4AkA49+71vQDbFWfzz2Tn2
xw1KXxsAlmvdM8+cTTltv1F8tvezoylygcgfFbMKOurVLcAJQHVvlmstigka1EFU
bAipbOX0ffGGHaenuhkuVcjeEVG0OrXbltmLH2gVvkpENymA6ay7XBBTYQfxew9l
y3L6niDDekmhfmEcZxKLxcp1YKRHbgX82Jb9mCyVTXBbZe9yNlOYkBI/16PlhmX1
ZEcmxwu2+QJXaiWCBVlp3ep7b+kbY7eP0wNnfKR9OW4FiSVHhsIo92Bj1v4Rg9sg
xAAisyqb0cbNfs2tkNmF6qQOwji8dR4GnAtsoJZANZHQGhQCxbEj9X9WYATob0qv
Uc6GjtdwX+B/+P7HDDYWY4Z7ehaaFVxZyl85Jp+qol7cok37dc7X2NUiQCKJtPWM
89Od8A5iwHTUnTp7oGyaHWnoQsCb8jVDjQ0JuC1IYSFfzG8plULue/bquGVdxQ+O
JQrpctgUdo6HcClVHkO0YMfWXY09ATgy7RNuEsqGNq9Jk70ANAQIfN08RRiXtZ8H
9Ea5ZqZzADJHZuAnammLKFcCgOQHfdF003v/1hglwETqvGZKPA8yz3e7WSZ70UP2
5vJMf+mXMXs7rfHhmmf+wcuJHQID0Z6nO/GfZyVrpKmnlCkcSpBvPmBwPHGNu1BD
ReJacRJjml/QbAkXniY1Q/M21ePV7uesA0oMchm59Fn28j9wTzs/73OGMfe03Nog
Ax22Xi6+jCWpFuiNNJSVYl+diGvuty4YqkLIU+WJYHCY6Ir4S/RUl1z3KCkEOVeD
DFxN923LDd38bnPPIZVCtb9vUKJ6AfkrtKTOTizdp8m+5p2vBeXYgrYVUqikXBHR
4/wAmEUXmVse3AOs9j0exoj6pIIa4E7Q3F9NENLXHeEcSvAfKY9M2eRdx0EShePC
lzyaSJt+PKfG/OkAOz7WSiKlfYCkj22kUwYKQytfpWZFQxRstE7IlJ0T3aK7RBCS
uUgcuH/LB20EOXy6o9cw7rgdbRSLz32lBV5Mucu0u30J/5soagd5cza9yIMk+Qgu
sbY7PaGdN6ncc2gmsDzirawOPW9Nv0oKswTqod+LgwCeelqRXWaYVo7ccs2ShVFx
ekxk1PNnGO2IIi18T9SSGpr9YgQGG6RhFWMnkEkwNPrBnZw/oFXiIk3Pi8QwdErb
1Rr28bv+gdyZ58KDfJky/xCt+sqR5mIniFyQw0JXifiUceXT1bnDeEvWO4azODrM
XiMAKv+bozw/sGldQTpnTsKpAJzZRgElFX+5ZyxULM7OoHupuaZCVceDVfObeD4G
rgZPKh4dZNR1UTWHte+9EpDPC9XX1+ymt8fW3UK3c6IHbUnCh7Cs/Q0MLyG97+1O
dL5ny8JlQE8hPrPhMRga7GUwLnSmyK0bJLIWwgifUjOGKPWix6riVFIYXU+vmhdR
9ckfMExp/FvtzPgnuNOiPqXUMaKq3Tw0dtLarjpcpK6ht1F91dSAcIZZR1V87aQ8
Xo/+36j19TFJ7G6YU/N+dgiCDvMTdY5cn14mBncU1omUou28ycnbqAH2vVAypyeC
kgYYyQeWsVsJq7UY9RrhJMm4Ub0o+VuLKQNdoApSSBHC+ttjyhUY98xwthWf9z8e
sk92ueE8m2Jjq5iI85CILO3w+WEI440Onf9QZsOBV0VCKfCq9SY46RtmsnLgKhM9
jYFcPrpsDPofmGQrjtqYQwzx1OwhdcI1b705gxkDXGQgQlGgJMZZcnT5ZlN/pu+b
DUcolOVgPsEVIYiczkaj7KD1D6a6bf0vt3t9PMqLpiseOcQ/zcl4p4gvh3TQpOlJ
AbFMugDEKjZmLfDEG/edzHI15EMf0dYyNuaQc9jGnOh5XhwQYGHQxWD2Uy88wupY
cDpWIAuUNB12k4u5UNuvwGGJltYV+t226pIMuW09Q1+1zES0/U797B2LFV9sULU/
B9sI9dTOEby6kvuI5s+nYDRGmeRREmNz6XpGOvclxtkUbxrkjDqq6axTJYl24hkK
mMyxVVand4Zls3050i4S8jsGBm5hZD1Ksm7RUnINLiAdo1SE1VPnSy5vkRGpahFz
3t7HYraPnMSZNaw6kMnru7ExZVaszrswFksMPpcze6Ti0wcp2TOmM63bmfr/BoS/
ImAs9mbpno12i16M8p+7LlWn7o40GD9cp+lxvfzmh3BqqxvM9JNIonW5XQmiAzvx
XWrf7Qyh840IW4np7/bE+O7cb5OvaklAIcH0jwV6E9ohEw8FGouZQjzZBtXihZzY
1UtyKGQcFge0+yZdtPoZT2Xxi6AKreGxeKgRsM5DCSQvJ23YMnlq0Q72seJLf06o
FJbQTMbuIQIlVXzITCVWOszSXF13IDTpic1WamD4bGqJv9mRp2vrGjAx0s1S6wbr
V1n6XF0UJyGZqe350t4+o7y858uO/bZBEkAkf5RWtaQINBkWYziFM46F7cwZ2QdK
V27uJnmKZBw0HJSQgrfslhq6BxYhvT/jwrPgNCoObM/N1g3lMAzH5krqqanJ1xe4
aHIQXNPo7oYh+YEpses+6cKPwA1trFfJM0LKvwksaAspuuy1aUeP7AQql9BIHRaK
ds8/NiWtSPxGxOm8Wurs1r5ZSFDmTNjVYSM6C//nzuSJSjVRZLzpalGZLOb+yrve
k+jwYDiuwZn+g1Gcp4rOIr5K/nSKbXUl6sOiVp5vbykvRUL8ICV/z8OKK1ME6i+H
RN/j+dm6TI9rWlps73DKBnQOjdfGacnJ0N4IdroT3vY5g7guYat8ng8rZoWmvkFn
UBeto1IZthLhTUpSoH/fkGOdnm7xTn2xQbpwWr7ryoyvLPgK2sA4euORwUOWG118
XZseHrCej4v/EIBDIGlnMkCMuiHifwqMzLdHHr9n2p3ZrT+2GlsRr7N9s9GuHa4E
Y48DQi2iwnaCvPqNqupNs3viNRTewLlEe6jNbxkH6YCeZ6yJaGwyE1OdBStF4dz5
l3Y/KQxEqGFx0OCCv/3C88Mb3bZ2XEbv5g4ceeIzK2p3aOG82tbR+QxJ12fIYAtJ
mxuD4jmPaw3THR3WgCkBydEjA8CCcPX+JYsnJ4a8nr+NLYpFnqp4XtC8EWWBL+G3
ylKBz7mVTG7SSWT6DI8aQ2PkrlSmLL4N8gIF5k7LMYSjYKLCSk3UplRIuZurHgVr
ld23V65BK5vLUHUc1pPfGQPmyzlgEieCacosvpn5dbYePE5ZoReHV5AGLqp72nBI
ySlun1FYjpOdx6qE2cZvqkqjRivIUP4drEUHWDsLmdozrEWyu4/AYcaMkw92o+TE
JLFQrj7cLfHEQNuJRMp+e2pqBrpdDQleZMh/dI52jesCOfvebXSejfeCqiPsCTbr
UFug/etqraQvvc8BTAbLWDibi14yTmeFBFD/iHrWXqrX7fA69rBcswUjznA1r0rn
+Hq5HxbuuKahU3gC9CmHJxIlPvRqiYm0rgU2U/YN+T+rvMKcIyIqmAq+NrLA5QGk
kcuP1awz7WBZ2vN0r+XLARHBCnCfwGw7GtPSm54K3e+GJGFu6yQbcmUWEpXa1oM7
PizVgRGdyGVWDwHsa4qC860bRjfmP38cc1uxOxnanHWVaIqy0IS/b9LwkH61u/Yp
5fJH9PFWwpCbaCMMMS8UZ2lEZdkMm3iBW9SGkKBQRWgWk5GTbdR4PjNY2XhhaJtv
/bbNLcpmAR6hgSMji5CJPZ/ipaA28VvOhtXcecsM4kS2fyBNGQECDahseEGRfOiq
jWL059wnsgcNrFbEyVIprr6WZyCCMe2Mv30gDZIWzxYUP/k80/eP6q7kBnmHQHf3
Z4Yd/0CaLM/0IVrhNLwFvh0HPvg3cMkI3A9bPpPE+tvr8XlcLw1PDf3g2MOVa/4R
qBCKitCJSbBKeHGoSFQkptcyXiQUPGJdlDkzEYHI7AqbSzlWlrlL1IJez1BkkS5m
7gpURpKDuusAwf8rfO0Olov3q7VlqGd2QQSkBOtzO4aLNtNiIlQo1PzcFPw2owaS
gEwoGAzxPkQlCiZQfqs3s+1B4Mmf6ag23eTM1d5mf73CqwAvx03y2DvumlDyz0IR
TxBUpI4ti/vvlYzDqR6GrV3hrVKjayBZjxnvJeTQPHiBpGuYZw3ykaaLynjPRHgi
1ebs8y3GAYsniBPXGft+QtWVS/c9meu0EJF8Vm9C1j77Fl0HKgQGrW3xTCwtX6m7
RR1mS+96X2wIqBUbaOSZ5XF6ddiNAOxsjjsNjFiIrZ3G5wZYM5YfL7s6NECIHIW2
Ydpg5itc+6Qas4Mq8ZiJNtVzUdVpsTYg2ArRU7VXWJ/4JaFAo/nzegHsJ0hZyYQH
DY9pblb5Fr77zd9u3WEWQguY4zymszkLLIyJRpUAOSM2oey8mzQLyaUjb5V/qX9k
6VEMEPDDLtjumCvJGDhw2UNbUfuNJ92OPgKi1aOhjByPYYWMwa5E1/c3hVFEUPhi
426Uq8ztEHpvUX1gdUxDeICiFxVJsXbSIxserOit0ayCI+TtUMQOlDy3iwGUPztn
nyVQe1Bni64PkdhS0lideBTPIzoYMWR5qD9bDXD5ajwB61SkECrarKuJZb+tpjeM
euAgJReQHMnCw6cx1XTcwHdeazmUOCsagUIyzyniI7WtCORiQuXNNLUnXYrx1Lzy
7MjRLAZDT3DDWK079gYmSCxuq1IhnT2TPv+84iuNOjJopKWp7QwmVn2Q5UGzl/e2
G7u/FpnR+/3TNg4yQfsX1REJvrc1T/6tmPMEWLddWXGyKiSMqEUM8CwVsguKBYaO
rSkW5oh5Pg9IVo2BIbe+n8yL56MmPP2SLgqN8dNvBAplHGo/RN3tDzg5gjEYi/Yi
wTmQD36qm/ldws/wxHDHWP1uy5c+PddZGmEs9p/O73NHvG5LzoQYvCQydWabHsJW
tH1FHWTLsCLLZOL7967V217c663/ZffKY9C2rLfZxg/yj1wtRZhZ2i8p2LIngIgD
pe/FFwqCcolnScaEcDdARygSJlVTz8ENW7+06HHgzQjzlUGBOdH+VfJpishu5vX+
5x9kQ1Rs1zHfFUbO7RVx3E/z/mnjjukcp4d8bvO6w8WUemU8j+ghAK0IUWKVuWZU
LZRgNPsohHdjBvlc5ZX09RReO4b0Iiuy3/Dkw24QhLsXaibTaEC0fzdk1fZhMDom
Z4lnUYjnt7byjmwvb1G4cnkox5MCcjwC+ZAWM0K3aayCNwglzYUUrRkp3ysGGvi5
hSrGJQGnpwJrvErksMpC4Rj+eCbEJ/AzIzJZAzEEaanL+lz9GCVzBCtNCsRU4W23
60vjGDnTZ2ZcCGR6hv/LfK7ZpH3AozTEyc3l1A4ZV8j3z03F09Qe5xI7h30zyflI
xTYny5nQ8l1ray2gR4WWAMjoYMkpVc7weiANN2wJ7CauF++pWN9u9TovxEEgcgjk
35I9wXlveNHvCunGSbMgWdihVutB0xuuiJlO4UU8SxiNREth0QLxb572Wi79DbiO
woyQ2Yb6BSUX6SLdYsMYONdc3ZLBdkoX5/PGucFfiZ8n+AyfNpJ4TepeK6ioSaII
7a8NdB8g/8GgsuiIGM+JwOd1d08NDUgzdxsazXRHBLcFoFQT7glL8iX0FobCv1Jc
aQjVcetxhk2fHnDzV5NjHdkGZcqeTwu5ohc+FoHNPG7lb6vMBX8i/z+DV0MxkdHt
FNHEOExByj5z8K4Qu0oQziD66fGsFYPMhAlurs21F1b6bIpZxoSIRJjSpgp8wlW5
toEPvrUz6VrC6Evh8B834ctvtkGw3vvEzAedEtZyn2Jel1Ox490E94WDjPvCD767
QNG9sBX4/kIA0vHr8gzubCfiOJ4nplR8qb/ihbtg1e2Wk3B/uXN/6gCthxnxzvDH
TFzzLlpvaVKinZJJaPpyC2bYfewKXeCVd0K2UV/WsryMRsYjytQu+B6r/dFkGrK7
GS5mUMUU/Ru6TxXl/z1er2quXpApao0bqo4JrVcjXH2kTniQDUGWDVd5pLXKJSCY
zhNxn93kwDkAInEyIoLnQ4H/4IHFItrtFZBXa7rscwdnPMYbHK1r9FuMUf3P6RAt
HyJQpxpwEq6BtNxUVkaUsXKgVkSOZYXFB26AYXOisqJkmoZ18S5IhSwPJKvrJDxP
9uvB2F3T5MaJfZyJZBOZVFbLyBwyuTZJsOF0ohXnobDpPLztd7To+BjfFIkACsKW
U/QW2+t3nhkJvNDR7ITJ1zwe9QwIHdmgczRIxSooxSF/Xh2THIlxhr3rEbo9XKZ+
/ZtIN0nju6tqQqjOvQc2N3cvIMVCtHBv4Njt/LOO3WxptBlqD9gOfdgT3+NNAY2t
X52FR/xHoK1r+hNDq3IfLH/noutyxFV5jJOyabtuCicivRWZjtDJreyZDOJ/qaVm
uE6sAHcYAw+HB7njW8Lo9yIUZXL8m5IN1EnI7bthgUnPzkDyloOvHCbsCWU89A7m
Fnnvkr0Crg7ghQDNZee0dW+5ziAAdDXNAmgyWN1dER7momxSLxMB1A927tVp6Bvx
X7GpGPjmBB0Vv+NUhHDGZ/XQdGVlsYnrf1VanCkG2iHF8j70K8b7LvgKESn0Rqj7
/hRWgbmV739K9TXlqGV4BurVpL5ZoCFAkzAvQugsyyyGVH5SSNWfo5IemY2Hkk3J
kko+CtgjfRnUN9ZJiT+wHljaqNgC0mFVgY3st6r567VO3bKKjInQPqmvXaeuDDSk
LYS/l77feH7YL5aULjqp21fxx9sbNuAgDKS9M9/NRRZs+gif7qd4NPW2/46NygWI
rKOz116b3QERImygGvjF97mzG5IlmCNEw9e1yEUdKkwMX5McKWLxVGETU2pqvKWW
/ucEccFyaSTbT0IKHK1gyh5O6czrD5xUTKwo8fseSKxnvY/cjKJaFyxp4h+ovOrL
BHGydf0ATerPM1r7RKR2vihHQvNBtXkaqIcnOmI628/IQ1uBdjJu1FYxbSt6fAnW
gzeL9UD62BQF0s3yT/6vMQfoIO+PifhJXwo5cOg+9c05B/tiyNyeYdREj+ng1UfB
7jcTETUQSrseOIaymyfdp3gDfbx0Zkz1bcjD9UyEU53S9f9GjrTwLfjmOONQBagr
9phWxKWMV2tmrVqhJpV47nrCIAfkcA/Ge5biAtBFDrSPnKPEqN+Y8GcTTXaH8ylp
H5GUamj7SNBvxIRCwpEk6qvHo3MRozgz3p0FM1toYKCeOT9aQhP5gdIPLcz8VEez
oxTtnqhmeb8U8TNE+0744ZwtkRm78AegXJSa0POFlnuhGbVw9z6ijf6vjnkYwPJd
8bIp3UZbSTq/jUXgidrXWLJ8fXkWEfK29h3xbTlHtMsWylEJKZPxIL7J5YdPvylL
RzWreq4Mzb8vgxU1WDPitMQahnYMsrVUwck25YizbCvVeF39KEURU9pjTvleKt4o
2829ADHMVF1IKxSS3Qf5oV07UkG1GuCdsBlFRCXExiPDuWOf5XMzEanYKU9qK66l
JO37oZ0+VOWbthAAq42PiH/ktTI9C6fzE9vWYd0OvjYCDdPdP5dTkL63RxDKa1gN
Wax8qPdopZqtrVoFhVcSe1nCsM1qLvQXe0WhtDsKVRioHFn5xtaE46l/FxtJTWZf
KCy83AK4d9eDJkyessZMAHqOTLaR4mZ38JNg6yPjrOH6wJtlRag25NHn44gxyRD5
R1vSntVGNMWQ31En/MY4OZBccUwTmA/JnZ4AgKR/hT0DcMznP1TBZ72iK4l8TWiI
mYVJFkNg3MEZNs2l4TEaanxA91omtQB+tGNftc0ZzGad4+UooLo9HLfvSi+YXQM+
PldHj2f5Pi5hRnoTJGpTyoNJZzQ0kquAelZy8OSC2p6rhDivYBeNsVgujEtXmctQ
HNKVb8yar+WLTXYAbxz08j1On08aNyoQ2MjckiIA3Pzac3kD03DT4QxmuCXETdF/
EkpAsgOgD6dkknO3jK2+VQJbFz79NgNeQF8rQTgzczbA/yY1QvC7WosGknDjOEOw
FaZRTJjP2HYvBbFS5/KKVpJUPamrIF2cEjxe5T7PVIQDFRda7Ik+J8rBIyLyYfLO
vO58pUGToNHZPkxhVa78x281sZ+NKc2UHHJ8/Izz1yz5XjxURourou/4RWS5lsdH
2+fT2qmveIC1bvXH+TNXlZ7/jm0Q1dmRIWLeoNIbVOjXbhshGweO4o5vTntRO3qP
7FYaM9PlEpNe+pVL+Cx8iLcGM4vqM1PXIttokLo2xZioMW/nQFJlqlgmrUlUVoK1
PpJys1Ll9pj2Zg0wYUtyGF2xlUcqSXA4+cQbnvIcfggqhJzQCJYTft+elb4qAZyC
dZFjkz6dYwWPtQDDH+zaZMHdaRUqmLSkfYjQM9r8N8frUhHKXorUQWiGTHQ5e3Ds
ohZGLsU8KrhRLDBo6dXs+UwhvGKGx+0WC5CsXGAZVDfbnyAb6TzahuK0P0c+J/s/
L3fr2f/12ZtfxRgJG9B32N6eCcgwLXIFHHV+XAB153IadzWU9/WFk0tZucuKJLe9
EV8u7iV3aMrnAwqpyhw/3Iu0RYDHJiQNM7ZtRs7iY9rwAdQkcUYJoKNAVGXoIAhY
xLIlM0quGDhonLBCKGjIIhQwoGzVgYIz0pu83hHvuQj/krTrfcq2Xf1lSAot9rxY
0d0mBcgMRZITZYyuQRe5ZDtYzFBJX2u43yXLtNlWFUnj5C4qeBy4Qq0zJWBh3OcO
AvfRPkXUg9pP+FCB5tx5AwH3eeUlu/sHmoNWQT9LJhWtYP755rVaOQb6KNU46qDt
zuDR4WjrBjYk0sRr9ybKqf726FmG3L/6fLYoLUrF69xYRWPRTV2Fvmg6d2hr4Gni
TuWcpamLEucd2r6rGZBlN5RhkmEGt35060zr2B3e2hKWJsTGj7i+xNctDzl3Ki9G
lOLCqt3mZ+qBJN4eyWUhgDIR1ULGhhrYKaqop1gib9x69Tp2O6R0+WxJmXi2IG+H
v/ONr49ETxMR99vQswvLNNrgmxMapEcT38oqJxZZwW5WLPmfXYuQNtewSPGL/Dpo
Mspi90HWIHmjZK8csqRSIcKklRTgS4rqCKdtbvZQ9A1MtYvvHNawBMW2po04nHGU
7866Pb09po5bcEAm5ObuexVyhRu9xfxuL/QZYa9MJ0HLdA114nhSm1tFV8SU1JsA
t6QmMjbDigzh0R80uAQxKrJPKVqH7BefUHfTeXw1YnM0J/6FykB0iuLl8HFIIvVW
Jw7ztztlRpKpJmn0cb/lotbYd3eKbwKXv3QbJjmg8Q3G/mSTx9V9kajMJ4QU9mIn
zIPFarjZBICEcxjSFFWAEZeIT1G4AVXUUGlqXOFVTxuieeFgOvobE7g302jzN3Qy
uRjEceGI3Zo5MWAK1w/Tn86NDN6HpV8tGX7pDKFQgIUywLZM1dLCqSINREGOYltE
FyDw+P9hfk9/P8DyUI7+nkkRWs+SJoa4RdIKlxW+ioNgLx1ouNB+G941f/mXeiQj
0tv2gyymSoO1flPumg8xH67eSXL4yzM+ikUWg6/2HhNkuDBww/FhyPwBW6M7hwpl
bYjEKg/5QujT8Tib5ObH7Nwjqeq2djQwgkq9yWbVjog/zWRgKOqvTG/RsF3UWwPQ
/B8iw2HtHnqXF+Oz32YHsOaObH/By1WNzTS8dm9SvnauWCJ7B+NQkcPWFGjr6eC+
m/8Pyelx30SJc4vqYc8Tc/K2g+q4ykvUbtaJ+AK6D9QE7oHJX0vc9ciJzjBTz9nj
3sB+xRc6fhNsmsETwlc7NNIp7B8XKQF51A3k9aWNEn6fBRoSpzx+QJPd4+sd3iks
Ldxl8e3TdUxoic0UCxy6UJS4amaLOUKocfT9EPXG67aSqFK17u1Lpbr3ExDA3Hog
xwEhyGMfJZbiXXs4j4n0+F4MZa0hNgDW14Ayui9N58ZTEpL6F1C3wRqIuVDJm8vP
bcIILcc1zeWZshIR8qemxLoxC8L4ryCrBj2c/kbRbiGnHe3YOJYq2b2AD+SblDdh
Ko/8agm2Dgl9jJZHon8NCgosFoa1OqnoRcu5ARQDoCheFFkNbbhvb0SAM+Zu2O5w
kcJFab7fNpw/ZoQYCsRP5ShyfddOf3oL4cBZWrSWzjQ2xsnq4wxZ6skLEdrcey8J
QGlkxMfj1/3ZNJkUjo+rzuNCCrxKrs2/r3pDrTCUm4FRaXZw49T3ryyQXzEmiENA
txT5CaU6rf5iNLuVQf1n0BxOcuimoOL2v474aJbBoGPLBay3ITbmVQqLNPzJT3RF
qqAx1MPTYhdjffVSY3Wp8+v+Q1wWZRFaTvuSqQzaKFLe5M4D0TgfL2XiiuYOxQQy
XWk4zqSqX+XGUjxdOJlHwrycgYBHTkiGp/uPSsJ+o43iZOOVdNl07MNMiSxd14+j
Ke4w70XHHtVveXuzH1xcY2C8BXKa7+vlRH3u6JB1KeulJddEQ06GwGBfJgDcL1Uo
UF0SJrkArsCpG4xDrh2KwO6uO+97fbgvA6Uv06HgL1HGHaEMH/Y1FTNOaLlM1/5n
9YYnnH3v1D/oUruFpDdrg9q94ozbZG6oNUeJbzOINfQYVXFmYvDjfnonDpyTGhYE
VKMuuODJYM5fLeD/79WpSXXh/76ZXAxBuv3szQmFjXDZuoojYFt95+7hETla3/Pn
fHH60Ztq04TSjue9OG1GyVZCegFp4lUe5ho99aBTMAgqyAi3ol6EiZXg5FXemEl2
zqwtV0VnNjcHGuAtGLU7Gcqx6iDZLPH6ZD80bGAHscdoXdYI8Cd+M2VYr2iVClkb
Qbgsj7Y4wBVjnz43XC7P6piNkjnJUmEvj6WvUOb0ORW0+hhsLYvtv7YCseNxLxfy
tRlLMPgO4aIRpU6umQ7TGF6gORCsx2LY633Df7M4z8fifrAV5Jn94q6DM5mxfd0B
g0w0gJYmhkaC13jJuU67G22Q8F6/bRVkuYzzH2cm8tq7wIaDBD5vXvrv7NtVnTGT
qsS/ExzfH8B8x+orjUh++I4LkgwcSYg9aeypk5uHHNHCWZXu25sNM8pV6qlAcaey
Gv64Ejm7f64UiLRpDnnM8YNuoUPCTUaeRSVixHEYTckrmqDgONgLjKxOyKxuro+h
oySJWKHfTkgKjryonPEoL/5uksoyyCb30Fr41l26p27DOf9PTSpKY18rM+Vka5Rl
mfR/eFBItWkqE8Sjhls9TFWYcAiHyf4wbL3D10ejQS6GljcFJt5onUBF8Xo9YYw1
Si4f3Q+7OY0MHs/iNFW8NDXwgnlrWHkHeOnRow4FDDtWvypFXxZJHvTy1ZYM6+s6
dnBElE+4+TRapvnvjVkO+Kowjyh7WhZNQAuMCtf0KKZmbHd+7v+7JNvLDQ8podl0
5q7uO93gM793gCMWF+yhqe71m1Yl8EsNLV6DwB+kON1JN0YaNE4IqFVYnQIiJcLS
Cda3Kupw5fcYX1kUwLcRiP+jIqXAW9e5c2LC/7BFh9eEuieQTMDXUsrOMtEU3Mks
7kGMOE3pVzlMNGEXxapOHvRzJEByzCbQK0K7vakZf49JsVzO5Nv6GKeoRmLH5wT2
MHqauJzhftuAX5cHcDE957FD4XUCOQPUwhQTcAGgpJQfg8j+5CsEbQDyXLJI95KI
5h3whpmwLYnMYwHYokIx4XgC2RawBTYCCGltw0+1XC3pMR+KW9oOpOoWG7QAyoFf
Wunujgrq2Cy9a6i34eQH5buDaBGFw9sBmfnCpkfihoLTaW8S1kxPlpvYrh7by9Ho
Jx0wtXoa4o5/GMzpawLvd1UunMagYWmLS6Ej1Ycl9BoLKxCy9cHB4TgecVsHtioz
RlP/hL4dSz9Mdl7q5Yyl4qYjJlhqthVnYg+eAzbFCy+HDIKG2dopFhw4XzAFVY7w
jOyAKTe9FdBPii+YwbEoQO/RE7xglCguAVS8Dyeg0Ni7dy+ECbrq6TC0ThrJ41yq
qNZ81xQ3HpgD4sCUFQA9OON2M5HGKIIB7iwop80ibwHjg9wh7ecfGxAx1uNxi/Ji
zwih81Nu2xKAe22hl6giYkdA6vy1uFVrHIxgJc3fpa7tAxtqLDBgOKxB4oyoihWX
cgpwZlx+sITjgQgio/JRJPJJFG/Y2AgwARLRUXZTMP9W2fT8Y1fu0hdJWoeA5PSZ
tWExBfjWzAWXRzOB5/Nhp7+UpsMMk2DQyrTys7QWMpnfw3A0k2KOTT1/kdEpH14j
V1e8vgZIEB1+DhFrSqStXKZ+Y2+7q15/uhtb8ErMFjcP2IDzAJMk386VklbhwJsp
HtXlfsrZjgBByr/uPQPKi2CVoUhN1+bx5gx5AIu0Bqzt8Tsu1Pzgbl1yvFuc+Dbs
sDfZy8aTdJxnF0p9B+r8IWsO5qEqqWmbkI7kN7efHht7OMKbPwttcawhsZ5UomH8
jZIs5gErnV/V9vGhNnD+CWXeTNcXNZKsK8R9/2CVibkvaO/I5Wa4cQytDXMHIkkn
sfTm3pBjJPgVx2fe6CE4AKQCJAz4lLdZ6odz8N5hEPF+09Ysi7bsRxMAMDTjAqxL
j3JL2JZWRD6hvHf0b+5k+4cB5JDZz128qgZBeB5AccyYP4gPVByYEvWoeIX1khwL
a4c10A47lF1REYrQuNdS5AqG7SYEb7ayUs4AQezv4tk06wS7RIyVynu2BdpMwq7X
d/wLUuVRh3Q8SCnCTTMt/0luBPjOxcRU9KVwWd58WokUnyj0DQ2M5M26pVJU0/wf
xKylb1w8Fg/KLCNFbUTRHanvMWOZumbn0Z8eb+uf4sUSwZAbUOTT6pOMq5alzRwm
zu2xbLd1Lm7dhiR949U8ma4zA+F3NF7wcxzIqdGtYkYz6uidGULy44ViZxccGJrI
hSQ1KGb6KbjyZvAexrcEKjQv6TTfw8RgU2iSEGK6QgDi5AyKzb3VToJSeuG7+ArE
357OgHXfU6ciokP6QB3vyOaFBFYlQ+F4zRjg7RXGmIYbBjXeqXbSeVrFNvflB1k5
sFhH74CHjtb0CKQCLgD8141zlcEKnhsgTUQIu839dtGsJdMTXbAQIohCOwGgKq/X
AC5W/XVg2BHWzEoIbnyzruADCp3cJrcAPdmQ0l0zNWE6y48XnPgcnoS4dyBUTUjZ
NW/EIeIIWOLSMpYUnqKpbBjpTW/At6AxeLEV6QNhiSdyK15V54KVs3yOr3AYGEBY
4RYPJIcz6DZnWu//eF1V2sCNmCt7tMVpsi6tLa8DsvbvUnez9+soK+2CKuyMy9Xn
vw+gZmTtBNClSEHLIPGWJk2lzCwVx9dssIWufpOonG/FBBreRpCUuxTEd1gbUar1
/FzvqHiHoox5X8lr1DqW9beYOVoTreROkGP8ovrl3QwxGjuqfkf/sDuaFPTg6duA
qTdGGAfYTcmzgfGhnRCnMCX3XxRzkrLWhCc/7MAQe8CEuwyBiZStFDbxiHenvEB/
NSp307ZdMkENeaVWz3UD+186jCm2TGDQUaBb8SC7g5m5GFCHJKfa0chayoCQn3gt
nelAx8GLdV4LklSlE3dxWELce4/0+M+G2lpbHpvruehQ6xdi9oMRw5NQZSMHpPI2
1VLrNhuOia56iEvIp+a2VwsHcMhSamtE+mgagvUxymfkfRghK1Xb7N5BT+wva9iA
EMoAtgu2x8qTjpcVdFbU/KgV7Cikb1QRIGef0byQ0oXoFm8+X271EaWZRu8iTuuf
XRctiM7nYfpPaabKy+9d54bZDWoImEyT0j6jdvNnhd8xhbJTOkjjU2Cgyc7UNKyy
zE9PxO8dyEFyQHQjvs07IotTj/LE8tIbjfsG46cRADSuY3fqkPdM+igwwySdkd4y
Kj/qX3pSKS013WO/P+IKksguKVufTPDseLk9Yb0hixiv8TeU/Un/hzxM2TD3tnI0
I0fgb35/DT5d+qdiSCoKzkNDF3UoT7muK0S1KuYV1H3ly4lBBuskF8wZ/8IBcoO3
I0vj/12eRKekLyHcnAZ0YeOEDstXlcV7q0fFLHgbz3bQAfq2dfk9Np2JsA2O6Sg9
+GRJ/iOr38fxJFNaq7MHqQgApNVCflQ24QevTC8oOHdTYb30xo5MW3lR79a5a3ZA
wCEc1CRXfygZZyrx6zprfgSDgAfaljC9GYQRDGlqxsmDlBgEwY3oL9inAc7GlE9P
qFeHToR6UzDecQDkBaNH/o32txJCrs0OqLYwxVt0awEJkdGJk8DLb4S55cw2EFiF
IivQ5lqbNIBoLPZVx7uGZEU17DiIe78ZtfN1SKpk1DJeRlzzA/LmU6T0/3CBVaU7
XacY2bcVGlh4/vTTCzE7XmPNgxp2qIe6MNBgPaaXNXUpExSqY4xYoK7VYhzJ0rii
4+igtT0gFZH06J3VemjRX3g9Me/sjKjBKMTBS43hbqdg+xNLBlW9JyVWHWwKAh+T
63jq2O8tLxTVp6B0Mv1OK8t9pV9RmR3GhwJl4uABJCzfAZinFMVWYNXI8ys40JUn
paifF9PWveKg0MGR4l6oLxc5CAOMLmZcOdfoenqMSr4tYLCIHn/S3M+bsA50vQfp
/1qql6J7WeRgp7wIioTdAcNGNvO+jtXmOK964Aog/sgzDlM3rXFknBs3aazgGkxt
m+mt9HSIMu6Edby/QarYNLTlDKG3sG4man+r92yB9U36disIhSD1Ls46tbzFVe7q
7zlClaGHJ0w3tG6ReQXwQ6hPOZU8k9OHN4HkGJ2yZBcC6CUPk4xazw4JctlGL14N
xysF/h1IvkbDgKu8miYoGBQiWVCKid1f5jczgyxCpXi/wiUhF7LGz/EFYmDEIRw/
koK7XJ4b75UnoIsc3FZWfaDbv1bBYgP9JZbZUiIJB9OfKon/xt5ZHQHMrGCDyx+Z
DMFDMnBc3QVyGk5nFPTKPbh4SbnJ1UI5x6KGEVSx986+tLaOdVOrhILlXHLfnYEc
8onI6m42sfLNBxz85aV3Uu4AnEhx2tVhBh75Rk5TmvSUV/u/Jj5UaWAoliE1Xkwc
d+qW2MTyocr9j42tXKV+gV6PXYhh7UX7iceS5dWFuNfrcfaB5Qh8Yle9Yu/OH3HB
4ppHETaRnjYllxIdaF4FUCv9VrXUKlSsyohkKbUBQM1vMMY7U2NN0caHIh//1pha
FzB8JfQI4cOn0YcNxKxJXYg4+ytNUpcZK4JTrROQQ/V426ozPDPwOrv1IhLr9DzN
nt6KvYBOvAAZLXYv4beCX2UyInC87lSCbt7tMD0tVe0J2MGuRPd7EtC9yW/uBYDN
/4jVhTdGwJnBdubLFEG1SJDxYo/xSVCbBQfWHZu42xWBO+ScTY2DJtmmUE93w9/C
GDDBTJpANzKA6QoKjZXCsnVeXarVSF844znswRkfC+Rmmuml0fQfdKcFeTWp4/bl
njJXJ1L1eGLiW853y6MH7h5UzyskZs5N9e5+Y5CydEBHiBvfhh3UJZ/ubnOVwIRt
DaEHyhTYU/XpI/YNrv+2Rl7+hbBvJmiTMfsgixq35kVIrA+ihTSwuWP3hr9UOyBQ
uNfuoN9StWCKbuPjCNr9Zr5uECJrsn3nJBOxJw6JYXgph0lDEvvHQ3NJA4mIiQ+U
g2dGjCuvBDNoyl+RFFtX1zaom506PBs6oPfG2Eh5Fhvfcul9N/0KKsBLq3nL7K33
fU8uJF7QSSvd5PvcRFPnLO5toDiSCjMyW/HkEtoX8A1q0SFU4WLrHmiKNPoKUNX4
T5m7ouIcjrtu/GMO0v0hoNXYLDChDUtH6K3/IlyxyC9Oy+zRsMc+KGAMc3FpJVgu
Ich+wV+JAB2quAtTyA+EE7RMI+FIiM/HI5Hpnr+nyNb/mZ4/fgQKbgyGVAjWaRri
fMdtkrKVQpGCTTHK4raqJbtnqQAIzsGBE6+sWdGuL9OxyoD/Sap1XxiZ6gclfF4i
XN3oi3JyOHSvrobApZyA519fr8hAkjwKgLg6z8YlFPC1ZHuRd9VJLAT1ESFWsY+E
D0r0pZev6sP9oowOSkkLaeMutNF53a6E11a9NAqj8uIx1neso2Jo/60Z2VWMS0Il
CSLUOYMI1eXWCGjvURWbpkcVn4w0np+poZVD2TmhwDiYtQG/8xC5vE72x/wFaYNm
I3qG+ke/cYfWXebOWCiNzz2HbM1AuIHCDqBKRp09RtOxL6IQEoN3wKwgvQbuekXt
tt8kx1n4lN+pXErdQVAd2tUSRaDJYIWv8PK88DcoWcRyk7Rx9AovZ2kqS6UoeLxo
cDIm7dPIiRTa5hwyZkkcXVO53DvgiTow6Pq5h1lTDIK6f/P4U6Su1JTY5PbRmPBK
DA5IxAi5NqgXKWbihvsWj9X2nSZWoIh3AxJbPZHjPlkaehW5aF6sSEBaGvSlWmkG
KVepuusSsdMsBhypR6odVeaxppiHgc7JFIecSLuFAWVzxAORoJiZuZlrT4ZSKzAe
7YTCRQjYrRqYZjA5fc0HeNC/3W/BdjrzDJn6MdqEWYJJTCvanaXYSP4pJ4jD5Lku
x53wIEXZaJHi13Mcpif/Gn8Q0O9miHcdqxZdmXqtlwIgAkgouOhFXxmDaCyYX5xh
LDYnX3pAg7T/ckNWA3wB0k7L1UYo4mOTAfbItML06lqEhIXt2eAodkKMKu5a1GJT
gQEifrUWKQJ307WrXZUdgkXi/GWVJBxPjlPJ2ZfnPKnHKDCLGQza61Cg4yqNN+T5
Sgx8IGpv7SrG0JjUpr+1lgC4gD/+EvWZTjHq7Pt+TFKqkJGAGJ63ortkGMKUDb8h
aaMqAr3qfs6ALVqgFVQout/+7EykSJsZ4rSPbDUFoGcH26LYv9BYw6+FxqRsBk6P
NeyEj8u11GoCK3X5ktI0qYv/EdrZyAO4mP2BpV8A20P5rL8KHSCfI3FyV9lRvYkA
9uLkUK4hgYBLQxFYyitm6VtSQ1sky3IwmJDiCZ2CrJD7Hx3KU+mMoUJ7mX+VaqYa
1i10rGeOkXTSiGvkmEWYgNpkhMQWqlPcty1FgFT3y/42vhNobc+tzgYRLGJGWjOr
6yqXnGq/i8JkqB8RSPQX9HcjiH/5quUUErcd2oglRJMo9g/b+0PojG46BxyTrKPx
+LZAHZ7H/mEarlOxvDrI56pCieN/TidXQwmYtJr8mpTkZLLTgT3HpXdTt6rAHqd6
YnGIQeLZVwfeqS57i2Jor0WGAhE8urfluCzkbU38vBiawrDPraxhPdM3iJ4Ei0mE
kE/4NcwGBUNEaZDGlMraaExD3rUjSvT2Cg+6l63/rMNH5m8odsR+hj3J/i0d6Ctr
ZzAN1sBz2PQ3PKdATThv68MkqFuqCQ8VrbwhGyMsL+haUrN0XqERJJweRQ14MUZu
SOBKHDCmIqpXdL7SUnTtrMqHjfqQ9SAAu3nFpIeTvU7nBLByEzoRMS+clsBt+nzL
eNZki0FfU8TWCY87Jlc4ewMI9/sSBwRM7MdLXWhWmuZNIkU+2tqD3lPi9pvSItK/
K7Iq+3cd3Z6YAM7S3rXOUITLCN5fgjP9H+FteUFiYEhwuaY9M0dtTE6cBgNl185v
OP84om+UdpCSJDD8DuDhp69A+hJqR4nmCCm4g/FIKOLtmRY9Medkq0B28qJgmaxm
mqgFAnP6ZLgKdcgdnBRefIhpktgj2vTFysuA/6Vz0hcqE9E0mIB55DHMzAy9lVfc
knh6chb+dLhJFu6NgjAW7T5Y/4aj3TzOB4qWjjjyonKq1+bpuzZg2cZxQ/fyHM9u
1qyAhvO39YL3lLeqiU159+Ei+ps0I+ZFibSgnm4yRhHrQ0+4ej0UaSh04+Q8V04G
mnGiACUUYuUpBqTsPt7kGvDaVqQDLe2IAcf4BOVU9HPZ4tJL8QTdAAn4CpTN4qO9
DcmCtASN6VAI9qmnHGmTyCjbOMRLusUTqDKeXJrqVLITjZt94us+kZEGNoHWJNZX
0GsLyFIv05U9n+xw73xN3HwuwAhYXAUE7+fU3TcwUETls31t822Zbl02oj1NE1B5
NckZaeoVFMK2I4VZ+DaqQR+QBwcfRTm45lip2TEgnK+8wLHpW07qsb1fXkS2+hrV
pW7sGBdlIuDm+tp9eH3HwyVjTSAyShmRr5/hm6+m8cicSiABpLwcPhKnPAlSBRuU
+qeckcSaA5oEQsEnEVul4tJ4bFK23p9RgMSquZH6aqIAl9teVp5aFt68asHi+Pf5
3YOChDLpz3EzoQ/w1Q+wupZAimLXgvsKVW5Y9+PxDwWcQ0eHKXIyE2dhpPCbpjHk
4t2ajtKavjHWU9Zs3aUfZbRjuMzNflOsj2NeBjVRA/hFxJXduucipcnp21GF4J5m
k4Vjjo/cLNbqZyBWsUqqLNmz/SroboSOVjnK0xOpaUgyQeuEpygqe1Y7hy1xDYNg
6sXtqVIB2Zcn3zB3Jqba3ZsNpSCDKQb+5mXZ6OqpxlEaFg3T2L2BO5NvVFPIs5fh
wKKe9g/BadtQvvtBnPNEzMYRw0V1CGJse5udgsvAvd2FlhUHqQWCr6ixqXCEhqOc
tml7JBf/huGO0R3/FhsuYzpO2aA7vpU69Hfu2imje4hDIRV4AYwQVoCmDrkOlg7M
l/A2QQOf/xKyclFxVter+LuXZ1eXU/cfMcEd/oDo5Hv9Qkt6cl1mQcESpp5QDCoY
DQjIMpNiD+3PkcnRi6S1UxTysgIfKljhDCREWKsC3VLOHabYo/gsCW8eyiHNm9oT
9/s4T3roIbzWkm496f297XCEgTVPuV4DDgpCBBBWmtTBsEScdYAvgdpgXaAIfSJ/
o3abpQZ0rLP2Uzebp5rZEzBWmzLYAe53QglbMjMToYEEanWY5kvhuxzOcOfabcZG
iky3uVGMGtwwrR3K8bAtUYsLsqc40She6LZwb0f18UwvHmGJZcW5o8ysGHzoJHDy
go1tBVpbHT2jEp6poe446ChL8ozv96T+Cy1TFLjW7PvZG3nH2/kjK3ScQ1fvGdNE
REhrAvzAQLIs1WmKKvmAfTxLqSEPUDVEF2owsSGYVViBg56aVHrPdqZd6a3AorhJ
vz/jvBuTP8Ah7gfJoDedPprQYov1V3dLZpz20cM5nsBbmdQdynh2je4GaYN9Kevr
gAq6zEFzsbzpjqP4vgxMr/E1IE44LC6+hmXNNhpcnMrOIC52BTVS43nq3SDV7whQ
RYyxf7dFBWDjEECJiZd/x/OVZ1j/WvnNBHHZ2lUYCQJn736QOCJE54o5qLPo8DMo
80zSTMl4yhMNUP1fVy+5HRNvF3IEwj4/+wpsVl7hq1t00X9bFRdiqi9UBX6V7pD3
6yr5OSxNv7Bsh7dvJDUSESwJjPesXFdhop/d2S19EKEAV+Ww7FKElAtxGZxDtStS
32aT0vecim4Pvug6NZB0+VyMHUbLHN2pkb7htfBJ965bF8X7bKSdNNwTErFb4V2J
B3f2JbGwcoSrbEZFpcXWIyGyNTZrBGAALqPbVlk1y6k1LqZyA5Ckxn8pj6n+WDbk
38XMfNCidj/y0oh/ZLPH1fJ/g2eMZZ0Jp7t2G8mzBJtfXxB+PZEQirhWoORMJxkm
3AJPvLwJVNf4Hz3R7Jv1Bs6XPCuAIbz3CbesfpdKdF12dHa+hw/SnLX7rtXVNAMT
ygM5k8Kfp/dAJNSPNJNZFlxYuPSAIKcz4bjrQShASKxyV2j1+quuWBabEtctPg5x
Hgn0qY6zqcSJX0NeEphKJpQJF/K/H+Xg2QK/CLnK7fQbbwWDqyHEiAKaDfGkG9qk
G2Mclxk6n0ckXgJWcSWB0c24fbUvQb4giBpSrJA+B7ewOF3/t4eENxkm59x5MX+j
lLLNLuUNB9s0N0IWqIQMPJKGPwrHbhCABWMaGSkbW5ocAn/DXKXIFyFG46iG/5ls
4R6MgoYgWNIgBYvQ56Kaagk8OvQWhrwaJLwX9sTTkxYcIgOj3LzgpP2Br+gdZs37
DJsVF8jKvmVDAuNUUaMJXDL5JUk0h0qf40eyu3BH0KD3cIVdjrDEweLAchZ45jsE
3ezx5koaSlzt6PitAGiUIwdsEKT7ASc4JI7AQaZ8q+40SduVhpgao5bBegEqXW4b
1604w8TNBI+aGpuxYCf5He4h7OieDyhEosviNi04OUqvU3vO5J9VXuagSUXnNcZZ
Ph8BKMz9Wdps0o1hDIfqtQCONe1oLt4yxnrT97zZlle+YtoUIcJeaJCK9pFtfa2n
vZH9iBbyeUN3Vn5+BnFlKV0w8Ro/D/rkbHaGQ/IpVy/USZGH5iRgkfv336+Gdk3W
4DKZ9dIPjApRhbxZLyQTeQJ98+iXo3W5/khgWJUk4EeTcv0nOhySoh1AUizPr74B
Xypx3UiougFevCr0yjeLSn+h30GY0bVj2mzW95pU5iHxycPbWVKwJrZ4gX0Vhapq
JT6WiHTUqbmoLQwoEEfIBUyTUObHMmBKr99amuDSCuTLkbhwSG/TXc5xIb4XJDPT
JMPesV5BMKoqSh6IyGIeCJdDvwqHjkwCgyc/d9Ez5ovbuReYN83X5bmhCu1KGQAl
njatGTRdPdiA0D15RUoO3dzYK0UdbGHjmY4mL0MAemkd2oQ0KpOldbummHfHw0ap
NZxB/7k+yArAULxNwflNnYEbuZWo0a5TXktVG2Wh/XngT4/DTfyy25gp3XIlCgiw
0psWNzM6JStFN2l7kuTX86MReF7rDmk8oEpV7znqtp7nHS6ey/IEAZ9e86Z1LcU1
f29/A5aaYtDirnGwL090aQ7e8JkoY50v3qZ41+/qiKGL1klJqStFkdj19TRJocyK
kGA/7ZDec2JBBbcTDceCQwlDTTbqUy1oAbZ+0/rU5w0z9243ey1UNm5/D5LZ17TE
NG8XwJEpQsKet3wHBZ35xkACD4QzRsYw60S1VrlERRVbvYOJof9fMNRwJnzVyrWJ
sCOEEwf69DO139pDc4AGfFFguSLWJyRFQxinyAuCOQ7n1GeNGLreXI0al7vgdMVI
A1ZVX+XJ9LPOItHJ9+w+QP90GXdF8Z2mCrcpTU2GuizvIBqmQ/BNzjQdVsANUhsm
HmfUSF6EPDKefXMulbydsjoRiiNZYZUGWbBLJabprteIqsJjpdZkNv+n4Dr2yinN
7LhQxALxA+QWTOOhViQspa0KqiIyVP0potZ1u7euWDt3/1u0GvoQpVdWQ8CoIbu5
lrwq1I6sYsiuOX07VYMp2RYUBS8fT6CUyX2Dze1mZ+qN2/Ge8hrrjZu88dW1czJh
HiQ72rC39s7blYOZxlTS61fGitmzrthDNGvbwY9PCdH1Ibjb+phyTcamG9qMCqjK
9/kdJEIuU3chA2A1Md2QX8Tgm+SRLGRefXYY2dY0coi4i0V5s320RndWjUtMkiL3
haW4bsmI5glzU/31zBI/kFn8JDjWsKd1wNN0ARnjUV8/ExhVNc+Ys0wLIrvy1R/o
5nRThtwCL3c7LghliKAHDTvixBl986+k3vRXyr2fOE4r5f5eFoLBz1rVCavjOMg+
gZb/KnS6FJfL13F2mkUSdLxQfkTNXK5y7ebXAXcvyCzpUIpltsSO48aAfM29lfGp
AWD4lOdLeLVLeTvCLdADWJwDox/Q+X6rAy09md0LjGuJxrkkaEbTg+GdHEPogW6B
AEcap43Kj8cgyN0IT+bwOsR4wBVCxnzVEm7pJz1YZnucObcN83pS7apKjrnKqDDk
X01+L+6gkeizVeI8lDdzg4nMfY+auTfFiuCfnKkOALDDcnNjJUmn45xmT+qHgYUX
I7ziVicKtf+P8ChdORH19nFj48RXfvS54e84/1Oc5UtZkHPRQArWn2u+TUDGDiS+
fUCA2cpND+7YCGXGt1i9Yamm1vaekV33RI6f+7lwQ7DRwdN4fsZFqotPTBUH4mG7
92Y7KrK7XK1x+XGzQMIgQEZMKcanN5mIzUvGLaRuEhMHja51z9A3hX53HslSi0E9
rRDXa0moQGN/JnUvWID5ENfE0f0AWmeiALNEfkh9JJuoGqmIStahTcSqt4wCi2tL
06ceObiu6HyDRWnQ2iqB0eqOGpuRrlpBcWs4GMQllYlVOwJcFoxzDNvDoWisP4a8
Cg1sOK04qmpu1iMnMA3bvEERw1lNzCwkGEDWpgx+GuVZg82QRKtNnWtSt7N7QKtl
CGrnOQGotp2xnHwyq8/5RQPWs+zHr6tODv4xEEarrKj5HEOJpAlexPYx/as+eJYG
TbhlotPo0YCyzeg0mW6uzAh8Wl8O2t2gRvDvpVriorEbkL00GoqN6FAQD/FpuTfZ
TpvhEMlSj2wu9BlIcH4F7mrzFcHG3Ew4wpikN4M/8jKOD32KjwtWWevjs3xIOTSd
PrBZJpSp5EYzEvdEBNiDnYJmzQjM+s90rHGg/YYukEO/9znFF1ufOh0GP+6MXj8H
Ajl3p0/9YXHXMLcEqVMB/gwEwCzQij7al4MV+EOfXdqBEG5Fh5gBg8VD4OegTL2Z
o5LYlla3agcF5rCNjf+PMUMZPGwsP4CTwsgBK8Hq9roeroQpBy73hJjPRWwZfJnD
u32+BVBqJwdTiu3tDsLLXR9YAsj6WlOeP/EVxEfUkBmZPfZ3XXsZOnqEvC3p3fnc
Ngx+EtDP982b1SH2Q3OQt53ng6ZADV/Zqx5o7Nw8hCZ2sElJtbO2fn5OkSzChMCa
AqbLWSZ0nPkXq2ZoiCWF+oYvjXrTEWLm1/QF+D6sK0j3Y2M0Mlt48PfvRX2Fdq/T
Sd/QrUxwe/CoceeIDehhPIamicuPwcuMLRyGY9Y8XRHWZuWaFPQldX4mMN03OWt+
Wx2DE3CCCPvFJDBBywvJjghKXhHGHmtP6wrYGDm2+wAA7zhC+JkqcLtDIW7lB5ej
MFozUcj2SCzW1db82zsWw6BgZ394NQg8kcrN474DL779tORqgLUEx6Mn93GkMuzQ
YKTwNyuQWDcDvZ9r2nHnn7AmsIXk4+vmywubUTbVYH25KbAUa3atJItaayv36s6Q
vbjAkmsvGHNH7fAsls71Q/jr1U7TViTZDpRQaYxozkWav//ZzuB20uh/vM8hq2Xb
GPj36b+bTEzhE8AsL5u2Q5sBfq5dviHGnx+OqtSe5MdigJQIQS97h+IjXYbSv9kD
rJx6gauLVmaQgFipFv1Xt68ISVEiHbRl85RoOctimrtAS8Frr9+hZrfst37VPf0Z
GuJd4JtJobsNQhWreRTILIiUh8nfyfx1Tp9SRaxREFBTcuTTfw9pl6c9YBRLkWh0
sgmnf7Okn0zJ/qrR3srFe24OD6SkZFlOyGifbdtLnFGNqEMaEPloDX+IyX1GaHqL
pBgBtzEI0Rd/4ZSBOckrw+XxSfHc8XltxjKtgFUw2BzWtHj5A8Vqe9f8UJ//kfoC
yXy1zGuj0n/hY/ZG4uei6oI5j+QMg8LWhij4j6KGKAEttPRUpShDb3fP+hRAk3Bo
x/h/J2Lpw1Ee5i2jSyhef1UE3o5pf4VmOyahbuLeeKhMkWE28ks0xsizxj6/ACHZ
Bm2nYULEMovIb2wgx8ZlqQGJP6hBDFCuXrBiRiYYOUMuC7aAy70lYjp79zvMN068
+891znwcvVZ9TV1sNMhgLFf0hOXbZ7x/OaixBfMu5lCkY6p9R9S6FloDptEVeJ1y
wW6iWZohjow+EIo9ryVLp7YtEiHI/OtZACQTZhFOWZhSMwchCWMibFUf8O3QavQQ
aTcGumZX8kXi+EIZG9qV4Q00QzlfcKrw3Ec+Unj9Eka8N5xOJ3r66dUm+VtRasZy
IP6sOEdgdFuW8re/T9dJSkoLYzapQoQGf+ukpfSIgk99XaN9D3XHqL0AA0H85W8Z
hJXLPXJ5/peYYqOD1Rb4EnE8p/49AAqWGyBSiGyUeP8S2d7Jjlj6h914SKDPCmz+
5BX/io0i28kN3LY0tXIfwo0WrwWf0sISznn8mRYLngBFam45Z9BpjXfeJqmJrmcJ
8zbRof3NlP9TmcJpFgc2+ZZXQDOHjkrsQG84mC1jmNcR+O2tg1VtoJ3MfPPgqDw9
pt51k4ZUlQRN0z+8d6wU4ybzCHAmFNgku5aX1sVQT6AI+X2ab0ZMwDwEUAZMZ2mm
x/tgtEHWILOLKnCHVSga7Cj+0FEaRj/xO/ezItp1DzRle1u/PuQb5hyrXxa8Yq/W
3utohmi8opG8wmipi7sMf1O9tP1sWNroC/YVdpA5ajgsmir8cYsjguBH68GcHXLO
lwa972oBNFyh4GXh46TkozNZJX/Tif0dNFehpMhy/+pFgPsghAhx/NTXLaU2lW5/
0YtrO1WBz5TqgF8AY3dJrIBr4ON3T7zem7vQps5TkBffq7c3uZmZ4r+eEeRXt1i/
qSZpxq2RjXMB/fatFQdk+E4F0rCMSZ+XPgUxoZV8yEKXZ8dKJL3Ga+UQWc+LONwT
3vI135AUiNtoa3RgwB4+0QpMo7RIx6hCEtJJ2EipLSAGsTP+j76oq8t+HPIZCCzT
M9DB+BvSwZx7HWp3GKyxEDvg2y4NoKTOZqHQLPdQCOnfE6Kkt5JkMCxm+78oPLWd
NA3UCf6VLNyH+4V5WRe0zK0Sd4/2EHnY8a4dMa1Fp9PVLigEEqNHPsJBWabjtEOG
Q1rxblFPapag7IC8c6pYXREX90Eez7oxB/4rVyJlTa4qqZGngL7g4DGNIhXqmfVD
PAfA3Q8Ov74iM2GXA2QsHI1SZ2bTSA0o9XQB33DSQu3Hr/VWvDLONPtOhgir3zcL
umiX73Jr8K02TZzUkZY9k/Pk/yu4NkLG109lS0tE8+4j0D7me3LA34Fu9oFkuyQt
36aWyK4h2aeRqr4AiQliVcV5pLouNyiyUd7zXFEbLMoe424ydctkt8yT8PRgNAOX
L8SGRDccqfH8ieKjlDX34OcSzWSuR0Yx7F9PnBrWrKrBXfC9a+0Ntn+PMMSU+d0D
BNfDxD8P2KvFOrhwzu3dd/ttfVwVZ3b9l4PyNKJM8KE/EaioEgydfsyeXrtWAo/i
ivICW3+J5sPTc5XINN20rR12IvZVkCeKuuQcIQuAVNxtQofS1PM7bZkUyWuPkWfL
v5w5xcHSCYtnS64fOFDj0Bi4jHZmgpnqa9QFfLM7OjHYfDrDbs2Vph2+XrfruBpD
11VHpLSXtmHTjzVxsv9M5M/glRaUzf6++3ULJNfNiZhHvJzbRo2PRWePa5WLiiFK
YNuaQwnoiyOExtfx1oEAjPnT3svdXDS7TyGfvwVuzwXj3rxyE6V8AvVhreQ8cj0D
EbDfUtFOPCOUQzZ21SWh+jc4GH1BQfFuDHUcP4hC50M5vv+hykp05+OsAXHCjWSP
oik8Ej+16SMhvr653FLExFQcooG7x2Wf5tDJL0lyOKPzgIGRp2aGgHGDCDGSkCmp
aNLT2sB/2kwE+QQcXm5ofISZCDs4vv5cxYUojK1lXfOYvDZci2RV7AX7USnIFPL9
9Ak9ZEK2rGPEafzNjqhv09uYLGJHat2cKwFBU71npEpGiU8/2ZxN5SihupFtzgvL
r8BoE8mBJY6AMK4yyiq9LMfT0mEmUNBwxpFxyzyCA3OndadkzqQ8fS1QDNcvtaa7
l0JYsL8qEiwUuXNR2FD935vTgzHGhoKHhAzD4zXHKFaStbColV7yN1og7+77D0Kt
DyHOhFwTIh6kPClcj8+kTspv7Sh2qmKMvAB7jgxV9kwxvvCXc/FhhU4xETUhqmz0
kbDvqIZ4+ojVWl7iBqXzj0szL0iYfiQ7w0FwOaYZ0BSqQwbIn2UVIo3GD8cX8wQe
G04m7i+iNtwp1fwX58j4YYszlWTE9PU0D020Kt+fGr62meBFxWRvRwzq1oQBRApX
ednLY+V8rCG0yF3rXsQn2Mlpfi9hUwK+RGusfDazfpO3ggSYoif3dFIekxjfCJyQ
wAlGfeEcqFOklp8O4wz/coNxIBsJUFUXgA6zZcsPk34NidW+g1x6qaQTBZ6ChhOt
0M7Upx1ecbZ05IXSjZreLkUT0vc4TWU2qJwrV09ZemYNde8mqm1nQIXGpKub8n3E
Q4TsSKzphxJzhfoju46cVepw2xY1aYJlLxMsEuQ/99VayvmNzV1lN3yIfqzP3ttk
ZPMypkaU8xSJDLBio9efVWVg3WGAfsCnRO2WehQtbqtkn7QcrjhaV6UZ03YI88Ne
Zh/jQFAPZWy3riINfadugHyf4n9E3B0COFLM2EicdQQeGxf7BiOVnhoKAAUCVxOh
ez2UNp1ilXtrz7WfqG+VXO1tPQI7MmtbNnYrlWokWZwJg5s26a2R9zS13f0AL3Xq
arCIGr9wRNhbgxAiotahuGXLspAmwo/lTpMx0gx5CpEVDvn6a7ULK1wUOPckwe1F
KkBrojSFGXy49bh05iy5kq3vdJ1P/EIzC1OGiWLY1J5BITQ208Xicu8UMLIUeQ3e
jKinVUFHV+TJ9/MYdnOlGfPQNzMLLeB3gY4OOsXFzZNCp/IPnVdlvIRc63Eew+La
qC38uwBCkxw2W1e6CeQHMID8hhbINUEvPzlSnCZplJE3JNoF4zVsHp9I1DXM12Lf
JOFlneDLqV4tA8hiQkiWbiC+z4V7VP2zvr79OtxZx5PxB/LA8veqWTx2g3iAo2E9
9kYyFVo+vc3tehbWo240/JqsfXwhY6OWwJ4TDJX7ZPMtnDcqAWqn5FjMdVrJoPnd
S0ZRPKxl/BW/kHQAzZtSrNA9V2I2ZP0jGo75kpcgew/QUOw2NEL4sMpHl96yjHRK
Z1HvAj2cweoppfV3p03Zaj/M0X/vGro/SpOOajevKU1oTjowPS9pXO2v1qkEkTkv
WnxQwOjSrYe1KeS4DG+EVOwz0tLG0+9u2U1FYNDfOedkLF78alQIBEIz4EAveHNU
OMHjFEeqUe0qhetXyR31GYy1lvdZs8E/pjHf4u0SsaDmRywNwLL+YAsbouyDAi7a
WObEg2Aa9BX0ki7fQVR4eb70dlK//uCDf3Y4r3gif8rH+oESbkmR7zi8U2UBomIq
hrG3CJzYClJls+DgEZyacKmMwQKQFyob/ZT5oNM6UBrY5oJs3rWaHIp7C6luayN9
RfmIdGPpZOl7BBNm9D7daotYyznirbU0wnA1QBEJJdFUbZpLvGuH+ZCN6ZmNmxa9
xMv5vOKB8NdPX1N+2A1G02Mz8IErz2OBOtEHwoKPAjEYQxsQVK4dzTZJ7Uz3iU1x
L+SKfZq/YxSD4rwkIuJmaddSoCdsfR6BkcIyGEl9fHvh96P6bf0wmGNona2YGN1P
306ghjsLd2hV3R7zFmYRNKKqSaePBKqGN/xJoTppsULQRERXm8bKaG4swn/E1HzX
txuxAq6780YzjC5/z+u57Oo9Ch+Y2Rt7sww3sEZFnvsiGb9iT0CdyKV8b1eF4MGW
tDxMDglnAS0FMyb1MTIBPAhh/nUQM+FnPLO3sSdfZOCaQRTV6IxA1YFfg6uNWhge
Q84TN/0nXQ5Zfl5eIcB37KgXsnXziaKA0lIoHKoKCm7sMeXYd7lFWhRgEAT00FXG
tQyrd6MQFHVAT6t+XyFCeeipnfAerDIQBWR1i3zWyG9FppRSfn0UuPpEFDO5kBvN
AxNZDfSXHcKKmqf87CtcJglLN9SAD0tfOlLY2m7OcGgUVH3oLg5qBsb6e47AXhaO
rcgoR1H3mv75Nw/IAQ9cemLBMgitI/bxLj8arjnc2U7pW682ERwExIMLam9vSutT
N3Jg4gqbD29qv4b6U9oLPFYARMgzN3b3PkhW7LC956Hg2jK00LuNRpuVW6v/CKmh
6vuXHOVkmJqRmT9QGEPnVmbFxEr/Z7GbIrFnrduwXxc3Es89cFcajpqJODDfdUHc
whR6YCTww/KcFCOAOxDCJnmGkJqUelDJVm8rsJ5Y5maaMlBbf13feDxZZuH2otip
3aQ3uTqIzQZQioOSVddx50LCHdFEp2kHdy1PjWIv/VKL0x8IB6TjSRajzO0VR0eg
7zhEF8qCz+ffjIUXLCYZZqtxkkukHJuti9qSpBIzY/6fZVDAfAwaRa+f0sOl3mLL
X/+VXxNnp5ZC1jBbHqKqf3QeKL9WiW+6Zx8M7M6/Lcs51wgRPaqlD6cUNcNWYbiw
ApuFEzMlRt0wTpJUjACTW14UFNEBkuGRFHHcsZPhgwTrHSAKv7Yvsomc177xw/kP
Ho4H7jEz8j2wEGDmAbeoHN54V196iDKMwOJkScJGApuPbCeEDUUxZH431QR6oDGo
t/hkdUUgPM3qT3XHYlE3hXKK/nUH0C88c/s/j3YmA2UEQfg3/9a/n4IViKIZxpkT
GGvjRV1U9L/L512xpg+DW6o5ZvRcoqkx77/MSvdh3DfjFTAnY6522lLiNcz5YAd8
UuG+gBomaP1cYRxs65utsmVhL/EJrEbL5C2GJN/7tCsgpfi0sdAnYTQfOUq+uJ1Y
S0BSBjBQq3tTvsCXwWzQt/z4qqirTpVR7nDrpnNdgl+N4KIe0YSZ3r6XaejjwRDz
nhnkSGHiYNJF8OVKvldJbxjsn3ZcSoShiAo4ShRcQd6Cd12RoRmgD4Hd4HPVszlC
1n0AgsyQ4euLzkl3LVfGxBYPu1bNe0XodBpgig/OvzoKgfBHo3jMCbPlE2Fqb4Js
fevkflbC7XY1E1aWHfUFw10X4AI94lACwjQxyIgh6dXkTysavAJIA+5IvRwcsnNj
ceV+N1BTxFpmSXVNcpB+GRzQaiYlSL58LzRvQZK/8iYUunyLABVxO6J0hhAZfQUG
1xWjSYwoEkLWydj4gKgIFJTMvUyvquL0bLRNztTsspfTyiEP1CYqsYs5ABsHtuyd
jCPumQ3Kx6Hlb17nRig9kVpCLLI+ut2yNtaijHpAiQMuQlonvYK38jTHPMtmAFcc
yKKrdISqgGTQLHw/i1DxawCJzlt9UuFNyfamCTzMYUdmH2WiO2Y/ciUsuKUOxgSp
kyfKaTKSm+BD7Km3OLcHKUi9pboO4PkUC/f+/YLcjYvVBmaDNlGlliqcaqeJI6sO
qxjR4oyJ9xemv4bIV/5BZO6cz3/YASKjNp5xl3/wN2IMIvbIAYffG5+maRMcocPD
01qfFf4j0pHQnGFpzkUf39xBsKjhk8tfHDz76hBaScZ5uTcAmaldtD22o3tutGfx
VfWTjYPK90ywwiocePOeuTmSt9zh3PibCCAcWwELw/wUqtZ4Y72Xf6eSDF0EvT5Q
OH+tHPc9PlTqoCujqRq+wbn3m0cp1kG59HZk9MlwbO8QPl2JhZQa4ugsgKlT0b6z
QgC7bYdYI3xn8llTA29k9g16gEKiVXsls4od7AIVgCTu64ppJgRy4ALB2cK4BnYv
80hI9xSpRGeFEf/Se+gX8iIHw39Lma49n96Bqd0zpd9DIvTGTzndxZ0QJOYHk+60
XdKR+2SwuM4p6M3hWQnxSE9w3JwN8tWQCA7en+gVky2pnzxXTOAaynfESaU2+IQn
soImSWZlyxoaWE35ZUgzltOFGWE3wKyLkTNKzguzwHFON7bAIQ3KSRxrHrU/9+45
7ZOwdt5rprguBjycTLJbblRsZVJEuXnRZGN0z6HmASXXr1wn7oZz7EqO5wIjp8L2
HIPt3ppDFXxEPH3EjibPUnon1ySIgRO+F+saUNaS011g6Lk5U+5ADJE7u0xrXPc0
JGDpmTi2t7789q2ITpzEO12ObgrUtWWd6MN41tBMvHR78lzi+kd/DBP88CfDE4o5
uFykqXrs4+lTDuf16k0WGCpkzfDiJvZGHjFkY94IgMmP3m+JNX7Ri2wMwngw6IpU
7H3/euo5Hld/m1xMhwCqMHN6GaTYlF6qKb6YDlpyeVOpILon/SGgz9hjhm9PJwm9
XM0HeVadguoEhHIvm5LxMwfVphKgaeACKy1wEGRhkomgWZG0Dc7E4zFgThCT/46z
t44ui4YssTPirQ7rwn8cQLrK8uNO+G4m2/epGUxSCwLA5DnONmGyjRm8R/oNLcrX
W1xvHmxeLYyts63xkVjoCCz1sGz/rlNRAKLkvkI0SSV/dmCrP+lMUvZQWexb+hAT
pfx/gJiGeCLgNuoYaH2wm6/OHgmyh1bEAKzdsL3skWDvhiXchwSn5tCuqp4YmykM
5yALwQgH0TJS34rfw8ej0hRiXFIQxkXK5vzSmT1ryUXV4L1mVTzK9bRn5Rr1CfiR
anHn/44CXUHk/bHP4AamfXERBZhBPqVvlD66jXCPj8GlA9YxDLmJpoMAn4Oh9JqG
rfQ6w5PhTdH0IDR4Go/FtvkWhvFzkZVNvogVXruhy7Lk4YWFmlvaEL326eZzk1XS
fPUITGCIPXlkBcjcuu4hsxHG4gvZ57TMg/UVv/3sf6AF4btGhzHacX8qUReEU5kZ
ynri7lniCoTxh3mRQlsN+qtwb03Z2l6I/CNZaL9lIyb49fMxWlEhTxmfFG/N3Ji5
QvmuVp97o2KYGotIRMWuTZp28O5T8DdRyWnbcYmQ19tz29gzs/Y9Le41SKt634CC
g5AofAE9yBVfU9ugJOHkYpzH9P+3BqWXZk+tunq9acNWADr9EHk1NHN73u0mYdqj
ObsidSlGMhWyTmKCJ4mZkp7hZy3rXtOWstQ8GBLP8L8pAuOuaN/2objpLkdAcPei
O0hJRnxx2XzoLQTeP78YxSLLnfOV1Apm38zjc749SIwRk5jqljAwBPjiLPpk097N
j28YrND1XYQBe6OhBhWrjwU5vonpufDIWCPkTx73xs4BdokygH3K7YgbGqeilPtF
dyBbdZgjzBnSWqo28kd/5gVWezFEiZQLKhvd7zRcitxgVUXx9N2TonLMkPm5IqXH
pEMI3k18u6SSLgBDfAnRZnrXbEmFDxvTmtwosXXHgJxT1rBMDd2BZ9NCv/IZU+pc
J4ZQvuIwleaDxi+lwZhy0yttH+2ZlsdYein5oNFC7en+WaiNBLkGbER2iBwXEqcC
dmnBQ89UqlpH4Jtb9E6H66/z503s97M2eSJFkva+I/7Hqq0x0OOjTx/yFtS73nG0
MnU0Q8XidMbO+K3kQkH9qZDpMIp37qc2kk1zqK5/lHAlWzh10WM0Yw5O7AMSZEcq
CMMZM115L70zLtqzot61l47gqZ8/wrb0uj5kIIn/pCX1W4g8c3KktWdfcrdG6IVN
CtFmqoBHFdp11Q9ioQ6ZIE4XGwBNAONpKM2VaSZ6a6bXvNugoWtcpqEvQQwJ1lgN
1zReKEq6VD/fYX00zPvwkMJdhIYMdsXVvBi1hIUtOsmRx7eliGqAXb/sjpkNDGeT
6VC+iMHV0kpqm/GnHX/nzgsVUiLw+hJb7jf4e4AibOnMjRlISwnG0OqaNZtUu+m9
WUv2R2QMazJEBcn6E0jFXeRDaQ+pId263GXWm41Atl3nmSnQ9e5iWjJQ5A2hqkfO
vAAl16oNGSwiYNCiqglKJpmQ50MTip0CvnVbQEPNwjbBmArKyOi3XlI8aRn7UW5c
Ozzfdjzw5NZWFVDU2NVC8hPZA3bJBubRV4uXzxfYYRgXWSzS2fGelUVdSqw+B0TE
6Bc1hiJCniAwQ7VzUHXXcEqyzyF1D9I+ugD5Wyh2+4ZNN87SGA1MKhwWZ5YNm9UR
2/979g92sNhDdSXoC+45oedPP8Sftm2hdARi6OAJ/A6i+MKfClhr04pAjNdqGhZR
fa3JS96cIOWZO3L0Ro63LhnZG+n3LEhLxe415WLHvPz387qc6nd3BvttkqB9+Vtl
NvsZZCc0Jtn3N3NWCz4h+dO/AB8VNCWngeXtI2oEuYoR1SDUudM2n2AKO8gdfAlX
ETBP0PNNYJgDEEb2BRhvlHFb84mi2UjtHFqIs7Lt3EQpvbnGJRUpmR7sP/ToQjTH
S7H1aD4D2ExfEDFtfWhORvc8Yk4YSHhXW4/OX7r+ayZ9QrmK/V4OEFxL8EiNujjH
OAT2yNowmyIeG2Hc+0uDv2n1W/vGI87n8RwOV6Q2gsDaby0E2Y7wdHosoMz6buF7
gsZi7Zu9WV9XRnnfPggJhAOGNbVMbzg9PEuhzn3k5NbrUV3FaQU3fw98ryLQ51k4
nTbnhsx6suJ7TLRRERF0hQ25I09vjax75F+vQXGEZVGGHr8VZAKKqswKYrCbHulB
ZWGDQ3eFTt44BPjothNAgmLOzuPkW/BQbFfa5z9yUDs6O/Tfy0BgVcJwWvlh51Yj
uXLunTJfP32mViZA9ErLTFNgNknCuxhCtuyR5JtipLpMKfDmSVoItPqDxkZzpEx2
2NWSuUIFp/ClWVVDp0AoBoPr/MVblOABvjC3uFEq5CfxF5d7ej9mNPk/iJ9yIBC4
mtcYMlMF7pZv8bFfeFF6uMYH7EmpP4P9r9g2tXmxPqvjY5PPt8nZzaQxb5IEnz9/
M9Ipl5MbLaYOHHewe/DU7nOKQlneNFoqptWraBGXuivdeimZdaLDilXDRQIQjvSr
IBp2fN+EC/fNaQMMOPzgMCjK5/yQa657DB29BQ1B1pngvkWiO7d79sJ1uXJyvqZi
eR1WyO1ewbi42yVPKuZWG6bP0+nK9fTwvlJH8hju+2l5qaMZ3BBFSo3weRW4QQS+
R4s0aKkOwPq9BvuZ8diCRlvrA5zY1l49NqfePClVCPP6fhGO1NYcqRJeXtvSaBhy
lbO5h66gGbBnMJC8UOIFhtzUvCIqmtsrJin+6Iq2bWfPXXv89GDoO/ZOUFBpLbPp
LKF5Jp1nmllS4SFM/RzxVcBsYKcfD5cqrVZ1j0bPvSnfR1HOQZpMljvLMibnnNrr
y22ZM6Wd0wSh+N5VBQxK1LekyoUNLcTuMiN5bCadXEfoI6U8CCio5Cvwc3E5BT2h
0aSrCV/TNyLjZqn8KB9F6cGDdsptetZd+mfEMdtDVO0+OJwwWpGShdzt7RcLNYFc
FLp8exi2HSH05QgI2fFiGGkR6ffMD4nYOoBDqn4kJsGBPAl9UdpwNE/EVAxuRuO/
6ON+35JMogmvMFnG1IcZiUQrrdJAEVYeUi72DOdh1JIlIVOBY3A01prgxK5Sv7fT
Cl3q32MHSW5HdcDsTzllk6l9BNY2uqmG3QuBW3BkFX1g16EGuGXYHwHZEnlhoYmn
+xZFoZ24Tvtmze42w2P4ydB9CzTdkmfMx+MGG9WqQXamO+xBRwwLwKaeqAosG+jp
0B/24qyGRKap9UJbuZ03jmEj/yHthfUwvvSrib0NkrTznQrtcDlpqVfz/nr/mUH2
MVkjplodfCNvQwHNVl+Jp00Zds4d8UBMX9dT9nqx21xO6qg2LNXx4MCKynZN3q+Z
CXzTxY0SiH6CXBhpMEdsUwFT7LFkFyUsMJxn4x033SBrYBzfSm0lenDcM9i18Hup
0pQT/hjWqWf+8Wyeo5lsWEWADOX/eHDPQyqTm47D1LA4Z+JhAdAKz8EVDt6DTJwy
Tep1LTD1wQ6zYf3U6jU3bhipRfRUmZVNVEK8OfdKLdURaRuLU4ZqFqFpE1Ul7Z50
8n+H99n5NL8efjmutYzAxaQT33J3alaaeDHgchIPABMlyoTwHNN/xLPjMIADqkFJ
B7tyFEJX+6bohtcft8EMHAea1pStMcfjwbIY6gPbUOedOiFXjsk763SUUNaug6gV
tQxird1M4QHp1Yfa1QRIhdx5/IxiyplwKdrxJzkpXahMmYFBcV4Ma+ZohD1jhF7o
6JHLCZD6yf+SFxEcB5UWtCOjbcfk/O6He5TyW9NVrAGdxzstSbwnuhp22FWXVrWF
Rr56htkuwVHJFMq20tKoAzrQstI2ahdEl/Fqv9KEhw7pLDzBIDRM23Al4CYO19hu
LRNiCj2AU1SEpgtjtbbpjWvPpJSkYijnpv/uKKiFrfz7rsP/iW8fVwMMqShppX56
GAB/u9CnBrNYt7mpwsMVGisERQw4uy0RHSZqtqpZN8hJheT7R1qlo7GpP0tFmCFn
koN0kVrLzu4dCjF/JlyCje01EBLz+2PZuq+tHofgyu865PUWbXRoDBc3srUe3irz
vENi2EwiqK/1O1X0a8uzEMCFvD9WIHKMWHIaBq+sZHeb2dsKRpJZAInmclRPAusk
PCiZLxQAV+Q/cSHSWeKXKusuJw3mZ6FDg8Z/VfdJeDEpuAkUv3b73zoI+pSIUMpQ
sYzIltFPPksKDPMj9IQ2cLpRdB1PDp7zUwRQqXrT8ACeRsCaL500BagaJFm1oPvq
0blDoiWN1Bq/p7Ztb/oB090Z3xvVEgbJkuIBl9SXStw3Mh9tJSiSrZ/KgYQse79A
R5oEGhgJjUKpahxQ/DdjR+07Ph6V9sHNlWufAyVgCz85shBUXOH/2zlM+OuDGKB3
k6OWrXaO8Gbtb1WdiFiNUz8ePr6DmnhnVJAFwQCNnuFhfBZgnk4vGJ8T/z9ulsB5
z46Zxog/cblfCDLsPFzQZnOUpnb50XV507QgVWF0ocLaZv7PDPR7UdU5d2BE6xaN
+MNw2phwyQ6eROWrhXWNTv8tNLQaBoiOcF7sXSkJmK4A/4NBXPoSrN4nDXpojxUF
2xxemI/Ot/7yN+gt/gMLVJQO9wSV37ExpN3LWBon08Zw7Ri0VgsMhRS3GwQaL9H5
F6XuOJAUen/cyyKw9RYXlEkDDjmBPvA8Wlfoz5Ka67JCpPjTO3FrQib/4gkpyN02
6DPzI1t4V5FtAtJiEoBdxU/lwCSQj41zSwK+YK1NsZKz3X46RHbp/A6JinJXacb5
Ubd9wqkkPrCQaP0itzVp+GnuR5Xe9PfWKldoZfxc0nP67IBsgEtzj2+AG8qc7hIY
9dT65SeSE6DFM5w1Z0/BShMGSyzRHhi+6eDcpHky94NZzoXvJYHDVUxf611AlnUt
9N2td5BXVJGVjlBQN3xc1PY/FoqUVP5ZOvSAcsY/klSpMhmZIImj3hvnKGAjqqZJ
UP9n3b7qb3pm2z79tpEqjnzuNE4Of0987e1yGDP2AiDVo2bF1LrBaaHGoFjV61xX
hlXUijDgI+r4d7TRpMoC/HzrnBYmMhOVzL74+9irYUd6csgE34kG/mmWL8q+Lne5
nopSjSQbUy0fmlREX/OTT/GSFChkQZk2os/9g9w/6RGQivP83ngGm/nZGAsjdbXU
RWtNGBCU9ABe3txn953hPl6fP3U6OY2yNwwkBMHbHBxWdLghzPIHqkE/Vps8rwbl
f9Uabwl31i8AHgF00q/uXZYeg6x8r9yIFI5lYmKKwuErnp4SPVlA5+P5A1wUxYYO
57VzSwRDH6KhX8g5XXOZ4lmsOTSXv6IE0cYNAhlfONnIOYq7Ga7vcU1PH+wjDTgv
9e4xiIATTiFqFx6x0f4cAEr7mGaNhMdVgdW0Tx75sPRxhhEJGfCMDlIKnc92d35U
rmxWRYnBnCLZaw8ANP4lmfQqdLsT8w4yNr+V2je9aD2XNQ7duK1uAFBBABa6AhxV
crXCkdBzR48A1oE8eDdh25AaVuqkOL10a22a5i5ROYKhpmK8MvVvSGTExSl8wVSY
MGI41UUcxt+Rw+sggXnf+AQ3h/jQNVgv40llS+KiWV9QZ/DHQjOtytmWolgJ9gKM
ihYDPEcXLfQCzxthXupxQ4UlVY6vRNNhJV0hA46EMAdc8jN8CJOTGUlHSbkr4m3i
XgosPN1yXUDorcDU/C+7+o/CX0xbFDydLgsrY9Lfbc1j7Pjk/jYKmfV1ouLnRBah
LbqrOFhOYyWCP9ZaM0kYEejQGyuzMltbfRImud7npQPG9CgWAJUHbaGVO7nCl9AW
0q4QS2M2WzfGokVBnW2SXvtfEj6vxGVYRQgiPxwNPCQcVZ7JlLeyHTw3EyM+jdGa
Uj687GoqNE2UmLP0tSyI+RuTiahU3qdnVuLmqe0n9PEhpxCySc8R5OQ3o5bzUsDD
qObPCig7vCJMCr20o3yWL/21enxn1aEiNfuxUk9i/uoQAdPJRcNgLFzKSWeY1pjO
cqBlaePF6KWloq9bxoWjkldBjDKF1XZ6ZqkIEIoVhtrggRUvUmZbQxV4zcC2rHfa
G7AceE7TKa8AwXlqS7rRW/+FuF8LS4HRxY6STqZDHSl9LTH7b1nQaTiynbvgSMlv
alEIXca3cpYFX+Pa4OKGLOgF5nRPMvlyXije6qlv7Iqj0Ecb/pDy1CJ9yQpJOln8
Qpv3HEtg69KRE2xuaB/7EykNWeYoU9fC4u7oldypwHSJGJDHQoPOvxycqIXNfGXz
YK6kqD8HY95q9W/NxoMSnDMF7wmBzMhyLFxn3a2l5IAf6a1EJIhK1l0d/Da4sTes
Da4h/C9tAoHTQE6hdHPqO/BGyqUh0tXVt3V/T6RyNtWi1SLk1DJUEVuyStHChoWA
JZ51BikmJKuSeSL7PsjB95/MwP8GJGqD9LgEe8fHE7NkCIGNH0EAzY8hDPDew59n
SGuE2qus6S5jwCITPygJVOobaHc+PtJQPBtFQlu7uSPAa2oiBkRQ5GLNrwarw+Sh
mAwXk4WAqEPD84caA7BdRvKRh767nerj1fSofNSTHq8vhrqZO5A5FE+u4vtVzBSY
v61lMGTqTtQqgGn9IgVZaLbInTPyOLYh4lYuNOvxgHfMGe/xQ6qj5RsMZ6avjcsP
lMgmTBd4IGXvDf/BIdymXdarfSVflxivLzF0EP0WHH0dWjzA8/TTpqZe90qX20Tr
eih5SES9+8ybpRruf17dAMaLOJycS/MH86RoiL9epXzY/xygr+8EOG9EBL4mxGZx
y2EXJqxzIXyP2dgwhKZTuKvbNEWYFNRcExElVjsGnhqyp3h1EBWCyhugbFCdMaMS
LRU/Qrjufu5eTiYckz3UyGUVQ8H7UFGVrSbtnJeibX0+96j+2SKIEOpoWr7p2yhP
yL5QQvbDDdqMuPghG1fxhhkhg05XQqdA2f/R+VDWabUeBOJEy+pbyR84/bVWYBsv
FzOaeyWOH/WDLdhxeXeM311tbVf4QjyvgPXsZUcNT3mYNUXs/7VB39FRje9P0Dhd
nPakGVC1XgHdPoQXGbIW9jOPuwHQ7xMvHflF90udv1U+RbkuQCy3JldZcVlp9yMj
LlVw4eE2DCxSqCbX6wcj56m1mMXX3cp0/dg/zq2PbvCu2B4hLH79SS79M/k5CNJ1
WJS/BVlETvBg333qSPrXBtG6StZuROQD1bDVntnKmhSm4wqC8iXhTCo2e2EG2UMf
8Zq6q06ehBEC1psDwhpSVojIYWFfAMC9W0YKC54zjo/6xOrIMx/DmQ7LOQzND8Wi
10H177e18WUEoPNiSwGKmZWzbVJuHBKUTrK8A11X5pPJIBrqeisi6JJ8OdrE8gGo
CkfhkmKLOnSGhnUUbPEZX5VypXaEdbInq0Jq0sqkwVhjbtHvlcuUYdTsWkZnK0fu
7BwDo4o8zgISMc8sdpRBtj5pKMt+9ym+jfjL8XUYj9qRN5aPDd66zW9Cm5mMKX+R
SBLxXHMxDQ4UDRqEIByYRT3owjtb3FJh3AIlLzh3lQvJmn5I4+BjVqyxPCuIocsL
IrEYCLfBCQv6Co/CwXdEG9WkN+5g/h6BGW2aqoymmhKngdYoeS/tnoE8a5Z4FPyD
WnLpGKfxuIh1V/0/u6F4vNT+FVhuMq+i1mfBkmdeWmKUVTrSaCGEFp2yBDGkk4L8
Cd/6cukeZ0Lu+39Ot2pmfTmYGFyQ5EHm5RCv2ZY0wlBFq7GKUcDlMEmeBNlpXUf6
4cLbpMncHVvieUYY82xCIXrD0TTboRc5ZcPibqBU6B7VH0H6HmN4L3OKsiQkph5M
838YZSdxGiKsyDrb/LF6gdqogX1HExxeXwt1syYverark/RoA5kz1ND4AVAwApFO
G86JITutnxc3la90spkLMhjzxQ+wFQpy7YP7dGSEcR6r3MbBwV9TExXa1IJVqeYm
o7utkwcyHmcXXkud6yeIftGDjbVCqHyR2wEyV7zDdzTh8UR2CD1E67IURbZ8dMpd
oZrv0kYzKltdu1w8SFf5TM6jIU0eIOxytD4Nr0ct15wTAxbezUZPl4ja8FiTY7o+
52VYhgRD2phJELZyGXtz3DB6hFoFLwXNfHw+QI+tF/9VyvxoC4bpDL3gPhV3SPgn
eZLlQDP9yO8yq6digNfFz0fykuNJRSw9sMxOUx+qJfPFcoXpIfuCHSerjr7U8YNw
fqdn4TfpNj5rb/e9N0J8MHSw9hizAtLrXfKuFmUAjQnH6opJRhS6k9QuMk9Jdyft
/ivfTpzqyj1/poEIzV/dkVYp0BV6+0al9MFpZ2tbyABaHIYuJFOoReaafDFKdBjT
5Gc59vBQLR0geiYHcsgkEDihh6I9VOwdwUKJKUsxGC5UGIGvZ3YuP4HiJ5YDwNNN
GPgybomh+9iXh4+pysj6WsQ21TL2nfjhR5w4RXVIKf+bDDvYVWq0DDhrAT27hWIn
1qTEf13tuO6XAAvrPIQ+234thSKu1JQrLbFbNUVieR5n2yVq97ncHsAXQVXcuLlp
PMgFfpNS84E25orov5ldH47EFlpTn0o25i2/A0t0e8QB9r6lC1WjSyZEskEa9r83
TUvKcEf/TAhFgE90meOXyZ7Sh4fCrcpray0T3/k2Q+hcUnH1ixwe6+x40glD0Uq/
VJDdjgo+zjU/RhfGsAPKotOqzvOei2Siy+LAvuU8OLm76n7aeZoNCsR6fyztysV0
QjKIH5JQji7DUiE/PLGbwAIpYrDetm0Jwo5lXWSe6sBZ6MYCYW/pPTbD0xPiKd9+
/nEML05kTnIYDMOqC5xgVYcz2y48BNQfeAvfZr8G+aMPtkrbGwhUC9hGx1O3MUYI
FoQ0rfP4D3WTzP/thwLKM5zE3EMefSKb1Ap6xBdEj1JBf/oAS7iJIbHhqSTgrqrs
648mQu+36bznx7MuW98nqxqeuXCUk2PYsVpxdi1IAxIcOMSIXEe6J7tve6+be72/
ex8uRtgUp9Pj1v/RaUKdJv6RnfOhwLER6wMJLsdZqE0AYjbtCWGE64yrQ8+GlSBA
h1bqb43Bpxq92CV1j0REpiggIwcPtS3dJIcohDbb9HCwZZtJqpOYNP3Nxv+u3dsY
9h2tr0m2OiQf8WvluAT3EfBHV28N1J0H3nisx/qzWclV2FahegBLHQS1L828XaA3
YUURclGQSrg6o2kBIbYsvsK0UyYtF6Y6BC2bDlq0U6DEBAsZtQGMUHJgtM2napmJ
icoiC06otSEZYBnff25GQISlXh+sIkiMGQGMAzQ0lztFy/y98kNHVBj90LNbrskl
WKTd3z8mn3brzeToVh8xJRSnb/tLLjMjZHcQd5HV0N7+PH1CxzrbXGHGTlOMavmN
qqNaqSLla4aYhqhsIO7VoOb110ipgpgJIOY7bBaXPbQRdZKOnACwM+u3TguyW7Pw
lR2/r2OlfFxLZfhIPVcsajja7zwFBs4iIV5kEMDxHJjYHCdhq+fd2KDNYK84QFP8
L2raaCQWI/EV/xuLMr4gYatKCUUNHi7PaOB0eIx01golGLprV8XaJpm7A112iYYX
I+FAoonnFuvjm8JrOHWO2FZ611Qh5uzhx8wxK5Nlsd1zSHaYgGBw+6lz6HT57L5d
eHiXvXfWc0VuA+bDejI28W1fEpE2CZsoZ+dZXXA5Xle+a60LR4W8crfVB4w5/saX
EeDl2h+1oT5PgjFUxHMQ58WHuQU4jeWTuwPtn7RBH4WAgJ10sNPm+ivRkxkinRHB
KF2Q4KzPgMOT22vJZkOIa1411bioJsvpzKhBlo2l3rMDLfeqLZHBrDOMuPgHDIbj
L+k8UGOGUxjUAuTGcFtqfF6PdJOw+6uynEb8MBiAiDeCJqF8fvK+Qx2AU3KhHqM/
21w6hAb/KmTaBgNDYPkFZDw7tASDCLXNDqbLTjGk60d/ctRcIOZxYcHa8yZCm+9l
vVu4IMnza7O6FkMP37+1gB9/B3p8ee1wciH+1x1gYyMJVi8th0k071n9Zew0g7P5
VfHgKo8tFnVjeJwjG6E1LtPl/q9rvJUO06aibfEicWlmDxVDdFdwWfz3x0xG7DZn
yOULXujvJZHW+HLE27peoN6vPhcMXwxeukKN5ozPmVBEp/Vzw0LL6yP+4jPYr+nY
6NhhiEz8HQujhrbydNN5AfjjV4X67umBXf9LE59Kg7Ky8GYatiCz3n16Z66K/LE2
BKoUFSFrMHfdB/su3Hyyjf6IDLVXWhtSOKORHVt5WakGTRwsneMJjJi/FqbEW19x
EeGrSXAmJrd6qpGBqdVtaVqbZvfpl+lPOUz2s34QgWy//TTs39Q0j40EIfp9BO1q
uZdwFL7KTkgVg8yac1Qu1gGyOV4Bb3QUY+hrH8/iGzPMHfR5l8ezewZet/FaTTxp
z8VSSwrjEluv05ye5BsAZ7AF7MkIXFXdkL/BEDZtfreQ1IzEpjOMQYxXPilDFalT
/aJihsVPk5NQkwBpiHejnD8x9Fs58ZETQ3X1Ek5VyQgtnVZIlUOzDEY7WexGn3gg
K51HlTKDRv89UffHH5IcAftx8M4QDF/WtwX/WPfOhThgo97ClLme3pVU3MCfHx9I
Aks97H3kIslcit4VDzQl+GcAJ8wBeh1vgfX8PGj8HeeqTgocTIjtPst6Xlpiu09h
QG3vIBYDA9gdnMV6o2ZTqGHCPLs+W+JraDbj8EFaCvunLQO5thRvvVYcju04ogsH
rkMyNFdJONMgbQBwSY0WOeOCaLcTqtIoldQG+FxA4/BaukQ3hwJ3RSjRkYFeOsG2
x8f3DrnJn6MgxkgtduuG3DEdwya586Lapt6F4aFw0oHr2Gw/lI8v2CYJxtBxkF+G
Aoy9a3K0rYVDpQOI/VbcBTGMC+kHKc3tR1TWAT0uQ/9CX45LQdcVDRtOidVP/lhJ
LcjUDQ37nCVfFK/gD8XmZD9nrKjMSZ0KYEN1naAJ3Mwcav/a1jWT8txJyXwTUytT
ReiCSjZucSSHx1Y7jPFEX05BORcakhP02lA/xrNYcw07kM68qXKpAy+EVj6cH+Hh
nMXqVEs5hVRnQzdJ4dAZOYosZFQwTl21XI/bXu0ZrIwrKOyFxYWWtpJP3pszgPZf
++0M+woI+5EpjW0IfD++8bIFBRIuFTcFezJrGmKQ3V5mrkZ7kIPlNl2AyyHi1WK+
nrSke5mElrhK625FfkTE0uqrHHP9gCNWV9RELHjA5swRelss8wuXyzQCBMI+necA
aeqIxX3zg6boaufbeAWb76w8W8pEVgoiBKYOfQvurMFQTaptdfE5BhlVUTnYvPeP
Ig4rzncN8B70l3caBdLWX1ucjgiZYSSyTntmADoitfupglvgd/AZ4dglHsP3tz5s
0Cv7duZaWpqjELNtQt3WIIJwWfcbz7ncVDR9uf9EhYhC1Q4kGQRbDNB+A2Koty3m
y2vGiyt+GygTG9fk0mDPjyTXpDyU8+3MSPGC56eJ6XUBoPGUbEo7+n3x8pOub8sZ
EcHYUrTNJGD41+9AxMND9HcfZGk8Z7eNyPY56ZuiJXJ2oFBFtC0TvWN+7hdkS6eq
HWbBfEVAtaDJ+rzxpQ3I4gG8dKBhv6cmYtKFBJVZjw6u2wzoWhtFd1u0x/uLRtcu
OOWiezqlwUYVitkjTd2F5YalygqKUYwTSv0IVEk9wgvDPPb83BYoz6Yo9KP2B3xF
L3C+S++IQ7rBeR1bxEsYyvIiS0eIUGywV31U6QDTBEPbhDm+mpCho/ICO+h6ByQq
x0JvPLBM0RD/W9b8ICfc7V8oLa99tVfsJlsLD7uG/+3Y1bgYkZ9kdku9TKKx+Tj2
cAmJyPs+H4b0LqeVf6DH1t7OdPMu01WBQ/9gyyaWjWMrGO6ngCdQNo9O64dxicS7
ZCyFeAlY4kIWsYuNwsU4XZOIVhd23iWIKTd6IKrHjzkauJVGxLzV1Ytk3cDAS975
M6Wfr3lIPTgN/tMbTjzC85f1rs1/Oim+7ye7mk6ehjfenvvwcvy0k13AtkTWXRqY
By5v+sDd21gRs7DxGsLpV8FvstUrVL9Wu0wqnM+st+unYcRopu8son/nHf9Z9Tzm
9PPUz/Y6Hl8BkyB4kaCfuAWCr/YmVbqdMtq+XuLzyaWUv6RCOniy7dElGew/ljA1
wnydulIpHW6l7PMVNrTzECI3PNRe8sEnpUJnth6mQk8iICGd7RNynAopWLm9FukA
VELmIroQR/eJqrydMNAStX203gjYyt9EOSSgIizIJ+qceheSTU+jbjW9m7dc6I2i
JUQnf3sCUa+ny6i0Dw3AlnsflzGHW/COLi/1WPrRbGT9naYZqgg781+T7Zf092w4
tUayFLlTTJmjLHApMuGspYL0m7kMVxkLX1xcRwpmPSVxI1tZ71WMaY8XKUeLIOYn
p6brGz++1djuWqiriGSR7ChqETUGAQ8oqsn9QvexRTuSBOBiUAf62ASQ5EimuDov
2qZS2ZG56xLxfGjjJVDweUnjz8KQVfRdAUD+3Z77kchCP/lB/z/oaBoBh4WRmKdw
h5eBz7QIVtLhaW1WCWJs5vj9EokplwrdaiBjjih279pq/iPms6/21tj5cbozqkAI
1o0MI9E+I8sdnf5b2xXX5Wz+ZHhDYq/RZKPkcID9qp1zvGFxh40yI7CVWNAjoBof
GJQfb2feRXS6Igvut286UmfGET+Kz63+UsFdPtZyGvYZXg35Jq/1+B3VaO1ikcAL
tlBaGNDi3VCjs9PuFyWSU3rHBT1AgJWDIp9WCyOYKJlOD7hNlI9+ornZCRh07Zc5
e+Ilny8VCEktYABlmRXofzB7aQs+LA7nnHkbVTkXj2KeaPI38suJh4xeg1sBBl4c
5+wdkWLIQrYb4da4qZcFOhSGGK9ji/btWIv5kQyh6eCIf/pXASWbl5qDFQobP+6C
l0SiReZ6uUhhKmE7oilS8dLXllH1QFL0rjuGS1mkN7XnRuMAKpjq+VmUnw3y4Em1
R0aFHxQt8KMoXOYNdhn/uQHAimQR8C3fsm34uKEGBdhzgKxQwIbjD+cnuaiHGOa2
g9lM9WeVgZbsMsGFXenLAkEOt4C1DlpJ6gJ0JY1yJjQTqpIKK2/fxqkd/6NzOIOs
IReRfbdtQHIFxxqHt+H7oMs3nes6uMHIvbzLuKnTR+GH3PtsREYrySx0kFrnxvx4
2ck+joVBWRFc08u+v78skBfL02WlI+8O9ij7gF8vU84RmROPsOHlkGCiQtjwQiit
5iJlzcUdKY+P8SXoFRPRP0R+hnAvbROp30hEs+ZBipqRnnZLh3XeNCwgC9eNwUz8
hj98TKd9PtJUPm7cvN8p1MyRp42bulr2v9fq/WldAhCEh271wohy4KZjVRvZNQRF
Q9/YsuxDOPqs9Eruww+oVYFejjxLpO4En5RwXKTaWWNyyzrKdT3b2+pAa3XVoPY5
sGMqlLr5Ibd4H0AZ8ujzC/lbm/YgFo0u6epBX/T62ciP8sc/QHH753ZrRAs7KDis
C/q2R3jSohT/9tTTZbIQXpXO7b8qbfrk5r8LmBWB9/uAQYlDTSrleRSBYqhD/cqz
aYD3M1uHU/RYVzrh+wsnv7djCp+qrF2OZ82KF18QwEjbn+tDRhYDsrHjmjE2Gfmr
uaBA3Xh6Tw/d6cK6mrE5ev/jEQ1mQ9k2wULf2bb5mWCJDNaaFcRY71iMM21DYRzu
18CvH1u57UbKaV8v+boP9JiFDkimwi7GC3cuQfhl6vgQvtxHphKJZVji3nAnhSxL
Wcagw3fCfR+dBoNeNvHUkPXFuMUDTPJ8ilxvtYcmHBQPCx9Z+JDXO88baBdVpnRP
fCertkNq2wn+3swAaw+d/sF+wUwpokv9GvjG6y6lgIV7JA4CAeUfpsGyF6D4zsP1
ZOkoOgAfdfHTkYAm1wFQZelxPAZxGeYFV0lQ/4J5xDuJkTy0zEGrWFlIyZ9hCMmc
R1csbshww/qX3ymbPpGGUbj9t+2/FqtdbihOWofBPOBxWjAJYBnKecwmiODmXTa5
NY/eE+yqqgVJHCPMRklJQLavnD1DjT1NZRqiWxiuLWUhAh5YtVr0yL0LGywgkizg
GXDxpoZSkGm7PzZjcmk/bI+M2cfm+g7l4qc34Vz7AFJjHM9u3UXO5m/dtqtuh4aY
DS3LBu4imnC7FiNyq/G9mTJW8nS2gL6yTKbr+sMFyKQ2MOlmpueaEMqebMrrPxQA
Lnosdj7rWEbMr4p459UMIQ1XgCpTsKBbNAD1JEDmsEbBOnA3iA1rrfbSAq5rtUDr
HwJL/DoAg0jyyT6Bt+B7VVSfvzSFE4Z0Sk/gRqAS0Uv+R2YthbdnE3D0EIUI8nVV
RnEEVZ6yDrHybqmxTt9iAED1F6LIdQSRHo4qysiYn4XmvrnfKZ2RMYFoBMdFWb6h
A0RxN0HVKi1FAj/FV0Xrj6IZTVK3FBsIAvjBQLe+tq8K/nXzDLf20WQ3m32vDupt
1+7KcjH9fubZWwBeLUNJ238dKZTMn4h+e/FvfQkeBJKk2UgqImChqq4q4lTmhLVB
R1fJnU/secbpjfRgVZqzyOItszsjr2k5N0mIyQEiSpND4//7T0XmufVnoE1PBcDz
ZmoNWJ9tHUZXHKCAhY5B/tw1Yn0Cubr2Tga8weAozgVYSGMZ59XDQrhWDsehFiSf
kctJwfYinkh4s0dQEeNKJYDiZmotBV2jS6Jbhjhf9bHUVfegYoJkk9mcmc6kcRZN
ssQtALh5AVmRSudW5OlMEzpYmWdP2dWFxZpU7eQJ21zuvl2bvjhY0ZUJZTjQnI6V
tjUdF/nRWeKc6rgRgIMiCa6PBqydDNAImq8abTigouly67wS66e1WyhXngLh07MG
wMAFHIBv4Rj9IkYDuP7ih6UVoCG+sukgtF69y7cFUObB443J+BGdLVAt8k6tD4DL
C7uTyDCNstETSAE7f7pFqAwVj3rHY0Yv7I2p7k3M8lWQD70K3EwPl0fNns6AHdNG
zX+2aB53L6bkM8wh0OricyvCrsuJeuneuMRm1teMracnnpPNVW3r15BKfK86n1Co
T2M5GfTS0zxV49fJqeQ0cbcP3/4mRAOXuk+XqqW808ZiFbLIvBAT1fPVKQWqp8q+
oGbjIcMik1ZbqU3bZDd0ijYML4PXfQTNUC2VV8RQcdupbl+sfkPRMlSuLyKVw568
f+ZrQQXIhDe9cxMsD2xr6EaSucg9uBjz05s7Y4M7ZxMAObBbVfWjp5izwq3wIu4N
U/Egf11fZ+6ca4Yr3klz3HCdAgmBrduC7JEX7XZNj6Nl0aCx8Vd1urnLicreiy3d
EqnWs4Q2/CT7AKfSzLWHmVZfViGWwYA1kd7XUQuhDcxjUpgz4CSo1ExF5XJUxvoA
qFdUtnPmWHv0c0643DCIayzxAxgZxwF2vgXCroVw4d/thFRAGRYGTEVjZXOabQpm
MD0/rE9EZ7lX2fIAiWqWsom9PUHDFx0a0VLUEDUdSnMo6QivZXUPyuzA0P0hEfnM
YyLfpjOEVezAH31/b3UBliPUNXet3Kkdl/M+OyDcrYI5isCPmrJL8Kh2AvtaIUyu
0v4Hh2E4JG8kbXXF1qoNro74jjYe+srD8GreAmfwInqcBi1kbwAmoXMrLDf2DX/i
eS2aXkMul/Rq9TFBAhbeDXh7OXpKpHlLZ5GGc+N6R3EZeEIBXgNoNaM5PZhL1C98
FGQ76hgblh/e0Xis/TDtpcsdBhK1BOOwJbRYfI+8DkOUmq8btp70vGTUnny2Wmg9
uz4uJ+khcpxVKLUrgLeFQnwHxVGytj5J4Qakfaejk/sA+wdHm34OKfdaMN16M9ma
4TB8yrLk9l1aMseshE6f1BiAE/6/l01kGNOErSxWsqKK8i8f3zvxOVuKO2SEJ1Ev
b81nTQMOYdW+U983rST5oON7STo8yzqxjD4EOb8q10OPaVA1spLDBcrLnBCupNCo
cd7mcsRx9f4BQntAlpWcfNZ00jKdgvFz8OHHT+RitXH5PFbJoratC1Uj2/o+NUpO
yfZFJfTNDWo6c2i0YNCCmFtV/3iWtK9Va4aYasW9oXjUpa8kzzK+fIlbgybFkwv9
ColW74hDroJekB28qH7LPu60uGHGIYyRIvTkGpMmmhui0EL2PHgs+AcKCkxAGtip
dJdzQFLQiRwPaMPUxx3g4atYpnUKRYdN+ERXlYlk5qTr9ureEoaSwVI/NqTd9ZJk
/CcqolAUnAp3FrNZSaoBE49U0VtO7u4WZpZRDkQXrGxB83XmwD+qAR37OHAE2zUC
+9O1MCpYTFcq6l5ikBRYgQOnbaSgQHBfNFoizsunbfg4kPfXIqV3lfXcz4ok4Wqd
vS1nv+10l5KQ3Xy5QK0wXECJIciCva9c5sN22URj998bZU6K7ecGvSGxO8csJTSn
JL7cEpqJdQfQKGKpGjxzZnpg4LIORYm5j9AgsnzqMl3jg1p0jOKbSkpBSgHAqdaz
EQ6xhxyYeAJEqbuK0LNINnzlFrgJ+BeKM6HkOnLBUa2XZD/m8Mi7Pg+QW7ae8IyF
h/QmB90OCwCt22hnHm8/hDM6QtqGuVM0kRhwAod/W06j6XMpAUlYIqy0sdcvTjKZ
Ff5hUPyicnWVJ7NJarochBz2/Nyd36EliYoiecg7PSefMfkzvReJRNvWgB7RzwSa
MaHpMr2IpW3f7WPT8RLN0oTsBnK1zh0qy25IJcST5FV6/++rQkWCaVs/6OrQ7Fbj
Ft2Vr2XBZ8oymxb9tn3aozCxrvLW1VP7gbpaRM72LGp+mcLVoRxbDDGiZGPm6bFi
7PvncwEQvP1ZQHfLPVjD08NCG4H6dC86f2/FFsKlZwgidNPQ054NXiNQDCSwXwwN
uww1OURBNW4sj3YZ2CYTjX/mlbSnip5lvWc/JQjrKu7fee+625YYlRID96rT/N9W
odLsXXdVOHLN9lXmLABUyM1gdjXIc4HXZbg4CD/zIDaTdGwf0nrLEvJZEYwdfbtd
DM+fM83Yt33mPfqiL/ZohvUYnbB0IJ14ggMJJss6EYwKq6saMe606GhWe2dabrQH
JblxgIrA1IfGJbLS1xRIUoqBUaVUxMA7dYMp+5zLv7xfJzLkfE5t2+TR7cz08KGJ
YfF7QZkJ31HB8U7inPGK3ymYLxUvtJek/cz8l/sOGNsp6vOWaD3IuwU8niK+70XI
NjLj62Ba/JV82nfP1a01/eimLu9ugLfr2BLcV57nwKmJklaafCYO7XVhwUSKqey0
OpU1Zou5WgWXVSU3VKChclQeMcYG+bHU00yRpPCCvnAN+ccTDcG/9GvndinPMXM8
MrlFf0AvM+ZFAh90Kf4mTCaswcxcFnOSuzT9Nggqp6gwiJlp6rUqsi1HpN7zUCFz
1XKMm5STmvet6iLno73K3BBY8Q8rE06kQgne0u+UYLiM5h7RUeVwK7CfaHZ+OVq+
d+ri4ge+sJDJSwIhju2+xyYXFfd1N+T7/1AJg7Ux3XAR8oOkcgy7CJHHaP0+0cXF
GJVgn9JYyows0CgnXU4vN5yuDMbxviEQzka/Hv0Yi3lqFsmzqGAJLpbKwFqUBPgi
GKmTmsGvLsLSjpVXCUPaPUMX+aTzOpW9YmiFRXL/ej4qKZMbkBpxA24UX2/d29BW
CF81zIB1FQlkdGYsvqVHW9ZQx+0NXzEYIC0rdFHJEa4pCkdtxLAqyeZgBvRJqA94
N0hJVb4J7NZE+ysUpVt6ZH0sUkDA6kkd2wG8VrMMslVL0iZFU8Hse8PNzOqnrq97
hD6IkclxF4fFpXBYUoNmsCyFIb6i12tPPd9RRR/IemAEXMk0u3oNul5YUwsdwQ/4
HPduN4RjnA32ZurWz0UxbVwUlsOxxMe9baWRZWFTNKKordyrZZIR6eTXcpK5rj5c
ETWSYqzq6bv4/8ZpGyxY+38SpmY5W5OzUBBgee2zWDdrEx46Tg8E2Tfgj9hKYxFG
U1ptsR3EOByDB8meVZHJp90s+1y6veaVjOL3ZlH5tD7rdhe4t+kVyNArK8FI9BBX
GbEBaVD8BMHQISWSOHz5F4bD/4BcLfkEo8XxZtYOBXFPM2HDcScflbPd2lLwHnI0
zUXBoCzp7wSoLMx+r6xvddFo3rVLdDEnvO5MFXqIiryhE73vKbkPAhPJgvYxwZ93
JBmlnlLWCHtnTa0tZYhOZiKDXeMGM3TWa60vRiJ5mAshgP+LD6yIuo8w9sTpxSxl
rk2YKGjjQ/xC6+lP8dHTb0NFKaucikDY/60UB6j5cT4JSLxSx5gPf2X+CHBIcVXP
5tGmli5cAp+/DP/J8Uf7B1luxD1FCVeA2zqfiEnymx7YKU5NIWQirRSZZX61HiWf
wYqnfh2c4hW57AyQihZmkPDjMSazSIganKXMRKpXLjMcfqHhJ73K37YCw8s/iveY
insSFYB5gTcEy1HGb9pCdLuvgw5A/2uUnQ1Qkh0IgqTrt1LyT8s25yg/N/8BD0lb
+j1Jh2+IS3DOFLPIgu0rN8ih6db1x1VQYKVYcjOo7lyd3Pbc4Bttyq6XEhGgnsGT
AtinhWABqvJGHkJZ3Q8ACYBlcmyUKNK0+lQzQzRLDKJ4Wn2K0j5SR2TXVTBXR8S3
DmN749K6n+NGOejo3Pbh5zf+ZPy1WscptwYp+ajYkiNoiPGhE0DJ/UsyKnaCSqXw
eL2O5c9eaR1nnljbSh0EPCLYYflIN4tvkLyiSIxEuLDfO932L1VXhzRdqRuUWuyH
E2kKSrd8K3e5KKE7mGCpED+eqEhVbfd7+f2bmljlW/tXhW+XOu+z45yFAlQX/adu
/I9jsDXQTqybgBTcR86K0n3GOAeOUg5opO1KMsNcp9ad9OCu8l3ElsuFGf5u8Cw0
jpofSNhwfgH/igNnNkQj7kG9TddNg3DHHJOduT+tyVI0HVi8QBqx8hdEwXouGGlk
+MzOOG0fC1ZZG71K5wpTn2yq1oTH/LeuVWwPOcPzuLsURJM+Bu1vvYqvolcHT89m
VEd4uw7awtuFmsj0CkhlHSu+ctm+hMOmzVAp/fREchvcTg0819mjq6etDoMMh/sJ
Mq+pHcunw0M3BP0lS/fyccv9YFDaJaRhdx2tTSAtNHgEf4oEZqv1Jaayx9K+57mK
f2C63zP9RWDLLyd+AiItY+pBjbF4t/GENgvEwo7ERQPbSoXUUsoHHHUifyHTLh5u
a9CzMuWMdANPDya4d0aZwklhC9b9Ss5bp48194q+j+Bsyd4p7zyffgzTyzcI7VBw
oI4p6Pk5Ce355dAO2t07INbUzMx48si/cqvYtI5dA867InnOVLyBbmPvK6fvjsf8
siWga9FYgUdhxWaDHFGaugR/UcI1Qccy0MUjHag045hnbUO5f33d2bHeCq63Y4hp
oBHhwuVv17rUxo7DRVEMgCyqpXOIvCkdwk1UF39lDRGJ8fjLAR3PSlH23qUwjkmb
q0m3ijggbCqtTaBH9Lk1mA6UmWYRAm8roV6uqVTm9KG2suPSlAHxOFY6U1h13ssX
ZWX5mVIhrimYOVTF+b6Nl8aI5LwNTRtdcFn6p17MEJ2uNuGAaFRlA/asUeX7pAlI
k6L4fOvdswE7Q4nsHD6mzVcPhttpy5ndad/bd1kK30fif8N6oOKxEq9CZzRnTV9l
s/KsQ/Rzaju4MyO8hcPBPtZjJOazvyCbbNLbzNnwMWExLuSB9JBSvbZW2MIl9DtE
CfEUA64P5gwyxSy0LKX8R5UAm+XgfjvH4Rasbg4E2xdVCnMSnQuSptb/HYtQRyZt
iSamS41MJueeWWsWfAcTYxAXZNBXgi4HapYk3YTN2OSWDtVPDJC6eojtf9kEn+Op
+CCjYjVq/qa0z9Cu801J7KDt0Fj0t+pcqcO9UvMbnOI0FFiyIPx1Px6agbqYzFiX
Nip+4WriQGW+h1ldg70sEw==
`pragma protect end_protected
