��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{j�X.;߅ţ3n�c[�w��o�z����kV��pN��Jb��әcS�{�ի��t�Hdf�/DFT�I�Q.�����g�k��qw9��"�\�P�9�����m�T2���**�f�����>ہ/�9؞��h��!�*�!oZ�?���
/A�vi�u�0�@*�M��Ӿ�z{S��*�\\}�5�/���ߞV{���;"�s\*��K�_�@��A�JuHD~��#[�O ��R�)3V(6͗׷v-;�%1�:���Sְ����Ȇ+?z|N:G��!�0-��S14�-ٵ�ӵ�Ygɭ�K�U�My�p�'�_�f��v�F�SJ�4Q��~�J�ˆx����I�6)X/�|9�S���^����A�[�+c�8������.5�)~��:ͨa����+�2'���m�&Fڒ)*�Y�eG-���^�>��J�Q�W�g���0~�ĀG�PB'cQ�>�r(�>�p��f�KnP�k� ��S��� *��ma5q^�ݓ���$m��Ă��8F|�L�	'�u�5T�_AQt4��ծ�r}���!R�O렋MM쁝�������z�ز��`��X��m���O�3%��qe㽿u+�9T��$�c�/)c������pT3#�$N�W����E��a�p��J�p$f���"�t�X\��6Čwװ���v��JS@L�ʱ�mʳ��R������q� k&6�:�m��l���kCM�w���gX��R����8X ���a���g��VN4��X5;���T�3�dr�|�&@�ڇǰ^���dB����C5���k�~G����O�V!\����{�������'�8��v�veB�_��g}=4)?�;���(�z&N�oF?_q:h��&��`{�ϪP�����6��v�z":ig��X�����٧�=v
���j�B��F��!�^%M����-0ZP��q��;؄f�03\��l�zSJeks�{!��Kr]�Y�k�&o,�eyH��ss��N��K�O#�8����t)4p!-�K��2F�vN�=��!HF?��t?b]������vܳ�զ�+9�kn*G��������$A� ��s�~EW�%^���c����b�`ը����JmX����y�;���q,�E������ܗ$��E1�3+2"�]pbw�A�h����?P\�wò����}/�e�{׿���	�u�^����y�1����0�s���b�M"�/��1T=�!��*2�(TL��A@���E���qk&�c(�L�4��g+�"��t�3���Zڎ�޷�e��g�- $��`���I\�c?�-GJ���\����?i4���Dpcp{1�h]�"��\E����P܇'w��bB�p����L�#�W�j��r��¨Q����W�X�Q��ݒ�G�_�ǲ����β�D���"�s^��o��]��h9��<�!�A'�����Z[��/�(o�^M����o��t�,|�i_HT���9�8̖���q/}&�I��A�_+#t#8I�����d�m D���
Pt*��`�q�\{��Ťf�K]C��YR�ܨe��$i�Nϒm��i�ZD�ly���kM
���(Sm�iuUS�����8�VsA�_3��|~*خh~p��(I���;�@����m%pA4�/��sI�*۹tA�aV��t]�n� ��NVތ)坴]���à�S�W5�����:�6�f���wfn�Eb���{��*���&���TA03�����$���'jUU��r+���p-�p�]�X����u����!��8H(�C�&�b�QVJ<��>�IH��=E�]f=�]��;�m�Qp�O�+v���s4u�/�M�1t���?̈́I�ڽ,'����,Zו�B��|�]������54���6�iLz���ܭl8E$�C�W`XD�X��(d:��O�Z*hT)�0H���Է��{(�U|���G�a&;!������.�@�����j�.��݅�&��UQ���(��[�r��O��y�r�IM?QI���������S�ӯ`Q�t�g�r�����Z#e�6T<��yA���*Kd�!P���F�;����:��u�GYo����t�c[�_�8��
O`ƥt���A7t��lJ怚�i�^+:C�%z�PTU�}��t��X�BTě%2,�_OD ���"1@2�c��c�U���K~}����D���x>L[������>A
\z�߀L�.��x4����n`�էq|8$���� Q���[�wZ��?B
x����&�����>"�j��$V�{A�����Y]��V��mޞ:���
�y��X�0��!�����V�{����i����U����h�Į�{y ~������q6l��J	�9��0_݌༵���円�׉��Q�ZM��\~��ϡD��zx��󊛀��#)A6A��K�o=�G�.�����=dU0|դܜ�z�Ƥ�])��&ŏ��sϜl\kIRSn��>��b$�)�΋_�?����[F�~M����ϻhZam�8�B��0$����q��7����� ��7}9�~'�ԙ��X;!{��ZW�݃+m폟Q^M:��L�1}��a��^ 8��k.yl�����)�秦��W��.3$�1����@�T ����������~�j\i��>p�6R�=���i3Ib��ç^��K_�yt�l;�w�����D���|��~��O6����R�m��!P��!�+ԑ�%�Uϖn[l���bƖ?5r����9�ey�#�V�`EXN�oGR� )�/�����J�O�pۮ(T���*�`�X�G��;ԃ���@n��III�p�G*Ʀ?ލ�����҇����P.+.���T}�������P�@}�UJ��V�1��Bۈ�}~�7M��2��-������ISC���M'�F=�8Ń�'}����e��n~�\��Z� 7�]�|���} ��#Z��A�L��O��X8�/�,gB+����EL���;8�no�g�P�߹-�m!rd���?�+%�7G��i'X@��"�rO�n������cPm	����jʸl�\�G��_�5�ϑB�l =cz	���m�@�>�G{�	*�m��u�;��塕�&�`j�X@���ywsb���n�X3���_p!�vG4;߉���@�R'�09*V�h��'_aՐ+2��XϒL�(�>��*�<�<�۹�D�R�*��F��eE�d�֘8�2�8U��5���Yv���]��JmB�V���+#��=5+n�X�)�4}1�b[G��ޤHV�T%ڭ�7ջ�����\���}���Jܧ3z��N�Y��^+�z�Fi�z`:\��#Ĩ��DyU?���T�%޷���:����Gk�v�W�I<���|��� �k؇��(r�w�̛v�8-�58���D��#�	ʔ��IO���[��[L� �p�Mш�)~ed��V��	�*7����@>䓿�W(�>\����hu��,���:=gs�Q;a�$��xۆ3f!��3Cb����{FiL���dK�/��c��Ӱ��H��ᢻ�Z���:�.xt_�ð?��N�(^1�����^C<I0�&�q�H��_��T��Lv�N`�p&���S/�c� x_�F�	�������b���K�=�z���с��@t�&���PP�J��Th�3�聣����,m�վ���i����"22��]��J$���Е�)k���35"nwKih�A\4���t��y��{�f��A�#i���+N���k=o�Iͼ<��A�/�i|�[���oܡ˦EC6z؀�F&�m�G�Z⠺��$���:�s �T��5Ġ�����3�<;~����hh|�i��S���j��)e��R��f�À+�܁��8��Y�}����0�����W����.<P�@R�)��}�Q3���%������(`)��sŠ�Bx�n� )��>1)�m4e]7�֨�] 8R�Ћ�E;�� 3�P�ﻪC>u��`^IjLkO|k�܆����t�Bxm�H�5̬��:}C�2#qHQ�$;��nx�D��O��k��C�6��hA�|&p��O�Qۃ�R�:���y�ZR���� p�+Ey���2�`E�c%��ty�����r�%��Fx�L��Ɇ0���:�+�Ȟ ��[b�u�ߐ^pO��(�����Bw��~���j�։�;P�\y��m�oH��zͳEm��M��7��(0,!>;0e��u��ʳ�<T�44o�+��T59�ͻ7FW�q���ff�X@C`5<D)�W\]�N�B�L�xg�M@��z$S�7y2!Q�ܳ�e��3Yd�f��(���y�})V�"w����:O!�n#�r2룂
r���V�#y$mULܕn�og�Cgx�N!�3�u�7��H�`Q��$�<oX�9���J���zKw�����˝��$N�C�.R7}�|ba�"�{��'x��l�%��ɣ��ǜܯ{+�Z�e�T�)u�^�W������@�*�^��ܐ�R���&�}�rtI��؍3/������tF�q��rQ�ʶ�J
�1-oVJSf��7�4Z@n�b�Dַ_�(�0��AAI�G{xG���[1~�SX�?���+�}
-��'�G5��EZ��ݩ�y�|��PZ���N�E��o�L�ZWҶ�d���V���&P��Z�La1��� *�}�6��:z)wk˯�*�\�QƎ����ʒa����g���9E�|l�yx`Mi�{���/H4J+BԘO�i��ګ4�cd����V��"��v;�GrDVo��T���E��q�g��O��R=
��灛��
c+fV\"� �G1���v�J>>�Go�x�{�ɥ��r��S��q3��f�BPBI��t����`����=U&P���5��g�u��n]�pQ!��.�lCA���BVW�Q	y	 ���1��3v}��,�ݱV�)R�E@2���2���E���p�W�d��%��!���2��'g<겁 �}���M@*B:��m�*�ʫ�1 ��nx�x�d5�w�7p��$����x���r�}� S�uh�Ͻ��tG�����U)�B=p�	/<xP�Y8u�c�A~�\�����ٯ�z���,��~�}�����p�f��Q������.�,�{�~"�~5�˲��y�����-B=zܫ�ahGU`�~R�ǫ����v���̵M��9,�T�<+�6�wȄڔ�8�,;�m�|pv!�ȥ����tx�S�sۖ/�
{L�~��Q��}��)�o�\�r'[�1�-�#��b�	���ED
rO�MAԝ:ޓ�z�SDk�А�KLe�D�����^��"Oe2��Y�xnH�i}%�!.��rb;��?��2ؕܘ�<���-�r>�'�6���E�se���� h�wWELoh�,/!rH)'}��X�R>���y�Í�䌩� �N��%��x����#²:5�q��~t��p5=�5�k ���#�л�|v�Tu�P�:ƂbU�Q�.�kC�#������9�X�Y�Dʡ�ssK�s���@�,v�@�3��^dN���_ݾ�:�Ăd����D�{~�P=~�U��?迮����:�S,û��	��Vm�쓶��K���E��!�
2�~z���Z�#![S{�V��>T��j'�!L+G�&��s�I��D��6I������fNS���@�����b���9��9��?�2�ba�4�ZuY����g�^y�%�XCi�(���,�p0Tb\���#���)�{��q�3�b۴��o��
mv]���Q-�]��V�����pRzr�T� (�Ě���<�5ň��ҋ��9T2�5��^Z��T�UXk��ΨS""H}�/�کg���)��#�����'$}��{�r�U�n�߈�kT�¾��x�ǎ�C1���2�J�2���}=2-��G��N�iN%3d�s(�(؂�s�{$�2:0#ps�줟�ݗ���Z�Tj)��t�~vK\���-/׏��4��|0�F�)ޮ�垇�K� �0�W�;��}�y���z�!86q7d���m <��Kw�
��ͦ���7SE1`�J#X<^�q��m
f&�& ߗ�	"�52��'،0S�K����m���\��\sn�F �,�4?i�V���c�
m�J}ͺ?�D���T�+�CA�ׂ�88lwr��=s�
��Z�Vֿڬs��"_�ݱ<6���m}�`p�q�0WzQ�)������0ܚ������!��5E��i���W@��{y���&���n��m� ����i�W$��x#�����*�D�49#gz�6�Ӵ&mX�%^FL���mP5l�c�)8�Lv�ЭƯ�c7�&xH�����
��L��u��h��*śg`����	�?�@?�O�E;X�v��Z��-,j�uc~�e����9�"~��V���S��u�ab�aEJ�!E��(A h���{��Vs��+��f�9W�D�SU����%�m4��B�F����!�8����:2�ŀC�^�o�·�X��;��뤤,U&A���ajP��<	���"����U���<u�&c�lV	N����Z�Ƞ��/��[���ғ��z-�f"<n����O�i0��L'�ATй~��HL��K/�'?+2!��8�fhq�lS���`����1G���Ql!�&�HZ:¸����<]�����#�Z�1���zh5X	�zM��Z)꠰�Q�7B�E4)jj�➋��̵��WY}��UU�K.������ug��Iq'��p�������g�7΍�����qd)k}��4R!Q��vGD�x��DHW�ĉ�UT
O8;h���Q�V� ���y�X��pB�-��������͜J�ܡ��/��t�ů�R�Z�v���zn�S�.� �	:� [Nn�}��fxc)a�ߔ��'�P�LU��B��)��e��h��9�g�3��Z�Z=^�ȴ�zI�R�zQO#>�����Cfz�_*�w|0N��M�*}���+�Z��D�|�D,�ɼ��2B��H�3�6`�w�Ќr���N#`�g�<��y˦��<��5�&�z��G����B7k��{KWP�f�o��A���2��Ez��PB�bi�!�|����������Ǘ1���Zxż��:KF,w���0�Z�v����<��`DX��	&<u�v`
���{�<�TT��Ee�{���`<����I3�y�'�ɕa����՚�ܟgo�7ח��"��U�W�g[h�Yv�e5�4��~P��Ŋ���3����,祐̇�h�L(�LU��Gf*7}H'�F ��bc�5�xeX��Ua*� z�в�܃��1��=:�-��T\��@���Ez£���x��Ae7�(�T�D��%b�n�@h@~4����+zݗ6�f�	t��n6�juh�� <>�i�V5�H�?y_QX㇉.\��"��x����)��r[�����k��uF�.��P �ܻ�������5�+(uTVC�!��d��#�<��&�d.�&��o�K����̯�H�hOR����xo�֊�n��)�����Ի�8�H�A��2�Z�v[���W�� ���aNž�h���۰�
�(yж��
v�]+�}�M�Em��$o��R�"�+J��k-@�
�=�ҟ��W ��I"��QG�m�ݦB��
5FpO�G�ĐF�NY�T��:�����V���b�X��Ҽ2u���g臋��<��N��k��Ǽ�Y�%6�
���"-О�߯���n���	-��X[���"7��M=EF��Ѵ��<'��l����w��Y���%e}F��)
�pI�����R[��42�-�����=T�uUt��1�ޟ{�Ak�H@�U�|%u)�,)d�=
�4G5�o��Ji!a1XG],���j����h^ې�?XM_���w��&I��ƨ1!��ڲ�ӵ/�j8C߅������t��� �xNݐL��gf��X2����m�2�Vi�G��P�s�jQ&�BK;�ro�� ����P���0�hpn��G�u�/c�U\Xñ�A��b�v�vG�y)�OU���R�9༽S����L��iT4@�U?�at�O�R����9�J ����<#^��S"~���"Y��<�o\Ef��.t�HZ��|��Ul	w��v<�\�y�tY�e^��=&xқT���V�6~`���?B���4�~���r��eSU�U�P�o���%��P�G�ݒ,��d�>�^*G7lje�.���H�U6����;/?~x��_F���o�5v���ӡLן��ߪ�6%�e#اS���X�pv��Rl�;� �|U�9������\�J{oE4�èk�#Ț�:YD�����<#S�7A)�A�2|ܒ�i�n0�FHr��.A��t7�����rJ����#N'���^�ŭJ"l?N�* �x��=]��C-��g�	�O�tcT�Fg)�*��o�����e��2���y�%dJ��2,�Ϣ���ZѠ䗙 F���B5���ݧNݞ)v��2G�/8~~�0$P��܋^�ȗ�4��f���啶=�X#�Km����\b�׿�U8��k�`���:�M2��K� q�*�5�k��q2�����-sRE�����[�C1`[mptI�U���\j+7�;�:=I�|g<���X���d�?W�D)1u�9�����8-9���x���,�SSRdkq�
ac�=����7���5���J\y.yc
��+qM�C����A���QY�}�]T�������J���]s�ٳ2��O���~S�h�"x�Ksb�ʨ!%�ܩk�ke���g�Ekx�I��u}/U�;��#�hf
C8,ܡ��w�=��R�!�_3�o��es�Sj"�P'��i������'�S^d�7��k=:�b?t����b��f�I�,ȫ�.E�2#>�����Q{v�toz�/v�z�C�D{b��[QZD�c���"啟ꆙ�D��sI4�X���gR�ߓ1�c��.v�>M�'C�En�;�P̼.��
W#p��[{��~���<΅�:YG�ll6�'6t��6�.�oK��b7θ���\��T	��B�t���5�:�l�N|k#�^\�6��}����Iע7��x�^T\�%V��9�22� rg'�j�y�QAA�Y;B��s��}�"�.����~��I@��[���~�Թc)���6Ǐa��C�iư�IZ�Pf�Uê2����1&�|����B.��������B�4���b�M����o�I�N�Gd��!%��r�#QM�����ׇR�a참�E�;@��*��>�Q�&.z���|ϒ��}8�ow��z�2�W��$�s[�9�$~�Zd�G�`��0x"�.^���r90�z�:O�h��r�������a�G5�R���v���R�E竇�ʕ��-�ھ�
U�"ر��	־B^	#,�T�|�@��ם��D=�I�
���!$�r[�_�i#��N$dyN�v�C�����R��%BLG�P��Ty(�	������:��~�hvn��ҝ�GVq��0���ÿm 
Rl��^i�x&��U�#bHK�N�3��[�b1�K V
��"�����?`�}�DB��#G�D q�#g�?{��u)!���Zo�E�}�uG�"����ș�S�Ix�3s) �=I	�3�+�S��[A��T�ߕ�7)�鶴�z���?�ƈ �Y�{Hl�=�������!�L��c��+��L���C�Ń��31���>��F�f<���T���h3��o�S-?��.U�<�T$8�j�(j����y:�R�īG!�(x�'ٗU쇩��,�:���O/	/:+��ο�+僩o��XD�;��v�Ȣ���h�9j��I:�;iv�*�����Z���f_V�=h�]�,��)mhf�E$�,wJ��5��������fc������CX�#����W8� *����tn��B'Y}|�l��T�� �-8h�G���i���:$�-�呼Ǉ0��1��H��e�Xu
S��&��I�T8v�t2w�������j�.�B� V�oI�(��]�S:&޴��ų���Z�s7;��2�it�$e�
i��@��ѣ�e��s��N@�MkAo�����q{H�L9�\s��z:�T����D���H�[�$"�I��+�*`���j"A����~�u�}]!2q�լ)斡�?��?�$ƃ��r�Z���f�1 ��?��AN:à��Ľ����2�%�{���t,�M���G�Ť21�~�J��>�B�;�_T�A�%�χ�O�*@�A�|Ä�v��[���PD����k������ЧwG���_�����4�ǵ�
�2-��#u�\8�~e3q'	�ш{�)Y399�!�k���Zzt�&�������"gb���(�?e�v4Sٍ�.��][�D�v,�q�YUl~0C�w�Q���w��~*��j��z�̔?��+]���e6l�(v��P�b�`l��vo��wr��i�T��R��n�ƧV�k��ux����"���J�r��.��"�K  k�`�~�1 �?B0�BV�~���X������d��"2���-���~��G�k|��2�S`_�O���<�A�L�����G�&2�E3r2T���l��\f��/�Gs�f��<����[�cC ??`���TTAC�ǁ'�i��#�/�#������$ԏ2]	ρ���p�W&A1��ů�)v�NH>�ԋʟɊ@��X9�eF O�b޼�x���R�D�v0�\����`iu��j����K���n-��L�NDNer�%��~vq�w��;�aX%����B��Ǣ<��]�ҍ��4D����ʊ�?�����2
�^��#_�Э��L�����T����Yc{$�ĺU��Q!��l)�GO֘mævw^Z4�C������fN��A0�qC�^,?�я�Θ���1scy"��F�ƴ��[�Z��q�mzJ�J��1��H]�5�5Ŕ8X��T�A!��#�8��c�hk��2Wrp�#`rտ{����@���Er0C��2;_~���?+��j� 4c���e�s�3ul�K�"#������0!Z%���6�x=���X%kr����3��%9�D%W��$�(�t[�CD��/ ��nE�;!C�C�?�̙�XCaH-dv�e�~M:;�wy����C���v����Zk��[���.{��5�;X�F�b�����+2��p���I�A9�Ox�9�LQݳ�϶vP��&�.�?�"*5Uc��eM#��Ui�H�zw~��G�~eS�K��%
 �����{T���!�8�_ʪ����ӕR��.G��ΣW-��� U����߯�~d�&yOϰO^!�h�����@� ���
@�ɸ`�j��Qv�4a r��ƺ ¹�e�7n��I�����j���O�r����7�a~߈et ���{��oKڊ.H)瘀oʫ�>�{�j�;Z6�_GDKj0k`�\�[����9�~蓳����a���Sy���Yk:�E�6�����b	�uZx�V8"�U���}J���p@ԚsJCB���x��j����͝��_C��
-
$�}`�(<�\�O��<45=�Æl����[��Tz�w�?�J���f�쿓�c�|ŝ.�E�'a?��0+L���Y�J$$��,VoGr%�`8|a�]	(l{������q@�qT�3,(ah��	.���I�1�M�腂-�+�ۭ�w�լ�C��Q����Jwg !����5s"�K(wc�f�TqAMW��8�a
��ͼ>6pa�o<3����[�����i����2�C!jdhO�HiF��ɓ���	
aV�U*��(�e6{ ��u\G�vi(�%8���kE�CptI�)�~G��>e�(߯�(�g��'�C6�����o�$�u�����_��c�xr�F�p2�ښf[r�����ÁF!L'A�M�9�������>��?�sΤ%�v<��>�og���Bb-^I mp"g4�<�^-Pw�a0�������sǱ.@�p&��I4�9&1k���pF��5�b��x�J!?X���߬!]Pn�D�5���U��9M�i<����;�.�3b��8�qnm��śܩ��r��߽�}ɣ�$2��-x��NGf���U�߬y�)w����$��>L��{l�1|+�d�����o4mO��/� |�Ew��*%T��粅a���}�Q֯��Bv��n����'�_��cm�s�ow���m����(�)�pN'}�J�BT�j^r=����p�m��͟�U7'�RV����0�0D/�š^&O�60HR S�ҺLf
�* �d��G�z����} �[#,��U'�Y���w���b�|k1z�G�4C�
29]oZ���,J�j#��[%���{�_\/:�xf*T3��0ѐ0-�JH�7fY�r����5g(�/�`���_&�ر*?®Q��Ull����'i .5��?|$��0[��P��X=��Eơ,J83 �e_��ޗ�����Zua��7�(b�ļ[<:�"ō�r�Q�
7s�"��5%2���bW`S��`>(��������48�}!VuR�Ӑ���ZQ�#�:���`n��6�7wl�8Q�ʛ�57e�)�9x(:���ύ"����4����	�b
)�����Du�9i��v��$`�x5\����U��X���No#.
����+�2�lK�3v'���x��C�Iv��2��̻�p�)JS�Sd�����XԔ%��Cc^��\��>zM��.W�$L�v�ӗ��mw�]F����,�ː�{ʺnQM6�NL|j�	N2l8������0ap��g�A�o%�J��L���k���ـ�Uږ�p�E����'�V���� љ�r����� �ݲ!�qe�5l�����U��4��~��-�X�0P���s���bJP��仑�hT5�EN䃉Y��QI�!J�1���N�v$^y������;g. ~e�@�>�0y�w=�F���
�V�i���D�y�������޹۞`B�)B�X���Ț��[F������L���ޢ���)�����P��U$'��Y�F��[��&7׎�5��c[����{_r9��"�x���z�]�5htYq���9zǨ˩��u��0a�~ľ��fKp�L@�G�C��E��nBX'ճ<m�)���CBM��M��o4��K�+߷w�K�D�?!���+_�0�m�"�k��{�@��L���)��V�j�a�U>Ji�t���2�cq�a���!ؽgX����T3�aF�N)�f�z`�"��>�xB���7�9����ud���r��n	h�9mfy�A/�X/tC���D�;����-�`��b��5n
\<)����a��ҭ��1�nAU�[���h�+�$P-�$Y����)��K���K�es��Q�-?M�@�tqo�җ���0)Ax-���F�Xe~���_W˒�ꄥ�X�����_��処T<6�#!z����>Z�{+��t�Ҿ��07)��0(�_�A!�AH9b���|)��}:ޠ-zrS&JN����'*��<MAԯk�2���R�p����p���8�d��Q8�<���G���͙$S��ֶ���SǕt��l⤈�	i<N��G6��y�UK��rm�9n�J�!��<L��}��z�`�����]�'��PU*�]4a��Q^ո�@O�f���"jvg)N*<�B��sbi|��bp%�Yd(b(�HF=A@<iZ�=�c�l�T����f�Q�Z�ş��� *���"������6�h��/ԗw_��{͞e-jO�98D�F8��)�/����D���E3-�\59̢R�Y�p6t3����&�
W��_@D�'����T5��w{_���{��&�;�5����}5[�z� \�9�hkG�`���;�&�����زt����.�Տ���<K-I�.���
����C�&�IjΊ�j#�\ew3�߇�����%-T��
Z�������~�v(<�5�qL/'��W���$�FwTn��S4%�dg�a����'���d������"��Γ�{�ۛB)8BxO=����!7�H�od������-��%M�z���O����F�zeN��S��%"?;����<�Ҷ)T79r�%u��'���s_i��nE��I;j�l5rіʵ��{����r&�c6�isZ7���!5���Ĕ(�N�I����긘([C�����d��XUٍcpL��l���_T�q$G��r`�Y�<Ea��$�O<PGD�#!�)`�Q�=|3�L�Q�z�l*=�]ƊD� ��(�+ɼp�>�ԅ��% �53d3VSN�J4�c�`=�㰧��T��a�FO}����;��O��μ����M{�}��K��H�?y�w��;8�f5m��m�/D'��t���̶�W��xjx�W(�0ѥc�j�L˼3MDm'�Y�GZ�V�86��b3�-�9� $�Z�R�4�e��S��h���p�G��8�����tX�S��N�Ǥ�,�k:<'Q�� �[D�[��Npkȗ�a�;+���ڴ�����=��A�����~K�^���1!E�\���֒ayv�0N�(�\?&�מ�m��j�"���i]�q$�d���؁%�R�����ҥ-�th=��b��QO'�0�������Ȥ�|��G4�Rx4 �b�B�$k�����ϋ8��r>_�
wb���E��PSz:���S$7�;�0Un�aڔUko�0�c�q|�]<���G9Y"��b�:}�+�\��f�W1� �&Դ��Bϭ"W�hh(#����q	��jX�_e[T��y"�ލ~; ӸUB�b'��WK�r�V�d����!��_|W4&Ƭʬu�,R��Ow�������KطйII	��b�A��C8�&g]�jT�]؁X"�4{����ש8dA�kuO�#CUUɂ#^-v=ꃽxr�$���z5񦧘K��]�������JI>�'�K�z�@^�z���qBGO#_�8S t�2�&�����M���"��4�}��%v��f��}�2��}�&X3�m��p10w���<���@�|
�u7Q�=E&������EQLplR����d������TV�N��gֽ&FMC����?����B�5G��ȵd���{�T�.�=�O��p��|3gI��{�x7QKa�B�ߴ���=�4ӧj/������ 1�ų_1�
I�Y��=E�UEU�D�z9H��F�G��Ɠɬ]��PԐ����Q5�pq�#�|*�9�/� jQϘrPK����ˉ�3}eq���A�pZu���T��8�	�s9�!���h=��j_��JM�o�)6�9�h�ʠ{�a)�&	+����!�xK��zNv��z��5/r��Zжy=����~A2�pc�i�)[e�qjJG%Aj�K�`��\��v���(JY̮���������<��|_�jw S�=��Q����
wY~�ĎDD-N�q`�X�msoW2��h
o��3Hojle��n}s����hԥD�T#;�i����|�2B%�0%<�^?M��MiP<�Ŧ������H+����֐��U�^�-��Df��;v���4�T��L�ϱ�?��f_Pz��K;d���*e����+�,�J�)�&\.�0:�V��Y�:y_>}&Ʌ�{���!l��dE���G64�U��S��,Փ�4yo��h��^g�B3q��6vN��4�̣K���ӄ�nL�4�r�V����I#�;��#{�%�1[΋�s��Z����Iʆr����4�?%��ᗦ�]���J�w�g{C�n�V�d0bY��n��s'zɅgd|gûl?A�3Ҩ���" ��6W�&�4w��MM��r=.�%Nl�b��b���ɔ�-������v���<���a�Hb	�3�ӿU��a��&�1�D�+�BK��F���;Q�KY
�ϼ��4%AU��׽��A�㘮�E��yq�>�e���hZu��*��0���#�4{6� �#c��������M1�
ˊ�<��Ǫ,Tğ#a	�@o����Gr�����]�DY�*.Q3_Sg"q�Tӱ��U�!������c�b�z%�A�]1���:�,Vw�Mqq�O���{�v*�?�{�m�k��/.��N�b��}֏��ι�����͋`g�p��-�� 8t�����v=Xs�!
i}S��_~�����{�Q)�*���� ��I�����^0[��P˄��rl��,��Vǣ	[�X�L��W�\��)<�����d��t,:b��[�Hz�5�4C�O�zS�J4q����=����w�_��^q���#^RE�K���w��N�>�%3�u����0:f�g��X�����N�5�{db���/�t���LcRi����}�E���g�%����Ŭ��yf�X���ɝD�n�G�/���p"Jwֿ#�pvSBc;����O;��{����N�"��([��6�E�DɡeFq� ���.Ů=�77
�2�%� �V�m7,Ļ���s�í��[�>�7�D�ۚ��_��o��A�T�0���k���O$٠
�	,�Z?^�,K��ֈ\`��&La���K����o? ����kQ��Mr!u�5�b��T�(F�v�) LO)'ɊsՖ,Qo�kW�Ţ�ځ�	<�-���C�QIu��(�"���� =.P��@ �����P�'��H擰`g ��	i��8!N�Pq$��:�χ����΄�#�ؽiiX��5/����`1���ϯ��=�T�W���t6��(~'ֲ`�ǣ�\\ �*p�s�~��C��r^
�e]!Ɂ؊L�"�Xĉ�����G�����Ê�Я����X��6r�m���#t��s�h�0=OB`�v"�����T�H���Q�����}�6�߉��[̊�e*�H2]��o�y�ST/��^t�q`�P�0I?:2�kM�G�v�ϒ���y�`,�5p�<��^�E��u�=��qD̀9��d�B8@�ܰ��MX�?��2V�(JT��R6����f�-�]w2*M���})[��C�=����ȯ)�:?4��h��uO���)@���=f�sA~�7��Β(�����=�k�uN_ٸ:rbS�f�T�c=�ִ�Ȋ��b{�u^�T(}�%3�-�`�G������)S�C�?JAo�.ń�;l^7
pxv��4�i���������wUD.��,i���[j|mپ91z�hG���P�@�qT6lb�
	x���y�J�mN����������PF{XY�`��}�<�(���Q�/��>iX�-|��!d&>˵�=3�D�],)2����h������/����"��k�DeMȈ2X{��&�ă56��9]-G�`ؖ��,c'p���S�� Z��)�`�`�1�rq.ǔ�tVqg>��2�`��v=7�jhF݉�~��r��r.6�8��w+�XU�����;�qHY_-):���RL�0 ���G���l��X/	5"b?S�6������=�t-��~�I��Qm�=Q�Vy��}��|ـ ��C�ϺO�g��*R!�ϑ������f1��,�#��	H���K���pL[dUI�4E^�	�~���G�^do�h�z�~*�C#�����Y͵n鈞0y���:A
H�V3S#W��X6���	�����q'��2�1l���@�`��_�,xf��!5&F	9�&�0vʽ��1�F������W$�	�=�B��v|�4+u'H�7c�fZ�X�	����Yˉ��Z��ͅ�Zr�,��jrA��^���ֻ1���c���+h}�ҏ=y���	�[�3d#)=qu��,w�I��t��=���"�Y������u�2��������p�@J9vA�P ��À(��0*����$�3��`G}7ga���F?W>x[E��&���BT�S�>?�V ]E`*�W����[��N�6�5�}@��5|����c)�����C�42�{�nǩF^ ��$�����ECݲ|d1���9�̽E��ɩ-m��MD����v�3W�l���.*��,tP�<C6��h������.���=�覗�i ����K��J�H�i���x]b�?sӏ��|g<��|�����VsZܓH�6ym�f!�4_�J}�l�5n�=d�`��1c3�g\o�[cLS~ϴ�XUǲՊ@.�%?i��9�\��b�(��跭p��GS0F�Q-M5��b�4�lj�OK 7�3m���Q»X�˼�����D���7����"�z.bOGG��}a�l����~'���)�;��mk�v1k4_+]^J���g�*M?{,��3?���l�V�vw_�)2��J�>Z��>2�H;�7����J1��+�uN-�뤂q�k�������>��lp_9���z,�G,�+�5������\s%��PÔ�S^!vjˀ�#�!�t�A����#6�Q����AAGгS�/�߼��d������o	&uQ��eI�P��Q­WT������p;��^�m�@t�a���o���ht��D�̣A,�3�w���7��^OA�I"$��!şK�܊{`�nQ�f����[�w[�*�0a#�j-j�T����s�����GG�Ei�pSz�"t��s%��2���߾�8��UP��ut��vL�<�[%�1M�H@��*Ƭ���.<b�쁒��H!ŦKh�?Ί;�6��8R!*v(�<���R��x��f5iC`�\��ı��ҴM��z��0��CBZ扣VO��Cv���z���/�$]��{�s�S���1��"����_֎a���Dc�a����@	.�i���=��Z"X�7��X��q)S��m8�[y
[��¿N*6I�;�d���%3< 1�~t��n�1�����I����rY+�u�~& �b$+4�Jx�Ŋ��gTHA_�s��[h�1ҁ����o��K^����ܫbMZ5���:��*�\-�T��'�52"j:�62�og��k	�4..��~C���q^�=�����e�z�L�A dB�������Z(�d��b�!��oH�?>2���]Ih\2�(��o��v�>$����m8��̥A.��B�<n�'�h}��7�}�,��k�Y�tW��_屠�*h2I=%?Id>)%�0]e�k��;r��3�V� �S����w-�,�M���M�s7]j� �"4�@�n���Kk�"��8>f�"��%��M2�w��(+=�A�c�R�����i��dj��"��Y9'�6���:U�BO�������º��X���&]J�횸�����  ۠��X1�.t?�����;���R2O�ث�ތT�G��"$���$P3�"FX]_���sh�U�X(��!F����t��#�U�OmV��W�K�C	�.c��u��.?��\���?E��;e1��uч�����q.�.A�T�L�]*�	����>1趿�&�U��0;�b����q�JQ��19��1��;�Pv�~Q�"���o�QW3����͘��_���{��f��(%灳�iŦCJI)�\�*��N��"(����<�]�Ė�HT�8��<�͹�Q��֟.Z���ݍ��r�@�QX9�"��������=}��1e׌�ϑ�5�Q%Z�<�獅�d�q�d�L�q����A󏾵cCD��������O^x�i+��kb�I�,��i����?x��XhՇ��&m��NtQ'������Ur]�xRr�isq���u]�8�y��<���3ܷ/��s��-�c���)u�D���x���s����G�NB{�� v�^D����"̚%_pdFIզp�x33�� uw�2��rN��vǒ��`�š a�cI�[!��\�$�x�ɽY�VW���`�D�ly;�,�պ��#A_p�GƜ���csQG���r����;���cܕ�����7��-O�	�i����q[O��K2��z7fH���U+�ޑ/��xDC�~Weu��@I�m l��X�W�z�xj�\���4k>n�[Bj�+��s��L�~D�?Af��`Q���6ք����c?���O�r8h�$�$��l�Ÿ��$����_+��\-0��#}��ܮ��1!��6e:۰��������(��^t҉��6����̸��)ԩ[�v����I�2a�a|�9�<���8�޳��t�ဋ �;�9�-!b1�n�N��9QK�'u 1��n����co��ճ�������|ǵ��@S���iC�_t<���`\ ����e�{�5�o�8�Bk�`w���Q�=�?`/��NS�2�����~O��X�Ԡ�E+n$�;w�/bc��ׄ��V��l�F����Tr��W!��D��1;�S�o�	�Ό3C�t���J7j���N�%(U�@�1D��A�2k��Jz#\�Q�Ɩ�ޤ���ls<#u'�r	�z�GʪzRj�+k���'"�Nh�eg����40 v}�����
��%��Rv0�~��=	;����d0��%��wWw�J���kv�<����\�9��� H��{L�)GV�֤�M���}��*�Ӝ��"��@_Ɂϰ��_f�N���d��L}��j第39h)ȗ��n4�9�3�Oh�<�B�����[��[�ѫ���'�?I��;5�fg���u��u��&a�h�e�G3/t�ǫ�a�%�n�}#�;aSI���ǿ\{s�JK̮�Ԯ��/�
E�^��*�m�@��vϤ|E3��c1f;��a��}��bز�������C�\��A"9���� �k��B�ܣ#������쮨k��&�J�C����Eb�O���x%�}J�Z
�:k�T튏5Byv��Z)�`�0�9�b0ʪD�f@�a��+��h�r+��bEd����
X�}��V��wV��s��-��5��ńL�4W�@@2�k�5$q�y1@4Vh>�*�oLlxz�髁���]s�i��X���V���1��fB��D%�eeS�~XL�e�󯼛�j	�Sw�l����^��Up
�}� mt"��7[���-5�5g��O�FoUU����%��7�F�eO���4�E�+�Md���5�����61��r��SP�+��'�'A{��Y�L�@��Ź�/ǎ���d&y�w���s\��,���ye�ىH)�'.�*J�(l;����]P�C!���@sE�E�L�0�ٹ �C�wеN��-|�-�Dַ���o'S)1Fs�2ED�<��j����DD�G=�[el�U�j(̧%����p�"��;��S����Գ�� �2�c��i�@��6�J���9��I0����ڈ[t0�;ҫ�� k�g&�]���
PzQ�(t�Cd�6\�s������b��A��]�tp4��{���'�e�p�l�(?�.�V����"���7h��~(+�hw��H�k��Z�U .e-�B7��Y+��c���^n�V�e�cR�onNr@��	�J�
P���Ar�u�k�{�z��6[�*lD�������|�%�d��u�������3X��X#�q�4�[>f������7Z�.?.�iS���_5]�5����d�M��e!6��7^��jv�N�ٔs��s}$ARP�LF{,� �bM��q�6U�O�Øx&sGs��~u*;U:�.����4_88��	�\�j!hL��{P�΅���6����B��ږ�tF�L�3�(G�H�3��Q��(E�����}�©�����`���sqÙ���V�gq)9@B,MW�|�e���+�cy�gg`T�A�\lg
��g�'��2��ۀq$���eJ	��\�� ux���1�_��^0m��JTxFGb���Fp��º��rχ�
d�ub�x��`�b3͏k�'�h�c}��X�8�C��rA�|&����4m���{��ɿ��^�i�LX����r9��Ew�����͑�m"�4��I�@��͛=B�O�p���$��#�����-[x~!���k��~��vHsC��H�u8��ߪ�5\U��7�;Xށk�"��A`#�"�%ꃛ9��j�C�&c�зy�ܹ�8
�$S%M��J��8�=�x
�hf�B��2�Yδ�� g�G�K��w#!�����?�?�]�	v�i��JY�=���S��+�ji����T�%v��0WM�)�%�a���'+�`�$���CC����3[3�y˭���\7�L)U�k�Y��cAZ-����"�Y!-�ơ��%�r�sJz�([U�+��X��U�3k�݌���#	��K�ZI,�ٍ9��:I�z�y��Q����|��-*��b����_k��vZ�կ�q�"\u�@.T���z >:�Z�U3zH�G�ݮi����mP<�^M�2y�W�U�Er�ۉ�݊۠H�]�sn�y�o��+�+}7��!�K{�c���_AK�Ƃ��e��ξ*�D%�W���<Gil��K&l�-Ѱ�酑�^����%ѝd��:sh�3R��!{�$�<R�+@=!�J:F���k?GI�������]���>��3T���`�7+D��{KY9�SD��N����i`Zs��wB4�0���k��V���(�P ��n*��Z�K�x����(��3fp6f�x�*�}����x�����[j����U��k�� ��L΢�nx>����U`#Q2S�!q́�^�:eS,*H�o�>JH���@_ͰM��F�Z�6�`M��v��{��KC40|	�	7%���Z���Y3�0�'`.�1"�Y��.� &���̩�+y|c�`�%_R�s�`�l�,]K]٬�e)�6�p�L~ϑVam$iɣ0�����[Q���B�h�u4%���#Aϖe�Z3���}r�R��yX����^�\ӊ�סq��Kٮ��������x����iD�3���=Nl����%���RҊ-��/{�l���t��{f��~ᇱp�kw�����ݰL�Y����}:S�����+��5$n����L��F��ȋ/��P���P}��� �3���0�s��>u���~E���]'�B��%�����g �Y��I3�D�-�r7��3�!ԙ��ݕA��f s.���g!�)���iM���"��Y�#�3r�$���9��g�p�ml������$� (�U`7�BŇ�n
_�¬��5!�#���&�������%��g�Z���K��ߧWs�	��j6c�� � ���ȉ�yVϪ���H�t�p6]Eqȭ�)�簾��X���ׂ]�ȡX���Tpl�����F�z�e[��<�^d4�
YM�|�QE��Q&zԱ��
[Dz��mw��P��!��>��-���x�XO`�u�yT+G���/���8!�M�q�����$e�����2=u��\Sz3�X��������4��y��}+"�M8 B
۵���FL�g��jF�)��K��ng>g�k'�:ę�=���6z�M��W�	Lt#�/�w������U��	��l�%k�l(��&̾b��Ʀ�}:7�~~�5��Rv�wN?�;1��F<�x�w�]��A.&ze׵S�S��K[��qM�(�vx�D��Mel,)���`'v��?\F9�ǿ���k����`K��i��?�z�Fne���t����/���|m�ҿx�:9��)�@��{�B�^e$<���k�V�k�TT�}�@��:��S��m�X�L��͵ ��K
&y!ȹ���uI:m�X�~�P�J80�'䜔d�t����?�̊n�?T]�PQR	l�G��g��aż�a:j�֧�ĭq�^S�>-���w6���s�b�t�D�,�L������Lx�3Ww�g�$��EH?'�bd��X�\as�������FE���!B�19��߬�%~���X����\��듴��4C!=������M�@�ݚ�rG��p1�U�s2�"U��������/�W��˗R �D.�Q�>��"��=����uZ��'5�D��T���o�X�ͤd��rӽ� ~���f���w?��D�}r�dݪ��,u���?%
>��\��jFpŰ�������YVz�F���#X9]��EW��ig}/vF�l�T}bU�C��'�-�pI�ho7=�0�s�.>�7�0��}�e�q�J8�c��""{q*S�"ܞ��sYڲ_�}*�P|�q�!H�d�Ѳ:T�њ�b��w`��e�!"���~t�/�ӗ�b�S^(�yp4Z�âg�ݲe���i9��j6O�l�!*hV�ͩ	�n��p>\i[m����`��y�Dm[����� 1�&�{k�+73������
���Ȥ7��,P�C�
��`6 ��¡����`��.��>s���4� o/��Pb.��{ M�V�T�V拏����c�1�wf-p��zMSb�3���hW�3]q�K�$���J�td�	G�]�����S��De��z�+pQ�Z����E�'𔗅�Y)�#�z��h����]�vX�f��rf����*��_�)���]�z��Ϭ�9�BtGKK������7���*~�/��F���m�c}m����ڗ�e+��)�	����,��E��vs����l�cNټ(Ӥ9���FKf�\,Z੓�_��!.�Q�w������'A_�v��
 �Z�4.��˸�؜���S�Y3�F}c�Osȗ-�D��#k$+h��
��i�lc$#�/pл7�+���/���GERi��i�@ץ��F&'jm�#��vd��c��QX�
wB�T�iU����*g���ф���(�*�,�bh>89}�mZ�YV#5�c1rtT�<�jX�ؓ?�KޱKxr��B3SXn^&��2Ʉh������O[ٛI���>�����c�GN�����s)�����h���v�t�g�ݛ���'o�Ù�g�s�{��5c�Y@q�G��m�2+t�k1�[���9�^%9���ӍXN�v$?��i�e�(�.�^O$0e��s� �����kQy���`�&�\w���*.�Y�5ٵ&�OxQ$��(ș4g:�Z|���k��j������+Zc)��o1��A%���wʱ���\��-��������2W��G	���\L�ʁ�:��}��S^}/i��������LR��`gM�f�����d�}c�l�q�0^1�P1��_�SI+J�S��b�^�x�,9���?�]�����EX,���w�a�ِ=?o�S{�>�[���?ƢZt�C����8go����F��:<�_n][���+�<dC�q[�k�ݲ���o�����������{I�]҂t�b�C������|j�98�D(���Vk�K��mfg�Ҙ�P��Jǖ63�jlSG��^��l����E���Mު��1@��7Q�w��[	y��Oؕ!NA(dps���{q�7���TqIF�]��R!a2��N��'�X�ֱuml#q�������%gn�n�1L핎tY�Q����݌�=�`�_P��)`%���)$OkM���p]�嫧�^(�ƑPx����K�1�@,�ݼd�~����,�R���q�v���4D��3�/jRs�sJ&v�K_�:��a�\���]H����p��rcΝm�րR�s��,,�B��o�P�8�1���u���+|��C��۠F�龦T�sݢK�.��q4&��Hv��TmjIs���t���}6�A�����ri�H:�o(y����}Q5|x���glm��6�g��䱥�b�s����lG�e��(�ӿ����Yc�^����=��_��u%`�HT-��\-j¨@��
�}�.U-<j�1�cfǛ�F����W�7�0jc<q��P"�L��Η��w��{���v��W�����?'�	k%�h\�O�`��r�5F)T���O9��i���������f���w_]��6�<SN��ƒn\��`1����y&U<O��iʰL���g1A����f�aZp�CH���{~��;Xǉ���=Y"푌���;&���Sl)�B�U���%��|�n�뷅[F�ٮ����M��w�oz[k�2���XK��LL�� ^u���mO���ڙ6>�66�h/�����}�=�"-U�yd��G� o����3�?��(�
�5�E�+�d��hD�ݗ$V��ï�C̚�W̚�!x� NmT�1��Z��+�p�J��$Q��7 $���"�w&���y	�ow�NW��謳��~2��-�"oY��y�P�݅ijiU$D�g�4S�����h�F,����U�O��]��;8LUi$?� ���/�Zc���3�)�Yo���	�[}i���L�_ǽ����굨D��e�|s�c&%�:EjA�`W�v��ț�Z��zC2�&a�R]9��b$ ��\!��[���BD�GH-�ʙМȥ�W��+��5�����B����%[4ΪQL�GP��� �Wq�b�=u�N�0��G�� TG-�X�x�ˬ�f�Y� ؔ��zI_K75ha������_�/���JzY���s�<TAik��~!�6��܁��p@-rG�h*�6G�T���}�Zb�8��Q�,��i#��8?�Ɋ�C{�]�doR7�1��ٶ^�)%�77�6�Jp�Y�������x�_�tw�]g�o����*�>���O�k����:��cD��N�o���S�