// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
BBp+BD3jIecisSN+oWyRaqgnyiJO7z46sU5asiESrC+4dOQwxRAnvchArtK/1hhQ
IV2kgii8tJ9U/XjOCWADMucj2UUx24DOzwwEJ3VzPE8YNLym6s8wDBBxjig/9NuY
1YSmvgVK2GdHjfNrgA6+z3lpZVhFQrNffbwp2EwUQ4M=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 23296 )
`pragma protect data_block
E1u4SLqbyc1gko++e3+GdG7pxv4/yLqKashbGn98Zn0PEPY62yCVhBVkvybEM1Jp
vxOnPRRoQvsjzKNOMbf8a08PwqPjYg3Y5MYDVm1mPYXl7WCdcQw5j28u0rxsvFwO
WlRSP+W26gF4z/GBgb3jYy/vlAy6IhWV4kl1IsNXLRouulyao+bjaS/+/hDg8meR
DARuuVmQEiPc9EoXI79mJnt5u5Z7qSC3TtVSrjgLRa1qudObjP1sTTK1vl+dayuW
Gbv08owEVOy7b1yiWtZvj3AL2PUTClUZ7fHpnlOPOFeZlVSEHydgiP3qsiydnNTn
Oy9S2UkMBBwO/LXYE+S4oQFNk1hE+o5cixGCTsjgeq9OzDXSnMft4iK/WFmfIWIa
rCa7sDOTy89nN3eBJCM4H2JBOTl2hr/WRoE4fkCP+xaOBpwcgLz2oh3Et2jhsILm
oeGQ9uLv62M++AiK6eHK/7qH7ehs0x84Qko4zJNzznI0LFYlaphXpLAkn5NRrLG4
nwueGytMvje9ZiQSrECKWnCeo6LrwZR4jFUi5MP8NFzZsQbg1ct6zDhrpKNyHdu+
W910XlpTwM2rYLDNDSi2ksNbTHw1WoZH7hN7Hp1cQKqbmhLCs9tvTXYx+xzJajkN
ZJ13WXBWy3fbmu41eKPSn0XBTI2zb94JXwBlT1oqjZE5VGTcpsLyD6tiJEYoy/Wa
/g1RlSn6y6eTY5Iyu4P23l39X0yDbg1dFrK5TWoTECsokHoH/1kAb/jrFC5hbJE/
3kuOHvYDY3p2sJidyCfEcQe9kx1BLUmOPkQZ++JhEnF02nPeFo7DkJtbDMEqBCvN
p/rVlZs07wRc4xGdM6p5qwI3qpCwRPce4TjFQ1VK1TUpzwPa37hvwRjJNBy3QrfJ
VRvnZHpfH6wQ12rpHOAKfJTut5wZvKxvnuBCy/g2DBnLJne+1E4kgla2PvfxWeAA
BOJ0yB3BHE8dmnav5QQ121EK7xIR3VsVhmJEoEK7t1fW8evRxYiHbIQaZA00ccaQ
0AZ3GqQ/SzmkHlTUzxg3uH0Is27rWVB8sqCP6a7u9wgbUuNDDD3S01PtovQIQV5R
5YGJP8p4IowBQjTF/y+Icv5Pjp4lrw2KHxSPM+BhD6NKoQRGBTxJTHBlwPHxO3D3
Y5m09lR9JDFOFV3yTOTnmpaIUFTINpbJEkuWp7PvCU142oGDASPvFX55qIB5xTaA
147KkExLg9mxyA1+anmSY/AfzIHYWwMrH72OfT6kOsGxjexgHbOlbVRsnQszeWMp
cSxX7712mAu36eNdgbj7qo/7qKzudM1HjlQNH8cCimbyC7yZjGEx3OLXfOHvXqma
FLqOg7fFSjAtGa/5zSFZb8lQd6s9Y/qre8GFFZCGCNCBez21SGru2hga0Z/n3XzG
w42qUD/uJTwxkT/cLi/xFIVwPyCEc8hbHJ4NydiGArEe8ah0DN2bhym4OyfSxVlF
ayT4NMtqHYb2kU24is7I7UFcsfTOh/9JbLYhYnYoLIX2unySb3e78ShZrIt1RjSP
sP/wzSFX3gbjiUHdx1ughasrI4h6OTvrGkHI0Kek7PRxPtQ4aIEtA1u/5U0I0ipv
l8vg0v8y/pxzOwoELDJeLroVf5dni8w8sLuH4FMcpj46k7eVT31CLt4IPNnAXsYp
PtV58FMpv6V4QrdaENGB2GdvN0RPxszJuZgSBmIbbPZaSfrKVLkBRrMlTfjaC5CV
BPlliSxa9pylIaimpnnsxwrxEpxELDO1omUh0Y7M3sNpLnlwIgzYExupIPq5Isbb
Hcml0dcv4yM8kytj2HCDTLDIK08hGc95NqyUvLJIA+7mM7oV6qtmU+h+w+iUBZgm
FcApBy8oW7DeEQ89vjd6kmqrCGFOZOsMpHMijmbxpVDjMgZ5MeEG62upScudOFHB
IkrNsBpbjx3aJfCcQUacx78OyrgGR1KXm2OM7I7S+NBkDCR/WbYcoW6V5LcXACrX
KqbnyNtxEYst6PJwMPUGpq45sm68AtC+/nTKpykHuxnS9EK+iDFYYnA43JrhlZbO
/zM7F5KEDeNzdWRyJ76UAuUUKfgMl86tC6ow66w4+TpYafr+yV1enORYOs1EVWTM
6QPYwXPcgjttORPKU1FdcTpReL0DUbz14xUmYLmq/gQXaftIKeZC2aDocdZQCTwq
509LbJemNo5567QgKheYRNXQxGvr/Qn246rCUzdYGOU81Oc6MrZIM/SsVl1ZLgNR
Zd4XFvdGb0hFTTFS1gCgx+SNd45baGdt0MwVQ1+FYcmduJOvTedMIV1ALa2L2tML
t24myxJIryrlX6NLRjut1zQKHvvjdq7iOcrAAr9/g7ypJDbNsipFhcR3RTJdbdJK
UE7ptHryDiXwccAkuuJBXsMySojozPz+A+AztTxxlnJ4Wcf4eeBJFr9GbNon8sGD
JqhqhxVQugUvxYkLf+7jsUPiiVQWHOhUbw0dLYD3oTXv6GlVoqtEIhyjdQ/T3LcJ
oiQHleQ75zaS6CURBftNDFVhDwLnK+gS1IN1SmvZCTqC25gJbQkAeyEmQg7bUeaX
8bT0NhWSoD60WUgxf/2RmLY9UbPTEV8iWBp+Cjn3qK1zDo+rmQR6I3MZb/t8XB9u
7tfGmMnLAq5vKr8pl+fBrf6zai44qGiRliTuIMQzNvmXGVkY3Q9Cm/5bL5KOZmkS
d0u1clrke5NtrDLkpIiho9aBRGtfyn87LUfd0mNyO6vE+2vxUIqSECw+lrQtmQml
EVis7oS2th2S1tFkcxIU2zPne2LXBwdM/8RLsWu9xoVHhTpnrMykPMkePxE6gmK5
9WTwUYK63ATGktm9f315xexaiXVkbETeZ/UDkJ+5hHNlyXg+Rnl+jkneUwlw8mIV
JXPOUd5FUHwyaeqEnIlcChylu+DRIH7HdFpSU0dxGze+KZ47XYYRFaUnSkHYDm28
uE/tIxGilnCwK0oXsYGDtuilLxtAqy33iOvS1Smee6k92dXlrleRRoji9o+JZ/GT
Ojp/2fxnmQN9WVK4d4icmLqUZvpRZypIGPMRaZgSm+DURNxm3k7M9mdEkV3dKiIT
xMyvgvpNpyw4HAcDbtUKD2cd3yzqq3TRi5eOk4asxGBu26KYgNz8UF3YZ5qJud2C
IJOktYbCL/glvU0PuRnWmGPdT9JH5qaJvXIYpgfd3+9pwB/CRCWX17uUHqlJnYNm
mT48pCQoMCu3lvAOLFzMwic2p3yLNv+As9hndowhIHhso0xGeg32G6QvDTv+5CKU
DCSQt2Tne3qMMMY5BjbUqZeLdhgeCMKWfGOTi11y0H8/GAfDF7ggvNJT5cYNMJVf
4zwZjItU/ct6VkcX1lYqkrqvOI46jsyaPEEMkk8RJkPCEmJDph6cIEdOHVYMEM3J
D0L9I0O8TxgMOxOwxSbTnu8fDryRYRhFr3HWYGv49Gb8F2iGzRDPuEupOgFpE49f
TegrH8997Vx7nKCXKv4nUVZLDrCNAgifzuBcsFMjrV6X3qL2KWfvDZqA7rkIVLKz
izp+QG7dj1UyB9KI9HHW9bxlS+FV8pAJkmeIFZ4n/uUocVriRC6rU18aM5W4gzy3
chFAQCVuWvZjncirjzdzmuGefBJeLbwNFN9MNCeLrASkuNgxl5eLIIrKepjCAF/W
+76QW4tp0n5RFl5im78LERtAk373ztwj/tmbqv1w13xBSBbazGCXDQYTD+mlothK
iKz2FbnjvN5Qji4rdeoPkrNbnE2Lnfz1Mg/NKIblAY4VfIXNYVWTnGmw8wGamwOA
/XxmAKsAeErVntyrqMEUE79Kx9o7xZ+cuPN5DY67u/zv8MVGmkFqqPN6af87Iwj2
6UZ5b1q45IVhANl5rA5YR2TL+sSdznSRxcg40KTEuNB8wubTqvCNFi2zs8f+1ih7
nnjTJOw6nIzC//PvX4TJoSrAUt7Q66rWbB3DvMZrgQoE9CjLmfUZjUF/0lnZ98Dy
pHMjUEH6a4D3H9m2LUjXik9V/hMhjlROucJEUftQklbeEO2R92moBvm3TRK7ExMS
E5KU9QgMwfFHelVZDYTIHVegPUsTE43G0vvwzIBaMQCNoPxbf4eK0M5ft7jp45hf
c9Bid+OSVJdP00W72B720VIGABr+b1k6aFhQqUvM8hfuGqA65Ziklnx2wm14bWnH
A/fWqBhuBOGIOR2aTf9MuYiB+nFUfu3qmuRiMhGSpL704c+euoWdesXgPMlBu7Xs
3jblNWhUcRyQXVu8nJQ+k92OiK9NHiAEcy2Ni0a7noQDmKVNf1/CyVW1keyjAIQ7
kHvFoWdLnsdCk7zONqp89iqlprtIBseswf303O4X9NZwF2QkznY0Pv7kpFGjFUTe
7d5BkNyvRI2Ml+mIWDwNY61I+zH/Gv21ReQ9cP0LhH0h89z8FTR29T3p3qDEvMbg
xTlDLXHZdyusLHJIViio1S6MT/h5sx4PifvXjzvyrkuiUiPZrtGrmPrBr+/PFhNc
P5qFbm+VqCuphRpDzqlpvtu1pqg5VJHv8H0jlt58RCDlVj6WaFAOgdc2fDy7RvDR
S3eBA5D2xcDiW9A0bwOz41ZyK1HSQPDSmsHBqOYBHgvAi0UEMQSHiiidh1GoU77U
l6I//Gr1iy+ppw6eROl4orTTV1bn3A8vPP08awjrCFxsmMwvu1zusLhebO/AVT2j
RMIfuSCTepq1Bd8n1x0MJxdoBPmBtHGufuUlIY0jNqhDcknBLyanKckiLjD4P7HM
y/WL/RPNl2p50rJtXs/3cDrpuQE+Oc0T9vJ5dLzIez2PjvVCwXCPskdRqL+8t723
n3s/RmBv6Yhg6nJxK2rKX9sKN0mGVO04BME7ovdtYUezn9BfNORdcfDGSZpXn7KV
3IgH1JIlpbHMuHniPE8mBzbZukJ9Pgzl0in6vi5Qe9kxYadwpKTPQMRK8W46w3hg
1+4pN4xsCdecOATjw8H0/juZ7edOZVQ7hPi99SE3idz3Yfu3aNcaJDzAzVYWBpC3
lMkXp6SoLvmIf25EZvEmG7hEBVYbu5teJeMe/It7pgnnSGJoRqasFttEu6gmZ/Yr
WF1/Rx8/8mFncVheyoSbUWggT7S4WHik5fD8zIy2hhv5vBYwrvva7P4Uw13wiD/r
a4rmIDaUxu0wH2rcjnuyNw2j68UBRXP2KqX5dGipyVhB1qR5AYhVRnkARN6sStB3
UWqJ95NLAO8cwZBP8+WQ/kHWxN4X2gHDpREGvQYY5xueFdAKKpdpHS2UGziGCKt+
6uKK9YOKUEPeQ4h/1E2KJZqS9tbHEuRrWRVNWMdTtwoirju8+5EK6y1JXU4rh77/
3oXOm+CjKf+mqiNm0kL0v2vvZd74eqejxfxk+8GNFV8hXwvlKDDc2KYlUceGoQhZ
duiB91oAgIp75EwYtVG59uIPm98ZQRE0Xcul+NqYAJv2LgUrYMKYQ5gVL85U3GdW
fEKQwnD5m5Th4P+qVmucVmE/yBb9g+P5HxbUT7W+XLEjim6bVYrSA+8UP9agkv+E
prMD1fDADwZ0vB/lhZLHSqiTgz7ZXKAP4I3L6kc3XOtuFvR0Y8BOunQbZ1wDedO1
4AkN5U3+6LFaBS8zOAOQXcBMXxB6giPxrJp1yBuK5M8/eCgc/5Ue++Fh1t2o37tn
I3argCJP8U/ipnGg2+KTrTsPWrFm5cANT/xa/0qo3/o7qt5dyscw7EoR8V2010u6
8yDirq6x1I2PPih0nm4dMTYOiq/lepgC9jZQDKz8aVAIwSJsG68exzNSK5sEJpd1
ipKQCsfjQTSqWyfyvnLTIGVNgORU0bkMB1d9eWISes10tEOUDM6ULAh8YCW/h5XW
afPZQnjotTpd7nFtvaZwxGO9Zs1N1hUFg7mSsHgyvNykMlGUtR5Nq+jil67iO5QQ
7AlFAFV8rsMeZ7n4QTwF9+H4aMXhH3G1d0em+5TmWqYc4MqkAaIh+C79xZpI9VXi
qa4+W6MKvR0SehFj2DlLT69VuNIAhn2ByN2pIzABmQNPUh+48X3cZvx6yiMiG99B
e7uv0f7W5RWWAqPLidS8+KygLWCUYlODlnIc9Apn28UZQyOJDsoQGvA/DZh6xOZx
ULuUZ6kS+nnAJXAqqFfBBaZjZx6LyvpeXyLmW9W9BkuFT9WJC9IUbog7J9E/muad
ooGnj7cdjeFpNXZHvNF3ywZGSUzMJ/ipWfU8prorVd76qg9rSRMoCNBe0NcOOxIa
4ZJmwwhhAV0XYHJKFCWuT/4upWMHAfkPPEka030jxNNUdRXzNL6bPMUbclCQo1Kj
mbFgq664/zT/zdXDGkRS3nyYK2zOtL9tZoQSImvRfzUeSr+/UBPxdWbbZvRumvl4
pj7sx2wbGl14cA8En8FTtsNayM12JgCSw9eR4kr1wYxJTWcy+rRDsb4Z/MqWvJlV
ch9tlrrfbh4jcxRVEuuf4Tc7rGUllZBvfAgFtFl0zYYBUHw9+0Ztr01sdF9o9qaR
3tX/twWo9+rJ2QdWFRka0QHtKuc8CK1di/Dzh1UIdN/8K9BV/0WZniqXtJC357NQ
pzzUYbCS9I445MdLcrYitrcfhF3AFY/3MQKDOivc9L9L4wQMX75o7/DSOCpggejd
uN7oTmYj1cj6eVu3BlxDHuJAL+cefHFx/TTsuLeN/uAGKLMoooMU2ayihJrPYlmi
jUziVpmWpBIq3FGnf7H6nN/76aEp04FmO3IUrSVlKzi67LGmje7tVNb36r+Y15s/
q20sH+/67JLaVTvSMUnlHvlZD/jOwqHZhy3pIZ4B+kwhkq1zZlOeEx8aZWM/cTQq
iwwQnFAVdfoQ+Vajxb+LGvkNpcTRSad+CMW5S0zcObWiJ5OS19YZjvI1+GuvVoJw
OqFwUawS7jBuh6es6G+AtEvNeg8OxIjL/U2AFCvI2UpjN02rbH1FyhZD1lswo1fQ
uAcka9OvZ9UUosT371OakeasxxZsXnE85Hf+HNb3AUywnupoi8rvKRF/bd9nSvAu
OWEeu4evlqn50umJ8L28o63Z4PvOfEflelleMbrZSJxw11g8mYNG8zB0wVRGLTft
Tj6WGIRNtnz65LWuUBRaZzHs40iALK+1Q06MJZufshPkVx1297NqwGMEHUbnIzSJ
HR4eloWO30GoLsDfkfg4svOfUQL2fKbgphtUx9Vcw6RKVykqC0ZAXMZgVMRe0e3Z
YhtyGRUENPoZio7KlEtV2wedncdKbfffWIfMr4UyFTuP5kTv1hZeHv2XJ7LAuyl/
9mFhfDXnnjY8HYvalZirBnvwsibsyBTU5SWc3q4t4Wf1443dQg5zuvoyxscU2ge9
fCNp62wbdG/P9nXj+/F3cUREQS6Fg6Dq9nTe5ZIOCLFcy1sOUBpeKea4lW4nlWEd
5bQnvzlXokZipG8qbul1YUpy3810GCj89ikK73c9Gux4m46oZaharDJ6p43J1pHt
SSwa3F1eDoFZzqOQo05iFfxR52PYd2PD9cIkxIUacD8wKb2lO+HIYaxLO3qdr/ND
rAN4hgB4l3BiSGTsmB4waVxwinebl8CHMOUsF5Lyyht12fwMQOgiC9jWtyRzhHB6
7bmsT7ikLMCAdPO+0E87gR5yJ/nHy0trjoz/ROZvSQc2pHAPS/godY5rqLt/xOrq
m/EQkjUGAEf3VrI11/tUXw526to/JlR4NWqQ1ZwUQQBc9a2nvNNWjxu5bOLUihEo
i6hf3m/du9J58+TyY0Thworq50dP9mG3sEta5DnwMMqiPuQ6kCBwv4Mlc0hICPjy
UfuaIBX1faaby1EZ3n3yTL9FPIBVD3cuZGfo1/Yw4K7qXeQ+Pr+VcpAAX/L0ZAr3
wOkQ7nHvIzE1wLvCZBc9M1t3xq+8WNympt2EXSc3UwhCIlHgixxadPZmJt3D3c0Q
mHwpSjV2khciHj563lgAX+sBkcrVusR9VPD/W/UyWdiQVh2ZkhpZIetXssTYjZuH
26dx0MgzWmHxu3JJTTug6jRKjPJIeXmc3V3/2/AlkXBeiyRuVQeNygB+SrwSifmz
n6ItIIvQvvoBT0eByRmdueNhgzjRmzdUFCi9kVKc1U0u2OG2+yR0BgszShh2iVky
n6/Uub3MKQamFscwQnuoL/LCaLFuRmxjrURM3Rb8HNB98knJ9XkDQnPbTBhDRZ4S
RIqrbbHIkVPatNRWnPk4Fv4FbfJzODjmqtO/70Ag1mL9LbsKSyhFRnFVwKeQRxo7
PIR/RUjV9TkjpGYRBN03XNY+fIXYg+jOl5fdqVFqD5NrgK3qOgPCBjieLF4DtNoP
ZfA4Xt2yazh/uvqWr5zYPDJdTPypzHu/aC/pkrdw7zOs+hry80zPgJPQL1cyxeSE
PyfiWtRJSyQDsceWsYx27ZTLp3bt4UoS2nhHEtTC2XpyrrotP1f6Z21a4RiVnbLT
2EMIbiVtFUI72Kh5NA/akQ8FmzdbolbhHwfb5oHRMRZ2IcdOO6E2kFL13obMIc78
UCi5ulc3pr+9EvN/PDANLmK1DDEeOIOmQpL+zqShD05C7wz/sw5f0qM5mdZ+VZMo
XWxDslCxPVF55TljNVJHYGGxy812CP2Abcjl5ocWn2OjM142APwE7V1rJqNJmJMj
fS3FIztbONEteKb+VfiME6KSsMe0AUyaXy3SSXfNMyUjuOUSTbLziWciEcobNLbc
v/8Y25g/0YdSzUTw1a5H73PyF5XoEIeYH8UUGifuhwrnd/q5rZ+g+aXh3aCiWiWJ
1TaWZSOH+nfBinp/7uKr16mpmfiAJxrVcA4qbUDyJOu9E/HK3+ZAG9xw6+s7WotT
G9leSu7frnpapXb9rTSdakZZ4rzF+t9uRi4AhVGoyuLX22sYKViyW+vsIMz7JuOT
Ddkez+9q2WuKN72svNkiIx8Df7g9kuGrn+usrooccICV9ZTmCxbHoaJswDK3EIOR
ls54Oe9cYc/EMlQzT+CvtmrnIfbX+P0iQi2W0OXw58pN6jgTQoiC88bOUy1fmxRt
EOpO4oTILRVqbFFcdPwQ4KdVS8omVDQppjJqukI6e7ycJzidvKXUB/D/nPQG2vIN
6rRV9fJrOKBmcJs0H2A2IoSoFaRsaXfGwfFxZsJ/dZgpOLMVgh67YF3qm+cbr8b/
Qj9nNa+Y6sXwqNVMmaXmsGIP/HKAatE/trNvsh+46df0Fi3icQUHIg8On7MuAf78
N6aa/UlQmUKzJNtGbMz5kFY8uOp07BHoq+xSROrcAUfBytoLqNYXm3RFzQIUV3lr
mtmUuQnOmKF6eK1zmU6rzsYoanNFtCgzp887gENfWCdE5tuV2it7514hBGiCKlg1
3Vy8ef/uqy9jom3Q/Iga8ZnOAREnjEhikz0qTEnKy9n7jv5NkivbcJjpKmBGmEp6
wFSEfQMA9TzMRbHARTx083tDjWspxK+POCHx2Jd+apaF23NfGmKFuLAgY/vqdxeO
AH0A2+E0X+TQWh5H1VVlOjXJm4TAPRR5HvWTV1nWqPtjoK+0U0rsrnvk5vXnQa1v
oddQu/TvMFjYwN8DKodtxGlSe09Hq5mS04bKhWjIwtlpeAfwJRklkntqjB5oKmey
BXk3pdFXuzjVs9Ypxv9qT6zIQobpe15njTWoKLw6+RAlohxrQZ2UNTXsUyQR3IsN
NT2FoVrb8B5fVQAuyNltFshvSrR5xIDAJtWWYbIDMBMmtPBLohz/oNSejoKP8sMR
ZLP+0o8ProB+DGRfWYReTEmyyxY8TbSf8x0OwOVYn0JITFML/tsn0A34N0wkzcEl
lDXRhPqCC1BCJvBfrN4u3Gz0fwexuGNIsoPXAg6+qUtZ3Lgf2Ng0dCStLB6GQjp8
m94gmPYlUbjOZp/6dZXOkChjOlSIs2n+rZPXaG1yCPR8qrK6yojSXdpFwwcOWvMB
ErVHnHyTZvIhguatU32xKWGnTeoY5xwcGBXtxM7nbe4QRyiOcyaK+1Gmbab+IWNd
qIkpZCQX9Vsp4XX9ppkY1BaHJ25lXybJ+jKGWuhmUPO8zlVHxn54jrjhL+qxgsVQ
Undp+b6o2n4/pTsTIRfsO7Z2BJ7xfdebMzzKHsurXtYaRf2uFpgNLfWxJXVhNPrq
n5iAHDRcu0obF1ET5eFzWbmgONTc4misSbTiuEPUQlRMExRznBD0pPTaW4cVWCN7
BYbe2kWIWl/+yvicCBRFqnJhGx+WGQRLrSaqdf8ChOXRAerNb7gzL4E5S0y+AbDk
J6BjAl+0PiVvgqehQWyQU1FVfa8vIz7s50ECtqSL6XjkxF6T9I8P8SFxw2B/K93I
qiyN47UwB6v+Wx55M1GuEpfPXCKobbxVseslJcM/YF4ml08FUJX6Ia/FKeH8vqxV
C7YBYI72ZVPmHgW7QfzCIdjLodw+bUH8gphqGvUCrJ4U7Kmie+9a6Ihphu3Vy+vu
7eo3ACy+DIupZ6Wxr5YH89CehjCKe+BDIvS5nbQY63Aox1wjWOiXuRjqnZOrVGOX
PGf+RrkPPlsNQww9kXWQymWiAZ2jiZ0YkenZATPP3+wib6MXAXEQjNSTZJyS+3Ru
LmWmICvPuLTdhLWpfjW7kgWDlym406bldCxIXHZPjyWfG2q82bQruG4PMRJV0TFD
5u2ekrq0q1HpMFwbtouRV4YeFmzZngA3BjZeJRhtP01IkyxG7G9QW27Ce1+J8xdR
sO0qAl0/BZUmgOAH/kgfroflD/jYmn3MdJWIIhQauHhhpOY+eGztxIhsTmY5OWsX
y4Ig+23zB/c7xlM7+WRZIctwmDDWAIIyxsQKkigMbHGO6fTTsMAiwaf+8vFPxbcR
B2GkmDKmBh22mzyNK/2SJ9WkXOSHfXbrXuF8u2DAaQzeiegZm9BButLb9/dzMJgR
df1T0fRA+CukjPXrE2s9kLELrDJbjD6qkJa7CxtAy2OasuEF2kZ6c0YpYhFolblr
jqxjs7HJEgzlcasN+DBcNblG9qFVvVbmGWM1qiN8qH2W3+YlWESxPbBta+3gefc8
/6mxO3CJ4M9lFlG1/ioe25XiFk/lbq0KX+Rtk4+XB5qloFRIhfVkdQVGh/WZcELn
4tlf2sYIpxfLRXzsr+Lej5CbsNfNM7f/qLGyY6VWZ1kMUGuA0HIlW0SCMxCTXRbU
C5pZ91dZhqmqiyG2GbuiXsJxRnSYwoXXBhMLqo3nxcXJsqTro4qS2jHDNndl/MRo
kcZM9zpMtac0l7kedRo2v9Tjmc5EYm21UU1rkLsG20DeAxIjSU2TFUoBV5iv5Vpt
3EgtkOUpEwekYkqhw1o8uE9lbJMqqNmqvQ9UWkdFL1P3lM7+G+dtdSTxVQn4Ovb6
t5B69t5y7oqaje40LT9VsRdX3wwAlcK+SipYMqvJn+1XL3N6KDClqYEtE3sycEKQ
fYEGrptCWRJ8xIpP5sbhfAz0npnLnLH2UzEJCPKwxzI6A3LgFIPOIpkqpXOKV3y3
akqSUohySpKOeF9ufVQGihIqIdqg2WuarF8Ezmo2FWJuaRxQ8IOIXgSGnUpYlYdp
16VRIkFCrAoM9pd5T6EfJdhFJxtbtWkL1bvbOrpAm19QwBekvGaLq4HTL/eeO6MT
etZMIHjUkQyjCq8F/jYlyseYdSjGC5fDZs+XS58MdnNSu1hjyOyIRVNxdKsurUSZ
X0klSnGldL5wFr1pXf0faRC1m9QHG4lkbYHKfFks37aRemHeX4HqwvC0xUc5YAUT
/um3GwiFA7/lacv0QlNr3OLE6YqnnAAA//Zx+4iHetwgxqp69Tkcs8fJOyJQ9amD
ljyjp9pff2/Kg08pdchFPHV0ENx9XCEKqLv+3f+UkpK57z7ZMq7lHRPkQ3YW3HNe
lx1TygoyzzZLLQoHhGnfS3P8hzA15AJzFfathayNRf4iju9+3n+g1NI0HAlxyzTd
Kxep5mKLfrvqK8yl3+PKf7osTft3Y1qKcPLuvGbfRO8y8O8o3y8peufmfD/FcGqC
vK+LjvYezRj6v2GhY53B9WlmQpGaFfe8HMahWMgCqazq/PR7WuH9yDPNDf4clQsK
fCfwYzXlH+qnlybduX5mTq9kX/hqHYl2ZVhy+9LRRMI5DtXYdNxyaXRBSPShqo2g
f05FO0qypP9fNrUnMqSzCocz7HV85bGkrGOl3YVDiVxD8fX4ynRkFZsMr557niXs
WdojLKqB5ROSRzZMvWjlJhO8/76z6NKQNINBUvrQi/rV1SbLYVBEippXEsSi+N2P
BLdyetRGbz2r6cjfuraURpUZWgYq6+XLJ73hgrxiI5xkNGSWP/o63EknJEvcfjtU
iphsVsgiG39s3iKxGeJshZwe2OaTGSUtCaiKdFMVHgPm/HmGOwccImdGlfiLTJy4
K6lbmxjr+ap+Ja7G/g2af4P1/+BqNX/+3iDfgk2oc50UUY7Wqv1dIktX+62rdwpG
0MlbWfUOI0dFtMdpsG9h24CgMlkCINAUlvmsSv5V8CaixVBNn0fKmkD2VwhRSUh5
Y0NPwoo8pOCfhGL562KYVSTdANnhiB/RpAXGpNsXs4p5Hll9xtYS9PbRkFhjoek3
biWjpRhI/hZgG1W2apWGP1cahvTZcL9Hbp0qx/VIFWnOA+Le1uxNMGHip+cl6S2A
UQxp2I+66Lp7qZ73qezVK5Y5Cmi2ppwWMrn743L7dWQsRo7Qdp9usloaevWkI+uK
qTH8nionmMtTsIxZ5E7aqEFFZ3M6iUKCAgFx+UjfRLrjNp9HwCTf6283Sn2h+8ii
A78zmaudjq2sV8thb21pxrmX36jUWco1yIo3kSo6/+f+nsoRMzgHFM/bRxpTCcqt
76L2VDAoJAC2y6NNav8UeBdSQFinG93DmOBldsayHR+iV0/5HPg9dxeQRACbWDv/
aELuFBACYEZaAVAE9XfwA9BPG5NeGOvO79E/DsDqOkZZ2+gCkrMbTZWWBEVQL9Bw
i6PkVLgaTGnj4oe1OCxpBc+ownTMVDjA/RUKUjPph1EVDkMfEZU4i7yomxWtZ8YK
kLuRmwrKvoeBr/Y2PV1o7dTjeE5vYAoKDRzcuyqOWuycqP/0Mxrkmc/Zonj2SZMQ
cj0USCeZtrH+fcVRScG0ED9D/r2GVBtmvBd+NBqJ0JrU/O261bVUrgCUKWupiZ0k
yxuuncyc60qUmQ1h4RifkiyCvyXUR2paX4lVB93GpIColT2zMSz7aTv+ZfU3MrPG
RuJCaXrnX2s61XZCyQJ0Q5X37+NNiA4x8Iihft3Q9LgYYR250ehRuWG5egoXBsw8
AutQqs+3V3BgAEVitjmY/u38HoYKAf0eZ4tyTxsSNUQIVQgkR4cS9RZi6C5MkKcH
tPjjlHjw3m3TU5wOe2RPrpFl8DPzsbaLaW9EgGyxqeEofyqTEi3mTil17YY4Z4xV
MA1fsdtJ+WriULnXnBTWDPvO7BvFoEKnkw31bmp8otTz9Q+qnJtix5kFeg+BU1Iq
Qx3JBpHMPvTjwvQALKhawm5M4NWn5qI5/UeIKYhz6tvhOfaNFggS95Q1Rf9b43NX
tWjKKMIW6RuRgawQlNuJ82Vw8/YRPEbWXRMAGvphkzzvCNIj9Q4E8ihOSjdpDwJp
lfBzWS1Srh7SwsWJmDGm6sxpJkkNQWF3X3TxoDPdA6eIyqoHS6/VsykQCnMBH6DI
Iq3l0xS3vTu/3kM8DmhZaIXePsV1OaAfLJmIeDYRM87McycCltPJaGAWSFYNpgko
DQckU6lLwyZ8CwsYulr6MIAa+0JEgS3XDiQlfelAnODURlsVfPczQaS/N+BzDDDR
HRJ4krflX256eRbbzte+qtpG4RnIKUUAMuv+wYzqzRk04pmPDIfiQXE+VpF0JU7L
AO7PFBtPFMiV1JUIjBHhMKw5nvxh8Ce+qOR53DLzL/fGKXY/nLMcmTQM5aFzRu5+
R31QhbfiUaLMgLm+cOm+ytMUHkl1kPICbkkcqer4O6i3wBkW24nXikAUf/HvLhkU
GcYrh2TMrN6L1sAitRQW9gQUqJxTKXlIWmIeB7VXs0RQfFoA022Z41Qerc2rzRmw
VVj6lRTQ0NldQTFKbYGXXJaXR2CqPvYw76ja8BbE+WaorA1oOhgbLz8idATofDEY
nn1isbts2r0BQc9II0jRkoZDsF9CWU28N/4fRqRI0Y2b0RXUG3Kabl+MjJkb8VGb
gja39Cp6jVdkoaDXNSI8aoe18UOi3V+SK4/crDdtvuz7dQkW2ip+VKjmhSneWXmI
E2yRbTBBQdHvvsNfvDOC8iZz3rxW64u8GFcRHzzVeUpzGhW1rfWfoq7dF97L6GKI
YpCttkzJi3MDEIs+CtCIuwQla81E5/r2JdqXbEkWQmfgUwY+AuCGIp6HvLS1sCIW
COHlee2k/qjQH2qdlg1Nbfz9GjlgI+rbRHiKa0ZmKvHWfhw18x22nZVDGN/DF3pn
eJI1j+SJpdS3v6+/Z5aUyLSgAxzNGxH3UgSb+oFS0OpSj4kzd8rvo4ad1wEP3Id4
Nt8phX3lY8qB+B13/4PFi+RTq175avLPRCAbZfoMAXMojnN1u3zNN2o9BLYN32mM
A0Yx7fqfM91BTkMGrVuPuzlzceIPjwxNR5dctWCrAvbG7Tcu6ytLC66vIftIamgK
90m9RHYEklru2iSAAEsMnUef7jtDTCWMqx9zAvsV7jlLoFdfvKITy2HqKBlQl6hg
6hOC4g2blxXE896nyCHA9ZB6IQ4KRCDKJMOeEuXDFyF8Ke0agzsGYvPir6UY7R+H
Do4si4aWNElyAsPRN0kfNZ85nNxLuVphug64B5u2Ar0bpUj8qHgjkRS9dJm2AyDB
evEOvNihGYfexTBExftwmyR2QqsgejPlRH0hW7G6KfwueoV2SIxJbvKLzKZhiYyd
H8iOwxZdCYHdSvdRVyaX0Pm2nVFgPNkbpNZfSjXwCEHSx8vYDLECWW2vXDzULXjU
XiLYP3KMKc86DkOqBYedfAbTrRS+LDNLkQqfMz/NrGazw1zEFAyoX68gVbMzORB/
JSK7yMcuoUGXHaHw72rXSDZAVrG80ikZroVuAJWzanMU2nne6FLW1lB2T67W9rdM
Ztgp803lUn22LgeOFT+JwqlRAqzzaIVqRzAb544H0KrmC4ZE3/RU0K14r8GBXyAx
H2kQYe39wsDgEHcG0TFJXchy0La3fipPwI5EJyZWFikwq4vzXVEDPydPdvW4SwnV
P4VcFnQtu5TMCwF8F3Dsg8nlKrSsskVbrCfDnUmuJXvXXgA1lDQNJPsi7uYZNIVu
6vQRNWA1qImtHtbg3hxE4XHGGQsikBP1imKeCatyemWMEhSHfKL2UNUU6WqV3x1K
EVZufcZAW3hpzBRMbO7Py75yP+SkY2yZO3el9ex2UMkQPIG0vg+rnlHdToLelADB
55Nbvn/1/AzCwahWsBMYXdswD0Ata9kqjen+NpUP/olnyoCCsfkbytWMnsMgAz88
OOChRI9ymOAtNq4IA6YFUlxad1NT5NYiYRl170GaQK5oKNH/OZ2sBgGtQ+YyUjKs
bTGiE1PA2NPSJ9fkCjF1TlKtYdz0vEz7bqgz3AJl9Ob26hIPBCf2NODnaBbg0qiP
MaeCMhqNyLJ6zfMSgboU2p0E5jd05y/ZXnrLyhD0nn8/0hzF04ZRX7E5hU/eCJWa
1D4GOthF3Dp742Ij06MXuN2kTBHueDLx8H1adLpCW1so/WVe5eF7cAS9DOdjOpD5
NmEDfz5EeYEVPcbNW1B8eAlIcJMm76UpDCcgrOYrCpOSfHb8MGXGY0jthWUk9N/f
PBur73x+5fW/2JnzFof8U4vzvGOpRmzOJ6s/M//76QIqlCxo+UHDBgFhWkjqsRiU
uhhUdhCzpwYPDSpuuBZ210dBLa9cbb11PvW0clwi0N0nuhlf2lxKl9DfUeaJVVx+
cr7sCfae94QtabLZ/bo5Dvnp/avqErRbq1lAPlBV7OXbHw8xfxt5W/w5NOQoeA5g
a2pB9WzvQetrUTZnay6y8/macK7RqiSC5KpvJRjsJZRjGCZModYeBjtpcFOS71En
2H3uhCbDRU44nquZAMNJr2zQJ105QuN35KPUouIEC4IYoSdXfxVS8IrwiOvVFixp
XvdPx0BaQnc+kiubeKAtkSg1uuD2ObOtUmz0vGuggyPnXcUA82Q2NUdXbTm6jCwJ
hUUu9Bmf12JGLsAlkFNLzg9vELUjmBf5ZwKIYF09lKKdrkdJ8XS38XKQce73pcwS
seUGifUUpY/uUjyzLzFLSYAQ7p2YyxoW5R41imMQYbK6d6CjXFPB9aqhSrenzjr+
czS2aGt4gVre8LLPf6VDplEpkNIEAfSWeKLue8seCMuLJoXlAezck/EyBBFa5SSh
ciPiKUAlKTU8TeerNNDlEHuGmAhy99npCm676KmfQJhIREUwyxdMuRLyYM+4l92m
GnTi3hZXMdS4ni0VtoDCU6MPHduMxLsjZBZ2R3WZLwckCy0LZCJ3AvDNlQKifNfj
JFC5dbedNvXh7Sq1Yxt+TDWr2J4kALL/ifVqmyUfcdSAZl9XQC8jpQCfsNLTJUws
J7bBfVS4cO/KG7Lz6Q642BvLDTV5S0KoaON4TWi2Kzq83WgSy9gdklkiBdAG7aZ9
yBF5znT0XftDdRgXkaT5mVNXzGK7eaSRQTVtXtYFiW99+K2PPrOteI2kvzP9d35G
JkTOpDnFZMlzSOAcpRKw8Rznn63KcYbyCmzDTB/4l6Q3qSGPliUL500+5XZNUYAK
Zi6meE01FQK6qGjeLfDICWypR5TaJ8FIjrPeeA/xnkDU4RTR8abXoXfQtUgPQNup
rkEUoMx/6C5LKNhC2aAugr0sSy7iWMXyk2NWMsWdW7XHWp/xE2Kz1BC3pUU8j7tt
UOJfcG9fKG0ZvXd2/S9y51m4asoiakHOlHj47cRSNwzA57Dp2qHlpDNxIe9SkI5y
yovwLQUPeRleH9N12Fmu7ZLlG5ttSleQd2DEHr8Ebli+7eSDTmlJrSe4BYIzk+wC
wGZ6H2tENXnK9GtizpaFDfpAUn5nRmwv/M+Wk4+5ogZ+0WpS1yqboQkEKFtQ0jcZ
8Uoi5ig+fju0pzxZJ3AaNCwBQ4JyFRq58YtaZOwssLRr/7jC8jga1b6L+n18Poqd
EldC+MhpvZn3ZmdCsLhk7WA4oXEM5c7CrH2ItLJM9Blk5L+B1qdfGeuJFl8PanAw
F/XXnrW/VW3qaQTYJHhV32i+bEuX2qcvGaCDMMY+Ig+wkyjj10itd4v8t8nwSu9R
5I+QBbFnNMJytnXwq2/Yd9DDD497QTxbtZT6n7inThImh/Twa8DZ4vNRxi5Gd38W
FxXMa2vuB1+Qa/bbeq2Cr5naRTCNhXQOEgj8FfGSTL5Mgv0F0D2aD8jxfQR93iG9
rhv3eHdGYKatDKAZWru5amw1VxVOOIUDJmbTw59MMPBUoPF0ZXZez1xQ5wi88cpN
Kil2f7WgoAUKdisCWz8ibjtwNKkLpUofdpdAbc1FvTld3rIf0KyzymQtGwWePpUQ
4H4aMJD1qurJ71MoSwzLUc2ptK4QCgnW0eCJcwxCNPUuNKQYk1R4g1on+q7mHBTZ
OSghBi1+ZYlvhnfopCdSHC40BtGa45lS6Qkz0jrBwE74Klj3Zto2foMUPvEWEFwk
a3aQJkclv5T1LOrRjy3GrAT3qx0OPPnD+iONiSHChUvDsxwXGYjW/W8Lno6KVYJp
HxwfK0xwBL7oo/di0cExQO7717zP3DE9DajVPMwkBgR0hNiVSUxy/L1g9jSG/KqR
GBxtDtr47IDwJxmfgS1FLQDpllycIit4AhM7Nl6TXzjJcMSy061ODRwd42MiNXFl
w6X8oXFCua4Q09EUavl6leA9P2X+Vd657a+upJHi+5T5fSrnOsk7VYkwloLeagRz
c/Vj19h22879V9jR7ShUFmQ51QZ8/kW7/5vpeUTJiA7au3wFOE+1HZZLFRaTyy6o
z2UUfC9KiBHw6xFD495ILvdtZ1qDRuTZUgttuIm6XAxpucvm2lwgmMTMJu0aKZGX
odt27ZWReYmist71oxbj0aA+/28QsV/gxzKv9UJsKSZ1VZJrblY5EScAyNYt2DFQ
rj8+Dk+ShXI7jBx7v64XQYRCFfOlJKIK1sZX8UtFZ5pDgERWaofgpmvWYI1U72c/
7Xfh36EgF/6BPIz0nSl8L09fcjUolVAQPUKpOawJDIw2gbcq41Q6FrJNtpet2bZH
zR9KO1bPI4w22Bahfdb1Nru2gmlMof5Fj/bbTzo42+e2+IaFiixl3iAt3int1Kcr
qrScmLpB6H9tEbv/V6zakx3rbyLj0EcALBNL1pCrxBoOH16UtHaYFRfVxDxZu+X5
zJ4qK97a5839/mg+Lpc8Z5mGZC3iQFqW/jdxe0+YN8norg+lqX+PXIrqtDEiNjZ4
W54Me/2gybnmJBuHosv5R1qmDhRkP6i5YMEQBT624xSzXGTXmOS9xYqepvefY++x
pOFwU36QTSHqa6Dq5UblhFC82yHTZIQZ2sLUz6/LiLlprX7mRf31xjvrkqSOQcn0
hdzzWdbT8iPeLPxzZw51A9mEpwm3DhfaXK6CF4xdAtPH39AtmVbX+1U4/4vfPWAj
Dboor0dwnUT8F48vUWQNT1Nkk7dXJIPYd5/VLKU0xwkybzgLWENSaRjYrLBjy+QZ
guh5tzpI4GScRdwxJh1CVYZSv6gjZps4O9giQA8z3vtzGth+ea+jCQTG0k+XM8hU
vKM+/jzQVtDE4C1kVtvXgrJIszEOxFfcIbrYtrd53kbpqxU2Y16s/uzJ6xKC/Soz
oC03/CZnN3odT6lI5Ro6OVNP6cEYSQl/acyPCDUjZLxnrY0I1QzKpQBhhaAIMJ/b
YiQzzxFwM9HhWGPhzQYprXTirRzWsjCryBFo6X0+/j9Wheo++EDx8pmYkfis+SA3
XXkUbho8gnQMVXM++ObERXxLNwAKD3ED3M+dJaHAuF6qc9IpHjHAPabw4RLMVKB1
HeVDn2rSUgDFVdbis94D3VqzRRV2IqjC/wbILgyN6AEDPJfYRkhYg/q+PTZaLiEu
nyw1jxbgMROOiezGMitBnLDjP0TGYBo0KxK9ZgD7+rq9X5dh9DSYkrD1Z/OleKAP
so42VWLopqjMj3sfkmwtY8Tb2cNGXmV06TLQfXGBxL6OAs46hrokAJn1pP1YcD+C
0S/09+MVsUkG98yBKIAODHmrotCAsryJT3yluYYvLyAXwdklYdUKcwfAMJpyTn8F
4h1wnHisNauAWP3Xjo5JgwdjvOBEcnxiN88XX0Hzkbamvt8onNzMyLHQ/d6EDY+C
iDbMh896ZhPWyjFcFtD/+cGGQ2vamsS1h2RCt2CGrsQvtkxawqTLER0nJ/bjB2hs
4UtBuSz6+zWO3h51yFtRR/ouNSAVVWLay8iJGmaWLeLAlzkupqZRDqZXFOUnFXvP
YhddP4a9dnzhGOaLlya9qhE9cdg/Q9iWFCWQR46tG3uAd4bq7jiK1AySdScBUql5
+Ytkdb5ASqW1NxiSLMm4MaqNftQBSlZL7mj4hj+2QeqKcZNX9SJoTX4Zeru5v0zr
d3gmszKONIERL2Gt/vxT0lwlZ8e+7goYbJgF8Ya4Lqrmy2BLLZVZ6VWvXqCxkBcS
pKWdB6BE8cBz8ni+h+HKdatiWdvVsXjxl6v6WYagC/nJRlyditx6c2AQyL1BCyjU
m1EBnmQTb3rIXt1moqL2v14bg+9nHedT1vn/IYyiRsGGN0OpkX/SoMihReznqVVR
FOfU5ml7yf7Qf0LxHmHnsYtZAAuRC0FQDjNDtn73k9TEjaS7Vj90BLSBdvrCP3qB
E2+bHfz75V7Ga/3xYu+ZPGeTXRroKeRTISNkiW737x0nBbDtdWyj9v+ZykwZttn7
pPv9+29J7lHMMD21Kxk2hiPWhVD8QLY+FP9cvb8f8wtkNvDMZiEJ8Em9+/3rjngX
nF6JIrn8WLjckefAUttQYgjR6peQHqe9pyOsWLgR/4y5IxYz4e9yDgAzZ5BHwz8P
YAgGuLTwSqp7+C2Uk2bTdmX63h00prg7ttsS9HjOhU/gjEMsv4xeWiElX4eHgwVo
bKcR52sQtxwRlZrf5t0KNsSb/k2iNVzceYrK1XrTFe+wMmVp7SPtv2vkIVMsh24i
G8rzQbh5ePXOECLh1K0zNnYf2/fena5MFVx2/xrl0v13qYEzgFsD1pQaSUem7m8N
dguI+hZf4QbzuRFAbqTT9xF4OgMSWSW1XtxMFkR9PIG9SzvVOyLZpiuMoWGjXfvd
f+qQ4lA6bNQeKX9f0dGgY6JX/F3CM/11FnN3ybUvYrm7QcE5pctN4rI3HSWtzthJ
63CS/EBjQoNMHhGx5GerA8OZjiIvXTXe0mJeKMD06xkk+afXFt/mF/65hX2rMUeO
6h/CRg7FuSeXNozKcS5P4fPQgLXlXXV5lNsmL1jciAbLiEuELpBESW18xYnWrdiU
F2xYNupggKDvUYNDigT1imF/sli2OS7/gIBmfFrKPblP2Cgnh+UurRb25pBznuGF
w2UxZBOcluwouEitDvppTp/GgfABL9j/jMLvcIrhm88j3KN9AZo16ZxlU6IgiLCw
Z5FAw+EPhPdB7eG6bqQRm0vCa9ZCL5yqpk5oHpVlX96pUnHfZqpwmuPOlBhJKMCK
YOf+SGPj33LT+9kWf0l+FwCaXJ43ABdbEYtGqX0mlE3QyVYRJ4wjFJu27dvjEggt
nsQhaF7WuteaHuooVo87uVTqkxa7UDhmQq7LDRCEOqjZWt65yMYiSvZFa/994KRv
GdtTN4Hpt00nowVmDZuof9oGOALi+WdpzLsGmSFZHJgC1SQFDch8AeAaBSuWOuT2
l6nunGtxtaQFXIDrouH95rMNJPePTLDQpZ7Cqm6yti7267jytip1YreA8O6jhRHD
rckPUHBXfP1kJBh5kMnNORuqSrGlmuwkGeeaoITx4uvykhzMummhJlKvYwCrKkdq
tB26JsOG521ijdm+T+HvHaVVC9p+hl+ONsNRGsUjf6ULpmmH0AEzdvSmqVvPyQ2C
Hyqbk0RumyLsRegjjbu2Ma9OIzWjEuyFK+LNOv5p+ujR851oQ622ctUGvBEa3Bve
JRGJ70yKkspXTOBMXoBa506a3d7yVgeYaAqegZ7xdgysM3rBDFiSQpI5AWpxI7cA
dl1CLHv7VJmvYI05Uln0hGlHgmxTr9YQBMsaN3NfOJXY9ami3c2F6WfDuebo3wSR
mEPWqUAvkY+zx7W8cFJUfXrvLXgNH9KzChBjgA0UkOlCTjzSz4LqF+UCfq01ywL7
zGIpYL9y2y6oRoY0k/rmva54/3vsS1K0fo/VgoP/Jt6ZFVum1XlLsX27YVn61NAk
4bm6P2/MCDbCk1zP1lHl3RbPSS8MazVgaFHaLYqeGWrQ9wWo7yKqh5ENCCOid1dd
U8lbKa6H+AaB7RNaPp5AFn0U2yw+yr/EbyyW2rru7bAYy/sGVQFrHgqfdNQQIZp0
spsIo7RoI6LhpZMaUadgv/yXPSRlmefTj9sSaSqr21k0aR9A4GoM2beCun0nctLY
nMd+r+YIeOsAdAzjpBSrZar87avhlaNheZhn13SVyI7dGKh/Pmue/IbX9pGsjhdP
WWNJhAkYGK34RzLpX+W1EwrrDkKH69QcDyHsAzw0ZFUA4saLmlk3IHJX6tMc39vu
vfLQ2NQHmIzt0pBQeJlpi8paQIsaLsxlSPfDgQOM/5jMn29JKQ8WUqebyA4U27Nd
itcEW70801fk0e0HQ0iYeoW0UgC7/sJRh8oo0xhtIm6LSRdtMBITXC8oXfQXEUyk
8NeGU9QjiCCDqqBQQkS3BgJHlRUVilCuCp4/XCsAA9b7Z9aumRa2ZVOTmPqps20b
YvZ82DmnmZ2tZBkgbcsNWiF8WpqAi2Bbjc1WlSPu7LQQ6GHlozuAcan559Byr99a
yzZ+yc9cuATZNtv5pQQoNDu9uACQ7VU4/Nxe9Cl4LxggeC2NiVK/NuMn+ofnubGS
2xOibbAAxZpfZR8nwVv7WoPytaRYHXHqvQjiCYLvMghlq0Y/Zvyh4uj6luyhYTxW
RBfD/WCWgeb35rb0fLIU1KNm4U9YynIErLbrRPlFnw68/vCrYvfPNyDq04ZQp9Kp
c65heCfB7YzEEvTAj7tM90jlRYSKC4k/YWe/l3lzy1DrMIbLZG5je7AzQunjdFi2
hhiqAgf+WXiqZgjb8Glw+wK3Rhyykcq0iIektLN2FC+5NPwoTD6cnr0E2yMQ5qBA
lmCVgn5O78KOPzZHZUz7bf3vqgnPn003VSbFZ1HHwTEuNSQHzSe5hW/35nD3HS8/
viEbUa9qvVUy7+NqWHZv64yIKL9FY3WNzSSlVFGLuY2glG278G1wixdBRBm2hdXJ
ZOkVkB+ft7PPIOkAVnwUDsy15zApA/S9QC5kEGzTuw8Zfd/KIag24OM/PIFSKAXq
A7ClS7pGLY0HEKpRAPTg+vL+zUrS7b/G3Prtwd8nqSZL9uCg8tstvi7bCrKqohLf
N+cz37Di1qtMzQ1+UeN8wyugcekkKjo+5tAc/IZsj1rYuLTYQjJtinm47fO+gicS
rkQ3FxXw2u0e/HhPq22bXc5a8pX/3yjiq/4+P826jo3HOOwYb0Bhndo7pgkQxYeE
W82hmF65piDR21XKRB9g3SS9Ui9GWFgydxMth5jA1itYPQ/e8nBenw+kj+UB0mY4
cCJJISQX8ZnO0Pj431a8i6HRhcNSFqtmgf7DaOsqMponQ0sDUcdy2/r8GD8JO1/r
7zG1InmEo5fY+iRMl1U3ut/jOIFRl4kR8iRvFDcBnh8mPWhn3AH4YQkXR9XQxMyY
yhoWU4alz1iP1cffuwdrfS7rEwXBXtxbHp1FmoOU9MXjucFQGnxu2lLW477bMaKX
vuft7jII7xQr2KvCQ1JtohQaq9tktT0wM3u5SkZve9JTRscSF98XW3zBbfKt3FcK
8K/VUxGXMRmSCYVsf+Aurai1OAnPP1OIwhsbsJ37HFutepyszuFEBQBr5j5D8IAA
YtvHdYYmdiUIzoUVXLr0x2J5J8lIx6Zvyp2QjuLy0tnHVG4gTeDvy+7+QScwfRl5
VnDZM8XUZbMCeKcsRJ23bbKXh+lnk9nRWPcEy6dEIOllUyhLFMFXcgdc/SpkCQH8
8TjErS8LO60SQHmGsKe8oCUtjryn6mp9ejpe6g4GNDaCgoi9K7AY+Sntfcz5Wo2i
KshIvH9ZpYVKunFePfS3qEOe0YkTXLZOHbLP2Ps6dEhcS9RYWvlFKXTY/+CmLVyg
xU27qYCIePGa0evR1UEUndl8Bph+MA/E3O2I1n3SZh8kG9PhxkazeFvFwIJ3gH9N
V1c+vlbOCCCgFPV6xCBRlfsQYjChr4oFbkElVYEG0NYiV1h4oN10iKb7+wTsvi53
BmiH986MD9uwok3aJ6JN5YxFZv0KRfmmJ+yqshIQjEYbgiRepPJ9UCgwivPblAcZ
Rnoq3+iL+iXCFOJRnYuXPAWrjX3z3AubZRB1KK20Jnyml3BWp41e8li633J5S53/
1bc870Wb8s87heaTRsCF2vZX6cNL0BgorIlyIJB9lWJq6s84C3fqrwS+dmLX7b5X
DzlQNniZgc9sn1HdHZk34111+s0cts7kmYZjaoWPkmaDOsvl/Rx+jf5eDWVNo7Ch
P4rtTE/DCNam9oLeK7l7m3nhYcUoKak1f0t0HsLVrrx3DUk7xKdbpAqQaV6YEITb
zd1NkRO1MZC60jwSD08A8LGxZGf1XDNPThBxO1WNIwODoQbFoKEEK9XyvJatMRQc
+bxcUMgxBYqi9KzswZHxt/vuk+NpqGth5mkgt/MZ2KurpsmObtdZNSJYyB6nTMZs
PfzpKtsnUwKH0wxBdZ4V1HjQAyNgYtULDHS2uWUNu3khcEV53UjNlTAMfof4cUXE
tzowqTyBqS40qP7rsPvXlOzh4Dy08vwqPru5vyxL1KrnP2ETify2rXFDlLlQam9i
aUtwHD8KOqkLqf/bMUEfugghx0VUi8ULwOczqcSCFSlHtSwOqszMt2eT2GeJpTZs
5RPUsDeK9StMXebB41ZdD7TRD7Rvfa0uUMTZQWl/ed/S1lxlYf6Jza1C9JZFhAE+
ejIJy6pCXqftUzpozcpHjyNsb1XmhIkF3uMh7ec7cNL6XG91lnXkiFaxKSrlctsP
zfq9sqQu7IE10kX4XNgMZEPxJRp5Svv8Qnkw98htLnru9IuFDBv8qs/VtzQfWbDQ
QIrcvVjEVCPqf28n+3gIZLYda8nm7ImSqH+c4Lbw/APIg9d+j9PheJFM7M2qJS4M
UMLZygK9JKMoGSRNZss/0PGxF7ss//1bVTWYTuJCLn1mPmKBx9es4roJoZNPutZJ
z2ilkZUo1I6PxRafkBYLo1088ON1Rkh7o7SYEP95yJHieUXgqBJX2Yqq3/TTwhpX
6kok8E/JvmnKK/wx1uomKi54XoXx5MWP21hjrtC2Sl0cJxH6TyVTtdzZvvTjlJF2
oj/dkeT/fxnhaATsuwT24EQ9RXHTupHs7wBGTyZqOIUEbjObkpMeW65KAjvOJraV
0KYAKZgZzfCeAaLKOm2NJbKRlZ3X42ezWDYO2ntrzOcHqVBx7gLrtYL4naicqOtm
KtWxLfqcsTslE+1xykhH1d3NR/AIeOPZDZlgiZ8WhE1UBZRLbpDRbSscTp3cy0ZU
czAV9u9ZU2Ey7VDtxtaM+bnKpAd1mu4vW5QxQWcef8YIE7RES612TaSpGsGGoWNd
bfS6NGnXgO/r8H04k3GG6Wna6OpBSV/jqX2LW0mb6TyUonUoBHpixVEtHkdYryM2
efKzDcMeHQEw2s9wWzUm9O9fLRJiXJ3G0QEkIK41rKRdIe/wuRAtH7TVBNOK5MM7
YD/YCm2k/uuk6aVr60etnXcM4+LD8tEFQbZ5JYw8V/hE6VeUSW//RI7ccxgPULcU
67hgiFUDS06R51T0lJPvV7k9vTq63J2HFZ99zsQZhEW5nMokH+DKqoXjvgzak+SM
3Ruv8lTfJEq5MU8MubWHsOlDhwAXvdxqgYkzwMCCaoqlgfaJE1T5JzNV3rGh2jt+
0aTvBTX2/TIboVZxsEClu/0I78+9mw0Zmjud3C1nRFLRRRSuR2PEljxC5b1wIWhH
s2MyWsaVbUxgokr662sHY7VDqAeqETqpZ6AoXA3y1a6gBB0oqUuH5Dag260ygQKc
bCWRKfh3cpaKR/yDq6gWrF2nyB4YEW+NIRyNUXKYEc3EqG2WnrVEWt8gWxDls3Yx
uVikg3UJRAM3qCSy4GwCK2WIBJdqk+GHh8o1PJlMFkqr9LisHv/Zrr8AufwLx3yO
nobXXlA5R2pkPJ3QXsa/o5y9bnxAjtAWr6B6JBKZVug0iSpRTI2P3GSbqSQF9+TL
RY0h3nQZGvTHuMys+PaForZUzlYs2+p5Ltrv7iyZsEJTWyGCcPsAG1c4ZJai1The
VvBDwhO8iZB5BmvOQMMd3eRiYZFo3jOGPQWBxekZ4LR8hQCWpFNZ1FV1WiUpRNLq
MKelH6Qraa9gH1/jORh39yXOU/ziQObiioXHJMgNTU2/m/JeqVxzW3gpTCEANyiW
vQV2FSwNahHhPG4FHi/avCN21b0i0aFs6fvNnKpiY/h0U7nUIRsMxIDhpelhGNTZ
d6MJ1npgX+yHz/2gwZ9qJbEdjHCSeJCUfWgiXwqNMVvoDSCcJDSnTmh6aXiV4O6x
CBPXz3X3ttcMQeAXFm3nCpkyvWunRySjOAgimSK3wc6tTxC0WKpFIK5i03ET8A2N
lcVyxg5VPOXCNGV8gPWx5zcmsesLAHYJvOjO+gNM0GaobnhyHcU6f9taKs2piKcS
nHQRCrEW4EqX32BTE4FDPI9HwHmbl+8gXjZK1BmTi+NMHmQuHT7TCYUWAb1761eZ
0OLPTz1U6n35SR7Z5u3z+vk/8GUt44ZwiekJBHFw7mIIa6pmIR1x9EpG5Ef7Fvei
XeirE2XsFS9NRZ1two90nliauhOoapxCaDQBDl78Bd09X/yMEtyVr8IUrImr6mIG
hy05P0Zdqss6X7GcftJAKPR+udb1xWDPRaxd4+CjHj3oZrVp/n+APfoEbr7uzRTF
YzFDRp6NA2CEuTOQ03NprQkMQEp/T5OPp/Rw0h2oaFQsOqaS+DPuNW0xiuS7Wvm7
na+X9EdseRCfWiZ/5WYqO6LgC0D9n3uftj+Vu35sObYScPjZXabwlkhZuKPHqflz
mQanpTZkNNK81UVE73QdBNgULgxIvAToHkSgogFEDf8zs+zZRut3VAmKAhFcv6VH
6o5Y+9I0r0AMbo2x2aPrIds5lXOLHPaVBp9Vh4W4sjoLqVPwYoLkInx+yBwZlTYf
ItpHkZxXT7J2pXKJl5xt5xmKQJUYn7Yzablzz9rIKcq9ZVojo4OTbSggvokoYRPO
yh1eOrm4kV7vX2xYqydnzAiB/iP6J2mGd14VkTBqyDk/ORk9191L10clj02mMUcA
KHlapOY/AAf5W1k8Lwql8A5gaMR05DBlS408ZsM4bxLhniunhIYLxEWS4kOLJ5x9
yx7pHX4Ts9+sj2C+Y9dgMQDnHAAW9dhvFr77eqAzc2hGcunqjBNfqpNwb+WLJOP3
MQMKVUItyPJ3b2qHzUxNp9P6ublEZfq5ucWW/xD8rpLMzatVLY7MGmQeDpf2aIZ/
eWumxUB+qnKlgEcl4B0W/GC6MSshUNpwIAuoPlpbEWyBsUl6a9KYz+PXQlIJOUZ3
Dvw6go/kCfVE/NUBiC1Y2soFic0FvTbS9kGn63KwmvZaHvgPIwoJCdFO58XYX8Ws
VlENy3oE/USaQOKs8f1IDYZNBEAXCyvflj9Ra7MQR3JM7wvsaBQBeEV5ovexFvtF
CbDtSCFVj26/XEUNt7xszk12N+uRODI3628H0G9ZUbx8ne/hsvTHWAXaNCk4D4np
Nw0VuTGC3tTAaADRwECmq+4yyTs7bs/sgzU7i6RgcTtUV/DleZ7ModeOsjkw8/GW
yYy8YdyU0/x5/+02uwgQY/16XlOKwZLNtv9hI9qln76mfbQxo239hk6JiISYtNx6
b06XD6ShlEEKvOmkjSv0DFevDo58Wub7/9hgR8aiKZTQw0SfHzcILZPH6rMcwrpU
bpNkCrL3pA6E2sJKuPGyG9OHzYAb3jiuE9Lb8+F/1PWLBlraz+G0H70sjJ6fbktE
HhOQxBFiVetEeI25BWVwo+HHOuDE2kMmrD4rwXZZ/gwfL6Y7U2JZBOKedlh0y/vE
REOQ4Dy5GXyKhOWaH/sU89iCalCDE9ghy2JbufVXV5wLRB5/OOdcLXHQ5Bo/FXVA
ttprEyVavLxJY/t7r+NIXV603gQGf5MHl4hu5T7JEsSOQmcJn3DGT7T+THutD4yh
kv1+MspPVltdOlsN4AxB7u95XurB9oizLDn59p/2IeJlPJuCu/SbZTXVIY4Vl1cA
R1h62Zu0kFKLVA1QHIh4mHm+LKN/jt+Hwe3uEJlkSRYyRoqLoHJtkX0Sr1hd7ppK
BVzirLbS6PyB9cNx6JKep3lrIKNi+kqElH4nAI1VnG2gEJp45yGOum/2juLN8mge
DQ/iBVixLd1D2shssDAyrxXLND0o4VabC8n0pJnr1irb+MlwGoei6uLaFN9+QbJs
ymg8l9T/mVwvV/Qfe/vfBA0J1+MaWEh8eFN6dDTUhw58uUICfup9IG2TvxFHe8Oj
/7jdyjzf8pHn9alFzx/Mc5lUhWbPvfl251LJhE5/4WeBXMmk5JfE915DmP391Drp
A/DZdoNnKhbo5b8LkgAmj8bTlpx7GI57TYrL/f3hFQF6QaHy6mrCxB+Vj9bQVRn+
YuTMwiE9AYhlNe7pLl9oROtkuUtuNtHf4m04mbog/VwKzeF9MFDN1kWfI2SDZd9I
zbQk/7DqF21wC19lErnvNcZmLxfS5fm1Ka6AkdFQXBacN2W2nA8D82aEbyAsOw7N
ZCCR9+Vu7aXcIptyk0+YZRJtwxrTKYD9jLF61Hrc+8CyRobW9R2HKn2Ybo1OY6UO
J2hzo4i4wp0B1swMnohiaa10ksHwzKXyRSKOPp7Eu8r9okTRr3tRBDXnf5gz8EXn
2dRePhxmYK6GrL3nxl/on0ptObWQd/8ci9Z3fuwQxg485KfkQMaxuJiJClCkZ92x
EEImMipq5iUyzXe3RL4FWLYbD2LQdoOoYom26oXpySB4+rV8aTVzMoe6N3gN/fpD
bk8TDKAGcQMy3bljwD18ucwlW//rMScNAGlnpUSY6XUw4hAXYBafRTalDloRo7Hd
vm4UBImLDLjTxkGzg0ufw/4k/KKLzLRso6Ex6D0LEuk8OLcbET+gfGLSHir3/ais
GPf7XlGMnpkt7NvANV00X4EXBNIY6sOQCuyDchjI2kqolgMsWfkUPt2WQjex8Lrm
z4C+6JNCyHjU07qABqCBiMDUPvrIkFs9kYJDvnmPDiW4cvcAXUt2a3a/3cXjcnA8
g+7vpQ0jCHtb3mjFdKet7GZtze+i/+nuhtytCA0oQMc7cSDsOm81Nxp7O8pCKgT2
qBLsYQnqscbtZhQ92xCCrCTdf8hhpAe8pGS/MYonU6Jfo2SgJf152b55TKuwL1V7
t5VWyyx8EEJ7eD6ZrEFviJbRU3gokZ9hKmeNtruxGXYiq7sbFAqPMUWXrDNbQQOI
HhejnzTwRHqFNf86Kj48fgdDpCGRdFA4NziwYArwpbOOV4zF1uHRJSAJSQk+MO4L
ANksAiA73nKbN7+F6e7z6eMyU1cw9mhu8ELH+Vw/HEXx846Hb7HiBB3KOXdemmni
YzvnjdK9MzDYWUNTybI4UmbgAPlnE31QJnx1+NZ7RGbpEecwFzUS5oL4MNWRGEO7
PCdFE/+9Fiej5R/7NO76A7IbBpqHcnjiTZ8wa+pJK71s2TSWzp1hdZ6riYJTvBE6
CVcyHzvV/sMLev1m2wvZMe+rAtQq7WhpaN6WL8cb4H6sxZcAHb1qIIjWgIgS+fWA
cbUAIwkD8BlEBLEEHk/p+JnrqlFNBDyUeQYWLND58Pn4FlfnnnHZuKVhXwGpmyJq
NYQ2tDqEqUb9ovhj3Ui8DF9QQur142tNCTnmiNwnqVslxjkUCO0Nt6UVfkFcY9RT
m08I+5vNofXd35geAVi8WAeC+NRK6lqg6cJFHr7e0E4bU7b5btU/kMmcvAJKbAor
QWT6C458dArTQUzqs0on4jZ2Zn+eYiAv/cfCZPzt3AbHQEh3z9uThCrPeGlMadbq
s2Dh7BSkefRof8NEn7XNhB9W+ENSB1QMIskzPpdKPblwbbI4unnhEUmPF7I0FSqw
gA6NTp41zkq1RvWk5jm7cmxLgyfQpP6NMgYS/zDlfmJX7xtRTVzfVJ8njT8qHa04
0sFGweJEbDhQNaPZctJe9sRruQ1dbTLNuhIcaYZ8a/QMzVwt81wHLfF+JMBiG/Lg
PAiBOC1f624Rajr7X83PI16h68mHSQCdO57RISFJkiVCG/Absx6xbDJGvXQV0+ci
7MXMMe0JT1BVDXkyISLu7pQ2APWfoPHNu4TfuUyCwmUHg6KEeS4hZXZYTSbb6o/S
5I24ZdVO8WTtmQ7gGAioVimXLy5gRQ3FInAIdE2I45/U2CiuUweLblD1C2kiMAjH
/BleFh6SxjPP7q0Ll7amwQekZuKAt2K2N+ontL7gRc70spIBqvSa+nVxYx8178vU
095GeglGW9zEhQ6H8JjrrTL/GS0wiPhkM1kYOY6AbmSHAJBYUI73gUnbYw2w1sjc
E8TS3N3CaNd7BnvqKhXpGGkO6aSUqBbXiUxUtgfJEgo4qQ7N9nHcJ3fkAMQenmn2
JBgIC737qSoMlpNtmFqaAmtbWwBR4Cb8r1DtCi/78ue2ghIiR/Dz+A+ouAYED9Cd
K81uMPKL74kBiwQe0OMJqczK1WzH7SGQfi8sQ1ZMumPUTFhBvap8EPUVJfNX00Rf
Hksp9BjtVu3aVOm1Mtb309erDIyDaEwaP135tzUNqsrcUSC1TMErq14W9/DzpTDO
sgu1TJzSTTzhqYgICTgayw2XmZLDC1Blx70joMG3twU+nrUBbttNM6yStybRHcDh
Xz367GSV4gPACBSx70sVR0eYae6SoUISbOXBUOSGe4PM/PjTBkryqu5E9Hs0Dyu9
mIOqRqltEmh2qvPDBvzPaPVVm9TT1eZnhRtVys1k9ZIBe8HXNrSZbo7QHfCRqGaw
JIjtKa/9/3BYxNR0jU38uzTW8bxWG1Uek7eI2CQNex+nwDbtmLJ9MTCTtGI9g29h
9Wpne4NU4FFJaJHttE5prg1vJ8sVRZeJJibGb8atMxFqmpkfNYTGCoEB0Jfll5EX
bjK3u9jHEjawVsdQppiCpnltmv54UKS8vQLM3RSGwLXCSaPJU4wxw1+iCdo7TPfy
2r0ARyVROp2yf+9TOqW6mK4sO9tEl7CvaXIOIgWdSuyumk/bA+hDABOV+eIox3Ym
DnQ5gpEB5eQ4iLWocdN+wuEMSd8JTBrmLdhzpJ5KWjmxFon8aZKj8Rwrao1IkrJ5
FxPREakelAAsIoMIdZFf2fyvO45rAJMg0nBtsCKxKDKw7tNfMZehPF6P23GjWTNV
HEbSQ20DNjJKC9kTxwin8JoVTHDf2oH9U5Z50LhsDDB9Uab9L0zWZTfybkaghyeM
S/uL3PylsWc1Vhw1ultoowy/IBLB1ZH9XQAtg66E7r3SnaI90oaSVpa83fKOMoF2
DSlLXtudXfqTQVT4nxqZkuAUuAPdjdrp55OnEHFXGOu+u2/6wRxENljzn64NDljI
kjPCzW6+BkXMdiiX7ZYg36NYRnsUvvSiOiozXJS5jNGtc13mcxffxBVWd5xjHRS1
vMSfcIUdT66WmdQ295vbnSfTf0bCcdDTlUaUdw8y9by21J/xIyvPGvoUy/fCLvxw
rdJNE80ZM7lkjBmB5mGKaCk/TmQDDESrsbR1m1a3rzeG9MBxrKL5GAFGibn4Lrb4
nBhZ7dXU6E/yJhubVNNfrFWhc7nI1znWXj9+P8bkXrSj90CGdooerN1PrIIHGjI7
Ohd4ohFc2bpYErdXWKzrkAKT6QoIw4TbPpBFFxAiHqs+MnaNICj+Cvyp44AVoCNY
PnSGqIW0lG8vco+ZgtZsYtfijrd543gQuYg5WDvfzP9dV/EvxV+hd3SwovTRO3Tz
cESSvGl2ao+kW+OwemZh3A==

`pragma protect end_protected
