// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
RYxp4aWEHlFG6cTvDWb6arKtUfkzS5nD4x+ISKjALjsLmFQHAzxSW8PAU99rtFs1
p/TCSB6GLbCXFwIxVyxBXXrxSnCzBxIYrvH4U8VCKGF1+pUbyICQenkitFuQ3pua
yK3fd+1NFZG/4gzyhAO6rp1pJOoIZTFFshX6iMSjA5U=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 13664 )
`pragma protect data_block
9UMQNwvqkHjIsU8gDEa1El6dOgubvMPlzJRp6T+A+IXdiAsbAXk878+5JAirBZPf
9p8Pv5AP1pzlmZn014BTOFHUEY6pMX2aCpbwF90Fe5kK1atGI+LY4qznhb0Ituu0
zj1siccOx+L8nL2aOiWF2cWWj7zA6PnqlLc5YbwzxvQ2SvFo7ceN3DCZALvTQ4n/
2ZxYS8xco2l3htNXlqtSWoY6jnqkGAVRhfdV81PLlHt6Eg8AaUHvJEPQPOMy0f1W
lkyF+MAnB8QsyIsow3+UBjlZQK8M5Y9eN+9iOyjTw5o5cOpi8MbWSYr/Smt8sbh2
bygQP40sdOqO/XkgMO1nTPs+qy+GVkEr0uTwTqcisbazvQEgrhtkSXQQBIICX48l
DCLQx5H6OPzegBWUFC8jyFaS4SN+8c00ZQQCokPJHeAQTs0A8l4lHMX0qupOhJWW
SYCFhTIWKfQaAizC2Mi7IIIygaju70j8XLhSjHFBBfrXLSlUT5q2l3+huSxd3H6M
mXW3wWfNxEqAGYYtFNj4lvhbeReGii4V5vbYlrSfeKSEIuF1RBSpjCkSHQSvsare
wOh6F11PApAWKghAUYnuUSH2P2TCRFhRtzqYTgkCpSQ2fea5KVL2PSs/+GEanuKs
A+VhVaspHQub7xGbxFIgdiKm9zncG4JDQxp1CG3ffgHqYoLA5dW8WGIe55kJqynk
9lQ5t8n4QEtqWBsI+hzN2UmA4KqmjW1ppFD01fcsVqt0eW2s6f9hJg2o8Hf+ZNXS
o+TEDsIW1eTIulAmTm7PivhLHv1QZeIBAd1vufCLM8Plb1dyDn8kFNB1ApDG6NO3
SfWKkD2SkWHyepeOPEOcXLy/WdEDwDrpRhvrwM/9dFuvCbBZBkzioHfsVpyGKVnu
n3E7o2rAXgYg7WzTHCKJuLhbTgMLP1Y0vImAnNnJtoTChRGkJ4YeKWhnAxlb9sRM
k9+Qwbl7gzllSq19atY8WmcRBSWeE7DzB/nuIOT1bAZBa/2XRF8aefJSJmFv71nV
1usqpfcAiVt9YBEMI/BcN498KRiWS9vtV1bTOOSFwZN7+bCxPUoLeL0o5vlTyuFO
k6A7OlDsNAAyA0vVe+dDrM87U6e0ZF/EqxD+9Slct1VC4TORQmH4cwNSKOdafcbf
yDcLTzMWFazGgVILz5LD2pA+XQinyAhz8bVDe4BJhaFn4zxsrCl05fJpeKKuP22F
1HMC1oBnf6WvVEpgysweUxEbCla3DDhJtpVrFkbMC4oCHuM8yFq4F/zUPslHLov8
K7ZcJUAULDR0PLmTs64l6NNq2ukIZlyAdR4m+9XJrSWz30W7vC+Fm3bvJiEVMbc0
BQ3VHSNcJ1tjPs4LdRSqTPZ+qTqf5almMLNoYygd4lIkQQCP8G1YIMad4bwglPxd
yRSgJ+H3kzfHtF0kPi0y8ZbkOptDAkX2C77LD3ALX/XEj4zKoCY3nTYsG4LOEpTE
jUVQmbtiGPBklo9I2wX7T4x6/XXJ2I54GsrQdtbSk2yljdxnasiPDGrPvF9nvrv8
4s3esoE2ijdJC2dChzLbDEHnE/L7xw0mv73FZQwCIq2bj5L+KRR1JXGfuCMe7aB5
sNSdvFFPeDGxuKd20pd0ccm4BatAeZaUnc/1PLz+LPaEN8nKHtwLPjW91Euib9rl
MizbnSyVBu4QhT1RTnbm9RKaMhndP6ljLAcZXCuasW3KHQBkj3awMWr8AkfcRmFI
+Bu/T2bnjV4ytjBMzUs98gb+kp0kxnT5GBtAPDZ+RaBNU3L6GFPkqbtopvcf82hA
CaVUyKkpUvIz6TmGuFO3K4H015UFIMejKKwzpIDIAWsm3TOSjPtTBKiet/U9J5Nz
Ut6FVdCCFNLe4d2QHia7pCKUgphk1G4oSZLDjeTxDg8JPNCw53FE28dJx08zhq2N
yHPxhzhCAQBhxUnUdY1veHE2rkE209oNNWIh156X7RAtyDLCvSD2G7VJentwYQ91
l4EsXZTawxvq6gsWCfM7TktXcbSRuAlr4v0AbYIjlBMDtcna8UmYSLhUV2cjopyv
rwYnEhkYK+xFUZVa640/BRT8fZ61hb6bYN07XHKP2mhEpAD2msb4DLpNa+uDpKhO
RTXshvootDO+wYwICEXk2lJHhc7hjZq69JQy2Ps/V0R42W4DwclYi1671/PmyHhF
1s5PB1UqF8z4+rZXZ6SqJkLFYvRhsXr2gZ8MFCjIpz8pAQBdB2x7RScSNJsPrmfi
BDAC9CwHcxZFTBLD3CDz7OyXUi3LBgE6Plm71XImZwbFFaYm6jRKqmlFMCyRrQYf
kMBnvX3DMLZK48BuTc4VAVpw+mf2vtKrGis7U+8MW/hkDs1wvw2ZV8PZs5CFo1Zj
3U75sFHqQkgednuxFtllhmQsU2C8TdZouCPrO1GhDkxzGap4/W2inYN2p2UYXvW/
QM3o71qQzYuZRLNeONj6klpma4vhG2ogEg4fhnqM1j4OZBunzp3aq7jAPv/mNc95
wMZnFPbWPCcbjhIaeVceHAdslw2QORqdOK16XHpjOKL1eM0bDP408Nd7H4kxfcHa
bqCzuDLk5VshenyzvXkGnRvS/D0yCnzBIg1PMOs1FpXvAJ941RzJ9PJeuaFKt16F
IdEPV8TuVX/kQ+PDcxsHBVGybE1sikjGJVHzwmDA/kKb97rgYhWH27QMUbbj/C+r
wxHNWXi0WfWZjz4v98LQAeHfxu+t3XOi/DfWy5YBNXBhCHddTptREberymCLE75Z
4uAHMstKrrIcLWPePwI9z/Ri+EaoJps2H47TbC1xu4Rvx2UOE4nfs3tA7MkgvRBz
NO2Eb0htwI7eWf9jQ+OJLUpfQM8jBrDzVyL5wx3YS7jEqobnZdvGCDsx2dqzOyLB
toY2gysIYvs4p/sQVDq2u78B4TMFjygmy0SUjYIsITGa9G6XGIcBNJRh4SpPxf+j
dcgl9olsJsZAJkKLCZMMlq2l4XIPxu8UIf+U68qdDAlYeIH70eOgvctQsFBidH2P
9kOFyZIRenxDLGxlrpn0lDmYUmTaQdTiDbYPCxplNCN/B3gOZl49mVhFfF1d6iui
GsCqrN6hFH92nyS75UTs7gLH4LK3zCSvH0AL38z41By5bTEOSaYDXE7/wORKEZfY
XpHJYjq27X4HINbEvbRYu2tZ8pa5Jvws9Zsw6B1tWPClkqUfFTAEA9MDh7W8xusE
dD3WBHrGAoMUP7PlPHCJCWhlumdW6nz41kwPfLWExQ8vlpIjPJQsD6Lu5KEjRZXF
WADA/71er2cmoiDkv2h2Ao1xYlCOX6T4NUTziI//+NbRPxnYCdzzVghvMQimjcCw
+Imnm2R1pO0N8Kk117nyAh86D041QrUV+nvXmgBsecwHjLmu9vymknlgKku84Iuh
l4x3e8FZjqy50fcEAyLnULcaf5DkhGvClYNjftaUCUds6rtHyGU4nsqpnnx1Va+O
hT7vA99AhYIM2cK93ZTdeSX2rvcCjnWErST3LC4xw303gQp8W8YQZoBvX9Yq4Q1G
1/52WlhAc2Qubq6+JYMLl0uRbR4F7KpckSsCc1uuquzz21mZ35lqdRaki1IFEGoS
FKwDA/xFLnKbtSnxd6+7DjcF1BScRAYO3FE7DThjy4M9FB5CNsYL4TCiegrrkT+C
fMWO1SftsblQxokFU9JfCBvdJ3e2s8ALSudIhiPRZh8kU4YFLK7IXZXKkflCIGtU
NHqLe0qriQzqiNIDyMq0P0+iCwgATRXCUQU63Tb3JcnEvQnTEQU6I91GgPMT2mKf
t+ebfoHHGZwuqI624eJ3pnatRXNH0/Lfv73u7gaNqiMtcLDs/GTgXWgcv1OcJ0jV
MWjRrXL/PhzcOCKM3tnRV4Wjc68ZZrNrDVmjJZTbYUTpjNU3KaxiZlRTDb/O02Yo
/IfKrkz/OCcPhDH8YYWU6RBKuSvcY7gX4c/UN03LeFUl3Orzk74sXCNK2UI44zLr
wZN7VUplJMVPkU+iKgSltTuAoH7F7XLtdrk8GBFY96SArImbYJ2H0CT71DV/n+Cx
5SST5BZjbeAKjC3XO6pztMYbm0Or1uGP/N5KNr/pHK1Yr+M8429voq+a9C1jKEuv
kx6jFIx9sMNdxx7aCqiTMTiZrIUM+LyWRVIMngk+WL8kiTo/vj/B1pmEll/tLWAT
ce25SjdW/9KpcrVpl4sX99HMToks5OnRTfChnpjO6N8RNWcoZww0Ru72n+zserfD
EYOD5qcIb5qQKWqCkHK9RCdznWj07B00Uz6jDzAsa1mSkybPcCyl/b45WAbI70vB
Nyas/Vc28J20n17TrdEYhWaqDPFv4wgwBoOAOxGwwcLUehTehW64RtuQHmZXwJUF
qKSmFrNy/hHTOUm9pnCr/XCkd+k4SORnkpl7vQnDEkycOiYlAyql8ayVhQWB7pjA
KeVL/jSIUY0ljXGSxBWudsM0tdHuKYy8UygqHGisWDyfTvdlhaeA4aLzrHLbKyQ/
nimZ6J33zt6vMGiItST40V4ZaxPkVZipooJBqEjRlElqYwe98V5/WzsAVRoKcz+/
fAVV4LKzCDUE1YxDTg2MT4b/IVIRFDmKBRlGPHuwMG50H+jjYI4zFrYCgTKuHeJK
WyKJZ0ygdlTewPIQz0tZp+FZMHfblAol7zAxLiqk1/A2VK0WqNQAj4tWq61smQZw
ZcAV6XSOB5mTEvaZoDOqk4523Hf6nScZEaRbBgNIxtV1paeB/b4bnVNmBFIsbFxC
EP+vYSSTJ3jF/NcwR7vu+VSVnylg6d4KUq5mW7Qx4feyEcZcM6P+nogkqsb9u3Ma
EOffGgNvgZ6vxWDaChffGcPD+r+g9K8mXeJZ+uWexiUums75T1PqZ5swQLdrRIJa
hdvd4BcE8tar4ZL6uGM7t6R9RZNevLNthrHLCuLCTbs1XGbfLJ51DwzA1mx2Tx2r
BvwFjfZDi9YG2nvrH/lk+gqY9GdyfVp1hT7sn2U1oNdNHFDoiMWDmVV+yg5w/b5S
pq3jjUbMLGiQ2f1S3bYevBXYhUj1/uIavfv+runY9MjFtGKzUB8dSgAN7Ed0kic5
sWUAcHKrhv68vbkAqxn+wQa0LqbLP6TVUqjyteAQplLHcKX5hQIJntQWMKE+mkJJ
3TBfSEfG0+aY9qAOH+vL3AhGYNRs1ltycP5KPZP3l2Wz1HwE0idbQLC2wcwr/MN3
0xAT1t8v2qb8QEU3iQc3iD2XKKZMZJs+upCM4fHvzVIeQVhWhuPzoZx3ulS4WmZf
OtyUDmqbBHPjvRWQEmOhWS42URpKlrQQxGApJDF8RLlMlur80q4IxZXsI40nfgVu
PsMg9z5lHVjEM5DkSf6SX8S/boRTg1RKMZdG8HHXefcApRuy720VKC9OyX4lPd56
v3jod9YicQjaLQbk9bn1UW9q6I4CsPCNHD85Lew1sy7Km/0rDPuOONRjCnLi6TNR
/XpFaQq5+5GXRlP/JnIS/xsijz1dy0kSBLSsowcr8pHukjRu6rk6y+N3s5p94HNm
eri7NpZV8eijQfFj/Vi9PgpnLdX5hEIhWNXGjL2hfeIp21AMtv1iiXONlAWJT23F
LQEdM1cxZjBfhLW77l13/PvRl1iZF9Zi/UyCyn+kOaPWX4iDl9ylNjPzhPLYN0Bl
554jnR9dGKWO9nI6K1s5zJ1PzohCKIY0Yh9B6BZKne1gRwNcWGfAxa3pPBbojidi
lcmazTozofHOvJrGDNlk4I68hmnZCXpFjM2TdchAjOeDHraPRN7EV9zTgcP1V9xq
a4SGPMvnAu1Y+6f7Pv7Asp3NvdQ4ws32j/oyTHqMucOnqG8R/zdpOMTeWxb1/0JM
gddByUCGF/CFtyYZqf1mY5y7r/pmzdsiYzjEf6CBxspit3iPbXoaifto1cK7D1i8
vyLeFHWt855vY7Hbx0iniQymClDotbih993ZYEvdOebZp7L4XY+3Dld4dZpBSv6O
YxoeS0T9kfx7cA8RjvzfiIqeZwE4t05Hz/Zwp0/Z9Jk6PDVQq13+0L3AYuaib/FV
wa8bDLpR4Yjl7T6MPlvQXJD9FDLuui2qN/EP02nKs0TEkLtfUS5zjK9NZBRWS4pN
mOEc3uzqkz6nbyWj6WMFJwkRNLRtgkZCYkR25u3PfZh5rD1ROGEoI1/ygIb61twp
HWSAEe8N5DH0MUcTpe1BPKqjK7W8H0gisfTRqyy2e2FpZPIC8bDSgnGdBWXh6q7c
4anhVR5Q7ugRT7SbFMEZQzUHSGNEiIITkJCHQZUplYWzaOaJV/rAV+pv1O+fp5RI
CdUndk10O5WOvMed6ZZty+I7+JSOFuox5ZHge/pyhC7hb34xcYlUZnXM6YC6GQ0W
zg9a/WMvAMSMo9vsQm77Hrat0emcJofNfjcvDoYz53uaXO9/BdfFpPX/2YbNrMba
VnA26dzqRfw3RWaFkLGmB+2YMJIqSrp13aLI21QD2Gvn9eIdqWfEUom1Qbe/WKwi
q8G920TWnweJJJ5HeM7goIkzOko9ASLK4fiPw5TdZBW4ukPJ19RxZdFATdraouK3
mWzHP/ahCCAFUdb+QVFvTqVOjsmcLbx5qO1pAP6w9YbGd5NURK3ktZwkYpJ+aLla
U1ENog2iRkWWOu3g6DpDCjxRVoz0iNmyX0Bb581F41S+WBB1QJUtsAGXUHjvcWh+
FSKz6/m4GTPU2ewe8dcGAVinBhUJTV8J6heAzsUrgxQT7Hx5V94fOIhoyf2cF7JJ
4mZMNUk/LW6lpg5KMHzO8OUhVroxn3TwJ5D0g3KTfByrdiA6ZSzlNSvp7FrJp+YL
bAwWqqMwzJnGbx4fYMp9dr5xPS+Tj6HBid4yh1m0sBxRmKiJDhr6hihlUCiaHrHD
RuHa6O/iSPmZHK2IcUbtPLN+MhqpnDPxMHvjpewz195VI2svmnR6glnUlhSQ1js0
GDJEjT7URx5+JbhDY2PoKYqR5XKkuOz/zwlPQ1KBg9bIDzkVANsdQEgNGMEDmnYv
lV45AnPlULOu+o+hCw/wrZT8dBE7AtRUXEnCy8EEQC9IBGEIfVQbl3C623dSIApi
UEdCfC2HwibvFlweRMZNcUtD93LpT5PTkuEjbEeI33ZdE5t/Lo0d9O4s5PWJlsGX
OWYHoAJikQRNMJo8Nfp/Rq/ObuAa8e8eapK2GIfRTr2ocLWHBId0AyzkAtgcEUqR
erkYjPxWH1dMhfjDNmX77yCYZ2f+83Y8CaGnrd1SMGUW4fIO20P2vQN1UWlgDFhD
7XNumMDbWhlJrGTJzLTUcwLohdPgERDG8KEyf9wLGgsAaQRqCyq+MuBLJXEcCMgt
O+4alu65k7oqW7eiZmaDXOaNX3ATN1dGPCssOQfjOInM1JY0ZCUAyv58BChN0oIn
BisBei+t60l6xQ1iBu+P1u/Px/SlwQaUOwMcBPf5SIBRXbO5Jv1eHEZyc7kC7RrR
ze7ymMQSUE9HUCK+1TgJXpqwTUSYFMeLbHbiwBJHcGOv3oSKFXHw8TY55zLQBFb6
MIf9C5q447rRsrvafXOkh64tdVgIGbit5Zl7ybvNReVWfQNCs/YDqhz/WFL0US4e
UjO8u8Hs5PpulgEAaxRxcakaUEYfs/OOd46I3cg4+unm+3iyh21s5aGMXFIoLCeT
S3an0SbtjdueOWBEfNaPZw4BwBNbBNCdI8Y6T8tY0XIst3BgQaE4SgMJZ/WqFMih
QvWWk6ahf2oYAXs+dRslumoSVhEfbQCXo3zZK3nfTsz3DFVbFjBYjqzhzPcbdzcW
RJvk7MOxq1zBiFUZD+1mp42vUnq/w/nXSoNo1EwyD1D8HHBVwgO+dKNQTn4g1B+7
5mReZaglWE0vbEoWEgx/1hpDxWiPfOoxlI5K/WR/SxTkb+9a7yP8TqTQud24mfeK
Th2uShPQYhYeNwS/v837nriEqSVOQaECNBYe/EtxkT2aLmhpAhon83zMcQE4RrZj
8MBxgMZiwZoldhAS4AAdDgsCcPeFgAIYaQnURz8UFt+39XUWte3e296kw/mKNK/c
WBNpPyCdtoJNEDagoOuWfW8/TG9xygKEgujyjheFeRlGCBk20G8+3gR1wNW6GH7p
Wa/Dy8aK0IWTNs6QAM6EDYu97kzfzvOyUpB6k2hy57O6khwtKS0ALGVm/ul8Sulj
6rJppa4k0N8caOUhLH7X0at/3XZ82TUEe0/OYw3bg8YMdaL9zsk5pdy6F9OnUPOu
ARcxFK1+lcLBGySlJf5aEZ6Zfl+peLrts6dYR5eEJ0VsfWPObJMAQkQ4Ghy/Ckf2
Ow2Snoeq1eXZZRkywVl0mHJ4wHca7Sp6dSTfwgTaC1XawoLuvCr/4E4JbTDHCnqW
h7V3agGkOPmyhiI+f3nx6Xb8FZfYRqOi0wDjr7+Zl3mzj570pTjyn1unMOvUR/qA
UaLT3WKP4LczcyeC4m8QeyC1UDib7/VXKvqEBXwURJsJDdsTzHL8E4bBDWfgDzch
ITeW8s313tm7QNEKVoI+WMhL3qcipuX9JbbrZnT800KWl4Gw/YJDg+uGxornZnkB
ycg/myhm1Z37f/6xNyqoCpxZL7T5YMz9Rj+TXAABzRzXz99mbGLU9tHS+ApDmYNg
FqWegSiuon6MwRQpw7smllWJlpgHeDJvH58xX2WvnlOu02US3qPrxiDKpmKIu5du
loRlrrgejxvGkgw5/wxH9anzNy5BVnupN4+65ej1D3SdCNSY1B4I5B2O1C7LyCSt
4kEY65mk/2m83VBiG9Pw5Xlduh7lGAkLl+ISXqX1fxCpkylDBRINnhQ/KzSlGaEL
jd5LdQlW9Objp5HzEJ1hkzhydM5w+DtD6gksToUnrvrvsDgtHCN57CifcVtvfshT
TaE0vZFFnfnw3o3DZ8SxjP8C37BYWPbBjrIYuoI9dTqo4bIhbYadujjO7vrs/Mm1
v5ukm+J00xked+OTmh5QXDOiuGh3CfNcO5QzXu34IGcacEnczyXLelO1fYfPG1VX
aNV5QNMcX0gdJobXcX5xr2/OSPKT+Q7tyIHdnq3Id4yb7rTEfkfXSHNjq6+cKDTc
/ToLiPx+Jp7tmQiRGQfT2dM8WhvNWke72AF6UjnthtG7qolFKleNevm6uC8HZrc3
mp8yFamAr8BZnAe8kyo/YEENOFPxCoH3D2QtPQJG0buAsWemfU9soqPuL/CC7hM+
uMCUO9ZKty/vFrN7HcWlVJ/+SD9gax0PtQW8m+XchP91dIxLxOD2RiNEWV/uiX1c
44UzUFcBjQiqHXJljz8lQpBamj1lw5khrNKP9XhZ55va4bxMJ3i4y1z4iA303yO7
tbEnebAbIL9CFxcIVrlGRcLHAs8smD9nEkMFzU4s8S6g6yKaq6FNpnOVVINfeeb7
WqdlVkcK18gMdhoJf2umJpnT4sKL/rYDMLiMf5Kt4zkoUGtc15N4yCw0jqqmd8Jc
GSu/rHRcy+VfUmO4RCmt9SWeAEZ3uK9Uq996O8x/Ey4U64ySRnUjkkUx3e+6cQgt
DNaOiIFR3QdAIIKX7kRg8dNlEj8dCdPdgPA5WMTZQkHZp7o6O+fDW8OF0Gk/l0oU
nkswK/JOskyaidqdGgevW1GePwp204hrY5HyzaKDRx6ncMXFMKLbNfYaWB2hd/JH
OjaD5ed+L3MJmkuvw3XEgZHGwt7Io6kzJx9yS0FlRoNTjMaUeX33pMaDzcfz6wqh
oVbe2RIPpOPqjBQrTGu8vQSjqtygc9DhzTPH1qx8vsZYQKQHvGZCtBeZyMwyUQKG
zmpDpB4RXsP6Ps1/c58L3CTDGKhU5Ya4KHitfg4UfIbIxJ1U11y0J2UrW69+gAGq
k6ndoGhsEVJ7Smt72eUC0VES+t0DWINhoi48JnlgN19DGt7ScCyyLexBgAkE9ggZ
4/iiinaSHSmu8HekA0+4O1SyFzMMBt/GgPVZQE777F2GAzKBQvzQk3NKy95onT7a
ffPjriZDHtTsbKbXJ3bEQlEBh97hrjDbxPsgka9qfYLAjJ0olN0pc5ETwvEhuD+y
N9Kzb3Zlfdeg+BnM3wdoYFdXRgDqpJnxp4cdDKiL1QhJW0/PwgYw4gG/SliEWcQ0
CQj9VVcPyS7j/aiPDTuNk6kDTvDoapk/wn32gwNUBOfJO1SbMPStRHeiLINKhYa3
dyLTGUdM5ZjOWdBcUqhaRsKYEZ1dfcYxDlmm+eFnGkcqqWf+w/GLt/sFKoTM8UzS
x6VJjiDqRehlJ1xb1/lTLGxUs0COTLZfqVTsW21cxVaO19t8Q9lxI1/xfzB2N6fc
33c7fctdx/oL0Yx3PC5NHP8/UU08za4oYwMw+4dxx2El134SM0QM/CgcYG8hNAT2
RsbKtXo/2BKd/g8CspfRKoYxEeFoTeZm98CmC72wo0a1ZmNBtzK28C+lHPTxjD9t
qMwGNGjTDXAjfJPD2zQHyps/LeYv1c3czQdUPjmnaddBX39BAcBa39wtORGAl8l8
hwnpED+dcq2mYA+tbxAfBmtrj4TazqhP4bwHF5vOUV6/u7pGMJki5l0w6zxVpMcd
Tv67t+/ZtetY/KCX7IEsI08keEg5n6mQvzpEm0Bzk1a+Vimo99H+q11PtrMJ3Wys
eiapSRbZbI95o8rUefhbJ7s/+vXPS2yXxF9rmLuUNZPaFrWxBfz5vh/P4eJ/qVqU
vwQVeKZoweldV2DwaUiH0b/mlqA2y8nib3rnTfDzUluT0saM9YZAMlz2g9Rdc/U6
Tv4weuA2dFGIfkTZ7TjLWjs+0dprU/QP4JChY6At2NRriRQRKjnEiJIZJ/yhDoi8
9c6QvrGf7XKK7i7JfRvXdpihDqrTqXg3lnRQH/nIiS0SZTK5B1p3mk0Z+0q38Fl0
1gSLcJSF8GXsQxGifbz3hdEEJ/FeH4b77fPB/o9A18dz0IAUgVOIRReWl+jMVriw
utqjdKVM6fZXvv4HkEgkF4Wn35XMK4kDqItFih+hCbj24zKtNr2oq79rUnZKUGbc
3wP+FCX7r2w2Pm0Bk5IUXFWisDJUEFJyFNj2HdL/mtj6FnI91Db+cHnCm4ffmcgv
U4QHvAwyLjoJVsmx2hwNdoLGej9owIEwApHZeuLQJ6wK+pf963nftlw25i3aF7WH
glmxMz3GT+a6Le0Gmkn6WncxkbXHOl8rPLU9hJNTHmPPLiNCEdkFNBABQs4jqtXh
FZFX6z1XeH6syjQz6zqr1krrySnyZVP6ELpHwhH2w4ftQ3gM/9QcjCqyJWWyBlh7
vfzhJV00nM5M55s4F9WYAcduDu0RrtDOL0sE1L3LTrvdV7UwyS0M1Z6PZ8LTIIRF
hfPYXSqtgIIR/A+jPUU1BmsByIfQHZmZsHYqnMcXISD+EYOPaNjY3SnpoPDf7pU4
uMgz9IDlPrVO4Cp+cAxUVZT+cr6Pvni9E3KdOpUoyMfXAdaJY9vRZ83ck6Z+sbFz
g/Ql2K+39CgGYqOk9lajMNI0XZ9cxfAN1azYgTr7eW+oBU/UxhWAByywzSEj6BA4
UZK/tqVFimsDIPLkYpXGpMD/3HWuReAVfq41y+dUIUKc6PWJWGIlwCVKrqBHRnHH
WeRSSQaFD6t5s0y/yGmvzDxBct7J9PtrfyYuRFImHrvD9Pj1i5aj7Z5jIkMk+v91
eLZHU07lC0h4jwSt2PyCDEXILDb3eq1WZnGBM05uLW8IctlRgMHi2yL6o/nxDKRc
+Yxi6Y71YCJfxjT+kl92p3Y/fQeS46XkQc0ImB6hv1d+EGyDWi/SpcKDJ4/yF6wl
7NjfOqHy8+TiN8d3mAPfKLV6y13B75fBCyPA/6Ttpomo398jHZ8bxP1icNd3taun
putX8XZORkqEQhOZdng69ko12ChGnnRaZKsZ55kcfZ8jf41BxLXAEknwzKXpsWzV
HzE0WrnBLLtjujf1RerIYg9sZ3peVB4tze2mVCVCSkRDpm6rLOzxSUaWiwo3+cor
HvYy9uMJ1SxLhUHNxuyktUtM3iHmyO5ush/Czb3a3sOEo3PwOkxHBLtFkjf9nM4C
ZANRqrOkvFnBqLVywNmzTMYWq3vX2X67AJjXQ2Y5HAPd75Bq1jpIq7qutM34OJOK
WtuScTNZi0PhxWz60YkvlUZaS9UKuvaYUFJTjol6b7XhVwizyhU/H7CK1O/vM1ct
hIKiUj+SWF6WMho7i+FyxPWpLOvH/wAxHZxVR0QzIAuMdO+RT8eU8qlSeo9TXj2O
GmWwLkmHDHaE/SXzsbROX+hoAL6VK4HVLx3rZu18HNJuDpxVCV8dONBZhiqS3/ca
eeekyMELRnQbVeHfGF/YDgAWs6o0j+9D1Vt7Ue/7K+1x2pBidaq0u9LO6l+/kzAF
e3V7BznRVNxAPoH4rA3pyfAZQ1JFQ2fs2p/fU/hPByBCEeoNQmoBBKVt6Ls92ozv
ywlwMsYRQpEYTL0QHaHseRDDMmEnxjhrtDbj7Jxu94FtLBTscI8kazaFlPDnN7WE
1FrgnN6X2F/2AR0oEUicRwNQOJO62gUecXjIn/NpfF85dbVSYaUqiLWurBjiRb/F
+kZr7u9+puZIE0wsJMXM0ykf4mizk/AqDP554W/peFBhIOBcuO2ep0GgE8ZYsXZg
CA7WjetCfgZZLpromPi7t6eGNhGK3XOpIGBL7w6pwlG35df2epnA7N5ii20j2L+M
gZFBD25kxDxoW4Mij78QtaCZQuodug0E0RZqk8/fGwmzo4jb1DOyNg/xeDiPH0pn
m2067aOlkHIkUAEGHZhwvOwxx1gtFB5r3LoUsxtUpMxmuc2LdSgR81bAm2XFoRLk
zcH7mrRGWiJAmdhwDwD4HTk4N2o398HiGgUsjyltA/qZ94NzfshEE3fjAXl/b5xe
5KY4kaW8d/AGhQmOPaZU5JayWdvVkPdudQ9JJMkot+jsvaokfkjrkjon2bPz9D3F
zLKdV5GzsCdgrTrOntGs7bXrAYS6p7BngkVllFK0mD2ZO1d1mXuPtTcD/puS6res
Vmg5uvCS13J/ITwHmX2d6Wf7awMu/VWoOko/9kjyBxnBAxrdQsB8W9knhU0FMVtM
kFNNsSHnc6BH39wBR58X9hOyi7GaksFLJCUAK7XFEU6j8ULRqk5ZbKfQ77VVBs+j
eAY9RLbWUdQZtgGzs8ru1nTw2EFgX6+UyGM71D37PRkrpIIe9NBfv90CxzkQg1j2
Icv//CGFfHIMVMZlnT03jrag4OCR8tx6/me3iCU4gjT4kSwAtmtONBrlDplrQHf6
cqpc7I/0wn3MvAkdkEnXsuSEl2NffvKT3YtFKS5t1Sj2eCtSuXKDoNqeukelMBEb
mnRPp69Q4y+jtaxhtiBiH0YNT9rTWlS87Tvp3y2Cv0AadQY2UPoqpv1m5vn9EzSw
YUdxRq8ng9icCj1SWdhWXXOPkSVKC+myM+52uZaSeqjb26WYvT1JwlJFP1bMElRb
PQ3IwupepBAVNE2DDn6QFnnaktbWzCzGkdnYPgz+RVTotE0cevn4epEZlgNcmWaz
uSuo/EjD1ZV0Br0sKcLAEweeDN5nnm2P9VFjyz5snT3CR2zUss6CXhF44NGLWQtB
9qGMcDrSS2Ybk8C+cqw3RQrulMB68PT2cn5KsssfW1xT2jxMJ2yAgL38iOwDY8t/
svMaaF1w0T1NwE4NsSJfqJHwU5aKh/hnpjb3sX4RgHvr/vF+uuX59lNzOP+cpE25
vP4atS35ljG5liVOBm+X3ibdW6lY3CC8rZF4vOUV6TkaZ0AZM4MDLdQO93cHNMMX
PnVpWjAM/RRHV3rZhs8mt/JP1h5U/CL/vj2G7c4LV7ZlyyY+Zm6LvNy+Tj7byTE0
WW/60zSfbcrk692d5K/hwIz1gc4HsQA2yc+NGIPFDhuBsHa9G3EQlODLRsCAqc5+
UZ9FTL7wIpwljqNVhiyUdwYxuEXLcqXOIwtLR0zil3WzkNKVQg6uB37npxk9nMGb
OZFjHVy2VMYufMR7Z6yH3fufhINslCWfXlM5MzIARtidlK1TxfAbX8pSewCRFC3k
4rhKxbGi/3qVQJlpcu4Svpd0hpfWbABdlPuCinV0CLpZv3hc6Xp5U63bx2d6cg8S
yX5SltFY9lB1/i0Fs7MgLip1hvKrHi1wvyy0VBbLnGDPwutV6Mc2JJHcU9+Kql7p
00HUZUhSbaoV+yK7L7MBaUf5ehSkxCy+apfaAl1YLlkw6Ux9OYh3k6qKPj0/lxYS
thKNJdV1EaWHMEnjbpD58XdvDKKPjwZsTM8M+lWtkPDogCAiomiNHsvHAEob9R4r
UnDE8Gck6ttr7whxlysGUss0F8ioti7bNILG+SmL1zBqiVZNNrGN7Co0zB6h9kB4
lOUtXggzinUUoUupkYOd7LxL6/lgFvWv3HP6bXKI2QB8IBhwZY2LjIypU4IFjLFT
Q1zrQRYya0MtNdf99HXeAWbckjfDFQr7cQ9lBmezGmFelkwUCcZ+7K2q2bb2q+rD
q9QVVcHU9mny2FK5eq01eGrO8eeV5ekqiISAgtZFTidyxUoZFDXKqb8iLN7ixdFL
uLevuVOqBemZkL3ucYp5YUPQ9Dmzeo34KLn5M3e16laGxRBXxmklaVPFhRdB7rHW
TKI0ktNiVEVhH6QX9AhgGt1/mnlu1wUe/FeHCPQvt0/jyTIw6xDdDHHw7llzal2C
nBRcry7XiUszRwOxYKtS4SMICiR/+1lFtxI6qkRD7CnHLl/mQnl4O55MUvBFRA8B
Ac0GGUeKyBGmEBcMb+7Rl8GgcNFyk02iPPpOL7EP3MkkPf5TAkvihBqHIkDE+2k3
3+Jk3zeoXiIp+n34288tzgLCkKPKzoIygCnPSr6uYUEgRgUfHGpsq4sGCDT5kiJb
l7CiTO6AWHlwFw6yJ8pT8QNizbkuwv9Gv9HDz/FkSIc2XpZqUt1mpyeAx0Bv3fKw
L3FjowdNTYDeeROglfOkPNKF51Wl2r5eDVjpFdvlHhWfClp32Fdfa2MI9fES7c8q
Hbhi7lFBRNFpjMsbA8Vem4EE0KJ3aRlYjw9t9iTjLTdZBmddypSBYjbR+pGaqN/1
p86+X0tN9QG8cGPFruHj2MSTfHigOL1/qek4vbbt1+DCQJumGcfz9EhV8Ae9ZCpy
IoIFhzCK7FEwQm13pCNvOwSeIk0AQaxbRDONBLCdRVuaOl4/yyok4jasCcuIFiBF
OTRy6NZp5MiC1q7q08dfClYfV0etP+125tb3lPIYoOd/ktIbrmCRn5EovBRps1zX
DXLnXjIo8PquSEuX7UPHLVvrEE5KNeUuDO3OyPa06wJZrelCqoLqLubYRVXBeUX+
i2Vk0ivgIbFc6yhZqOIeFb5PvaGrOTVnSzyLfdD8THPDd9xkENbY0Z7G8Nek7WKj
rtUjTcvD3R1MwA3zrYdW2GApKhYna2P2ssekIj1bGp/5TLYGFaIaJR+gm4p+oVag
77RS/Qcfjo9NdIrvaSH+dCgSfN6FBrNjTjjsn2/vHYLWeeHn4hbx+qrRIfb7Gx6N
TKOE5mRBzqBboLobvf4wubPE8GyhVPO1LsOBXHF/NQFMXTMPp1fWr+yVDgZZwu/M
cUFL77B2BCutkcNNHvdjMKe01YFJZhoKR9ysxY9SAe9A+MiWxQAjItO+oY41zMBw
bsM3R9Bd3GbPFXTVBVKAIhVqsW4uNRSMR9fsMSBQz7lOjAdYz99bJmxF3Mg0VLeq
Zga3E9w8/zApFUZwBfsiSXP0VDh9MiTjiEX5c8tSvt6G326wS14XrsWFlLm9SQkm
k4CKetKrfCl08ebvsCJK1BzEYge3mRUrj8sW4befCz/3kqMBVn3ediQzblP5gXH5
zlZVG4tZRQwce16g412iqOfxGHWwJCbLN+b7iUNNWHrnMNUWWbyDqV3C9jmaepl+
6toiKskgKuhMrZqpyWqmNx3hC2xkfHQwEDqbI7YNuBrpLTxVpC8E4KJ6hQDtIynn
qP1579OodTskCWDP+JXcpF8yryC2JVcp0bk0EkRKzo2Bf4hPRkhF1tvxC3/tywda
fQZQFCbcjiR/DPN5tcTwAUVqOSpTjs9QW7YecJ7BVTomdkPYbQBWIG3pYjGB5RIx
kA/cUf7mMsskXVtKCTU7BPUSEBHUfTKZbBnZIAUD2SKHXWbHrBAvqVBatXVCOJY+
ZimWbUXEh5t3/S1uZaHPkn9lI3tL0LCFHjmjp483H045aitsMYwz9rp127cZHXbS
e3dGgn9YKtqfzNPeetLDQn+put4M2+Z6lgEjqXzuw9Qglw8i5TT3nIkapdW45gFw
QWFkt1siL4eut14FLOwe8fkDVhPtzLRKWEPCo6u8eCDLFnrp1LSZmb1bFbMCRAQn
mNxfxenfgNUsZ3bmnrMij7vzVKWIcJ9UYIwwzf4zIiscLS3d3dSGFb9/K/pTsU51
emG+NvwckFM5rMSAqkCi5ZcLwGAumyksji1AkUOBA3t6ZEd85vEYuMyV0ll8K5xC
MpcaX1B/N8crB8bsZKCDjlwYUNRdfrHaOAEBpNlOzhVV501jA3uLlKHJZy03eaWP
t3Siu7ApIbuvNEIlIKHcvwSp2WfqB5O86laSHC/FOLntd3unhuAncCtoSteQW9oC
fUIsCIuVl9yEnCx7t2CNk5Y+JYqFhtLocdMoyWPLnf6G0ywEDFxfCTbrYUNNWE6+
2oBfcUXwtc2oNDxianA4Hzyzx5DxkrXwMQwFQgp4cpBuS+Ef+brEgqbCAjXXJ7v5
1pPwTzrBvLBc74v0ZdcweWXl1j1YBgMfrgPjF3tD44WMXzzob5Bl2QHQK+LXVygy
I3wL3Y9jksrClahEBaeS0GoviO3QknW3M0YhlpTbbAFl0AJBdXQi6jEJA7bQrvNe
xZoyPl8FqFXBQZkXwNKsS8S4MsHBu18MzaxjzLXreHzJZlRMWxgoCy1kYGwwOAIP
OZbyczUVo1HK+a2+BAutvMP8EVn5jGBtR6uLo+Io0IdTNG9brJPqXycc4FRCRaZg
lJnMvlowOaeoCbiYp+HlEGklNn1Lms6LyCRxXm5QKJgW+pqrTR18D0KJsA5PhOxk
ZRMvWl2QHsBRxkS5UDmVKXCM9EEFAguee3APTSKlAfeVas7i0T+DV+kdBAJfC4Cv
UX66nac7IClijM97y8aHUoaAZNqCRUPOMV7wv/gvugzlIu0vEU2JgNW3yWZmCFl1
rfmmStxNwqrxa/ku55tYEVpRASvT/DqtfsUyxd+iCobphFS+qGZ+DZ673DiPttw/
xyNiHexXutFGBBiw02VmolzHWoukibYozm7oaV0dl4DMf2uG54juK3LqBK+xkk/+
TwMJMrrTWEK1os/n9LMvbopCLGPuJqXis9D2x2B+3EwVyylTizd1ycBXZAL7I+Mv
C5tlEhTXFPfIno37c/GSlSyh1j1SPeTZUHzhMpqurj2FlLyxQSUyfzwijb5rmZyT
a1cmLAs7zwJkzen+8HBL7Pzq8GHsZJ6Fxo1r7r7e06afYRM3I4qU0dG8Ojta/uga
yYhK+WjDM/nqzG958pzMoaszTWoALSyxWkDnO8Hxm00ctperAV7VrhlnpqiZ6ITi
Kh1pxn0SIbyT4I94ogVrbis79nJpoDHEm0+4wFk/WZW8FW6IxhTlVmMgZvCbxple
vkhbXEgzNkOP2RXd7quXZl84pBUnVGjmnk97t8EnhtFh6aPTMrHDxmCuCt8m+wLX
PPKF0tjhubg4Z/JQW/NbD2P+63qSzNrOjShW9c1xjjVdwQTtvGGSw4HYdK1OmcSg
WE3wIdPmPRH4ZEWPBYJ5sfUJ90Sd50gm2sQZNOSBTuqW72xJomeAM58StUOFfXYG
kf1Gfgav6SG27VaTn1QQGbfcS1Fln9kD5t4WUJVrIr3qoiDjsYY9u1yU2kPu9PjV
Xt5sbA4Gc0Xj7xuwdDwmC4dIwjuxJ8GbMQdgJS5v8EWRwEvEp/Jt6qGb5a9/L9cf
/17xZKVJ3+IR2Ly6+vmpVe3UuVq+ki5HrvVaRABNqYaIbSAxvgNQmxPbvO9X2IpY
71+PKsGpBKIT8GMAeHkoZD84XC8GYzAX7HCs3j7jPwMiqfc+wTET1AJibJVstKsC
sSch+7jyMQeQLI/gUJXd89LK4GkDGrE0snCh5PLUH3LeEXsY7U2pwwjRz1OlLcfk
g7L/cpD44G1bKbzmhCAgB+qOzhh1uGU+KvJkjkxB3sTvuAJg8hScanwwBERYS5qm
gwZKVpXpLIedc5XE5GeqU1bN88ysLqR0Hzz5AXpiZpZ4C4uFaH+jvL1mw3NTbH/W
9fTz8fFXW+EqN1D84sHCZD2hxQcd/z+B/4OVRDByASg=

`pragma protect end_protected
