// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
zCBYvSTMupQmLW9DRrYGHeUGid2uxnX+oDlXQct0catLhKhfoonIyinfyIVqywLJ
5AAEKzK7drP7nK+DX6vEurlcCFdWgwFTEsrXWVwDSV2Ok2oDaoeOWlEgGXCCPnxf
lBam7ZPvnUI+iTLfF7gVZxCiGE9usQH6zQxs5ZiuSHfBLiYzh5EpzA==
//pragma protect end_key_block
//pragma protect digest_block
FYGVdwrpo8oewxcbzEoHXKZTO8I=
//pragma protect end_digest_block
//pragma protect data_block
+6pztuzqVl29F9mHTQPx3uj+D/NByDFuBRAtpE85tN0SIETm5MsT8NoX8nSj7M95
HYPr8GauLZZi/cs7FgPjbDpT6pvvZt2MF1OeXnkmYf9XtoQFOI6JJu5U6FYIcbXY
+9eiOzMjV+nfsND7W/EgAJHVRBTuHIGeMn5CxVu/nhjlOgSbBgcNCH+HbJ//7P3w
9+t1NM/AFhC/TQEgLSdiHx3Ec8s+lrq0fltdYEACi8i1lYUBmdjr/m5uF4LfFFvU
CMQlCpmHBdhWT8nb6omjaldCNA01Zj5HHEL3PN5L0Y5j8ijQ+6ln0fgFaZlJFesA
s4PA+4a1qZ+W2QL8E6Cpr/yyTDwmeVtqZ8ndedkBoTeMB/zkVk/uYh7i117me2aP
RFlR5X3H7lDKYkvxg+rXmR1VDxdrX0UzPbuM/J+IoSSfBXuUpY9lgGmdyBctF1IL
B9WkThcnYjqDuzGurnW5JEhb1FtRRpTgibNT0T9sHdm7tUdZEzx6hYTQbXdItrR7
kIJymq4yBScNLhWvFhPHtkRaOLNmsPg68IiIOgEWaDB/K1W4PQwghtXZzoEZzWQZ
DQkYpIe/1EU0RIbvy+8M9NS60p9+xY585GeNkQVyut56eKZHleUrvMifcHpMoMv+
Qk7xc7Jhc+veCaKU6Nxtk6oB/vdymps4uA/u4ysM8jSLlzOjKZHUye+BJiMNaMB1
SHJLwgHFhr7yR9n8K81eB7jwVIYaWdGywI5Lzb/XYKhn9y4HeYpnVBZKB9x+LV00
eijPjT0ARckyuIcfv9/RSlxuPE8WM2Igxt91khNlFG8QDE5NgVbLPsmK0cOyGkPC
AygIjIYsWiR3rZVJqVsB/lPv5Z7jbmYeTt7lZBz0oawDxFBNwoHnySp13o/1SQVj
CinQ3lLhZ+6CUOoGcECGia4yAjxmr/hBtKsM61TzVOoRft4uH2i7U5Y+FaKZJb0i
kGbX0LgC8UjRnyHHoghFv424mdShPKLh4IpceK8I4wAYuHCQWvxArfImRkJwg5Vx
k0bJcP/O+/DDgFk0w8eCkRfdiDjOWpTfTtqpUoR5YZTNBpkZclUuhDARoaqQ8JD7
0g8DPsSM9V1p8vdng5/IJIyWMd/8AdmP5EmhRkNJA0SYadODyFffevo2nvfhMI3Q
gLR7+dfhRZuLJbbmO+hsuaHlCl+s3x8g8h1Zspuk2/yVQVCfZLmC2KOdwSADHsHX
RUi2fpMCCK+MNGR8WLImEkuyTUj7i+Yl+OCVxTZLaZGgXSUjtv/V6GFK1dOKu35q
fAuZqQ1VtvYttl2QkaWsiy+31I6nLkOhwmGPUuvr20N6KSI0mPXZF6qB3EYTDdHc
lvFAB0tDro4cqgRvmMJMgFmfuyQSyBf0PE4FZCb5guc3ZY8+psDwJPvJETrfcngP
pmbd3c+fXDbtSZGPJSXzNBiItFQjBdYTAb7vKXugOGD+mcuit0kPw9e+7qZBGdzE
0lfVrg8WFG+YzDECGq3TfgZywxsk/t6i00/gPycli+qR2ne/6mjeDaL9gJPQW5Ak
EF3o3UG7J9o5joEWgZJSMxqPYthQjirHgAt8KuDIKlOUS+fyvPDCHflvpWHCseLE
Xgv15MTpFLIXzxpuGfTZYmPiidTqebANNs4Gd/2/04kj8PAmxwEfIippCT6Cud76
XZwrfJb4B9ES1jNU1hoGnxtQGp8/062apE8J9XhP8C+N98g63dxJRrU3F1KmBszA
PfKILP+8K9fm05ZfHfGeTZQiFHNOGJzSpNJ42XGz4AQuf+S0K2zMrwIwx7LcYEDN
OiVEzCJsSJ8ch7bn5zrEgHDQ7xhWVeWuto3BzUd4jmYCiLrQSGDCQGFLZ1Y6kfXO
mD+MJjaT+66Lw7d9YZhhLBc5o3GBmQFH0HxSIr+QiGOaeuHA42DeaA5M3vdPLT8n
NJHqJTQz7Yq5Xcz66/5k4BE9zA59Mjwyt+sJBgmir74XZl6JHwnIDgg/0EMlw36X
HaWCAwZjvcRIeMgxXkDmUtOYgPcIQ3R4dKzesp0MCYGjmWioAGUSHaS8bf0Jgu5t
67G7c6iQpcnZoQGzyc7cqoLOPk21/kMdawJYEhsvZpZAxZVVLnzdD6LZrcNSgzC0
2TTcEDszwzLW3hrGQF1S6Hpk/OoeQYdi8q1ZC7F1jXa4feP4+M6Uv8Ki+tG5PaF+
yWI8AoLxLfxNlh124I2DzY7gk1mxzmkhYNI4W6bpPtTzTuWuXAT9NvMLhwcDk1yO
VY5R24SGGrp6WDJ3ZwSlkO6MM/NcrQ8F+RPM3HsLMPdwqOICk7ToSGgvL6uUT9IH
WC/FjVpDiU11fFESkPncLstxB0YFkdDse6o26iz1JnVQuRZ2LiQLxTw5yZSoGQ7L
ny9m99PQlusqnTlNIcYgsuXN5O2Wlftu46lP/NGbw6fxOL5DWUjl7FUwF2OYoMR5
Ft+97BjHvP8rmDTiNXDHS4q4febRVo+EHcnWlpnkX5YUYeLKqnJuJcs09rN1RXBm
OqieC3y1A0LZEa5IGz4YDLtTluBkd+OtDxb4fl78d9IdjWD48r+sV0313Ke0Jdzf
vim1lo0okmvI3o9TW/+pioqIr3S/vOH/pvrhoirku8ozQIz3ml3dJFwF918BqqJK
qaHT6fg8xNXL27oYvq62GFgRHgjx5zlcc8Hf7kgn7+geEJNUR17xJtZymgfVYmFp
tE6Lb4TZCDqbTSyKlWCDzQQycha0TiSEfnHcvnSfYDBsbEqxDVevU+10OlenMXzN
gOU+GVgu0GfZ5/iq0RfcW1X8zNETD/yLo2Xu5zAXlP0U0q0az2CCCbavA3gi2q0B
t0i6AC00Ev7Dw+de9KKBTtV5ArzlyZcJgh3SuCog2Vp8pnep9pgCy8N/VG7yNuG4
+4vdH7qerh96PBI+EQ36uLNuia6Fzj9M3ckYoZx5GjKF3PkmQCfMRF63FJicCyyN
LGIqJonmprTbII3cW66E0gr0uaMnPBLOSIoAOvc5SYilAU0kH15y0iFTWMCcmreP
0FxlgxLCILl02x9L3ZiSXnwnt3lnJGXfc44IYluYSVvA6xCbKsBdHJ/yrMUGnjdo
dXi813WnBRCni0wLpncOTp0JhY7f/8xlQara+9VHgDUifv0nnVp6rI1qNEL2XoGz
j/sFKbyvC7OYq6JMdsCn5Xs29WRKT8iQmATedpiGiJXopIsx0mN8NjSn+d3aSU38
Eo38xopBJkMHaoBS5Y8V8K4dXP1b7HTKL9wJ1H1R94UcIsmWl2u9mF4snjVGPc0W
Q7f3dLnE6GmuJxkmvk9hmFmIYXOzA2g+LPlTfnw69WEH2AB48oIsMxCkDOfJ9t7O
RlQsGkSWyDgi5CMluiuK0kdZpnGM47U+YfiNHw8DN+KtDBZHBZS8t8jGo8igyLnk
JHLISeK3oPhY3elXFJ8ao6R0kA1Gp01mWpGbjwARu9HlN7FkXLoywfDQx77G8bWP
uYizJwVSNTgqgQxM7F5duy75ijPEaoJkO5G78yUwshCwpuMVOgM4F3y3cbCCq08L
mMlBKj+FY5xTSo+YHrmnxkgbV44pPXxD2ERl9uBvYOaNCSD1HGmxrtoJIoieLMdd
geBmdU1TfpQWSJEKIqYHIttutzWDPuB16MoXkzj4iJQtwTz6BBtsbGnNDO1dR8zu
fAghIFbLYaOF9e81Ii8Y6Ysdh7QZJcDxK4YzYznaWKy8BC4CGAvTiy5wQzZgqZjH
io2LgovkdOCeZqHQQ9keGKqQUJrStxkQfwilcI1jQOsZ0k+NGErZCUzyoaZKC17Z
wtS4kQGNtsGtXNCXs3egylyRVqVzEnSt9yqMj6k3ctvM5WEHGSEQCvipordZUUyi
FbtgFqWzw9OSVygXQ22/5uNLTtyxNSHXdVjmb+jsAXjyI5b8MI9MQlihFlK47R95
leSQLVYkORYjS4tk3kijAR2fjGA8cH5Ugt29oOKjjlKc7NbjXKDQ5TYRLVpaBHiH
GV/oWUvHlq1xtPlFb6iyDW/bKkhunQ2PQY90gMac1jDC7rLySehyowG/X/QDd4WZ
FcM6Q2g3jfrwJ5Zrf9MOZD+CxhTIAQdarZZLzDftsDw3fxvPoOY6laJaj9KJcM3h
9Jtz7R6t/4ag8Pqevzo5dTnjPsafdz2YOKMvMFpNS5kj5SeWQXcBIuvjOYT3qPX3
PIOIHle7CyHuZXQt0SZU6AxmPCVKK/2XpeU/Gh2LB1I42Lzf03BgIB/D2qIyz4Dk
E1TqIq+7nQWN48jHOd01ZkVpGSVfsmO2d+ej/nQuu+DbsOooB0XFQxOkiu4DqEmt
Z7M2i2heemdNUr1JfszLn2uM9XQab6/SbyIQc5F2+o1Grhqp4GQKZ49gWXEoY8U7
JAebAMHHCELg3wypsxO69z0VJSZy8hyNnNMhJp9rIhIKjrJC47UyErNfG/5nGLPs
u/ir2nVZwT4skBeoWBiEh1Pq36S1sRXsp8kFXQuTby4KnO75XvNMnAS5rjvJMwVZ
YHfSFlGTdgVyhrrvW47SYSMKKwjzA5I6W8tMCAz/OkYoJDnfQqshyV/g6JiT4a0i
ezi+a6otMn6HNP8ffw7UYQN+l955QDNdzO8vWIJMuFSdmetRyVpT1NkHqJ3t3cIu
z1gUFEmUytcrt3MblckRfUUeMUrH3d6vnRLr4fPcTAf6B0/Kc4y/KwbVNQbeAUiB
kp6qFhXX3D1//R8V7yvtDnSdJpJm2yfr1Zhsiph2KuOvmIK1eRW2WqARlLZukXRG
bowTLjQdqoSss9oG8WsK+Ey9JkKX+e+kIGYPm7+08mbZCXrMI2vPNulLDHaCghW6
Lf+mEA+BJUK0JVH0Z6BQxUCnHhrobOBAZ0jas7EPKUvglnrfx8/VzDFnfah2Nn8i
xfNnZCsrdJaGkgl8t4CKD808SLAzG+N9S7S8dmdbI6xargL9eSjtSIJdAvGMtpEg
sKHPH4Yhy6A0p1gbeooikG621ffEuMyCmyG0hvgYbm04P7TaVRuGUEy7oxU2C4S/
E7Rf3TG6lqGlv2TVQeFzG95isWb68MCRJnaXrtcszwQW0BzmKDFF3501z8pRHYoE
7KqKGvKEFViYEgbKfFGHgkX4xvdy8YhBpFK44eeTwkpja1Z+bRP5sHVCcXYB3LIP
655gYxCSmWkVk0HsWXiy9ZzXXVlz3WxOEZEGuQqCF3pS4xjxRGfHYgmEpv0eBrtZ
9IkGukhrBkVQHAWevGhP4thRWP/e/dEHeBwhS6+OMTWxyTPpcZ7nU9vMV2j4sRXs
0F0/2bbf1ahJ+zJTc4uW411PmR0jR2ubVe2x6f50cYPelZY0IPtuHMHBUWWU3bm/
gil7eE1RwyC696UMKMmMPoddY1qvWHLXFZ1lZnBWlv519Aw4nMDP/OxMNiQJWtKd
QutbdAdOfowFV/v//W5io8EjDlsJuHL3C1TZ3CF8Fu9yLuB/pkuVzJo9s/CF359P
VF99CjKvO5TDVdnTroP7lIPA5UK9oHwXzsgtASC5YcBQeveecxvu3pnuqHJfuC4f
ylfh7hvgx8BrWMMgLqEpqJmO4ydva2EdAks1Zce1fCxCaqcN5pPw4r5EzCTpEAXz
vIVan/guZrrtA2S50OlaRh955q4QYe98ZSquO9b6hf5mUBX8df06Gd+R5EvzNioJ
8pGD2lpfEcLoUVxNXZc5h+wjFcJy7X/mkLstBOEpgsohh/8SRg5NCakkrI/sR1hU
gxTgMFYh0Z6YdXWfGia3NkR3RmJBjDH6TnuZt/JxK/qGtHHXIB06OuBkoRuWkqGG
UKi2RQhq79Zav7ZCiU+Ptjw07YiFgFxXD9g9f4kLhsm7JzIoqTN7+PKQYYpUapF3
0sLc13UDEk979F6huiCvxkwS6b/fRAchGz16vDeTuAiPL1zDu51lKwnoF1Ew1vDU
s0R9wlHS3O8QBYYNC+UO/NcC9/QkVg1cxOi9GsH0C3BruOTZ8jXgUWFQxpjCsa1t
kTiIgBiiMkn848gBvO2VF9uPa3AN71SQ/dC0FEx9tchodFaDfmhQAWHlk3lZoT3d
jcXRXQomLVqvsrhFE/iPcmx7RX5JmNFcr7bncrexHxWOElzW35ZTQW6tWAn+jqyR
KbRZrzuK7rYhBJu+jjsZJofJ+hG16TEehXqM564ylUFsZbJpDjXRpfAOnKPV2/FI
lNLNx169eAcy0GGWVcdF0eR/p+9tkpoBWlmVu8kv3JkRmvyFxs7EXmZr8nTRgYdQ
LBtSpU6sYuBYN2kafk055t4lLkVk+DWIbMbQV48khs3Smb5xUHaaJ3FQqmfpJ5Ya
cC1LXEL5uQU9DRg0Nz2iq+WI32juWXaMaJ7YnsXPjBqgJNSP8EvqU3HDRyvVX/Gs
nNzcyqdGu7mqan/kxk5DZA0I00FZdYzmGDgMK+FAe87h5uNnDhzSbnh/RV0DDPEf
uvwhOa24QpF1Thj4XAlEmVaLKdjLvJOvvqJu2nThWafmpC8nYK1dYNUsKGuCm8Ma
+13WNd5jhQ26tLd9m7MAH/wo6iV5szOIVdLiEwvl0Qm2Y3FH/fXrizefFd0KUGWl
KasPlSMWRJUZ4MgIKNVLPc57xuhegIuIzyriQXL0kds7GxqJH5gMU/k9ZlCFR6wN
y8DqYiplEGVaX3KcXK9VErMeKgHXF/yMTG75sOqKWa9FPAJ51Hjk9z1LtBDcTp9D
W5IqTjTUI97/97Z6RjfaHf5nHANzrw4wbgH7C0/w9aDR9eWqGOUPoy7/DXrLcs3w
fic0UmH1Kpk/PWMaXdZPtUYWzcoffHQviagX/NMlJk9YJT4DP9NPubg61S0SUHbp
mwBXtEeYAQaNA4HwK9AsSxLIJHYxxqkE+RvOR5kmmXx1Mh1cE6+MzukazBg7oGA6
ii8+gZHYHzcISI7bGG/CEiNuiV0jYaeieohGM7IjDsfuuISfou0Pbo9L+TRkAs4N
H7FBtc35NOQYLHidW9I64I72764NsU0VLLTQNS53OHoG5H4VDSEpl7zUB6Jb3pSU
GD6JKpbiYqj581QTFwOHob+/Mhxfzi9mjeHAcH6+FqOwbInBS5Rf7V/IiY+0gd1t
7bVWqkY5f/DTNKV4dGW9TKGciLnWf2iMCVR62/V7tIEnAVHVUPUXOoLR+6ToQSeu
b4gF/kMx48WwIFslbZklNW5WnRLKEjwddJgPhSCB+M2UqP4AXQBRDHVUFWk6N4Re
2bUFp6OCIfRKvglb88jTCnFH2VcLyi0l0sZ5EiWY/261ZvLAhCXaMvoU3Bmd2VfD
EGR5sw9gT2T6/Lcp5JTX5NBNNNm9crjmWkJlbnGvv5MnutDFULzRUc46vi8macbi
LOtKtEIMq1i4DeDq/efOjmstnUrRwHkALGECod9zmMAul9YSUAYDpL+O86I3NxVl
o4gaTyNIbXqQDi02fz3cjaAy484amOCSOyM5tWmhw+yvVfltEHtM5+WJLyR8yxop
OnfohJ8O1GxuXkQq7lAO9SzRWp/g2fBAzduSMl/ZIbdk6F8DQ/+VLJhhQ4tWR36n
rIt2bVijTN92KFCFqx134Vblv+jDEgbc/B0UacmDdNmS0+wgMSOtnyQAM0KDtVDe
UOuPoXdOCWwOKrAyM2lPTui9ryzqEppoAHY7AEnO4ro/hhxok8hYU8yt7bHueu9l
+EIkcRXhkmIrOKUy7D5WU38LximFxbclC5LpeJoKhhdqeV2oV6LRt6uwDdwXct90
vQhAmHG6gj6kI4RtY/XIDbbLzI1HYlS0Nvd72tbqiXOxg/TKD4aIX7Jg138/B2kk
3UF5zkX7CQjRwz80/KEN9eJuUwXeyLLX4QQPE7vRsIQ8G1HLc/IesopNha/KUAMd
bfjS6TdwdrwiQkMv/85HeXSggU3xWofj6UIT6zGH9lB0HzHsHYfXByjeRypIqDlL
DG0sdxqLZnr5vdKEhVj1l8JQh9zsIv2/WxL1iwqWhSPVB+zY75w4fi0+T7vvhvR0
cr+wYcBIcT2bD2MAxSsMR3QjwLyWjkUms3zDHhOcBRZCGX7965CyLF1IfWris+Hi
KqkbXkpkd89+U4CthzohQcOCf6jmn3MZHLmI1ok4lGxeLsr6BAJsDbev1rjuGLt9
P3DeUUKe1sV/so768Zifqc1kJTtoDob5kNvBAr440FB8R3LwAk2+WThMkdUhkylU
5K0zwDyIpB5ah0vi9mmtHjsAEEUF47BF6GtgwfgOHFJGTwSKY1covDAGQuBF9djW
xP8gPid7rLt9Ya8Zt4rQvBWeyaNPUkilnVHnZpE9l8tpFPN1Yaidt+aOcUtHo3zQ
uxZ9kmoS9Icg4mPv3AUw3M8e3/tRk+4JU9jdP/okfsIGW16pzoALbdH0RzwS62qS
WjRZGNXRqBR26N/2t008JAyA0bftp36MW65VHOvszj12Ivz3CZuLSOS0EDITHlcf
ZnNoWHXwlvS5vMpaR4nBFC60tdO1GTulULvk3ufRqPiBf3/ITrD43zsaTZsvrRjS
14KXjGXi0F8jYJHoDx2YwRGeUGbwCHOMS/FjUsvovfDN25/lr+UwnuiOmeQKGhrM
RY1OJRX4PE93VovSIB/UPbRXQbpRjdXrw1U8hhxwGj9YVO0XkqPDF8U0yiRWMC0/
GwtWi6vVIFAlZSHeIu6QrBndeHqBMFh44z3vUtOfWvPvtZs0Bs33AG7Q4SWlSaWe
8oA/uWz/Y4xvXw2q5HQHBwgguSDai01zFn4z1FDYvdvwrEbUm2JV4GuptFbautji
dFuyjpL7BfbV4wXvaZTzJLRoNFN1mLY0WAjo90CNFqTeiIADH6JEmi1X4hF3GANx
R/9VAa/bMPygs9VYnen/e3ulP1UEeMIdtZA/igBxbKGzJ5QM59ieEOfwO4pAySHT
5ybLjmmZIjSgmmOGh1wE0bwHqTarntZKFwmSNmK64vTrFSfuOm3xj9x+Q2zuoZVK
8VauBC2E3BlI2iR+QQsTAOZ7CCVL/yXcXWU/Nr34HTmP7IJHWihXQExe8Nm8CRE3
3n6zFFJvtMoZG/g3UR9bir1DqEmkmCniPQd6xTcelcXKPSQY1V48sLMCnWIEuI2d
ADLUzP3M/4pNq9HIhoKvoeI5DhZVWklistdmTXcn/7hPu7I6GPOFIEp4PPfC1PrR
cqOoCA0VMOHBwtkeGPq2OGxA8J9OW6EnROgAtmjkhWGl9W4gDDEegNDhaaoHxY0b
V6nKK0gklX/UGmYqrcHhFX6zkBT0B819PYEMP4F0XMUpa43j16nPf9PEs19mKM9V
3dTwORqgO/YmfWzDSg6J2Axr5VSSN09+uFxYN1Ri3CG83TsfhV2ulSw2RXm7+5N4
2QNZlrgDNAHpU3AO4zu5fXFxHUiXsMI5nrhYgnRtAo3UUOXdVbhF0Y4r3yM3E2Ae
v3MgpsW+Rx0DqGx45YM8fFvhLlboKadw+YsAbWfmW5MLnT6tafNoTI5tHD2utPPa
THXnAvvn+C6c+QPAKkB2ub8pVJ7DhZlFTnc0SG6wIamdNQ0DEqIqKy9Ewb9yTgqm
RZsYOmiE4osYpCXcO5R1bu1CD2B90Lagdd0Ezi57gl64Q+UvRFdx31m0CZ9jlSby
ZlT/CQ4c3G3oUHtHm74sHHNEx5r1pej2ASKn96HjMgT8A3gsqU9cvGeleHRToUfA
/jB+dJgKtRuNXbZyXVyRITpqHIioYYOenmpRUhAThXssVgn8CbXR6tCJrkBJyIRU
y4P4us3Us4t6mdHfISmWyYCcuAtSjZTpQzzyUlJQdgJqu92vCEhJAoyGATKtPlxA
ijvSGlI57ob4TBGfFEgVXKywKNTVH6JSOLC3RwLlrXcWCedjtd5EjKxSIvmiBMRO
jMqOhL0jh+evfATByIv3aWtD2XmRvjt6nCpZdy4GCB41i4I2nmbcMAmFhIzMbSy2
sT2W2+NrT7MdzEPRDDjWrNsB7J/skHXb8vCYCggCF+WsydeCRTwNioykX4dSz6wI
CCpacQ3LPGFRzlYGd1PSkds9pI92wGt/D2D7RfKS3O5m4jBAIQ2ip0sXdzt1HTl3
NDDEPcG3u3WUEQlZ0592heT1qImvf/Kj/06krhrmU9EymbUtfR5vQX4IKyVBB0/Q
PmYoGdu3oO0MwmU86yBggHgRZwyf/5UleJC6fNWY+RZs1yDYTbiYM71ugoqtFVm7
hUrUiWFRU7BB57jC+7vX1uN1y/zEpNqz1HtjnaV8GD1YOlu8JITl41nDpDm0AM7U
wWIdVdnobecWJO0QDkEsqH1+7RNOVEihuIHpRaGnFHOl5IRzyqDj86lQcEU2YC8r
a3ssRIiVChW6JYlCqpWr/zil4mKATXUqGbeBUleiWGXC88Z1QdtNSf608G8piVvE
hMNy5IGRWvQRpDbF+zSseaEE8N/vFF2sff+5kRc/qT4ssRxTlIw6BVIit4PlIiLR
r8/Dqi19qoolpiPzgD+xIs/ML+My7yGlFcKNHP9SKKKjNK8XYUvZIMQgymit92X6
BCSnrqpi7fTkHN/E3tGhgz27m/9NDr3wDgoz8KRsaNNclsSBBoBW7USAL375FWSY
HySAI8Si31lnK9bvh6W7vN5eoVkaCbYUaXNUEYsy+/F+PMhcaGR9ZBGyibVGQ5CP
5wEOvNNTrn5n6VXk3VK6VSBAcXjo5JQHVSdm9C7Q8C/4zwpl3fKRJqjHLJnAA6yP
CMX8cSTNpH0m+aAal6MO7H1sSkYpDwaDketrCbZsEN5xO9LifJQEarDsZKK3ZJBw
QZMPgq8zOcNQnqojomI4Cq6U0wsYMEjtBtUjMx/kyyL4uThZLe9MhWxo3yBlaK7M
aWoAHrOH9U81muC4LaJmEeuFRamjZutr7UhgdkAvDHKLmfgG8DA/3SKe5flC8D/d
Lw7aNFYZGW//UWuFkbpGtoyvEHFhQBOtVj5x4Imv0luCyCkXexHr/8gulgZBzHQC
QkeXNfNTt4fuc3gYPMAfhko0Qbg0SaixEirHDqQvU98rwmiv11bSWiWWT4IMpd3l
/eqm0qde4xWgLzWTUIaQ6DG3ImJt6e0MOK5aIPvfAkHR7LxgdsDPPq11xvgXmhmu
x3+ZB1fOcE2MrgWJPJijgZdxf5szwnk0zfjYZmpHLgleNGcsJDrdkLmVzfP+GigS
I4aMRG6m/tJpwTcVgs2A4og5OSD8xDsqnpR0IDRn54hJQ5otflwQ7jkF6QrCMS+7
H3k2VElq5uyIUVvHJrnYqwu25qOwzZX+2xzWsvynhqNWK61CmomDG0MTaGuOuP9+
oDQ6VZ/Q4bFVchuWMGQzC03fQAEt3JzK88++K0JyG/qG0Gl6x2JtpUn2ck9rzdu5
y+CduVlhOY9m+kD3Ox/tVgbj125yS2YjLmbT7ikkRWc4IVtiwhkgJS8+EoW2grkK
ybNHdXueUindkeZ8AvKf2nGzRpBCppj4ogZmBdWpI+yxC0zhn8upWTCwmTZnjPc4
+RYjLZPZBrOAedT8HoXadafYNF35Ad/EEU2HU8f+iB0YHqbpJUyqImQ0WDUSf2Vq
/dVh8/BV+TJZZxAnpvoIGESFDSCCjDO7aw03GaVG5llR2jIi/KWS0lcvQsaSS/Nr
ezyPfT0gtMpN6FrStWmfQchjhaIpsXVDyd6bJFwS3MKmyNpsHwlBaLIjIxQxTtid
qHaRYD7TQvOYo3YjezxqmhJCSdFrkNYX8MC/2ZMWAOvjkVKLDZ+ZX57NbOknVQ8f
qdKq5WtiiUuP0teENDWGUbZznEr+qijncKebvuvEI7naYBUpSYMsWT08zbxV8EWt
VG1h7tVPQnC1hTgugmnKlWvKixQc06NvrLY7+WHC/RDav5RaWhVxLwUEHrj7EkAz
obQ3MLx/S1wRXqFEVqWkIsdV2v0p6sdhDVsC9PeT8KVxNMcAcgzyLZG/LoY5bJB3
7Vr5rMJ9Aan9vdvbcg2odX9WhfPkkz3h5a23VXWY6Zr30CmI8Umfliwndsha7rDA
anG9fGdLF8T4+pPiN0QgHhDryXtm7WmXsWTtpw271FTzL7VpqgisruCe4jOf8bhM
tgQv+1frxJLyu2UF24MTerQ2RH5Kv6TQXOBfy8sUGs4IL7cnVFcT4INYsSpFkh+G
cuWCgHKnQ4N2zQwcjfKlRto14hERavbnPEp+94dWh2LeyOdwrlCl7hY1SsjRaFb8
2QpmbkOUT1wlSnG+QwD2CDjQrEDKZkZezljFFkKhzWRjFSfwV1DuTGlTqPRBI+R1
PHZ8Jpu8nuQ43qMWGpD8wCLRWuWnB5JWAjEdgKAhbWf1c/mB/yQgEOp+aIIA8vUH
1KViX7wY5KJ4By0t32Ft3/BE+wZ+cckeQ90myLP6Gt1v2eALx6Wv3mU1aYTgjtMV
rt3WjdWqvgRz8nqhRzZx9oXtrJ4N9mSDQcSRbBkf+HQeDsWPoIEKJfaNyiqMQRBU
bHyQMwhyrXG3vNQ5VT44L9LRdQdL5k7th6Ht8YLRAsi3/t+vaNURq4ihUWE0FFd+
YElBaCT2Le2xMDjiln+8gL8zVVntITrPzujtfWqVjj/pgoXDq8wjFnmvsUrrAKoM
OXKH77FoJeSC1x3L97eg7a9qRcYLh638rSYGhbIugwZkJ41cEdR4yzlVX0e+IONm
It7TBlQlNf7QbKfZNWkcsF/rQkWAJD87Z/lCWEytWwwQdzYTDYVeBV804rOQbAPs
LHqLl5GakOA5AKaq/0oF22vCfu5nlyH5dfadcPuu/YMvVugRtQm/b9nM1qJ4t5I6
EWM8nLIRlAuaOKX19/amNYeFZsxbTPYPQrdGRF3tGFaVnMCznUnZ538MSshsujeR
Gcn9Tgc/DcVKhirxVMM2J9Nuku1rxzjAenqPbZCVYpXK5+lX31MIzahFZOUMqM4/
VmUDHJ9l7dR8Jt0tl5I+VQVwCl0ngdPW8HqWDzxZ6gqotLYjxG3cmkQdNJrrsVM1
+ohfPaknLoB2/34dbCUtJuIvZIzv1wDjoJHuOwVe52holmAj9qofJs2fRGtjdmem
Ez4tipwHGD9/bKbx1KcpZ/z1BVsJa1zJcNiX6cW3zQ6Rtj6aJIUpTA4PrktB4bfO
RC+t/+GZ0u1FV8eS0J4VnYszlYxQpuVqb4D7Xhg1VP7IAVPKYlraGB3WpZ8FD9m3
TZIkJFc29eyY0kWdXD13UnfKsRNebJAID4DAWlmv4TunfPxfVI0y+hzIjFGY+xb4
bmf76jSvK1BmVCnGPn8dK/w8EXreksWQwJhl4TaC+17BIondYnLz0iQWgpsrmZN1
NOpYVdH+E7R/6awBa7suTCs0xDajANHo74wQlkQvnSOtRasVuvr/FtTNNYmhnnPk
3qfRtMsHg9n7R90pd+JWXYDthpop3t9lGpFTXr8SGg36uxAWLPT7JwViWSeA7+SW
7IaENHhOu4u98JdDOgkAtndURksnmtivmUp0UgcKIavBgKDSsoifSaoHERZG6v6b
M2Rmb0eQY5pRwfbBOw0OE3+mSSIGsnnYb5E8hZHS5KUQxNYoS4BvomqIguf6BI1e
IexczJFprfkFX8pBcr/fw2D5It/KjdC9ldF1AJqITCQdBNZtBSltXV/GiPEGbi9c
j1Qtx8XjnKnrVGsaw+DdVEFHjqeFgkWPncP5VrkmO5Wq/dGWbydHV9AnoAVncIaq
8yue8EBiNL0Ksfyt25skOqT/AxT0Z6H14q7SMvHssjUO5SmmkOkxTZM/Xa3IpTL+
Qn+NFptJxq8chk19tJ2uWZtIx8v7in2ktyin9L/bMTOo3b2nVJo8q5cTf6OnsD41
SylNAh93GIKT56vdTiMwCVt8ZJkVe/Fal5QtDmt6wF1wa7+CrRuB/lmcCbuEYyWH
87zteCY8vajsRmDYd7fX9vCL772DCsKHF6dI82GIEDSiSSSIIjkHQ1oy9OFRfg9l
QEXOGv9uvZ0xA2l43+aKd7s3QyCHMZNkc+cy26i9bLrM3PXUkbOrOH9Xmz/fQI4d
6W7esD1aSFhXj4+ssC1ugXw33TgxJAe/V+zcYK56ru2HIpueXW2XMT5D/ED/k8UZ
15Y/YCwQ/TZIvVIJ7DWtimZH9BrbShGmp4qilSVxCabqK+75kajmLZ7hAWVd/j3L
ek8Ip9MCcHRgj4UjUA+lqB59V9qj3q92ns1tJN3umuFqWvmUcWjmWi1wKGl+/yFV
4yDEq3v0wt6iNQ1ws/J3pTMUaf9uizrxOV5ZTWKZ2AaOFwOfZOsxnohS5VFhhQjK
5MgCqvbkl4aSFoINfLvKHLEqbcA/I9DsbrXeWmDqVJJ9spNc45wu/89QojxNiJ+X
mFauZmO8P4LV+0UI1YSCg3PzpNeGFGeiVHmhksF5Rkn86bf0j6lCGkS6GM4LRFXb
P2VSxtJNBzFz1wl13imj+ORmp0kpLkZJ8Wpd1tb1uHmCMEKNlLBW1zHHfoQIX8Gm
uik5CBWMvDgoTfhQ8EzZBGeqwKLbhu4n3Bn5CAfCbaVNnmIUtk5PHQYMB4jv2M4H
ly4v1IqlTukfFCoG0gNy5e7Gf87bZXOqSyjSDueTiwvV9gmJW6TxMO1KA/n+MBrg
pLad1MKwtXEOpzq34Gz7uVh6I4JSCuG/jv4V5D/Iq0jsz7lztHvk2xdHcagsP8yV
2qOS+8PW1JVgORnIEjUmn8CBGNOTolqByq1FjpwrZD64CIoa+xJKrtVpd0r4UfoW
PhehuilrxLEWXucVbrkelNTOokXFcEfWVvM72/ijfGrbnV1uV3QCs6mT2TT+PqER
eCcmvIzKRvdWPpIHuFzOZSF4B9mGgbIjGpwQKtrm6fM8wNyWqScCFKgYtnylrv7M
ZnPHjDK6jGOWsS9zIkIbi2hpAqUsLnwcFMr+aqnBccSWqmKiBlQ4ssyThYaZyxOa
djGGTrvXYsjKQkc5JbqhY5lDeP6vEM2Z7RMr5AZU8SKXb2WFiLUhlSK+sEeEaoSJ
dJsgDhHHK6aQGzf7pWwwkTaxrwcMSmAz9NHtbBK/sdoC2+k9Pv5fyery4b0HkVSk
eoDdOOt0IQgw2mLU0GmvQWdtXXZUfQzCbxMVpvy3DKHCucyA4stf/rAhaViyaKKI
NxCwNCF7IOUdjd/qxdANCSKOSxvwIZksNyzNNixdYldHE4ZEyNeFB16XRb6YP3sn
pFGZKN0r6enJDlQF3GDcBFlFTvoUQSO2L9mThNIFL+IGMR2ln8BK8ayQ2a6umhnL
3arLK4bLOFYpgPHAupOYQxDNAkekSQPHxsuc2Ka3AnNIYkBIUbBGEe+2PkF11b2+
VeNIenTmJ3KczNAgWKLN6eByhc6+etNHHs9XDbyJFL2b0Vrisk2KIWTZJo3k8WmL
TvjqYZEOMaAi2wxXuIjJ6vWJVwW8lSNvfHcjLrWswY5YKQ1RtWT6PyCf3fktM5WR
2JhqHYf8J3MHPD0FPfOBVZ/5WKvRdyQOeWgugfIA+XF266QW9L2ecyhfo8UGRvsm
a76rw0g1QVbGGlzk561RavCM8GpNYwo1kD6cGQIv6KkYN04bku3XzV/5amgmuymI
y36AXcO8MwHudbgj0Vi0bdu3HpBMtPvctJ5edsps490lBpNezCC5lCfkPm2kg7Ar
+grFDaMMKQmt/TIP4g58L5/OCRLu1j2ftFogIUJMx3QLKiSjtF5kahB+7kyreQG2
uT4ZVXmxUGfENA7o1xTqmLlk64vZqkJR2mI1aY8XpqH5TZNkF0Wj57JVwT7kHtaY
MN2BXuHVYJ7ownTYjpEdRBi4fIdszkfe6nNT62e/Ncq+cR9YCWnuGcnssmK1FQ5Z
2u1zDM2szd8b+LAuZL903Op7kq/QzHS1tiAg5PjoMOqsFP/ZKj0O57lwryOvoaPo
VegkIKFICepAGewdEaMz1uZymsm+5jcvN38smJPWImO51Lrxxl29TDhu0ZlR0pOT
AUM+WXCyVhP40I7ABGodS+uMcnI/FZZXYeQ2v3IiXCiYeJpPEBeBLVQUM0y6n1gL
4aGf9rVuFd8Jn6ey0+H7jqx3mMOoLHH4GuS5i4QE+SXXF48bXIJQI/5f0dQ2L6jm
ggJRabYiZEb5W7YpzMwK2tbtm6QyckdnJAjk+epYTwY0sENrmSPoe/805nxM3DBh
K3A5BUfxppyBq2YEVMg3aajdaUtrT83veqtxs2W+/D8/kBXUhUY8IgIUY/7yaNmq
uXnnUxmsNPQ4xEb7h/r+EtbBuyJpiQPyIORJ2DwQFGqh3QVMZDf9Rj7sB0qX/3XC
Mnqp722krNwlAq0WAisF9qnpG7JtFBDd7YPrj8Thn9EYluouRJk4rF10StRFKMRf
j+9x+40i4zj8JVXEAI+dl0JQE+umtZx+h4sEXQh9uK7n3mXp0C7JEpH2+sDJtltG
q+3WC/SPB80Ho0hxDRhXXSJj2yiuhNcjFOmOjDw4C1ys8mEkXecqOqCJwxCoLFDw
dmY2INDN1zSt2UTbdDRuKHcTL7tlL3oE6OCl0htP13X6EJbWDGbJwP9wd3ljVAV8
CHJgo69tnTXps783Syabv9SQYhI/1K2cLHkcbwo8Sl6m7BT7SGAXQ/BkD08WKVxO
DhcdyG3GpIn615/L/9aSnVzSOT2mCMwTVivB2UMsS+oTwr9OJ8FOzzOjfQDDXyr0
hWxmWK6Ni+lTb9X1C48B2WiJMlbfRszJUkX/cvGwU2LMxOBED6LFBKIRT+TwIN1y
jFElXt+2UDFjJSfRkzqdCLH8OkMsiQ1fDWTCMJ6Wd896obCzNYlg/KKP7i0x0ezx
TlXFfu9lUPY81Y5bv9ArEOhuFi7xo8F88Y10YkIJ2e3yzQbXJeFEkQ+dXFNQXwd0
5obEFyjKOjtS7q1UXlG+8n9357bXag8PraDnq0wbfeSkQ+yjS9RvxxpQ9n8EGn+r
li84PY0IEWfiMTqCkJHBB48vn0JUzhV2f7vSN1ZocY3YlOR6nqV8qD3n7j0gpjR3
63D0qTDhrn6S5lKiGdTkJaREIPgEHb45unz9FTW5Jq1DmAvOC4glGyR6Ikl0wZ5L
OVMJ3d9GLUudEtS47AC4su/F/37oUUVeljemRn/13O6SF+baTSXhb1shGCZSZwWA
F9QVSVa6b4o+dTxdcevfZXTooh0y9prxLTQHvMKXFAsTucO7jn5JWWG5PwJhUEqU
kFS33ezyam6UmFYgL5OBSGan1CtmGYRBwmm5uUGTV0O9A5DQzQsq/ZT7Sg53kxZr
cQDFE2KBZGVp1TVE+mhoL7wJW8InbcdjiRvlR2q/OXqBR7gtv//3y77njOOO7vKf
yJNlRMs0TSHOamARgamhiDi4kOfSKapJ7+bDzdA4SnYqUd6IuC5mAVA87R2U9lYN
hCKrB8cfP4QqM+qujpkmdHPntw56e0Q70hcEFCHh4exaZ+ZBM0QfBWDDIzMYwatx
dM4FAUZ2HnCdvbdYXNRY6Dix9vUwSFJyivfNIw8GG5DUSSy07J+TIIaogK98HeHv
9RR8QoN1Ae0EKDrnL22mQR2TeVtZqhDlPc/fNuDNAGUORGNmurUm//ibtnpzipQB
cnGdcJjIYffs6bf47sku1UsgKsAw643WxNqhs9AiPw2Bo6GrXpAAwfqp+glV8O/n
eVn6hXYcK8owDVXtlIQNyC02osQhmkdspfIELTlGPHlX+U0of6XZY/0yWIBT+Pf1
tNcDtMgFbep/OV82fnA4dsBsS0XhH7Gl88mXsFmA5asGhe6j6I2GuETdpRm2nScB
Ovj6/Aklu4K6ZZqEioAmAzEPx61evH4uXuzReatNGYLhHY3Ppq0WYGvusjV/D9NP
LQpuIBf89LowlEtWPFHGyswvO7DW5XuQTzWdKgI2x0ggxig0Ppr8QBYmZkypoMo5
nOf+Tktqmtnq2NMVwSn+RrmjoLu2Y3KL9EalvPgRSceZmPIdWX/4LybWm9ivNUXe
meIHGpzvc+/41UDvxJDRG400LrPM7rZDzzLRa6oQcdFVU1Vx9/6nAQWCeWao2po8
L74dNeECs7Hs/YubjDd0mHKEpNCJknWwaZsLvSsu/166zwb45ZUYQe35qXZB2zZH
IHOmpuRkkPj71+lsFTnvzV1WJqYhjysaD5fd3XZ09OsCdFyzEnFE0KquNEShFKNi
qrTi1sUv/5OxKzxhoLruwbk9lrQ9MLUqDI26IBNf1TB4BLdqbuAa+oCxyzLUzPgT
HuPVIAmJ+JJAcTzSfeN+y4RrQMvohyDo0eoiE0oKEmtA9B3cEYaVt8jelNp5i2BF
ErwqXqO7jYdlQ3pvfYKsl2J9q5Q8Ykk1wz6eLtNB5Bm4E9rPlq8+6bAM4FGmWnq4
hQsuBaL3tzbpd5HooAvvzLkB+ZiejFKS+loOOuv7r0hh92TbPIlBHQQuFchZdsFp
sdzcAk1mDF2JtfNnA58pYcap7Y/s2VGmO9zcQ3L0l5gJtO398qVr0E20sWrSp6Pi
NaSdhwaV9qjRAeoHkKSpnfurcDLz5f+fwI7R7bmjIL9Bby31n8PlG5d4JpaWyVEc
apt/uB6SbykEcprLGA4bO1CsbMql8+tgzT58qiL4mj3Ig5iMWDiS+iTRgovJVctf
zNkwtTmRbnzPO+ELySekmBF5tI6tqjCrpIOgN63JIikzqS04MO71V3fCoHGhwweR
3xB1UecdbMcHWOat9085dhIZ/DVsXtuRP1Q/8HNZ5nqMRTOW9Oxv3HFTEBQHDfTV
ET+GQ0LfskxJfhulgB84ES8Xc4e9ZWejFPRz5c381VF90jUTWmMAc3/SDDJ+ePU0
AOrNdTwASyHDaECFm4U+xexiV4BFOD8WRsLcnpLIrx3AlNuRXModL+M1BQIDGT59
BCQaT13/gDzlgMDG1khts9xHMSj67/ln0TNaSx6dvDIPLZPjQwg8XBHrbEz+SKzv
a5ha8arzFsil4qb/YoxFlp/lpmA0XyUdvdMjMwMBGec1EoWVu6nSf7MwxhlR0CsF
lbdKdysvxKnlSDVqzjz+wauenybpwk2Ro5QbNf85ur63d6OgR9voYcEYCiAUPHyD
CIlllnEKhnm1LqNmlUWtJMp3pcOxArHyaKmOv6UevPE2U6bunDfSWYB8E4jNpvdT
t0R5+QSazwPeIeQLyOcEU6I1ER0y6PPVx/gA+3vX3isIPmw3XzSI3IoMlsuFMuLh
LdIYbG4Y5tv+5V0VTFFGZyObrdzK6b4X+MUEqe5WwvhNhjEv2V6o7mFn01S+hzF+
xTOaqOu2U5F4fVUMLz1b4p1tWI7OMeoVwzPJGZncEYY2G3AtiD7hsqg6I1coq/Jw
aCfr2YFlA6ySl1OCaanSJkj4X3f7Ml6+vcyOYH0ireQkl8iylgxcvfbyl9noCdqI
d+u7WzBLMqxxF0JNZ7Ncec1RQ1y3EQqpupdAwXvldihLKcjhxtv5z5Ajsl7vJqys
4N6JllGKUkbAqaiPrkX4qeRoKxQ2F0+3wPHrw2MwNDW+B9QGu9Udd9S68GPzV4kH
U+MNabSHC3Kj+eJdV7mJ6KC0ZJLsjWD1f0O6yzCpTGUhgJFBvRdesybJPzaFOP1a
7ViTABiL4KuPmvyRMl1D3uvUsp9xdgKRES0qCkrgehsthJQfqK4MNmpVx8wWDlB2
urU9I3u1ehe2mBWdbw00m3WVPIn5lzFTPes1rTzQQh/0u9RyTxImy4cWxcbKDWpK
0dYjABCxW7IFWTaTysJimyJICFAA3nduqSSe4fUUpN8qMVw4/v1Mt2/Oir0L+60y
ktfQw+qXP0Ems3UsjAKTxJjt4tTOWoaadv/9sb2Qt4LQO0PmR3hVgvPhxYLI3wGU
PL80vqqIPC/UH3ep/beYMcTHLR71r7aKt1Kfjp0jDs5V/NGEVbi48HRN2DHEuSXR
8FBD35+HY3+paJoQ3HdhMBPR9Xb4ZYE4X8Y1ij3doI8xKz+/4YsQVznES9cLDx3K
5/EzqXpLs4HPbiHMtkJc0lkAsJIJUkGbgldVvoC7Pd6MVWeL9QorOQ8CUUIMBI43
e7TsdZEWKKapzU25RGuo9pj9dh809GCrGuIFyzXlMJab2LrRna/Q63tU9x8912Gy
9Me57NezyRkvaNkbXl1OvRQ1/3P8tHvohkfzK8BLKPMzN09YhtFOBpgZIcb3/0Xh
MWKoeVg5q3Wv3NQag101osQnAoI6KJu7AbuPTNigk13eZzeUMhch3M0o7C/g46eB
ujziPI+x5+BQoW56JgaVrwUpLUmu2XlquMCxv2f6VU6mWUGOGmAAHa9v/ik88xF6
OM8GXspRIxtacSzGJ5aZ+etWwMTADdS8wiAxg8GBRnATjlYcZznR/8ix7hWl9mbC
owhvboahKyPcXZBI7wir5nxlzXp3M11NW0VyyGdqHiP2R0I47fkaEzCxKMwM1AUK
imGRM36BeHkXRvx1yGpzJTa2TvOKpTExHuE2bYZFL+mbzHhI3iTEbzOD2ro+k/i0
JvDnxnw0J7IC6r2WC19F9e4JJkdvTJebsVFatOGuorvmP4govgRgPWWvzy2A8B40
PBGZvetSS6s37aVKZgm0BsL96rg62cNS41lhkvIA8a+fjiGsMBaDVQT36Dx4g3ZB
hcKU+/KQKj9aiH6i0gZmF3DWxT4K6P7GFKndY1DSUdlOR6qUcJKuOtwOv1OQkw/+
6ytryYFXmqQ+MTlCGQdTOXJviJ2g7RkocLkGECeFpGdiGrGZOBrUP0NgYguT5yXO
FFRZXqg86CVVzgSlyQP16gIKTPPpNou3ENIIOtmBAhEOGE9f2A39bi7+PDyrvqOR
KW9+UCzqteK4O6ix5qEaOpLskZXo6gRjduldphZPmr197clgjs4U/NdEqLZWXrKo
3fGgC5zCJcIH006rzXnXWRexF2w//2gA6S2utPT+Qp53TWGM9NSBOVCp9KLqCTyI
lIFCu9sJ0IyLNCGE6ilDiQmT+MkVBUZEx+TPB6+Z+/yslS1VFRNQLKEicOXjN+wS
ojqRooSHI8d39I6L0floHI65RcMbpHQZywejmbApYsDGH7p2tNnecWFXPEpajDr5
UBlqZjq/7gMukTSESPjCYSCix737yykgxi0D4OIcpAZbmo9KBbls27sdCNtgSsUY
7mrWwoNVC66aD7XutrgtmsYlPtc6LDV9i7AXQsX9NWS+tybQBAil5sxB4S5z17Ei
2iQSJ40IrWfdpnjhIRVm2gtscvFo/suQW/YMoWdVHusXp1iw9Y7TXb1aFnf+ExbG
USp/6l7I7Na2SsmIl4Bsu0wiUDdsJdL+/D6BBd+X32lY90UrkwZmq+hcNm9E1h+P
92YHCU33ZWrqjsyt+JoF7Rxin7Vd2lplik5pM6dGQREICQNLPBFFR4LQT8YMvJA2
/Eaj4dFDhF7qWOp0Qf7Y106k9VsHqRoZ01aUcYSnoyzv2mmiq7Y7xz1cx0cfPKpE
8p2QwIouRrXRaSHKtN0RerzQdXpvUKjudT16GtbPuNLQ/skhJ4lfsXFKX3hWMXfr
jeRpgtmw06Ev+jA4gdSKlzarj55pDDXTX9CGA5Pf/luqC4+iIfAsOkfAoV/u8GI+
k/mFf8YoKdnYqdfGson/QMGXHaTyGHnBId/iufBVoFywtDjmaxcP1zUVns4mIdok
x+GGQQrik167qgKRlEHl6YJHURBO05jAFVKC1Wy4Z08UK7jpnZaIRQk44qBmesgP
clWTA1boyBxWn6/ujjr/mtNSJ5Si2rtE9wwp2cg5ws+FF+6O9lLDahTcrTKIZfSr
hveUO8FzAdsBG5ZGbVMZbmOBX+OwCCRBZRBnbafMdXcrFTO6iO68Ijhp+Ig8xkeg
G0bD7gSftGIxxHl4nd6sa1GzX9sI1Di/FOPFFexec0gWNVGS6RbC8G2XzN30VvI9
p6GedVZzWgBz/LDLPpaT4eMgFqZml832hUFKoROOsR23KIP9cCm3yOmGGy1S7Hjv
iQg8LVHD5VaTvkgZY/2DNSIrj1iQmXf1+IWU1C1kHBFswEqinDKXPiXlfr8gJXoE
6KWpMk6IqL1KkDhau1X5adUzo2ZIC35oZKTcVdGf6Nj+N6rI+GvYYQk71OUFHD4A
BoquvlDlkrbTvmmODX9NR/eY4N5liNOTn+bXBESMNdgLaS/PDvaNhSTE51/fG9mA
qXXwajZVMlkUn7g9dnjQbbSUP50xekZe31SBqRebAu6m1g58CqSJX04FUE0itAD0
KopuehTTasXhDlB7demJSwu+9yNIIZjzkOdvHmLM3l7Jjchpc1AmZMLIvmfaEVfg
/yWAWslSr5lgC4NcFKCWWCXHfCutO1SmhWWGx/H0XxYfQare9mb/9e2g4dVFdX0a
quiQwRQX8tH+lYLHe0GlOy6rbNEfGLE0/GiRDLgjdF/WwI2CfxyD5/sVTla15jsT
JMEv8gcRG6oenNUxGRv2w0ZSEVJwuxWAZQhOLPV4nYqhpyy1uqBrQ+z641rW5Y+p
1AAYjoN1yrANyyY0+2TfMPGN33Njglor2kwNXn4jxE7SzNm0Iy5k/lgtwWhykX75
clgxqHyPm3PiBsIO5iiv9bU+snosvGNaE6t6NRvaffM03yc/65Viwwu26zpxhPw2
+pEnV3gnn0v2TvpQMYeX66XEUx0lpijd9mGfZvvX0/omWyOzm03rrr+aZyKgsVD+
EPvIpSP7BXB3eFpITM8bml4ZpUmk0j0SALVZPnzehlaVKRg8ipA+BfdXKEi90BtP
QF7isfbx565gaoZXzn9R/ebupkTR/wkE5bHSlFBG94utDxftdYOZXeYMUPIknDeJ
SX8Msi5EqSGKUQLc6k1J77+03n6+/OENidc7SXgU0QG4L8eZaAbTZfCsAcYX4xNL
8cxip88edKkCS3HP5E+LrvNIOwbBU8upOtpqOPdHiy+i3jsHG24YB0u0jP2jlktz
+LEP6D3eeq2y8Ek38ok2M9aQDKchf4Ik/YBgyGqbFcnKvzEJeFw4UQTMnzY1ZB7j
5lvMSO2GbKsD2FwfmwtzDq57eC8DdzxdHi9UqbWpWYCGtErSaTxDCjaieMa5Fcdp
hHGxnx8uF2NzdzFYh2XWIBCvnmlX7Icfck7bBqsjNQ+Y/auqYhSw2bHoGTbxu+lL
zZVxIxbGhD3xJFfIKRmO+9WifuCnLrO81F+oZlzOzbmX8SpC0DCdmScX5ZC1f+th
UgOIw5DJKDCF6RcluI5Rz0KfQMwXxnTEMqnP5k+7KkZoTqXtbF7KaGtYbkuF6YZ+
HIKl+mkbDt9QgctkUNuYUJuKsAxGT9w/fyzLWghcDiVQXly8oL2uEhR2yAgtalNX
XLpBUl7e4Z5orb9h97RBKq3IiHrczmo+6lvpg+J4+C20k9riqHKr2p3lZqs1z8u6
JaOFWGK7p4H+R9qKHxV3TsJBgd+lHje2wVIA9Un0UsaaYrlDicMz2besni+D+l3G
gj3fgCvk2X3EsQP5/rNMLNMiziJjbBk0lrgkQqwXVL9MwZKlVQOVyiOLVb/Ipb8/
dcEMPvHdbIfSrPr3AvJ84SBGgFuXNodmHF0s/Z3nd+UQ37nhZi8CwMayGAYL/JpO
r/ERvvBoyfcfE8bx8td+Fk28o1MRrxrxspIMo9pj5F+O4fWkCTUJGmqT9ye3WMZ1
mOtF07i5Aci5xu7h+IA8NVEc2ANVnXnalyZh75hv+nd/aXFxTOuvopTNGIn1NV5n
h2BAHcm8Fs8kvXOsKYGkk/XPHP14Xj32HiNrFQmk5s4BHy587W2OxHncHXbV5Zn3
JZXyGYpWTU3Z9+4TdPxY7Ub1hRxmOUoDwq6kE4F9iic+gejVv6NVPgFqHLuIaOaL
LtoYlIRqfelQXbpQLPdwEhmlaniqcSUEMrn2TV9pVqp04w439wt5mXVAQdsF74zE
eF5Y+L3rlj+XVpG10jg3VW6X7q40j2+Z8TdeShFRisJeBwz/VhZ5/N0ilHCQMNXY
MhCLMnkDpJrwOYVPahILASHCAczoQ62zLNNSesP1Rnpq9FbUObWMkZUrGESFPgT8
ufXr7wYnBwhnKPGdX3EzQINMf1DNCGQoMqyAjHWeqe2vNcKEhMXvypkT8d4jy7No
z4ZP2/Fl4l14z7WGiZ2EdUyfZJir+JP/2yfPLJQNYm7Mwedts2fipof08Inegjmn
lE7yXojgTuZATLdS+TDvBOt/hGLv950PWyVZDLw3PomcA7tmZZ1FLJwhqZbFXOcU
kVAzyImxDsKIB5+4SdfxpyCTQWPL7lzVIWPt3O3ezm2w0KLaTykp7s6o/EiDbkR6
8sHIcZNo2mr5xUKqaaEaa+TT1Q7T+ihUS8aOPDSsPFNmtmkmicboEDEdz2OyEdjj
tMAnRrdJOM4rHjRHfOZsOZN/eBmMqmd5T+djxR7fn43GSwqAVqVQjciPLROFzzOK
vGYAni9iSuwp8CGDhElPoWQpTBuQ/e+mWoxCrHnzHSDIfev03H3NEbwuVbVj2MAK
+0ljVnVJg8wCaQRzvI9kXNzPSz8vbak7qGh1DN3NmjfyRUcgLoBb6LadOOBKZDvV
uvMzDDmq15fvxG+QuM9nf3+GPZ1eU/ZZxQB1kQ0MWxnJ4FK26+tc+Fbhq85gIUOM
qQamE2qP0cBdwcnc3NlwJ8EVVID9FxLEA6/AdRXCK8R9bH2JdzkT7nS1O2pt7htH
TvAeTLSAdw/+nz1WXxi2sCdSJdiOfaQ3ITtQ6810t1dB+mCErEFLPl12wusbWmHu
hMRdboGXkeNPCoLg+sqAqWmz9sECXu+B2MYFxJf2IK1hvvTQyd7+h7GDyKMtVrbr
alUXh3RkJh1lNqanCZnXGDG5Yfv/F2Yt4cTifd33kE+p71T18ZHtIOjp3nbvhj68
Le7R45k01kN/RApZHOF2xDlbZA9yET5EKPq7QtPRfIBZcTdjQPLia8ZVdiqr2LiQ
4RWeNBG9dLjqgqZILlCUkmAoUTZLMOhDla0JpuLnT7tjhSj8ueNWg0uFle9zgd1P
yx9JFK6aWfFw7sh2c6KxuAjni2ygi+xZsi6+BqDPfxfxniNghbnjBVLcpAZGvNG6
zDmeu9AFQy8PaKAUV0C07AXN6D4hWyJAF+Wq3v4YKGf9by+jQfIy+vsXDrlZWS1n
TSwdKchTNjpzcDyF/W9et0lnSPqGfhtCTaj4NTTK3AA6GCahzZ3Y5xlC3wEfHjhl
PM1V3N2FcJ0w9JNaNcnE1Mq8vseKm+tMHyvGkzURw8HxyB1QouGE0IjdlsCNDARd
NmWcywysZZAnFIw+s6J+LkfRIAq4Iz8C3Az9XxCe2uY/hmBrDkkSGWc7CN3Io9LK
faaLSo4YnuSENRvNK1RRuSdFyW4ZbHCereIHhp2xd5bqWeWjqTxjtPsQT/a7p0z3
aV6i9V5O2v79aJNJF4ZmPswjR8kPFXJWYp0dc+N4HE/VKKF7t2de21ZJh2FhHLbZ
d7aQfftyLOTmRNVOfJm2yPqMU6mwmachRIgVsOT5QYKQtN4jUH/G2A9whm5jm6Mc
jzY7wc3yTTkS2do5jGUtaKpiPfm9GIb3koFfeFFM006wFNMCr9CkDmXSPYRuD8l7
XZ5Zr3XHupYSgWCaJo1Jyi45OKc7P2IQPmQrQtwMDp6tvY8JLksDMHL1nS1pAB+L
gHStHhrLMERdhMvpJiLowzpvcsbnGRx+wwJE/urwRXQ3IaCzPxAVIoRk5MkiBIgo
fiySG7aAXTwFXpCQAS7H3RwUeyO/W4dcS5Zi4U4riziaOlXx9YNJ66PbC1tyAVKp
2ehBMKGt8wPU1T88Ryv2DPzD3FMfzscQyS9MN15jkZ4yrlWnda+o4DQVHSBJJGlT
dGY1AOaJcls8gsEuMXw6oQLrYlK/+30bwNpOSfMjW7sPbmpZBlE28H3xA0aGC0gY
qIYcmT1tL0mFr7GvEQvEcHU9/Sv7gvrnQ9aN2eHgTKI/aGwi7v+3AAw9A45hcNSX
FxKLjQ7uQ+GnW9c2cL5XofQBc25vilMS6JE+eqiC8tUN+Kwb+1/Nc3i58XEXYAD7
JWaSeE3B/Lg+tbxNugl/rFqF/+4zKNDBOKrI0unuhpRE832sk/hF40rkU4B+XgGC
T2CIdKLuG3yhhUY+p5X1zaVy5Q76Sauq0KKGs3UHmG5jIJO7feyeexdB3RqAkza8
ogSpZMgwm+AihBNG8M7aJKnGw4p2aGaAn5TJVxeaBtGtZI+LqNTvxoxxwD/eBVbl
qZKiMkknNRMROhHnERsPoqyIZkiZqa2DFNT0Wp/gFpKFn695voMfp9USnZHaFGAc
Jk0zP7RsWd5jmAv+3vWhIm01Lq7pIDczvOe72pVtt8G+24x9OB/VRriOaPNjDFnl
S1D4mbftNcbAu7yWMlyZAbPEvbrmJgr9OT/nJBcFQF6LHpIoramYcMlH3NIzbbra
kaNOz5ouaa/HBhEECw+hoION0O9N3g/tI8t6u5Z+s+WtmJLyv5lwqUZprb6xubSz
BP+Ta3Bb1zTbuIM98gjSeUDIjhtcGa7N5m3d6Z7rR96qI+swJxgBofrbCDrQwXXy
uvK7yQAMYkZpdiMmu5IS7muYdGE3GhYb3HAR2HJMXdw8R7ID/yEX9AloHjjnYq4H
lq+waox8oa5IDxNdh5sg2Nk/w6liGYSsWWigHq2F2Tjsb5cvwGuct96ZYDhyvtDj
x50Lxz88GHb6c/MCXNpZs7MVvO4/frViDnqeFNTBdTrGBa90bXh8G22B4ui/PzUt
ySQYpebCBeizBykceh9VOI/CcGHIjnrCDgOPgcMbZx/Kwp0jHN21xzihNiZwmyoi
tzjHLT16fdPh4KQMRNdANiI4UZQtMnxWglmAugRjOG4mnuK/9HQoSNxBQdHdIH5r
9Ec8dKvvZKLsefP/78DresYMbsln0P9UM4rXHHaqCSdHBqtZqvCO7URAt6nKzRuM
9GpVXZhszXkNEzOg5iePmN4PfX1TXNVw6HQPndvAE5ZgOKVKR9/MI3VVs3KeBx87
r8PXPqxY0euOc+E7y5wbLqWvyA1HapstdXUzjs0ygusR+huovT1OpNfvEYhFzehR
pNelUFzikysEOumnhTn8jRYCOBuCAeTJSZa9CqFq4mxD21d4uONMCNgEBesmH8kl
q2Pc08f3YMZUo8ZW+YLr/HiDPR+XCmDcuxbCYJ1IZqvCITuD4mY4URiuKfUC/4hw
wDLrBcP6d0f1bm11rwu1J11VYs50ghoYxJfdEjIrlAAp6noQKlpU2Z5UZI4H7Fxl
cmsoOBqSBzuRDw31j+PRVy7A3s/34a45qIQWdMTJHB0xaDbucWOOmo2Mk3M6j2T6
i3C4zt1CItsHtO666kE4Kct3cs9bJY24KY4MzS2tUq9kKO6zjs5zz7me0UGiYW4c
o2xAU2rtNRdiU/7Lff1dscnOBg7AygKZYymoevwKgXqYExALYG2pbSo6Y7ZP1LOk
QLkVPiQlJcSusykSa1nIojFY00pyHlmTO4fNtjXcdlcysi19U2TAX7T1NqZFbjO9
OVTR5mkx7OKelbCcI2LVQgCcsDKmJlXr5cQqvh0NY3MUbe7LA7kjgGI0v0v9icVP
MD0w/cppqv9s7MWeP3HahH4+W+8rxNrrwBi1OFxxm3rDrnyradhewAmFfIKycnXf
bRux6RT1Xmgl+4ULjsNSo/EkVbULdFmzAQnEZvtclMU/xwmzQCP4SDi16uCzgV0C
rmjebTblTm2FPKJsPXK7lr9FwoZmAkf8V/uPFX9T3uzzK6mijt4TED/gYtGhkx20
SJ9rLBDgEOw0SehFFPPLSnlzCn9esCBVSTKIas6pAquBhLrT4C2r3o7sGvwgMesB
sKIY0dOkastB0lCLlnsGSI/LiHTXND3+DkY8pKb93fa1DMhaHJGghE3kEe7hk2Sw
hBE1+mb6QW0enuMv1SZ9/3AUycRCUXwReRmVLaujMnptyAF92UfWf/JodnIJ7vLa
MU/mXOV9IPqmMctkXm6l6fownmzQ8AerS9arqC9Cv6SGQJQUOyh6wXyLfeNnMw8o
Xz58rtXNjWqzVmugta9F95G2xwr1hyarkzLwunduaNhD1JIqZ1XaaJ7TKntZlDGw
LrwGhuERBcaTwqhns4veLTdGpfG90nHK5ulRVm4U5a2U3JIy719FaZ5QxKIKbi66
12hJlE5QabY8bh/e5KzjM3chEOyLMpn5OmONSGx2BBM8umemTiFyXx8LnBE94SnN
ghUP+ovH3A4/GF/Q8bSqDC32sBbhiQbz1i6HLft8J8Ha8MDLBtJRp1N68DhhQoGu
fefZ7c1XOimnxPDEn95gIqOTFEhP5DepW94mSTyqlwoWMQQVfZwMtKwfmw7k9JOw
0ciBmSDoze0WNh5g+xL4P8AeICX8/jUe9zMOF53HoBKDytJuYUtU6QtbKCzzCUzm
INpQXBwMW+dw34Uncy1Bj/YsBwGM/wy9t5j88MMDh+S4e0b1StNBwhENWK0nmK+C
Zfu3J6THi0meg96/+svqEYyw4H4B71InQG/U6RNdSR6/993LbDfwZFf+GGeZiidI
og87Snz/Y22rHfZTYt3b/ZvmoYa22clc+gWH3NOGe56VXjDBExh1ueQHTdKaBXjM
mFIANkF8u0gIFc5e9NYPn7/9sPTMMxfOEdhhpu8X1l5eXj7A94DBCEXF4i90qNVP
lby5lJLVL8ME1vm/xgNQhg7V1vE+pr6cnVyhuZvOzbuGeYLqzIJtLgFoeygGqkW4
1U6ghkTJprH4MgLUePV2Wkep8800XEc1cJD8kBMubvhNGqWY0d5xovO3ewNxYFtX
vjwJg2PtHuRr/rsxyxnZvlUO6iR+qKvNIueLCdjmsRusN8vEQy9vkjLR1uaVi5Ui
aPG4rvlRzD8S8hrFCmz7AnNs7Ojb4uQvT4zppO0Beig35BddS95yc4C4fBaloy+X
RIv11IMNruXThvKMQYqFcfegBhg80fPDsN5VsAWXEwi7MCNlLTGWrxCEQakmYJ/g
87wkA0fCk8bebKovSz/VbCfEXsf0dCFJXvqLAMO1UV5jAbknbgILVfN0lhblvI5G
ET+i1LJ5dkyH8Cv1j5ThaDoiqxY6seuvwIbOQwgVfCMUSRrjkg7IqmkRWoHVPrwr
+L38IqAF+m9xny3f2LxSCQt5AiGJHpgw8BbJT1hAQtnEvGaSRVfkjfsMN8HFa5Rz
02Zw3qEDGPgWUE5bdeF1aP8w7Z47rpxPvdYcQ7jDqF6O165ATJeSnx3H0nvC+y5+
/6Fw/6ZkhvrDD9f9TsljdWUrA/f0abTJ7Dvmp0lFvUnIkaDOpApzaMEcgcrpXglk
12N7B1baLdQqcJJbXHrSlFRUHmMm1vCVDqt2q66tasHdLvZgZm2nnTuftb5IHE2+
iWVHxYZFbBkVdMhPkyT6Ra1k6HLlVGO++fGgpLG8NMzbtWZ+WcRnVZpukei7h0mW
Y7068vB2nmDySGd1cpWwOZnW0PPljIlkoolr9W3pBcB4WzYsEMeMLMMygDhyFGR0
c2BR5vXlwUgVRBswyGoiK9ScDmHRmYe5o13lNc6VmgonuoJ536IR+f/D7LFCF4Tk
+p/nmKorl92hIXx5pzm9y2P6L9HdYYBdMPJ7MlbxamawPXZwmE4O/NFmry2y7bzT
UiOk/0OWCaWj/llyr3M4N8puiw8cfar/L75Bng4oFoF7vL+oC1MtEZDQyQvq88HX
Mm027/ggZouTAtabSYn2BY5eHpdkZn62Zz+BKBbVvlSwTTTtk43kwHe0v+S/sXHy
BlHncFXtDG4YJlPUQBWTQYXO0dgjmEZG1rtFe1JULHq8JKbwNiiu3DkD7qEpwizU
SBqlG97Du3lRADBi6grUT+N0kvl5geKOiGIhn0JCwHTkvWfy0Ce/h0XOmlYLmWVq
4CxyTukFC9MuYwTFt+QV+JcX1LwLlb7aEpBI9K8QGneC3Ad14+xHUlGAZwWJJeQ4
nwYP+jhglHC1QvFTrBLXylbbxxf4wU47ZvIHbeseEY1i2FMMb/WW0auKYMKia44D
Iks+HyzYtJqEmV7Lav+LtXk4/PUGhZ/t8LbQjxIU0zIxnuak+JMM/6f3dnzRqpvS
qhHxMyFs+yLUGQALgtFBdpb11q14sC8vvKY4ueFcnLpPtpDVXKrBPHG07n1vJdmX
zdLk4+oiH87E/bgZwkm1bCOj0qOeB/pz6uILGqzcvCIbH4br3x1F+EvMg/j/NTFz
aunXPB77FHjuSozthmzCQFnFjG+RA3kxS1WV2pjLWQgiiZIBHzHQw0oonNrlw2b4
QU8NFNWdor2Qx0gU/Heu5qmWxl4S87tXlqHy3QBmiRZnm+1e7KZzG5dmwSZfDwTD
cGNU8TrCS13eNIeredVU0iqrPDzej/aN0XH5p32MoQBsDBKsw8pvs3jNbGPPqD1H
PSzy9NzHvf+W5pyatmacOGYd3Df+7ICkunHzUmmOGkF0O3hK5k8j2zxTUT8kdmJS
yHmIYEY5j90gipmLQvIQ6wkw//OW6TCXG2OOku7xi0LSK5/qoAvbHjVO5kW9/fTH
1gEnKY+zRpoKReU+IasMl1M73+8kN6cLyjImWnDjQcsQoiYGcr/cMTLQ/O+MLFbG
qmeSlTVbgpsSPRY0WniB/+LBNN6BM4bpWMrjRMUBWXssh3X5b2UWmvVoahmlneQR
HyuW7Wf0uAWYPq83C+JS8Ow+2jqAmK8gHVLncVYou9rE83Vm+jyZfV/kVQkQxbOZ
W9hSo02hqC0C0bdZyEui5wIXZEHJZcNRVQYASi/iRcbthQiyeZODcEray85BbBLh
8WnovN+Zjn9tDho3ETxr6RldBs7qfrBoHVCzi2J+AXF7yVDIIkzXEhfaj1zHKpyK
1+vItsmKL6PvENA5mZSxHph7nOzquGZJ9iWIn4zCnfNTshSSW0Sgn5d/sjWw7Jav
VVnrjlxSMSYJpjwmWmGYfzx/kfqPyn3uqs/aEuL9SCM2uJlrBdyWy/Kud4auxr17
Vn34pgMqeEDOfza/H//n7S82T7cvuhlHez1veFyyNDDrEV36qq0SjeYRoNxgqhkh
w/eUA0VRajIh87uTlmNlfrfjjPZ/D6tfDzO43WpGB3NF6eZGvRaaka/f5xhj5LOH
EQZp7kfCSmmZfH1Ila/XtWKmv7lo65jQXgqgV9uKoPoVDBAuL42JboaGS9IDfNFH
i97RhwrJE8DCQIV6Kw/UfWOMCIevnzKyLLOe5NbPxhPuPhuGe8NPdYwKELGGgqnx
KQqnJsgGd4dsWf4mIqqoWyvl/LYlz2SSKh1wtIWoVXu6pQKj91q7KePQHYR1GfYQ
AGJiEnKFoZ7QVyNO5yU/8CLafE4CM7toYoVqXyWDxPCGRR7akS1eLJse5Ex7Mlxu
M2i4Ai3UgnXFKX4zzoxLSvnFv4YjT/cTbU3i1FfmVXIXiLD1Dofn35dbeHauzlmT
ILovnopG9U31WR/RWARw+DAct0TGnaIgYfV0rbi40eutzmCSTNOLoQ6yeadm/dHo
BRB+3J990pNao9xdD0poGyOkFw5/6i6LVm8fYPNKO+dxPx1zLM6P4GITdDp56lBq
KIgcVGRj+wo0OwQ4MGyGSqyEgPgPQATW1BCToPwP5ysCqZz9YKBsCZJMSrPqYYma
V6YGASvwmJs6CtssGAPBbec5wJDSJnbZl0Xp4P4CQ80nA5X7slgpY7fPeaDF0Rjc
YVgO8fqM5MpA8nRodRda0gR+Y/H+bC6Vro4ixP0lewZ0iOj9Su+Y9EJA5/I3wnZ5
/F4GLY1DJ25bqXKw4wTA/VdV9hdaawN2/Xk4shiUZUroQJz5nwyn9GWWKZzyhSSR
1Fqj7p6XGwtnu1hzEh5fnAXITVSseqEjr6+FJ8yqrsINCwZrWNVVk65k9fXgukUZ
TXmErJKj+MRDfQ1ru1mJiDTPY2KhKvhHOQeye0KNYNoWxs+G5E8kFvmrpsezmj7V
wG2gniLmvj66iK3SYCl5EPyQVExTL7QOjj+2n5c508PYrl/E7t9FbLxqYIfzJbvE
OfroweE6m/pGJ0XctuVpgG0rmxkTFF859XJS/ObJ54YO7VbSHI5gb+07vcVD0yqG
c5mDnrhWEIpkL3t0erkGlL4so8wBnAOJPWgOOtrfnZ4NcfHRYPUWbmgxte1HhTo7
bJ9twNaDWSDrTIkqhYNj8vFunxyQ2nxwIyjsnUFshVTVwmV7K5G01NrEsGVk02EC
yXDehPVbvkjQQyUHnx5HrhGKrtmKoanX4knq4zcl8ecuOMuR715yWoAhD7daFXhu
H+W4njIeDNQHwQ//qR97z3plkt20mWe617eQyT10BSmHuLgSUSPI1ib6Ne46aKsK
I6mZNK7/Ir4kDe3gluksxZ6CI2ePFfxHKEnIBcgh+dnjEf9TJxF5AgMMpTmrsngm
rVXt7nyBUdPtXFVumKhOg++Cyw9VTy9MkcVBsGZwPB4UtF0aNqD+v0aeEDQhozNQ
pU/rbG1Jv57ngO2HRpZqvonxx5h/IWsPcvEWlnPLIGlE3+h9g4+mjyRoVDVCUpP1
j96LZm6TyRzlej+vz/1qKQz/y68a0OcYbQaI/2Y9ZDaydEIvDz+odC/xcm0qWTxz
DSN3RqvIAQpq1Zm5JEjDfzPH2L5Ao90NkjQGkywxe4WLmorI93IIzRNdRayMvp9Y
ZWWpIoNUIKjCTOT4eaHyVkXBgXpEgPjLZ/NOAFx/D5xmFNUh1dBYjMG662wARrP8
c8pLp3hGY2/9/lfo+p8XZXPTdcZ06eZ93Vex6xwTmd/OCLic4TZVBkH5sGfzKtBo
xsEZMfVMV6n8fOXfc6nyhWbXSpYuEi0QkQNdNZxYYzjY0ZtZhEEqmQ3Ng/wyQoJe
iKz297E5IDMfH33HZ9xqHfdmuTNyRTtzJAEDv2TJuYpWAk+OE0SBS8L+8CaRrV1C
pRuKS4oXn/9sYOat4cj0WARi05YzElJGuwBkSHo0CJiB/00CJP9DBoOwEEDY4OhS
T//UPjEXcr2CnDbwySXQa2KM0IyXnvQFQWtCFakXc1F3/Bmp6qu/Wd0FdG0llK0K
TZg8s81DwKh/EZyPwZFffWU2ROvS06KaYcFlZAs4U/qyrhSouQ154Mux/ZlAouOj
uKEwhDhL3neE1nMoVsnx+UOV2w0pu+Td3QhLcCcASn1tjfvO4OmTke6Ttz5RBZrc
mAhpy2s/4E46FPspHl9wwl5ynJTgY2WVbq0foD+Kg/mnJGCoYdz0AajUd5HeUOvI
U6HeOsUDFF7WsrC+GF9I3HwFMxM7YdZ0xRLQdrCa8UB9NmypvMwdY7ymjohsvNgS
i4+tRl/QuXNbsH2sw8esvX3RJDR/xYmIYwy8EuDZlo1ZpizuQZFuIJTlfcSMlKP5
FxkduF8tpySzvKUJ/t+oJx3yrdpDGalKwsi9zhQpCRGCuluNS3l+yublBGlhvp3/
BWELbON1qnvaQV5lYlzifyF4CWqNh2kZk+r47xddFQ9DA0CMtkpzgA8gFIOi/Pg9
h7PlBLJ1ypDFewNREwdPrZjCUz3z1br8B8blslpdAXVv7ghmYTVpaThCNPZn8ps6
wgzWpA7tsBPs1GuXDfLVWx7+Y6K6xL2bRNJG2HT2kLL9d/3p7et0SHQZ5AD95Wzk
fKRuk37/QhPwueNX4OGqrygE7WKDX5nQB7Ie04z/AYawxbpknjP6oNMAvFHK1+y6
VGy6E6TnmSI6usbQQ9ker8eSqJcnplQowncLM68LfYJ2FYYHHy/foaSDsWjSCjoO
4l5NOFjs52pzImJcp9wogwNbWaUpMazZpjcvWzgvjdcX02tdace7vIxzI4QfsWIJ
0o/p4YiidFbGc3LwlagJAhpoTVTNLvi77r44Ss4fwRJkRn+hOerLbPfVGJUdXY/Y
xZE1xPwDFIB0F+oFaAE22fkqt8L9KL0qDKkLg7W30MsNWO8XKN3Uby+/sudk/xXB
W5meIOo8by+n+X8m2LEpivVmi5ZWxCeC0pqc2thrtMBwA/wuBEw53iwv/KuZo9nV
DjZhGhbuaGRDqKwXzfeCphran0LA1viT70QJOqBiaK8mnCejHfD6HNO0KmwVHzUc
nfKxLTjpr0pmq+vvbJFNNVBJURgbLzvXV+pwMUeLi6+Xl4rTHUO+C+f5cTjD7cM1
wFqZ3Nas+DrmpsbyCT/Q5AnLeU89KmdFJtXg2sXgbH/PQ/+albiEfYYJ+3sReKzF
xi883YaxMOEqutHQT62DiMGjDNXcvZOUtD9yNeW6o1npCjHuhyx49enc03sFSPOL
BPuQ3B8WBaSiEmguzWv6S3fGeX8dSkxFG6YVUWBMnNtQBV/WDkDdXqY0r4hXEASx
Xj+E/1/2AJHnqHfya8zdnFUubKA3j2EtH7nN4h5suZNhrqg5IRhMl/CurNBq3l/7
PTOhuTJltpjgloEknDv8u/sJOT6l8Q435FRypuTpVhu9PaLgtpWraA7oaI04chse
bwPWHq789b0fox1wjJ+DDuEFWN6yxRxutr0XsubaEUJFEzWqX0s5+3ly++VGaa5G
vRx5c2f6OUlyjaimp5xb32sSkierSBqlsNm/hl3TirdW9riDjNmSRAA3WRAuk2R5
QPyhNkxkV/0l/IR3VZQGi6MemM+R6PULNmS3w+Jbh3nHzhWxbvDqFD+pINtOho0/
OsviySegWrBEJ4L2hMBRWJV0G5Lbem9lTVPuy19ytEMKiy7yZxQvJ3rmzAAsnM9x
fSkPCS9pNkl/m52pgch2XKhL3XlH3dnCypOhWgYASWRQNtaNaV4Rc+Us1eyGzrjR
GSfpzhTbRxDQgn64CT8ni7Bud8jqlimSUwO2iIvSDxizpEeOZGxLHz+IVNYnox6I
9YQnFxipO3pPri7WYtumvnxPPHoDruaJSaED6OtvwlNjYmBx153ySefdMXBAGsJR
wRMss+0dlYSY9ngzm4hTCozGX2HErRznwqfeQi8BCwluitfS25+0ZKXb8+Iq53s3
XC+u8CPZHeVTcttS4TARUDOE20yc0pciTW64EkkkpVgnlHdarKEiFdueyetHE5AU
P9xCJ3RkH2lRHpQqgeFAY3a2sfgdfZyc/Isgy219J8Q9/cBK9UsQPADFLdpXG2uh
zEIeGualtMpMekH61amw0eESx2HC3QrX0KJmI8fBgEdY9lRmu/VArVwTg5DYQUPj
GLgI3rW8BixDJiEF0qf+S/14fjRB0Izrc2S+yfs+MzlCNxwtXkroEeHOL34RLcAj
KTel/VP9OgQRfHJmgpp0qFoUKMXolVeKaiKYsTgm1mxcbgC53OIFFt7s8YiHrV1k
beBh5FXV0/piBCVFYaLdRBPPc8pNnb9WBq+dKlBMh9qP9NMrmtPPBlNbSOsW4yqk
DK7EZXYChn+OltYvglcl75KTHx8a+AZn8t5s96StA90k6pWoHe0Oi6HXv03Ti29r
Mk3/Tmf8NVcN+N4ZF+HYF77YMa1kj7YBCb7NccKvsoBZtSkjnZXN4dn5OREyOp/g
PbKKNOZiWQ2uDjIWOWm+3Iwh+99nCvlMCuKHfrfTNhvuw0T2rECeanizy7Kwq3xX
wXjQZIPei1SDarziRmIiz37BDXp2pA4YupRGLJTnla2kx2ORB3wP0yJK2gsO1Goe
JzWUt1e5drtF080edR9ENHSLJQh4aidMB/Qtg2Q4R3M2QPpm/vGh+wdusApJeBH1
dtY6aWYV0OG6xLMDwLC/+IHaSAmKHxv42LJMi8UnBB7kyIqI8pVhIcTqis6Z19+f
8tQjG4KUTiQPHbO0rJO4II5o5aqFhAWnAh7kPulUhI1frt4MfNNcaptAtXNBsGYw
n44GV+PfekMqXDbO6XZWsN9js+tH533xAV769Ew2BQ7QIdqprRc4u2N4g37FIO0f
irJScmbaaEd80WdiNxVzDYt1tAwKfQEccJTvRCi40S1B5hTT6UlAoOXwc/ZXfSkB
lvf49uzhGV2GqnqTwJOCYqzdLD24AOjNVG8GENPYi9O8WSTPoXt74Vy9FmH0XWFn
hqoW7SW/R4w3qxVw4HW1rLR/4H9D5xfaOYvvOPb0vPgGd7vJVdWs/ktUwJ+RhZym
i3M3EqHTTWEBv4DxQbtFZusR1U5zsveflqKdS6kFXMAoegQH5+IY+vX6Ub/f/4Ao

//pragma protect end_data_block
//pragma protect digest_block
xk70naGcLfzh5xmV16T78feK8rM=
//pragma protect end_digest_block
//pragma protect end_protected
