��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�a�ȝ���,��p4���,�	G���L�1��t(��N�|}	"5�1����kަ4zf�HF^U���^Dqk��sr��RH*���
�D��;�<�0'�Xť]�5i���Ri7ڸ��s�`.�i�"��N�(E���!5J����k�`Gt�C@0��-�NQ'�d�t�C`a4�y�T��<�GU��L"��I������r���&��U�qp�Z�;�uZ��4�zv?��e�Y
i|ٱ�q9��L�-���%��=F����c&*f��,̟,�ު%��$]ש�9��[�&�!��Ypu�O+H�Q�Q(ZVB��3�+*����,�O�H������זu��KmM5~ABOה��?���,"U/[���2��䩵.�۲r��z�ݟ��tC����zެ���A@�ɀᔮ�\9��7ӳߌ��\�td�����ײm0طIMW*��ɟ��������~�t	(���&����'�z�MTX�&wP�(�~�9�.zbr�A�<pv�K��"#wu3��R�%�9�֕�%�Z����!In>�-G�Ftv�vZ&����gD���)S�<)�?�ǌ��XOp5r߄sn���u���]���leP�ю1��	R�Ql��PN�/zf䩭��#����*��I-�e����j�{�~�S�[h�\��j��Ezkw�[��ɭ�r�.��L��ri6K�����ۿof0�<I'�_u6�A�W�1��#F}������<rF��/Y���OÍ�7�v�W8��wZd��p��Y�4�Vl���:�`�z�:����`0�O�u^�vY�{t��Ja�u1���8�o_[A����6��j��/-U �>�u�Z��ɲ����mm�y���s02x\c=����*�j�%�V/g)��'��-�΅���`�T��Ī8��+]l~��I�=e���Ҍ{���H �?7�����I��ޟ�(�:8;1n�l�=������H�󱏿��>�;��d�3ͷ��T�4Q�g��Q9�[�����	����0��YY^9�"�T!9@'���u�4k����<�mu�H]v�N���.C0MZÞA�~,�\p9�x�5$"X�)2��y�����a�{�K���B�J��ꍒV�n�?��N 2bz�����Ks�{�k��dW*��ќ^��Ydk/�M�2�:i
���$�z2����T�E'�ޘ@2-���~#����e4�a���ʩ�f0@B9�|�d�#HYV}'�x?���>q3f�d}��[����h~���&���M/�/�HB��9��z�J�~��@w����Sq���fE�R��v���׉ů�M��l�av����7��?�{�팗&�WUf6h���[�5�6���D�Jj�����U�/K���rn�ij'����t_b�mγS#%$_hq2=�h�j�
��M������ݰq�����u H�d�[�Q*�%г��ɒ9��y������&����]3+s��b6�����'��<���gI���Я�3s��@m�)��\ C�=�\`�U�+ @�a8�$���2B��zv�V!�0X�VB�Y�*�U�܍�������F1���pk�[;��A�}P}�8��{�K׃VxJ�ˍySۢ��FM�.rZ"�؛�R4�}nm�uݶ�$�;�ஸw� ��	�1����z�:���T�PW/s
�bI�r��JU��;���x:?�~}Ve}-�S��6�&��#�n44������5�]oJ�)�H�����gR6UCo�Ԍ�&� �S+P"�7��"7�9oU;���K�t�D�՞��C ��[��O.'1�s��9��0�s<��n�1e܃��ii%U�OR���*�8�ёb1���B�,�"�4*���t�#����ڙ*Y��C�c�ɥ��}�<������C�@��*��2�H���Oi(N���k�2�^��B�PP��)�ъ .�`ȏ|�SC��9^�H���l��f4K�����ɲ�1uQ��Ysz�Y)]g
"�
G��õ�I��kX�s�#��K]�oE���X3%�S�q+�8�����J<:�l���"<@"[�^�Vroy��ͭ��nA��֖�]}��zdr
W�%��?ۆ��C��W3�~@�v�%�"�B��Z�%h��� ��������5