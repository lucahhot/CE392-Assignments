`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V2Wbh9Wie5muavXiWMv7fGhjExGvjB9b77T5yksgOArsN06IClcxbuVyA/FhZ09i
jLavMNmPRn40KnCkwRZpmVd0xmBQrg31PlpL9+Xb35+HRRvjTMng+0Rrq6y4I/ui
AMod2IES/tPNsUZ9qszFudK1Qr35zsjXvDZ9Lq9RKpU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6416)
jWzKOlIKxl8OfEmO9syB0pAH/Nr/71GvIeZCyoj/ivYlLjbT/3L2ki3sxC+grFL6
+mFbCgV1A193pJdzc8huTKuGfxASw1pxgI3EGviL0vx8unP9pvLxHS0FQd4SmJvB
w7kn/gQ0U04J2+TNYPEGw9Fr5ABgpUiCD8QtphwOqIiHClI4cImMsdiuEGRoghxR
dJCdVHkOqlf/nA2A05rG0Fmu9uFmvrV4bMeFux0kqvHBl9qeh7N6uigMrnVneEN8
zId5PpIqDMs/nBx+EcPTz+vK1iGOKGi8rbcXq2YYoMsFh7bZAoWKTrpzxmXRT3CH
XBzMtescOZlyHEIK8XXfLnVgQaZdSPFT69SQAUuBRpPVhiqpRcw9XKGYKZ+1EZwj
reTdMgtMQhR6pGEIHJZqFfLYgZ3csYHFztQv9hSXeZeGgH+Kk6NZSVBJJgLfO5BI
9lJ8k2yYpxQF5g2i1IS+94JC+u+O+35c0T+3E0yaqDmhADrMzr8WhTqNWudoRQQ8
erBDCfH0mPvONelbcA7Xf1fFtPpjx8WtqYPJvYmgdrv1pLm0Bzl3xKnUcImhJapY
ZMp2n3QkSMg8AuYj7F9JeIlEoak9Htrt2P1t0WTi0x2cdcBL+z78qGyqNei/H3RR
yQ0gix9C5AI2hz22qqEYjwkcquhh/p9Wq7Cl8PknmaXO/m7i+ysEoDMwerrHL446
2p0t/olJmmZcIW9Hhp7sB0Pse8Gb6JbXovh2KdTn98bGapekz5ukQRmsgRTnY4Sg
UBrL2JbqvGuH1nZrfBQaxwQrrl9ljxXesYyQ0fyQLxgHoiqYu0vKzHkVeYQPv7x3
i3UEALJt8V3tnEs4DufcKumz9IEQZ5HPp3EqhnNZfzvbx0jvAxXKiDIbhD1B1mnW
4f1EcvSfTO6e/p/gcbkRuG1+h/cYJ5M10gDn5vqaft34WM5L42rnDozKxKWif37c
CAEn/4FLrAhvD9NWOeU+BQZX0xvXuT1cbOdI08P+KcXtoFiyzaIumYHT8HVTvQ0g
J+2IZiXfMhs7pfRkezGwjN3hbHn/wc7ONzdzs6vfYMLr4gs3PIggerHYtV5z1ZHa
04XvBrL4EJNE/Zc9KFBDp9lYykufowoTXugblgzXMiq+4TBdYgDJnIpZIpwhc8kV
4YhFQUPolrG/BweX8IK56kUz9gIFB37msEqoXzqbOt1OsEcAGP8zlvCoyW5WV+m4
i9pGSq0nnzQMkdOOtSLfSO1hwzNwZ7jL0lbeRE1T/nudu71j/C+7O3Uzc7IXayVk
OtKS+jWJHEzzMELbwB+UDSppJ9WXJHXctFcnXGCfrg+w05eaBziLOvxJxDviIuEC
j3qUV3U7PzeJBR/NZnxtDOAta8AlpeyPKmcavLYpUtqmiyFq/RbSLK4XF7j4BwWl
bn03kKLnQGu65bNWHIgHkBj+5gKJKT5oExqFTbZ89W7sxCDtdmvZ0ElOEKzudGX0
t9cUMC1fXZN+wXv2XWHKR+B7CTaJSOgGme+9US/L5DvfX87uLLy6Q/KDkPRjo/9n
eI1NJ5D4kjcKLhFl9LsuXLJdkrOJKsoy5U4T0SL3xWcxdoKgO9GDgIr7Sb3KcDNW
A0707iJkhvDO0YeWwi5JkNlNptQu6Dw0fhLlzenTFKuos0Az8rA4mh5sZBjait16
IiJMhOCkMHbPwI7kYV85qr5GKNsv6uX8d3t/BKNlbqhoKQ3FyFcXSx3McCGLV8hC
jxOs3zpne44d5h25+JZmOCB/xm3Q2yuyAbH7sn7CWfp63PGWeOFxfr3yxNDbWpTx
/3Gdvj9+IUV1n6YvVEziEv9SibqbRxLIlDLgHYCGFFsJ4XFZf4pbjmm56zBlwJbr
io3FuXqf/sBwMJq5PbUvhNvtCiGFqxfBja5psZbWwNgpzDY0UyjNRNDb7QM2/vG3
x/xpiNiIj/wbwbS2MmKzItj30a0uTP9d5PTzfpdGO2N0DuiXQO8Kg6un1qM9FViE
FCVVNHF9lUGEuAUDFdHJV4sr/0Ybh/Z4WJuuKjVDJz3nXbSXH9wOMrU80XDAsxRt
VxXNgIuf0f/zX4OB16GrM0rv8OrnZnBbVSsmN6x0pLNAyFYczFd/hsB3BbcFqc9D
zvTFGdm2HQu8vlhvLGmUyN6ZUq6JpYYu7uN/iO2WsVH3qoGXVPzks/tS1/ZcIDwg
q53PskGZ48ZZZnR508QTux250C2KrA4QNdDQaPKjKn4yMxdDPj3R9gxPTq7mgbGb
ISIKoDSoxN83VDPcGqRC3quh+3RUz2KX9Ypc/2FluT8P6tgHBQA3F1DXnmJuHQL0
PU3MOAcyhQ2eZIuzBo57enqOFbYVaIYA+2nufHibOCwClSgVZGkG8u2FgL1fbgCW
2kd5Brylplhznz14UBGiKtA4TGN98IotxZKBKx9rDcQ78qZSNBxf1CuQ2oQW9JtE
tVKHxPsRwCWjREOq/+AjtuWMcedO2fMbYd92EC8UuowFg3WhuZ1/Ic7nbA0ED5Ey
dUP6YKlvqIgwnCypePlig+VlOSDX61qfn8AfFeBrEd+5R1HwXiQWGmpw1yT58niV
n+cewR1CYzLZ2J4KGAMUsxEVc/nTB/dhFEZPqMJsfAuJ5ZMGMohTVPytFmpXBbOU
E4Zd40ETIhLne4o/FDkM//cmmNw7+8033zwmt9LOJWuA3CTXv3lHyoFXakZJ6qQE
4Lb/W7ZqXto2rHRR3q7V+pphit79D7bp1EjpT5ftJBpm2ZDFKibLsSwEqqQqzQle
vPdLqwY6RLSISjNS/2DeTb0lcAghbKFvya+VnL0pc1B45cbr/QdlCuu+jtXIsgee
fJKicvEHWUGMDhAEABHSUogSRsiZTiLWWpZF74v+t5jsBAVVzPAzBAJtjPUdoalQ
z6NbpGdBN3dNz31g+cPjTIbQ8lfttmWHc1x6+n6YhmDxs1TpQmxgRg+LrK3Orfo2
tYO2wSH2mtEHPfShm7rskGheng0+4+xYL0Fq1hsiLKjJR1qff6wWFQbq+HQ34hha
O3rTWQ+vt0NmUHaBRQ39x6FZ6VNtl9K25gA0aZBaqVEu0kQMEEIgdfyIcDcansjQ
RIaOyZCowGhZHdTkW4VFTZcdRKz/vpU5tDMJWAoxGCBtpimgaPUYUrLfy4eNmynq
8SpHAPkzdjvV2igEjqDdln5itvej4BmSD8Y12wa/IFFBMrZCYYbQLERAjiDfWp6w
cMAMtSqpo+/2FWsnpG+rHH1mnnmlKU1BA6+0C7TCaTJ/tm47dItFcAF/SiPAjaHO
v6WJCTPXsK1Cn8LJvtuE9Faqn7EEiCT42tS9Yls1KZ8CBMlMURtPVNuZkvNf+3O9
eFfKxIr/Gc4zTI6adIoZn+Yv+egcDdo+xD+otTbyMtXQDNpuGg3G+qo7g7wNAELM
f/WnZw/O79a7MXL+l+fIP/NfRL/BtF1TcFFwAMio3CQVI+Pp+F0rIQYwloTgWBNq
/m+c6VG0xW3/yjr+IWXT3H342HemR6s0Re9eyUnzluobYmj0i31dBWkfyyP4oZU+
zcFKC3JIMfw3z2vEF1fGWA5LO8YjU9ZWLUojirielb7xOi1aSuqlJg/xw2DU6g6l
cdK0h3dGdVfdG/2UR5cFe4dK8VAm2R0pc/5AgjGFTxhDZP6LURtOiujyX/gdRb1S
NjO8JuQ6XkJdB9dfVeWZIAhAG2pBPoNWCiCPTkCmcMADiMgt3SUMW6205kNS1+na
6Z7pfTP7uPtb6z+1TNEm+VUArzQ1k9+uSA6iM/6TEntmz9DyGXDU7z620K9Jarfd
ngJwLWtMgWIjqC8+dMI3+Uu8aZib9CNwMOI4uIRBAsWYdm/232NB5umscYjxTx8t
OR4sqOCJb9XaMjXl53LJRcEGiIYvj21KaKg7MjTiPIe/WuT2Recpy8baojvekBED
JxJno7i8G7iZMqrdWBe4INVwGVJI3REuXP73TQfiXO2DmTvB4B1ln4whwVHVIyM6
2Oqmle1e+GYaBUa5V/IL0paPRLm9zcTChFEsPHRvKRhOnEFoyUV5b1vSSwu6zrSo
1ZfCV7fsLyPDu0MRfpIFCwsbusfUcFXgCfBNUPdu10IE7mDriZQo1UJ6OGYEfOh0
wgv9QrEJBO3Kza3kPMTVTcsVLWNaHRtTTsQP+L8bp1+/PwBUymQN/XEY9asFP953
MMH2PSWADWhmAPS36MaYYa+H9ZKVhyeV8ME1GqfU5CdU6apENYULVDc+dpmQ/CSI
XdhSpfzZaG2SmWSwM4F9luezQ4jmwm6eLhzwvKKbEmHbwFZ7fTqcy4Q9c4YYRlfD
b5dC2Wv6Gq5QIZZRuad1JuRbqp6NV7C7MsjHOZQz/++sIh3NDWsP0xDR2ENxmvXd
4MIjcbBnUAN1Y9N3EuTTNhUE4DbRn8r/Brx9hVY5NF26jVvl+NAaiO4lmh+YyD74
YTtVjMGMvanFrSOxDRgLGBcHV56+3+ud4ZlVloKcOJXdTM/YkBVGTUUjmJ5MSSzm
TYZzWo9Si2rselaJzHMCQWsw8cVHt3MQxvL8jzKQh7QoYDC4hmE597pN9c03Xnei
KkFIE03JhE0xo0mT3XgAQi+01ox4oFStza8qMvwfe8+RtXuybDIJBkAazV2lgLtD
p/5VidvIsOJTGRA7i8gO0SOxpf8ZzwPaf3T7XtA+k1upgdbiEIjtX23Qd9CZuiRi
tnZNb8Jvv50ZxHQRsaNFutXjRCbKMgxwEoe/47j3LX7QLRkSsxyrSYD1ciIDDlHJ
bEPDq8WNsc9++OQUBGhObikqezGJtZzI9QEoGL6bmjs9YDCpJExo8NZhVwwNJJLX
F4+k/kMMmRgnynNEv90FQDm1kQ7s6obUnrTgREj5z+04Mh89yTQITfyyKUmwOvIQ
OhdhSn5yB7923F6GcfQ+4tzo9hIEx/4xm6QrlzZ/iEGUCmVDfuh8TzXHb3kWSNko
whN1bJhij5R6LvFTjnfp2K73aP73WCUBia9py3xHzhHGLdPdRd3xJzeRb2+dl6RO
ylU/WkH1SBxZI6r+WUXKS2JCWJ3kmcRjinS8hAZNftQrh6aFL79fIPg/4Af9qj67
1w0enyLvI+7P4E6Lq6uoXizB8p2WljQ73CU9lRq/yg97Fe4We8cmlsOlNKhPFATd
5y0LuA68V5NPIVzVW8mJKcr7crYid/hXyxGjgz11OAQiTC9kfDVOCa/yEi9CwE7c
596QkRI71c0SzgnmRHFDgQ3DKkNU5NVNXRQKi3QolXVwgOitK/BL8SZ6D0Lr6FUX
JzmRwyFYSSEMGM5qGP9Vo6ys0ePKlOKRPX8q87bT7TYBiJNV+XQYYqi+AxylXivG
mu11GEsqMlod0SOPuvugHnHpZeIqp2b3BEIWg8/SEd6sWk2T15hrSz2eARepym1L
3KhtjICu6Kisc+MIJPc0tJmQJkibF4FStLwT+Tf+P/yFKHYld7qdQ/JGPcT+uE8I
V0OhMl5VcWLLOGdFVa7mV1rQ6E8m/xnWOFaubCBN8rnEdt7n7dL0llkCOggv/t7n
RUy3lApjYUyyg7vTQtF783Dj7I8zhzrGQIox027HjL65V7hK9ph49fEQyjRDsqaO
ierIlzrEsKat8UeVhf+mupXxftFljQFbZ9vMWqVzbslHyKbf/Eh4EHRc88OTUACh
/o+vl+iUsrhr3PLbjYmJC9KHK6Q3gp9SN5DTdNpUzmtAiTAjdmIhSrPHoc0AXK0a
4Qyl3ObJg4bZfhfGruICgkZ7BVgfOO99Ud72mOZsCIEycmUboa4KwcE6EOWs1ZzV
s0m8H+xhC7B7hK1iJhEjdUwHOLrhVzYjSrlBQdvuNbex2N8EZPFtF9ZluqOltuBh
ASz/Ue585Jw9vGUVHeswerYgpsJ3TZ8+6gNoh+oU/2aRm6Yk6q1ylPYRnrRtqoMO
SQysVgikBXUaE5MWkZtj9rT2VBmlhxoftBCrC6nyzKJQsVxuwfnD3JYVv9yLykbE
U+vL+IIezEPB4GizEDvnM85NcioH7//cC+yW0Im52mTyA7F+vRagGkrJuM9Q9gBQ
FP1pO7oYIou1PbrBOMAPmcIOV7y1jO9RV5GpKxmzjyiSjaFY5RefFK+IQw/8/xBg
X38WYQQA5dYofjxmrElxmDHyvoq3HoTXIFQmoOTCguo4T13QSYCoqrK3Qfk7JK72
H5FS8CDdX00qKEUiyJ9zsrI8OFP0NrmKMYwhW92zC3MjBB54q2CA2YB1T0zRakcy
viFMmYUdp6bbqJpZpQMpex55j0PlNqYn3FXR6fdMWx1gba+j6uUpVwf8lI0uHTc6
tYHZGuIk8KoX8RCNTPHlk4A5K5bj+0EI1dtIR57jvIWgzwsylxXDtdFLtEVNSkB+
QWfup2XpBCjOja2+Dozih2MLzYWZRWG+n64uLMxYqZ0DqqIYXymHyWFQRzq1AxEc
CdM2nKKJJBRZpecylHH05i8ZSGhj/N2/QwmwkBd2sC3fF/kkvi01Sn1DLNbFGbVy
VsyuWdInxa2UYsPhIg9JJLJdeHEB60+VXquyBPzkzuw3N/094c6vC9s8XfUO6EdS
rcM7zydBtezY0h2IPTNeR3TCV7/fSdVYoKEczuwWg4UDOfCIek6CSESsMdQuEXSU
3IGF5D38Z/WBpH9oteHdmqE1etvgSW/bmu8tW7adV4Cr/PLygt9+m1U2kkG2Q44m
x+CDWw7e4RqDhOr84AZlI5AKFLuTRovkr8IL2tTnj7iFDcpD5HUN6zVOUKBh72AB
v3MS/+WarHH1aPLVXw7qLZa+iVJ8SxszWd7DOj9xcZtevP+GDsMOKhq0ALHGtSgT
GZ9oMh/T25blC02xlMe8eTj3zJFpwO+267Fk4Z0vZeqcWT/CJORpxC+kfZk2qq7b
y8+du4RBI3kLDEoFIcECBPwnV2yOqp4lfcd1QN4HrTH+j+j5b449Y0HqdBcvxlco
ZSErW/72E70RVR2B6dBeUtHdHILSYtP+Y8T8RtLQ3M3my6ogmL6nVvzTJHNswq8O
2z0CLLC6iLYC7K/MbAvfjb7KXTmddKA2I0FOV8fTUN/PM6/9WZNWO0GlMH+IbTE/
Yzo03rE5gc53oq6U4dUvZKug4DkXqc49LbjkKKl28mqXXqEGkWGLF44Qux6NNSpK
FQXy9F8p+E+9CAd9Shr7KJS278SSmLhrq3TlL00BX9ZGodFQE0JCSDvpxHISYnv9
2X/o9YNMM+MQ43cLrk67caYdOe6BQndP3Wp8Wjr1X0X7Rl5PmTs9ULgvJ+9F6DCT
inVl3hBBA0MmVSjGvz8LBpepv+mCLDc0ryKQOMKL3HKBr4nGLRHxijiC8RTh1PWT
SipJIlbc3zZ3rc7EKXFDKHCM6sufi/M9m6JfsRBgN3gyP17XU4KPwVtbeZ+TMOWB
clhEjDJw+FtzrFHFq0nuH3wB5pNwYeLdHv7LK/g7DsE2rW4ErL7P4Kl5yu+b/CXU
hhWsmE27RnojrRKB0yxp5j3BxUI1lIY5EqQkAa/gykaH5JV5XfoR9RE1M/pLpzUn
fbDwzRHrcunWZ/KeuxIIKi2Riu9QH9c9A2nEKactvX+PROQGA/Ksokj2Gcg2LLGt
aDsQBW6X3i2nXALOLZrUyj7rWpTQj4x2qYA1XVcPseESBU3HPfrc9Hk0rOknjfUd
mm+OaIPcbuRxXGDdVy3Oy/TKF522CwItJNObjWGrnpJMkh5AZ6kUAQsYOqKZoSBb
DwrBvC5u4kLDOYFajeZ3v5SFKtI1zP32ZpxjfQBSE9QKSrcn7Uc0vHb99yMJ09KJ
75bwaJ3g+M0u1ym8J05B/jOqxbbRZK3t1jnNVjRNf/A/O9sG4v5UQYEKcR3rTjdT
tibyM2U3J0EOqyK6e0mWDYD9zB8e4XZ8sJm4bx7vvwpDkw389hN06uS3D7BKrcSy
1VVM+GCHmYShnIHCi4E+v5NH3YW1DJ8NWfRQgUmON3iBMQd700T4bp5c8GqL5cvH
B20bpY3CcSrvtuoWD0ZSe47YNQLofN3d3aoNSZWPuXIek/oObdnGebuudhnzWzzp
XAsOzQtjpAsKdLNfoiE0Ppr2uYdd2vMbQ11DCOUTcdXbpfxTjnmxxV6Z+/lXhgty
RaBa6CFYgqqXMdbVx/nmnnM+5JYnyFdgMvSUe5QUk/F30La373Jg9NXXOrg/CLPA
QJss+xIVOaaab4M0mlqrVm/RFuIn2aspW+zpysy+Wz9/BDHC+Ifv8LLMeobcQZKd
tgcHvk7N/nThy8fx8+11UKmnOjdP6kQBd5drlfFTgfr4SB76GGwQ36EZ0lNAs4Dy
ICReY1EjK7ywMp3afMB6MtZcSasiMgdYE0FonzEGgjjmJIjosO6m00mE8sF4RH69
dpxjfS8mMcGqvTqritjsCSCqcK4EuUkKxLRhSpqdKI1VKdnd/DfodHSxWk++ePRO
VBQH0+lrkI5CXCRmmbW3vFfh5K67T5/ROdzwbAkOdD0pLqHc/LVvmNYCJyi8AEA/
Ti918/jLk6RHNLok9OotfHbiE3hwj5yFJ/aYWscYNoNdb6pMqMDkuQmKWrNoHDZR
AJ5lDog5F9NndeUneS+H4SX1OqC+S2/LkXPQLI24v+o=
`pragma protect end_protected
