// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
szGM89be3C9lvv4XH0sV+Fltkm3Mq9mJz9aOXBgrk4eVIpCrhlMBIh+xtTBVqfwWP2g+j1DekxTF
MG93Tgifm6LpfvNsPHOBmpJGHKnrOP3MdyKHk65XvABl9a67nD0mF5/t3a+r7I5Y8h1xIGVJ6iLS
HNj3AS/qBNc/E9YAJVoEb0Tm7jfm9gtwuIRhYAlo/W4BDW9/d9aacoKQRCSpWvfPv/j7gt3At4jY
vVXZra7brkM6/ebOCTuXPCeF3A5BoBxSsNnKw08O7S0j0GYubiEPkUcDqHthrwI/D2inR6fvkakm
NwnDsVBfrXQgH1nvRGB38nmQ2fylvZReS+ITnw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 34352)
tWg4VR23K4eVPn6NE9JSwcDjzyNAGGL/86SOClwp4cL7x3O65f+Z+MqDr9IKONqTmjfEHbQIN7Z2
fwfSauP+yfshZFZwbdngU/eOUKUa/OGcOgBg3BQY9Ei9pmXMjktBAU3CTTPs+E/2ti/H6HFA7E4C
cbtDy0QCqeGb3foznqaot8JrqIAjzqhdW+pzzjH16nc3/e8FMk4Lsqmkfq2y24o7Oh8idys2K4JL
8NWZe/6vpMLo5HsfBTF9mv8tWrV7eryl2H68KINIc7pHun1KQ36fbUhX6CXpiaKPZFACeSC14COC
2fr1+3zTp/BVEBZ5x5VGO7YrbnveNcNt83AVciqHknvC8kJwFonc2124pld9LUGzQBKYDv8CSddd
btcFlNZFk11hFXF3FFhP+znQOJKh8rvdDA9+GvP+ioVuuPHKNEn3xj6LPz4uBS+AQQBUxmPfOluz
AIfX1N7Hv/cRvPJ+0gMoGOEEjKK1V3yx2RD1d8qepJ70NN99t7tnPlUI1a3wXi6lfj5gf/PQ/7zR
xYaYVidy9dHT7LQHmKV3g2Hff7koD1Z5/xqoWS1ic2q3Byk+atEGvkSASOCf5OUeEjHrNAmuBzvG
vAdqhEn1D29LR8fEgvXO0tBsKcFtD2NOj7lJM78BG9Rx4XY26R3EyWSSdabzzJAfsAQrt+GKYuAP
LBXsJKbsxYfIcYVZbV3Elyv6rnS49aZxCDW58IrJ9NLmQzjW/RM3+HUn8/Thr+11ThihuB6MCJPr
U0ySiq8rSCnso8xk11JScIc++j2EQ5tOU5DLLYnqB+E++b8rjgCcYWUCweCKNVBegkqb1GyCJFmw
BecOue3R9lEqDpFjB1RBH7WSGBJbimX8nEMl6qe+oI3eW59krzC7Fibuk6QT2CV8cPg5gmmk6b6E
Pu0/lEqYztVSEVPP4WWHjZ5tqRV/qob/SnpnZKiex+nzZrfHI6AcUC9C+R1cHjVOB1XLrFSqSSS0
fAzhVihA6kINs54LuhYW2oeSwXnqRzPHHZIOCgvaZJwXj9WPf6wcqMS0U3DlXL2lFkKqXdtdb3pb
VIaPUZ0VoKNtz6N3TdSKJ7B+JjSMun/y55Oohvv8Kojvo6ifk+2vH3RcZzt13IUavUxmJVRsFcg0
CjAnfqN58lXtMFggBNFvqDE+EozEMpfv7EOod35XNH2ShN9KShMztp9CJiFJ67G1JDrPt7k2bOqN
xpkeC0oejK/rb4fE0iOjsFiP9kvVXIR8SzGuFrQ/weLwolSlx7CHavltn/eV8xgx3iFQIJbksVWE
Z0N8ezgHGrhGY4qzHLW8M0ReegMc4f5oMEyD9Tbaao93chmkzknq/60Yvuz9QzDKQJDP6L219mXl
LwYGge6eQSHL029X4ArNntscZim+N/U86VMruLqDAhWng6HGDdURyFpyVxS5QDrfOfFq9NdKoH7R
O7QHobRqmEOsKuxQwbXClA1nK6wiT2iTI30MoolI8y+VunG8ZQveeMA/p3DUN4Ss2YYvGZDBdLvp
swoE3p/qD780OJpP2+vdMLlk6AIx47oOoB1a/69Wx65qz2zth5DnPAb6hrA7PqqrIHLdT+KVxDb3
NdKBSDHUa7xQ6z92o41urqbXPgXBGyR5qbznbgOlKfOBWliakYLhPBDffd4EqERzBiL3yVM6h5T9
zZscBqH6F2qHnbKKESSf2jg1qxMpioLxr1+DQt9/88FDAOlDCi/KKKNSIQVeQGGbsXzjc/1hepxU
Yp/7H+S6mPH3sa7LIObXofEDYiNgvnXuBU8jPgAp9WF5lGFufzeAvP7LyDIArMA+cryI4BLMRxu1
AMnRm7KSvEJWr9ue1flE9ugy3+gnRxZV7oD9ZfpuRc8EUXN/EU9Fu1q/GueUivEvFYFU8le0RHYu
DKZWRaah+Oj8xLk6SFw6Fw+wNJD05smh8BWscA8oUPmGDrymXOn4OeTsyqdDSkQUYo85ZQjcBTS0
bb/iUq7Xczh6iTHPlRmYyjnZ0mq02OBgP9uq+zq/ZGRjY0wN49McSoty4z64Rdmr09gQ3fama2gE
qFRjXsFEFypkjDcQujQURAVaTBIX0PaGvlect24WN53el3mrWlTDO7liM9USYG/gLHsyXw88m1iQ
5Zz2Bdm+9krvObf8tfrCIfDUxnjtJg8qUCODqI2P0/waaHAKoLafULFe8IO0G0ySytI2tZdiYflh
RUNHKMb0bQNz8Y4YOOtLra/JvygW+C5RihmOtzMjN/IrfRSlk5Se5K+MBVT9+7qeHw23ZmM2NSRe
gyktPTimicJ872t3qUgZd3C01lEKwV7DRL0MOZ2GlQr9apiPqR9c1OHOU4QfpV7yyDp0nvW/Sk0n
9jJvZP0Fqjq3oXiTkPtTI0QGpzB9eMjwsXehZS6K7BS+FUc+fIb6Wl4+loPZKXZzkljXAUqUrQcJ
eucn+DHatOFexhCxXgMNUQ0sbnZl+oS7iTZDYejbqu22bdKF1lwwVlczwEI+iG3/4aZLeQkeg0QE
gsZtgGXA1TQkp40QB7KpsQDPFXDtuv4IKxfG8bwsgJcU6SLPTP0q5ff4GpH1snPoc9QWEBGN1bHn
CdJ+2hkiUeETW+3WUAxSrJ/X2Y+Ifp34QQn532KhLh/F8+WdrujJ/W+4lMaLUNRzu0cppt+he5Bu
d3ISBfcVgmnDr+w/DP/qLvhB+AISHxwXkK54WgRm1R7vk2U0vHS83JoL6jo2F+Z/i/Ef8RCCpDLZ
JD3lr0xTXYrEXtjkWBkYyAyPzD2cE7kipJW/eVlhWYkg92PcrzVsFoNiIfm01LQ+pT/+j++0BuEx
fN8A/XSgGMnB9QnEyxfwPr1b6FgzjjAvP6TThnuG1f+XOUsPAyx0donthcygcn+8NYIJ75s+Zy6q
Ofi0jZHAea6bNvDyzELlXl8XZTOqOMFzIwZmhnm22xMOfg5hevkY1JPoa22I2h5OWUAUDkBsf5nW
I5gYwOk75Fv5Dy422AhKoOTwRyFkyBE19Hmwa3lays967U0CEYIqkTodl4QurQ0u/l0RPlY4hJn2
Luf4zuBlBSUkWV8yO0TkT2fXdVJb1n0M5dRkLi0aWZuT3b40qvyLRiN1OSCk88tFk4gg63hxMA1Y
bFO2lm/cwfYw4CcXqBopdXA4YSga6MBhd5QEJS+XqgT5qM4XDK3i6JwbTIgr9elrsnEqER+Sks8+
OCZA4oWO38XzUrxz+Nof8Z3hLAhwnnTtYFNuMXPTpg7h8fVFxhha8LYIZ9IF2Y5dhq6C4yg1hZC1
lBO+lElTyVibawaF6+WQJU7+4DzdUhJ+Wym5xP+uRPZXIbZ6yL0IRd1nBjz3NLEKANLMq5rckx+F
J+LJt2YEkU7YS8a2hG2qzw6qB/7PWQwYkAAgx9sJq3p8l/NNWiGeqtOxkJBhwOfbYJC8jW4oL5BF
DyvJ1KZIX2KRTDF89oL8Lns7rtR4dVejlpLeLcb7VbMrXsaVdm/KKG57xhzQCPQGpRsjTvfjiq8e
HAjP0Daaiqkliy+A5Aq8OAG56K621kGf0CPX6KBGbEoGvjp0WANWqtWtZKv8cVs+DnmENb6fmPn/
r60PhQ8a3qZbJY4+9nNIVrnieNmkpF5nII2bcDlxOAQF2qWHpItTrRAgpkD/SI6yC+kiIEKmY/6F
LfvhclkV6HwhZ7aGr1V2fmOkxqySYkPmEGStCyn9kQfrWToCiAFsF1gtX8cz6YDGmrHFyvjCT5P8
GItoGIqZY2mutYNuJEgDJHLfSGVvVoKYllAve29hkAsYhhz1OfYmHI7q9rXNzLWjAB7krI+0uXNz
PidAExj0RYTTY6y15S8Sx7N75D8uKPxk7M7x7UO6X6qoXp0PUGnxuCBqjgyjFInWaaZwovDe6hzh
NU+cQRQ8TU1IAMbubbJjq6VWPz6MRKJPIbw1Tadpmtplc6tm22/3KuXulLwdWR3TZvw4rqQzNql1
B9IMzEOqIg5nQfUGvcYksHsbu1bF2fY3TfBvn09WpD2CMDXSrzerkWOINGawDETl8K88PPNmw5jr
a3oZbE+tSbeG64kGfmUSiCkXj2+blgr0lgdLJrZl+nEcgUIVaq1TD627/gnWmyj9pG1XfqakktkW
40g5KHnQ7ly2KdIdF4etJfHCk7scaWGjByOwzrVwPWu7zjY5+YXUfdI/GVKfYoimf4tuuaN5Epui
0ugmlhRVp51kBs3VFKUT9buH5yoIbeHunR5KEGfKkz/IsvQCpveVrrEwkXoO3QLWqtfgkKmobqnI
8mULuvhKuLZmGOWZ2D1APe51K+g33sBn032q34Z/4se4uRHsMiO7Zijy4+Sl3dCW3FqkTvDiE+Iw
5+r0ibHo8kw9DWmb10JdEIaAvb/cZ64hiSVh+qM8/J+IUTUvTnjIMT9+mAbOUwUJXHK5ZxelZ0xJ
cAM028Y9pZ2Vu26FT84+o03QKF6+GlimwZKC4uawkTq5Zs7HBUYB/MQJDwUDntQWRk27Q9xPgPul
lXU8pc3fWMACy/gjdDX0YFZCk/gmPJ/OsRwn0XerGKGw9oPv5M76hy3TRSeLq9gD3KvyogUCcNqv
b15gnTwDWD+m+8r+ir7Su1paTNfOutWgegFNB8WxWE0gq8oQYyggANUYns8dARP6WcPQkEG8Wjq8
FS9MADi+c6jDIrr7Z/NFJwq54x0T1P4vFevL/9qi8lJkayeil8AMwm1etSHmUp7yu06HHLLi+J8E
Xqq4u3tQ2PLaeyu1Fcdl82KQ5N+jWKqObvt4j/rfiyGVYMyfbsOtCoMovQ728/Z1ywFTU1+GWxAj
JXhbuSFcAcWTa9uhitwlCfP/5juyA4Q0oifWqvVTUpbFZGBiywFV+g99OrLjrS9WQ2QUKRi0K6t2
hefOxmkNp0i2pgGRUn7J79jxgHcYPbH4f3tr6GyxQy7DC0BpzQtLBm6XBiMLkEuxXRblgVwLWee1
lgkWz0WXwNfGTuFtcHOiiIN/bO3jByihN20hCwP1o935iCzg16g0gc9RmxDhywstjFmQpz3VM/Pv
cUKlKD8O/PgbkPjEtw3aUH9pbIjqXaVPY+Y4uz5AF5vL5uLadqNMtAkDLV8G5ztqexi3f34GfozX
hgOgJUslqujCdSfXOdlGj2y20EX6ORdJAooe39uP7+oox9zNKIML+nSeyoyWhuexncfZaTxlmJfc
DZR7ZGNTG5suTzZ1Q4/X/QrvCePHsh5wsatMuaEoExVo3PpVaEUcx8QaG5Ei3xx0WjyxoVYgk49x
qnZg4Ut6lGeOcvPLrx7r/ehT5P/k+ODMWGpEjmAIE24ZMhc7s3MWy+Xgs8ACV1h+iuDqjutknQbj
XP0qGVkO0H7t+YJla0uLkDZdBKQgv0RlxhHUp0CtbhQMyG3379LQskivBPWZx6xfAvCYqn/sl6YH
CZPbaPUkV5vvQyT6GOP2w5nGa5VP3BwbgofhfNgkruZ9gQKikHymVzKYy5T8yXSsCexSlT2Ningh
+Bu3IKZX070u75hAcauqjT1JEhaz6wlCp2Fcpyt9Duzj/GDM7oXa0tjioqyrWqkUpBQsBFB5jFEi
fu61visKXpgp5L77QU7xgJKlgWE6n7axokJc0lZjPtP3bS+wju+wL5yBVHPwjqeAlNQIBO0WI6ji
Qm3wmbWTZB8TeBkSqFlLpJLz020eyUIt80gu9JzvOk6dJiuVisY7tohHmwNXRG/USVAklEIpJLko
QOzRW4gjjTMcHob1fS/DwfWRk6YQfpxpENw4SQOWhINNgNyIbHanpbx+oLFBQR0EAALmTBYuFPL2
YyYSdSFDuBujAiLOzNtDTwwCzmr+FbzuVE76enWENMCAA17Ro/WOzy/u0zZsh06CDlkQA7Gt650d
JgjGE5FIsF0Jwt5v1TsJMYwcWYQ9JPwqtqW0dEuwffYwPAcnRjLa3vAtlbVIO5aLJtby2YVjsowO
0gFE6cixO36WG4dwp/lVvrOmQqYGVcwY/nRuIxUJiZJC+bJhIc5Ylmrts1GPEnpi26UUzEQDS0gD
l79TgrgSAQYGssZA1TJ+ZLOml4n5HrdJVaWXhWMeDzkhyuD9g9+OxDtdz3z4TV24sW98uzy1e1Dx
98MrmyEBK84djXH5z0dzjzF9qP5cSlq4U//j9W/tVD50H3Vmco8l6NCPHb4GKZ4dxnm5G2UrrhQy
kr68FxyCj8GZilKdXw4zCJ91uH9Qxz6bq3aaB7YC/Za0w14jjBeMzbnkLpd0QuBrTb1f7T+IQ/wW
DW4o2QUxXjxZ8W/jb0aOhWyicEOhQJ1j/AOHOyvzYVLYoxd8ZEi/jHjLhnBfo+iSd6Oa4rxaI7E1
SGVsEDX+Dtcg3un4wxRNwLVsqt1nd/BWxiALA+m4Qku5CgVOigWvxMiDqEd7ua+0HUXAyoLle4Dn
Cg21CfUcsDW1NpVJxmyI6h9wSoIY5X277Wdi8U6iTKcPdixtfNQ7BOLruTLKL9zV1Ndz/4eenUGV
7QlQvWvZRpcqDNXbBYdCdo7tuKOTl6cQ6dr+8Jwl/3pejwTl8bKFOBB0ZchVQpdt4GW90IgVZEFZ
6uayGlcHKOQSFLTyVj+WVFQjDwnY9Yzfcy7TXvMyCi1jLeUpEMOXxqgH4vbboEtvRKuYIVBKRn/b
HXF3w7/swtJVCH25QUajk0Bfa6rY4fFVwXqC1jdO/DYq86vtWkgf9g3PmmWNGzLR8ToBjjzpQNAZ
sX5eE9A4teptWR13DOFlZBbKlMve/onkNmSIjK/YqYQoHnAVk2T/k+GCzgPJzu9eKlFPCVQ35ACy
jj90CGnI0v4cMcalKYrGgcrgFk/5WbuMcBVI/TbJvKhX3r51Xy4Tk3UqzSjqctwQDilDF+3G5+j8
GGPDZYGMaB5StiqsBR92KJOsXMfDzmTfNxeFjJZBDNx8UxmuljuSSzXkleE4ohjvnO9SbuE6Gw4K
bRyQgJGuBNZ3J+swdITi6fQwNORIF6vU0EVEiSNuKX+8qx2v3M+kYCY9TfiVw58NyJIL0IYTSj+5
e6JHChUMLquS0EWQaqVjQ8uAzM34FDwOVWywXi08VX4boPIf8IXwMYGjiHVdIZENrUuzU7e+wI1l
h6ElEHAw60IGSx+WQJ6mM+Mq3LaTH6SN4eHW0aciz9JQpZTinmRAzaWvyB3/+NOF2WjhMU+ME38A
hEQ7Fx9qJKff8ZT5BDj7O8HdyMiUGmhE3Jjv5sSldho38FvWFp9BCIbEftsgrvDZQ+9OVXsirGf1
X4jmEMSyElJeFn8B5tylT0wF8D3yCv4XuWSZKWRrKSOm1wgAZsvZjBMqMGG6BqTmbG8isQQXPDDg
Xy7v3M+P+qr14BrqCvIk1cu5kufSHQTeQqlBUKRliae2A0Wc/B3iVmVPsz9EGlisnzXG9V+tXVgo
azW2rPwAMWk4x/bJDGGX2hXbh9NejymKHGlwqz4i4Mqigtbr3n/lRfv+t0pkPZ9MK6PHl7sZP2sI
hfkJG8nrUNZII3qnfOm5p4TuC7A5bRamVnJJmIIDUzdQX7PkymirKJo4QXS2OsEsCC1PoRo0HDJb
rGBadluykefPitW1yT+BiKZ9NDoH56Oxdcd56XXqe90zWqiub5qv/X4EGopmuHTRVLFdvFa2WNDR
MYpRit9HJQ4dq3D2uI3kpQorNllJYYX4uFks4Ssx6lxCamQU4XtMTPdWtPOf0jVCmsFBdPP+/umO
cYTgnMnHQmOb/NAlfr67dhhwkeIFz4kgnLBj5IQrkSQb2QC/wRSlFjD68i/eIDhHhtV8JHm/71qj
ur0CWWeYnaYyi2DE3CwxfacwLFq4MF9Sq6gNdRRS/zzItlmRzz6MOIm4+tDHkkg80FQGezbZEbVI
0+cQf5G5E+TA+ZK1wA8M/pweMdPgvJoDzz43Go5dhSkeMbvvrYQRtHL9ixAmE1wITvfFHzBNkpGj
7foekP821OtHVSGF4R38kNybb+LqyxBVQnLPJYkSaaMREuxV5GC52hkJiDsbGOasST6EzJF8xtNW
/7A7ws3SrXy1fVOfUI302rMT42aNsaQYBZAehgNTDWYFdylEPH/8wPvFdKoLTi5XnHUnSCKIgD4f
EbTUaYEq7cfZUZoCfvUr8vZvwi7yhlj8rJ9rvBf4GBASSAjPrSf2tBm1Qss1LEgh/I1VLEzBhuTJ
pyWQqO7sL5BroeY6BQhdejhaxsp4mzuAAkp4xu4FFxD0SARPak6NmDmlRB5D0p+XRfC3DEaLWxV5
eyEq9DEsT7Q54nSyp7nJAK02OKYgmMa192Gt2zFATiTvjMVNvaPJ2a+3cZ3lVd0B0kbQQ5ZCjnbu
gPaBC8TErmUIMhDdZUfOA/WVeSzitVbqXo8I1Rzrk2PLPQcFjo7F+gHcJfgc7obH9OK9VQcN8Y/7
TVrfzgL3AsrB+FNtNFj2bokTf/lvXONOyN2IjbtcMx2WHf4YeRK74sK+iKmW8IFDPFQE49GhhLq+
TDnclMUeFIDyy2q5wrZsV6ey1Fhxcg2MEDA5HBJnrQNWEDk/0QzXQVDO2yUUf+fiVpjOV7GzAfPt
5qI6xlHwKO+X5e3Xcln0UUHYHXoEThSbkAquwEgmwlycptcBjlzWrfauW8eu+Vrf8g9F+YJEtMrD
gge2uuruENLCFPHDaHi28ogjprlw5AS01qldYY9TwihvimL96sSD18wu0TYGGlNTTV/Hm5zFJ8ah
2YOueyV2LLOex7s/Ncvh+Pxoh3S2RjBeTNC/V5KLCr6Dh6dWFJljKcPbB2+JR2pEpwSvv8IqBHY2
VYv+ZQnUh2lYhWRt4xKAfRd4b4T7jPqSetpFITLwJnRDA2ErGcewrIz7/SEvuPMFYro34ZOqdZeH
wUvhMUxemRvDOJHvJLyGNL6uyKXjt3ktKQP/FAHhrI4K4sIyrW30+od02FUkP1udpegXRRlu7EwO
S0xOt0CAcwx4REz3mKBI3VOl3iFcaM/0YHVP0h7lXsYwRG3v2PGyUBViYQnzz6nLlwPe1MPsWATs
A2xcXKu5fsojisT6ts0i8MupAnp3Y0y+YqvUe4zlhLcpexIa2FeMkkHlkJtLoRgzM0o/wN0HyX9p
mDf7T26fgXfawqD3Hfk0piQKGTy0tJnPS1O4RHmNld1xOI+D8T/6oqDbhw5GF7vq3zXplN+PatG+
oNwpqUiALM3s7hKsI3XPx7Xb95ry968nKM61EZcOR049yW7RJMXYnShSXyV4Xk3ljRTe8Fgr6R/2
wji6yglBiPjvSqpDcvdd86AUCJKi4syKzkwFERnGpqHgqc4DPbOY1qfu48iJNa3lN8RG4BkJP5Ek
ETcv42SqR8QfO6njFXgrLyEAMhI3NLCTEe8VEx/u6kqf2OucY45JaKY/dPvC0Rp4ANqNpLPJqoMf
eYdp7iC2AyFgVG8v4ZP2w5YvH8yH8SpX6z2Hw9fwxOYKJYo4zVJIjosMhrIw59V10jIAlvQFftyv
V/IQwoomn8RCM23n1JP+55I7jgddqscjYdZM2b5SsFo4x8nX2SjPL0mqQGoysKDepcz9cyhVnWT8
NTQ6CNMnY8HWtT5YYU9r4im98I7qBrgfU/4pX8isigtpv32AH03EErFQqRJWsOIGjmJLCdS3e29g
Bdd1EjJGiRDXz66Uzv/sAucfVxiqn2GQ2PYSnUnvS2t/udBYcuC5z61qom1x8Q5kf5ZEKlV7vZBy
srouVhO+xBLY3Hy6esMx0e/lI+cS1mSoShk6YXof23mw2QqUYYkknESJcLzTe74+WYVozSRAzHC+
HimQWrZRn7mRUCnURxgRQKoJDPdlDYVYILBE9FA7+xHoedUQWrkzbhMfCNUwhgtG28CClCMShg2Z
H6VXN1DhGL0XXapEkjrPXprrfvKI7WSR6AHUUaIn7q+NWfWmJ/F9wuQzKLnS28xcNUd8XoS++GO3
QvONc91sQfizmd+UvVwTVjNup46zs4AQasxiqDmvgO133HTzr4YCx2QkyVFdPis7Ln3Rdz9sU39T
aBRrpgOW7yU3JkQgVlTPTkEldmGKZw+I5m7tervpJLf6LDbLF0A/Ik/sqRYZ+OyBjhfFzkQMLMLo
rUOETwFA2IzpKdNNsgtMktFEng7kLqrOTa78LhBYxBaFTj+BhJVUDQgvUf8KZ55pVwxkpIrQjyb6
3jmqjnKKHoeinxsM0sNOHz0kkNF38HT+FSRS9u5zoUv7W2/3gtanBvjIDvCXzPrOS3nTvX4za6G8
DaMpIqedefewAgOZcAF3muVwAnY31IcMBoZGCS4j7vlJbLVqPwaDy4W8HQ/Hf7+26/4CqJ67ng+Q
uaVWret6ch6DFblJfZHZ0BSzKyfV714FL95uHTvqnFSntU9R903ThWBxVAzpaC4mkox7jbt6Ja3U
5ltLJP+Lc4iBRz5UzY7cPOcj0DwzEAN4uSuNjQK3+MZLKH6CeDmSzw8HtW2mRdqKS60A5I3qXB5c
xliH0Lk1L8zowH4B82ddtz/XraScT8ukNoS4aFwvHakbSn3YeGlO+xZ9hzdPAaPxt4156+LzfWP9
kCU4KfSqSXIXIHvlju3nyOlVd1KCf41orGUVLFoNhB5rsxHonofGKz9F+IxxL0dQtHza01oaTBzx
43sFmLf7++QULO8zjyOHXQXqfcjmUNWiFJD2hPbGedX045kikKQ7h8DriDSoniWq3QvlSZGieN/9
aYAk2+AjmU8vv8Q3O8Rvo6dU3DIIkXWwErPXWBYkFbVi57r/vzZsgWVpJkb4XW3Kjio6aPpZ/teH
UoYWg4KICLRCN+QPdQpKOAs7vmsGZ8kKf5ryr8lD712ED82ZwzhnJTg+LgaaCH9wEiJ7Ji1t70V0
fWUGutB2mwNHVl2PfC9UbIqYWkCtXXuln7oIDg+zFkfGvsJofM69higU507zRRjcAm75nqozCQSK
on709e+pUTUllSols6Ho9D/YF9OHc2Ot/Gp55qmZgkX9oCyA62Mt667tGthduKu2PCddwhC3UEgT
larNawXtUo6QU3VtNYNqbCQG0hoYzKVQIxlIXE49LLEeQWDaa4u357l4cnskVQUTNFt3O/YOm4kS
oaa+sDHF4Jzhe43bZWJo/ICcGzaXo5yFLBNMNHc+Vn5OHF9Cy0fv2mlIrc9zGdjOrntScJ4gbom+
QKHc0uQcjCWWxH9BRAsSgCfKeoPFwe6QZBZXIiDog8VcM5oBGIrSgMVubqOtApPRoTR93JplWZPf
Z0h2kwd5pxYGEGAzastfnNHSsNVnq0/bGsfxeuWzLuGBkJjwQGKmTFLBU1Vz38z95ukMBwfh9YE3
gBwXYXG4fAmt1Fci8NtCTGII8paH9oQD14WS637z4e0ulZKovmmFZ0s3PTMZS0/FuUdpctOpGZBy
EVYLFsQ1PAW1gO5k2klpr8vWvSk8sHja2bMHj0A0GyeRsm77ONH9hd+yRpUjxXFGNYA7j+DQ3xlI
9vNK4kvlDBuH4exqIsjwaZ3eYLusoKI+kKDXAramXQTtKCdomf/Ta3tEC9c5ArZX2H58ujusK/wx
8U6zqltWVC+Xnj50UcdwGXFhXTG+L+c4xTL2Gx1pUWEOX9E9yDStkADvCNYK5NRgItXysWLrgdpV
6vDs+7POD1TI/eCuyp6+6XsHtlOCRKpdMXIJXK4ux8NjJZWvY7c9vtZf0uIutMBPXR543uZ2CGJE
68OW9c4V3uwYHyNtfJHUj9hSJBCAPbFFJK3Y9q51AjsQ5pdjxS4jMeERHEeVAvGf1HO1rXA3IJl9
lkuCgG6on66fmu+PwdpsJS27qIzKru+hgbMxCiMuu+aVYh/xbgGAPk/n5JJkmF0EVZ1iYl5d0Owx
V1mEtWdCqJXd1gxG4SeH6iCpFOW6mRge7rnzHpp3MQb1wqNfxqFbcrPpj9jajUygf4AEYCYo0eft
D+mWtukF8DfbzKn2Zy2yNTHJotfvyAMrY90VuKBSmCKQJjl5OipnhXagSPy00JGwl1dsd4NFR3XO
F2OEZJTPu6j/49o3SYipJMzxGE3VKWXr4zsYgkz3iHQF03gPIeZSWraXc6egswMjiYAjJjlHVGdx
wC8uZvUo7PIyrUAa4Z5XSH1+eZEUpsG+Gfpv9I8rJctXqxF2eUO6rezmZQ1elKD2xwyiqRMsUigm
L4RMPko6Aj0b3eBb6X4I2UQ+1dhQitSLbeunGAGsWabezJb2CiS60oa/hzvDK+3g7Uuik0mMhFx5
U0Q6LeJKkFaLo68+JwSsJ5M1AJsLcanGYINgTa5FuMx44NBD+zmtJWcN+64g2x4EzHjI56d0UTt1
0xyZrbhB0BYL09bQYEDiXeF0hcLFqP3X+y7CDtwim4zJMl8OUbLKIyEZ0wRxFkk/hixrNkBZ3COP
ew4UO0rvufVQwfImkdCNdZKt7xXPC9ISRDYUNdospsZnvdj4S2FVjulpb/lRpLF1MVWuxkZa4c6b
46z5BSEeMn9QYjt9UOF8epI2Zeb3Y0J2rCBqy/qEkIiDRoSZ3TCyD6kAxqmZVtxp/IQIT1n88494
iWoZKEXzCAMoUCl87idnDxzMJCWG4JeM6GIXUd40XVDK5YWzzWCHHt0BGCF6CtSwmPpP4H5jYy99
phMofAi7eHHJB92ooCpBcPLAjxCtlK5N8K+UsFrHtlO1dajk6jgoiMEVvQoTeYB9Tz/Tw8uskaQd
e1riQS1tjSehSaeQk1fw4qY6/Y0SUR3bL6XQ9kOi9w67MLPMggcjyICQFJSYXEr9OXO8VDj/Pt84
7UQbtY4WnqPtIUjPme0RF7qMbJa3DPeR4Dv7iODXOutA+rwbW1FD9DAI9bQigOmduKBQAoniTWxG
0Ai6acunwx4r4yp5aEaEeERnB/xg6ftB3cdbEG8lzsd5LXt5iKWfHzxZqcYkDLOH4a3js0RtEWIs
6jTXPuGB0aViSmdXtNJtkkVs5xAW1Pji1xm2B4MmRyvSA1JMfCpRDsdeYk/7iX3pBhy/nx/88YUW
HAEkh0U/2kWNJoVElnnB6d2B5eL8zhHsxVQQx3QbB1Wf2XSCwbueGJNvSFDNl3cJrTqxvRKr9zL9
5QQOyVfB8SlrvtJKYsG6GGKAJjJyaryuhOU1YFAJyKKzqRYsYRC+dkdTbFjEqqDwj3+GbsHQhRUP
o9/Js2VjCCINcH/5RWeV8X1GPEAXUvTvyOrXNg9x0a+KJIW6fPaEFa0RKGzBnABkks+c7jyPCw9g
rAR/AYCGi8Q8G7sdQgOkSRUg7O6eJx85a7phCFP2d7ZOYnHZGkq3Ezb4OivyMHxjy38cssWFxdPX
vnodbi80R+macc/vmbBrA/jwmcz2gEvER8flpnMB7HWRGNKCcVa2P2mF8R/z52Mh3ul6fh7c/9VK
gN2oMfUuzjkpM0Yg0UKflFP/f1V/rCh3nrrItPpcQkFMOIVK4emBWYQcBU8+h51FFSkzRJ8simgf
zqIx8TPlA2rN6IYEpHsW8MWjvzhTO25ARQ7KEYELh2qYYiRQP3Ow026I7scCod2Q/EuXe/djp/4M
ZlEBZ0XS5XzpzJMkK3LAY7M/AKd0Xf3Jmz+KwWUjCOxCrlNhisPhKb64AoQxpnDl3RJxP7Tq8nko
ws8L+Ty7ClmZcpsB8SNHcHZ1mIIjckUJYhp+ACC/4xOU9xv2gT0k0AADzAV5PY0H5skNfJQlOhCN
VQbWgwdQLle7JO5UND8i9YE72J12ePZjIfTPU5QXN1JWJTrUVxhhnm/weNSAajOK6PSOWB5gNlyc
4JpjBBb8ex44loST4kmvgUHZEMWB3onPHY1QL3vFVsBDldJGsp05pUCCSjZAnG5O1e9JX6F6k3jx
1GKDG6FpAx3FjrzUYg8Et66l5UZwkB1+bHeMgkIdpI4whUx/30+2Ja06CprBYVdQtqMvwd3cTGgN
qMCNgcOHkPr48wLVAvsu4W1F9fUTEzbg8TLZFSxg0dnh8DwNp7tGBa4SqYu0u7GGKAiSYc+Xziuq
yNvz5MsmCuMNCDNzBZRvnd79SfB55eXVI2VCMqMSvI93/8rVY2rHoEmm9tIWfhKZuRAvsnLdy8/B
FylivW+P17Z3pa2DfIXZHi6bmotkOtXy1rcYKDj43pbScej6xZPG4mWyj/K4ghlcMQ+WnaBpF3CG
I38dL2pv05EiH0u21hSaYYgj6aDapimWI9cLL3YgR/uNYGCsExjZzkkGCOs8P7kqF0etgyTm2PJs
jBXNW+Yybr9tiwn9ZXl5suB1gkSSeJSABxxjiTq9drt5db2IH2P516+1Uf14ieBscc6kf2xJF+QV
t7spLzaeNWFbMxRkGXTcv8TTgrHl2p4EPG0OuN8IMCIPdAHX6thNPzAT/y2TN+EWKmqWV+0ixj4D
R1Qcze1R4vX1cAV0Osqj9lqoRfc14XhhPdTu2fN4KomRTOQ52wktUfnlu+PQEqtsFDjusvZfzUWr
h7mhu0OerLqen0MQTd0vjvFwL28j46orWnhEyzRyRCXhyhpTQbPWdZodw/pTbBzpfwkqi9C6IDt6
qGoTpwI9Z/MucDYHx+ChSiQf2ELtxQcvXEo3AtklJozyeKUMA91akMG+wmMhnV8jgX7PiEyIzGHT
LFe0YlDxztc+h6gi69KVQ704K4hjH+3P5QHOA8znR5bA8qOBfPKb9kYO2V98c7LG31fFpMvBssup
OecP8MYRa9QKPKtitLhehq6ASCk/07B5eUGf04GmXYwGok+Pq5tZbI7gMrXL5aFKjlX08F7dLLqL
P/6iPq3b7gd218PvE1W7QkWOpchlucxyNjM/hX1VsUo4/ujERh+x3v+hr1kVqdWViqLOFM/Cn48z
cs5kvcK9oQP7FXhlGH7ZiXT/7JmTfcSpqKb28OlEiGQjP4UW3dz6zj/l7p08u/HHJjHK+L8ss4VG
q0ckO+SLkzYF7C8aAHpwJ8VopuEnsGXfGXiVGd5OUPVp2JRwTlV6diN3wdUWN1w+nrTPUr/DdhQY
610KvjkyUDaUvQt+NwgF2jPFBzLFbrrhfoi+AiA1/D7zwGHHfE1rY/Vo/4bX5hiGdNWveiscEqaO
R2JY4GQomZcrGwhez6hLDiSgUrJPdTM43g7bcUDKmFX9ez6NJPEcjO/M3BkMXMANM5nk5WKrLonO
zjMma5UTocadJ2HXD0D6L72SoTG/0XQkw69PP/cQ7Gkr8PtlDainSVIa+Jya0EVsVvIaCIOkPopX
qaNrWaOTaCGhYzfmFzJOo6pdjn1U59ockloUaI+P/cl053NaRA4yzGopzOU7+srMO3XQwHtbf5Gb
KJ0plCKoei0LQfRMkygpDwcmAdmbJs/rzbR9K547XZ16AAyzHROo5cc9it9FFTSBJtx1D9gSeWgj
CoKQgeCgKTpS8gU2pJNv1P59csnfIsl1uJyLfMpBAZlGwq+eeGumLKswlI0TbV7IuVOw5qxeyhqX
K2bNmeFFJ6/n8T/OYszl0BpF9EFcX3TBo/FM21VroeNxI9BaEMIJbwEQ8gqEUu6fcztalT7OsDoD
mY37MArhcNwfOHqahSnP9BdZw3Ivno11LUauLYsE27c7bA+aANG/J3pJNr9WwHEOa4XC0pAmqIEb
YQP9GSZtvy0JEe9iZP47aB7yahxu9lOIBAbaf8713pzDEH/T91/Orn5C5GRu+BLmvMQxAkfYPvLJ
NTLlGZke1jyb+5/l3DsLY/cg1ZHM7wAVqWhYwfSNepxJ0v+UgXI+la03OvhRvBhv0ew1TMV8K4xm
a2+m9J/nTYVRsvz8ZLdtcBFB/keaLFFudhjXfy4gfRDpmVRzwveOyf+wQcDxVKqhlJT0f9O9DbJH
LdOrKM+fwQ5sNsNp2nwTKkTSBpMSWrIiPFZu//9c7FvGpJ43o4WMp3U88fxGleJ48riCm/xJpr30
D0GZNTYCjyW6Y/j79+IVi4wWsYUn4flWtwIbKszQViQvTwcmn4ahT9o85Mw7az2+G8mEQHcjTIbp
WCe+oosHubs3kWkikAadJ/GZlckVmaETGnW+acFpKmWSnYLwI8f/7BX81OeqKxoQ+cmrmtVeM5z2
Vwi3SCa+TGc4lI5VA/RvBYZ4fJbJRLzsizpCgQUBa4OG2L61I73NQFt1VBEGj5K7i9xYFwEjusNw
1iWL5ANuCYn2ZG9kHc4mrc+PEeMih2o3Y6enn14a+WMGGlIl+ZQnPD58p5OwGmQ/heTRJTBlXepq
nPJfq+Uxt2hHhgt/yqEAummKSNgnp8Nvun47KZaCXgrvKetORlxNCKFKFd3KYlQ+k8G4kzSTU+5z
uw06VWzw7xD/gBdLWKfUjK8u0W0MXqwAZNzoWb8IdpHDi8jJsJxbAl5LuBdDXLSbuK2+TcN88WZJ
mdRCSZN08sJHX+c1m++bahvRNfSm7xLVuCcaBilSOGXJfhRC0BKH+isFbiq2sMbOPuAL1R08Upec
iEmIEbvE8Jj0d4J4ymVgczUH2neq7dbBr637fWEqqtfKEXZZBCDS1UIepA7uddP9tnp/JJqSmbCn
9SNN/2zrfMp6Jz4dqOVOMERp9G55AmSye8pUlinLKQVajirQ5+cIlm4TZ2uYog6zGOXvkpdurXFW
tj/Fs3AHG97cwXFGI0OAiwaukniaTZ38P1TbMROOGb04XCRTlZpgKUgHgJXkUnlpECShreU2NwJf
iQwglkWWRlzeU5tqZJUAWK5SwvivUZK+WV0wG7PZIZYF61ImvWFrxthOkQ76I7fHkFngHrl8WvSX
NgSigY1lIrFLLD8ltq+7ZkMF30BSMSnRsWvK78GK/KUbHpmeyk+dQ0a83+h1YBk2Zr0+YvgLdLpj
pqBBTv4ura++ErvnI4idWRIFUcS9YsBcFRswwcyFL0oX3zKCKWxsvIaOYurc+d9Q3v+zZGWKN/i9
aqQ98ppEKzdZG44KsZDAHGLgsekUmiNZLNldKm1Qiv4Yt/s7/CwwITflUkrcULBN800iYUzOL6U9
zKMu3Z51tCC4bLwfhBW4IokY0yIKDpCuW03YPxANii0mNcLljkWcM3cYXPjv3XdSpOAXC0xLpMPN
pDNssQJtOiePWqVZfGl/WiGWoTSV+q379FeupRV+OEHt2Ypq+DgeuxNqoFj5ShdYPYcEgYHZCIBX
r0WcQo8qo5/la+HicGTTFK3VvKYJLIn3ExW7TVXisTNlfMOrgdd1+kUI/Z9axz7QAamOIIUE0Vzj
Hxf7dNfemk3IddHhTQzSkBgZHc9pLBGZXWMWMafT0Vb0+MV4DiJNOotbxXV0Nskj0ofJiYlBcbUj
GzfLhgXwXH/te27V68loF5xqB3FZ6DgYIRUpuJCQ+IdmONeXwLWDgOkQXKv2ZfHXYABoPA75LydA
pVxjojG9ql5qalgKloAHFyGMbTK9e9uq6LtiAApny0JicaJes53emgsfxewuNSx8QbWwNPIYC2nu
dGNtBYxQI9ypyZmI+LxAVuJxxWZsA1MKZAS63+EZpLZnmJBIzOy8rQw7/jNp1kbZEMLOIigAFNY6
P5duFPYi/foKIs7085/yed3cPZW5s/AHmDGsUJGPG3U6Yvv8x8MMN6g8nmdHT3Lt4Fxw41uvxn3d
xsxL8hAt/OCuav53YVdt1QNMI4+68StqIMUO0tr1nr2KGg6uwEwSwRrG9Z1nrZozO9f8xqXE7AGA
8nDu1k3/u6tN1KOHlKhrTP5QDEa3HDn6O7MeuFmDbQ1t0kzCrFlDxcEDIngI1/sYOENvs0mQdoeX
RcXsX4YfaPsOSjNOkAeVy4TUuqCSzY9K0Bpm4UrT7QqWJ+kSAWDT3CE5S8g5mR/eUfptWlj9xBx+
PJ6lL/0OavQqFMLnWaVma/Ml1VxEdDZ+CHZEXewjKn24ajiRNZ+pRmypZ2Cfvh2jXjN9nAYG++SL
0WU+RbPPKzWnVLnWt7KrqOeYPPO6Efh1VtAsOtbEkrIRclmXYHcWS5YHDJmvl6s50FCIXVu6cnlq
7B04YuNtC0QJrshwKTgelR5gKFgs8D9jDw/F5Tp2fg47dzKQ7/xSpUxT71tB8CRR9b1W6xxFVaQd
O/HfEKzh7P6U796vgEiVtZgUuRStUariKffORb3zF32Wm6lVLbZu16BPMPf2MKpyhg7BguR5Zq92
14CJ88fxKXqSv6ElhKtk+9OOlAQe34xi32XCP0oWpm1QUiwjnU6yocHnW2pniFCKzVPpFlQdqHbA
gvBfqrFndEkKii04S6V8pXjiLokEGTTbhPTq30ZqrOR9Ve5bv88QIHx3lcsvG6Z9r3yKJPDNyxW3
/ujyx+gjottflnINw6k55VwYQ1MHYrNDDApEfCXneN8IF4ItG4+I6tDkK4W6ti38RlPn92mbvjcH
do+oY65SNsw7RR94LYN/UyRtDKD4/c8g0zmjMYHLWGY5g3EZY8w2psHb07rumd3aPX9bsW4UHu97
357OZAdN6+2daKPUvSYeaxcVPpgKsoJzkLkDAFBk3SIrJQALq9XawVGgpGLylsZrWawRagNGngOb
NyUY67Rk6SxLnfJTZtUHotF1JG6/vDk5g/c8kaKuqtfbbEaRHT1qNzqQEaienD6n2CFBd9KfQinR
EGLJa/ySxCkfHk9Rbh4KK7RxVMHn6fCSOehyW2UKz19LNP/C4y43VpN3WNOk/k5eplCinFG6xRJi
QqDiZAdX477Oio+3GZ3DWn8OwWL/CRNd5KgQ/CUA508S6ycZnZYNUAKiCN/ArQyawhKb//zVYoWu
tmURrT0gYhwWOpYUFcqngdmRyGFU6vj0MtiDqXo5f/fsWgz/smyKUzMSunIytzHmNuiyRwMN9xsO
w7Zpv0fbyGrFR6bKfQWn64usp6XRJQPY1Z32prbvUnriw+JkPjdUrJ/JSxLwiwoIXMan3vkxbXA1
GSNj3THO7Cr8M5DoZQK8dJErRMpsZR2U0SkixXyUqqZ9TO7/7a75vY8H7Qs5NstR5i4AcP/KdkoN
lnOPNeNl3qHFuMBRuaSVknx3hCyHelJXE4oau9VN6guVmRLaueX+a/wSvVl2uzbN/4Aqqa12850o
fb7FF4kUwqNhrPn1/TYua/T1hQn3qzD0ewEqd49NYwXb2MrJxB2hzZTPwPXohE23lpxOkOLtjP+7
hldp8wkBfyVKnpknSSRjsoJW33IEeyvUMXXAiUQTZNmnWtB01tZ17FBdiY+IeRKwYNGLbsB2YmnQ
bZevgOZ2Z/SpEU0Jqsv5k8zYgMMFt6ei/yop5u+yieKEuqdS2pzpwrApOTIW3dKdlNDFBR2+RCSj
1tmzLo0+9m7jWO95Oh2201rvq3W4vjWoZE4TMEcxQucLyp/MFQhaRN4MULRwXmqHHo47ilmwHCSg
aN3FQRRj/ieFFSMV5VCFevYmKPKwhQn28DZAf1Xt1f23s4OGtyTaUV/WTxPYLpPgsRovlZ9dwlvA
2l72mw21vZpb1Voibx/EWF+g171zs9wV+rPljmluUDdhdq5MW+bd/p2Jth2gRQdjyExxadKlDYPL
tdUaBIcPCSWvvuMl7lAMvYQWRrioY/zEgXMXFJqj+D6ydJ415/fXSG2YQLy366cC6yKQ5JxXvoJZ
fzj5hwyw0gWbdsaP9rTU1dhsvNi+qQcYjLx7N588RpNs8hunWr2e35mgEmmgu3VS1jQxh81wXYus
tXbQJRLjESotxoYg/H65b/3Uprkv7PnOJ0HeGdIkOxzRLD1RjqrwjVgxN6O5RT2tIyXYOD+gfYRV
6z7wVQwvUHz423fcPOWZxQXbC/oEwliiZ8r+j36wPOSKiBU0EnTe7gueWzTzl49lj8m9MMaTQKw0
VuWmoxQF9lkZr8yI9DiQO2ngLMWmPDXsrmVqTEqJv7VyjCL11I7rO7ytslow9lseOFpu+GVYpJpk
c3g/uJ3N9+lsUmmExTMjNUqO94fMqXuEfCZ23k9t3vJQX/s8Ex4GBoN1v53VrL9+/WwiYt2+Mz5Y
2jAgs8A7kpvige0QnqfF14p2mjn/Tfcf9DYw7uJo+TZZVHbGTVl3zwTBj4986DtEbbXpVbYO/PKC
5g80ZIs9sZ3KD6R5/0eod8F5yrOsCzctByE4JYM2l1065Ce1gztusDF7kxDG/5NApfOITsIUrZCE
8gTB+8e4tPksLeboLaGbCEm5+M9LWxzE12to9Q6sURfKWHgiFrNHhj//OcpBb5AW0gFjwyvHKXqY
NXOHyZhOGTS8C8v1PI2q2KGDM7MS4HKpfWG0rDEmFLmyOS3yop1V8rnK3TPI368+nUKTTWwXDXy3
Eo6sqxX+E/KNt+2zemfYqIegiqSacsw/Mz2o1UkWB4EipHucfTqbMElhGEWZlPIVmql0gLcinygR
+gRLK3yvKd+LKlOvex1YdX4tHfmSjr7bBji+GE8LQHTldr3Ud0BrYAB4PnBx9VNymeGepq8wXfJa
9FuRH7SM9Wm/gDeHN4RIgWPoT6YwK0cmpTMWWHN9HiulZc091VnjvQAFm1PuIJnSa+kLl7hurEwU
Fxlh6x8dPIhimzFiiBNOjEYHhVne5gPinbWUKNgZOudWvptfAAIYeDA246zgpO1ysQNaMxd8BTZZ
Io0DhjLy/I4qoWsFGu7OTOldk2NkYb3URMjdfcXin6V4tL6M5I0ioepIiDL8Poktg2AQqV1MhV5A
JA51QkNvDG0FUCCVsklrmu4dzg59Gn4jRpNamHE2EiBExO+MW8BrAld3ThvC5ckHNuylhau01yaP
r9ko2jDAAPJ45T6FFgFJ3X5ZmftFaw2+31zqHPUwMGAU4PGbuVbM3GgT4he0I5N5e1hDMn0cMEuh
RX1/+N+5Wdm4u4fwjs0wq3xWRLBPsyThrsJ22FqpnUsHpMOUmb4XvjOKn3IXiM5oA5SdxCJARTm+
4iDAO9w3CKBhHgYjmt7ssu9yot7dm7SF9FgMbiv3JYNymKvrhixzdpXQjdm4Exabd0YHHLqGQIJx
t8ZlJh45G+nzkgwoNm5q4zqW3Uxvf5lLoMpJWEjegGyayPTUmWMPDAG35f0PvkmqfYrpIVYzD4oZ
We8VB9i6XxvBQOHYNFLNiM73ryhg7D/n5mQdVz6AlJ3MugRtLIXNASqYcRarnG+rfhIZExEjcwKC
+7ABfF+fcsxc9TKVdBflFhcl7DgLk7ZuVUeyFgCjiYrSZQmsZaKHZq0GVZxYWt/jslnouLD6GVWY
p0ngWlIB0pbQ7jt85814eRtzuCIrQggMeeZ9aFowM5ciXXi0p/DdTGzG4oKkXe1Gi03RYjkCLBJP
5BjOBBBaOqB8FZ7dM1xiqXuKPWYI++90ZpEQYAkam2WXYvtru8RPgDL8rQm24n+e4GgjQrVk+AvV
+cPnkiHpilFJucEggwgkzc53B+XxWeubmBwhNQGCnPQ8Jo0gwrtvztaTaEU6JcgzBwhLHhSUGydI
87//RJ2GzD2Loz+PP2gfYGy7akb+qDc+kbUfdWE0cwi9TUhDR/r7D5MK33OCO2n30zmou3a76rff
Imok7CqXmaMwjz1bK2G6YSLsZJzDjJnvP2T2DuG6pJGo3Wlx1FY7CZVSrhWk253iWeguVOy5lifP
3tP42sDLYXKy0AK/UxkfGCK5iZEBxjBtDsuYD2i8zPSLzY1hwUg+3Hz7eC7RyuAEVrMsm58M3xYj
nbtPZm16M2TjGHD9fk2VjIKnb8fvUAwNLVe9XyqWEL6DrkZnHqvHAYKvGmo4uUdkgXf7DauzXjOf
mbu0rVMTkUIvqbbCiVqIOXzC7z5FwyCjn5BXQdWy2StMidlyuMeuSiSBfQ9isHX8p6tW/LPKP8nQ
k7b85CWI2Kv+biFU9gXpa1RQSuRbEplC2LBMELXwFuUlGjRdvCbDzv0PmC25KXf8e82/EBlMDaPa
HzhJwLkjH73oPJM82qU7VvSVybeDefFyhfXFF7lav1yu3f7pCMOAqPIkHArqGKSHBl1Ybr42Ute+
vGo8Xpg2vGll7zi5FJvfpofK9Q+jK+h0Xzq3sOP0hFPoy7JsOU3yhSV36wpZCc02OGIB0+poI8Tz
4iHVCmmDbufOHqCCMbGKF4ZoMYAzyMLZZNAYFqoi7nfBA7MKjQIDB2sOOtZOx94DNVD6oGXpezE7
q07sT7iHWwv9aUutuVV3kZzTWsjG3eydnqVyr4ZWKAbaQs+26pA8xJ76kKMRi+iR+sfK7yFnfKuj
gOrChVtA0X3PWw5+390XTJGuTAF++hE9fQD0KWkN994r4WiyN3z3vmJLVSN0lnGEOtboDduuHXuD
w9Px6Rh2Z4wLfExfdtMSYjDZllkP9HAjhkfS0hrkX2ecmEDzG1/R6l7bhQ0R5dAxaxkrM9MAJEGb
80ZfwcvYk6bGuLbtURi/hFvmylSWxBNxUdVOeR0oTA3T6wu2q5kQUlhlSzkJMX01uc0NfshsdlGA
yFBDEdEAw8WfO99BRRvhbiVgzYKVoxa7qeg1MleRlflT67FiqLDQ+t8ZSYACP/GKfNnHu/yrROmC
H6LkEAlmwl5N6409Oz3FQ50zn3653HNeXEx5NnqrgYKs0imEYXxQ0pzNMunEsYdR/eFkfDl76NKp
YGHhqW1WPUNmpAFYmeUpTKmp38JYFZHo8yTUMBmrP4EeUZPmlBKmV/lqxCOwIb0exnEf+hk6VXQF
8kDN7KrKqtiGuXd8IAWswPUm63xai0lQiSNh0EtimU/4Vd82EE7EBuPWH6cJDd5TW8g2x0NMsvLx
mLX3ROn6yz3PqScWR0eujq3RcMHON86LbiYRfmrc/b+KxY8Ial4/YnKcjyDyN6WqI6Jw83L8/I9t
9m0WIpsS1vyKDxhrjAchoa/Sl8ViTOaC7kf2iFsFkewQzcf3mKopLRh/Nr2z53zuYUvr41khOa6m
vhihShfriIftyz9E+E9UhzjfJAR4dSmMcY3NAuPRQCWPzEyrJpnSlWZvodQyo9rOTlDT9/3BRqYi
u15Rl/u2y40E2qI3Qh2um7EJETOlis9qRmouTxNOzSRXv71o2TDa0FNFkgrKNuYJVYFqCqf231Kj
8Ez4ybWCJ7pw55pAwfLExeG1BXJYzYrs+fL9xXcnji8IJQpAu+zhaXPAi5q3HcwflRS5WDlktYrb
AzxmIBjR2pter0SRcfKmKZvRHIaN98B++GxaviRBF2jRXDRzXjmc/2eVqeHcfnBA08P/2aoFjM6S
e/oAAMTNlZaD+/OQDRp0roZxUn4VWwjNxqUbjdwNTSdHD8BxGJJaxfIkeS0IKwMgYt/b90mqwLnm
FsBBS0sqIr4yx9MbKa0+oP3ZnQMAGWnjs2ilEc+nA7HL1UQn9pSsiw9hW5OlnU/5upR7InwL87YU
CadQQ+WPFajSn5OsAJXwUIhXJ3JB1eo1bNgRfWR6jc7Jfuj8yUygIe96wFJu5QiTbzGVx0EJNF4w
gbWKbPSOa7SRebiwno769VifygDqnB7AMt8BDCyby01WBmZTTAKfyf18QTIz3M8AGY1OJKIuT+nq
ZeezHVRR/npT55JVZkQWGemUwhGoyf2BvCQXyvJis6FXhL3hxJJEOZPHrrnhAWFsahS+mpqa9tMl
Ic/rjtZdrnygG9a/kPmPvSq0xPGBje5Y8aeA6UZCeYJOcCmIHXXd/EqiNQceNdJ5NcJxR1gpenDB
0TCV809+VSl6mf18X5pup0dXz51n0FX/vgpwWTjF10G9sRWZB2BnRC1+clQRnbok4avqg5ylRK30
yyWKYpdSHzbsbZk0c6mNohQuysILUIJV7Km3GwkhVUQRzIHMMlSk0Enk1vx2T7tW7unWII2tjMXH
do3MPlH+19FLmv1V/pMi1KrFYqfh6ide06Hhg+G8ilTqN1eenoLkOLHvdyX7ew2qwoBB+DjB88x+
/hIQiC1ElOdq+98t4te0BPuyHalaDCCq1Q0b7GBHLvdlL0K7LkJIPs8C7k11YdHTJix8ifjnTazu
ygTGon8zq5Kqa8rBRWWdmTfbauu5ufA0FnT/HIofLTVt35yOt80AHYjqR7tlotlxqCLqAeetmgCE
RblQTt+qjJEWeMmRzakz73Cvv3TrSE3ixS4aRqgg+aZkt4knoyu3C7Yo9+UvtWnSVkGLaPViWy4c
5lqRK9EoiyOcLVn5yzeM90R7e9rawycWivU4SYp1bigq4CzThIWiABbB4KHKMhJ44V0fH5/HFEum
CTOmsVryj5kIK9+8KcElw6mWT7kbIOfY3Vj7ArIexskNC+mHIOLDoHLGKSyd7maJ5XvEUEREjDDO
3ur/dVAUeWNWJfSD8l1CTUktiGAc7MaRh/9v25xrjOoEXwr6ZQGLu9kvgL2mCda7pW/t6H8mNu4T
Pkp9eH02Tc66fs8GpWMp6dvLk1L4BBB84wnhGDumVtTJ2S8VGhGtmCWORohc97jd0xctEqQ4fMMT
hHYrLnKVhk7YxZWFfeY2RpSQgIjMRXYmociqyl4uu5n5r7jGEmfd+SFealjtpwiUcINbT109fxmh
Zta+VafL3i8FhVFqO8qwE0zmXu2kTu17tearCpsl5S5TMmKMJQ7abUmd2qZcUy2f5UKIaxOhcctH
cbvQ3TG+VbI4zgoXEa9/Sd5h2GtGCJTfSNju4ubCPaETHh+llcFZrUsmwWfTH0/I0uzJBa7mNI4L
2ySeLVDifLOK7hl+qMHvJPHviSDbrrQBYTDD4X42I1A+fd78eOvePKO3x94Vo3oiEXPu22vDKSL2
0pGICrUPyzhZdP8iMAdAWZA996iasRpW+mTvbQled5KU3ynWlFHG3JR6BgI+93pRaYszsC6S4l9S
VxPkdPZh4tRSk6q9LDV2v5IN7ybXvRJNoojFT/dapByoZ5gjVssLngQFLNajhp6OnUB5pantLb2b
VMpGH6Q3zcQUBSen77ePthBpuvyx78t+IK6z7IVbayKVtvpz79vtKRgucCXcGe86E/QPLTYhBLRl
nHoVlubLj2VAU8DL1ZHyDd2xTOAo8zV9y9N6y0wzqdEiAoO+7/3PnWckWkGgB/w20Bm+hAB0PnGk
W2/pD3QTQpC3it+4eCtAHNbPvjrfe7wbKaCFl87xiiUHos/8zL81knBa0iVxFoOWdvK7lNkK1Cdk
/hZNYTQfQEwebAuvj+EJ01CaEyjGNvhuK5uS8pxh/e7dHU7GGPHyrunQfqrAfB3l9krXA29ehKgw
XHn7lQlITk75sMMelotAjrN3o/GpGLkHj+ds6A+2V6D0TMGQKjnd0HMD9FXgtR8CAKvCV8DaHncO
dnLeNUXLP0yZoTiIi9Y+cKS977VnrUC3TDfCz5sOjUvyLIppCOGcYzSroLYhlEYQgPd8Qg1qABVM
rZOeC+BGTn2Z5ymc2i0a9T6QBUBWN+Raw5/TITg1qAVjENQ0JASstrLTaWGqdbA/FH9E4Z0UjV0H
yzhxifhZ8ya81/hvx7bQIAKIGKw+zOzadSR+AJb42HZ8qVc3SU2hTSEwHlW1dfDLMKK0QhkUfc83
uoyXw5te6/ZEEyFWzZEwkTYWXO1vWNAPTyWVIDm5zU8i07cEWWN+Io85MYhGMIQpQbhPDNk5sRd0
hu7c89EucKAAQFMBi9UE4RjXUB36dkVCCyAhIV+N5MdCh3xxqvijArfGf52CArPvdt1A3CEP8Hkl
UB3StX7+4mvBub5XgZO2KCFjzVQMfIgpqkV+Aw0/DHI0bEMMaC4ZVYh2/ksB3EtZsq+T6Ss4JG38
sDA9IbmAuMKWFjNvejzlOiOBEqNH597mLNCEdo8/LvEhjijtyJ4mBvfiiX0UfxM5X1o+r8SIgVtK
ztUx79RcO7dELIqLkxwI7UdaJh1NuDvh056s1DQW4EsdxpnrBJnOCs77+W0m10xR1L6levNKKsKN
bHCheTIn0UO0RdF5y2W8p0w749ZISznchW2cbxzPEeE/Xy/0ShpuVa9ENn4DiJ9Xkl9ikT2UKsoj
G0333ZTIBt1X9GALh7PRCcc/7svjCpAa/DDssjb2DuMvyOOT/Ys6+YGY+5EkMO9OnnJaDBKtRVlF
v9WxuvvdwfUBy0lDdb4rRNhyzjopbxxbhOSfMilNivRXMNujxTZ5G6pKE5WFP8yf+XnMCepwVIip
QgYh1JrlRZuhFayaQjNzpbL9xS891xy2lztmeCWGKD9Nz1+UKX/aO96R1Jofmzu8Hcrh3hfGBUmN
Ju05s2nE7n9qCOaKT1Z3HV+TE86bZCjCRH7EOXXMtHrZfmBu5tQdZLc8gIuMkHRdH0ncA/B5Wgc9
iBSlSyM5ucJ52cHA5TnesNkiK/klU4gdT5Psk+NQ5ggzfsK86pYDWmmeXcaevaXnrTo603GcMP4F
b2Oo962HWVd5Oqp2cLAurBqJCAX/jD9ATAeUF6wY9wUEfWr8d72nL4nVV/6ml6fCFpyWvDGhRyo2
IXXoRrqs4UpXKRPIGGDgZpTi+LGh+5lxlXAYUpvdeyITJMsbelHYOSqam++uJ0Gc4NKXyNO2IaFU
VexPEVmqi7otfRhsfOlj4Bl9eHAgrV6GQRI+tXj3HFSBaqQCfBdAOIL5bAgAQN+efdJDpzRe00jL
dcdSqxozVBsZkKgJNZxJ4fxYXX8yFiQsXWnvjE9MTQIRqQ7gH73ALuwhw2HBu3ook292kp8zRK1V
3+pB4ZtUO1gb1rpQSxmuw0oWlCA2qroViapxElcVpU69pib66KMN15Qz3+lmgQYJdS8xP/94W5H9
ask4pMq8giO9xSfmVv6ldl29Gc17qOKIxT1c0CI/J94ehTtP2913HDUK2OLu8VgvPRJaXmeFf606
MC5ABgaMtcmXTZJQ9OSUxSstGZ9z2rbVMAp39D/puHNFTCIo/FU1qrxcSucUB+4s2LkZGC27ta29
FDwsukFQq1JNjJ+mTvSF7Rg13tBk0lmq63oBrIAiTM0IMUudLrsnImFzkdA6L5azcbQEL2o7knf2
svIMsl1o3uFLBxgI63Gzxo5apY2OD+4N523UpBmCVoucGtdaKmHGTMLDihDo/KfWf3UOqJYDUuqv
ks3Y8lERjU7IOwQ7OW5tfGNnCGWShd7fG/murahMPYtZUSf4zXbHSScwSAvm7oAOfEx5hN3TBrjG
ed14xDg4WQXTSaWDK2t1FLOZWeem7JQBwp+mmettr/x9xGecLBV6TUefqcTOnZ2meERFGaLx86s4
q5GcGywASdTn4DyGA+HOtf6QunsnOHs0p9RO67GXxt3WkIk4RzH8VXkSTqpcA2RpuYvgeGX8rGzt
FYCzb2h9v3hadNcXw2Ou7OSamSAKGTsWc3iTDv4sYPLXJ2ceSw1L240LdSrQcwDG5Gukez2ujoY1
679Oo9QfURVpVEF36erMy4TXosxdD76iu981XMx+bFpX21Wh0F4v0+ve2oAeRlNhwK09fwxwqPIR
gAOlHn6y9ib+ZtYEKCtGh4O/wBZ8PAzbPKTs8LaeIQTYwoM3lygr6pISRJK7wtoPsDSkmnvEF1Jp
d3o9cbW/gm4SoQbFcQhBzcCnh0XWN/M4foQEh5HBTZIcplNDXZ85qpYBffqlxibMF00ttLi15ZOi
pUTOetZ/JcM0672irD28opTGnfWyckly2gNhKeaqx2oJv41OKO5TTRH8bhB9ot9pE+Qyx+yoC+oF
BoAWn0TI2yQwLczq3ZX9KMm91jCpRzEuY3LlNlyuPziuXjzHcrdyH8v1anxzoLJm3XQJAhUu3R1P
ikzNPakfUdEGpsCVGGGmF+yYW1uyvHX9lYVilBEIBhlfz1jxRYkJjtoAYSLMQJFjEYKLf6Gxg2yN
B7OFzwIBCFZ2dT7XO3VWmis2ZpKxivn4lOd0VZRBzPjXcGf9EPTHOU61zeFDXF4W8cNQAPNbbqQF
uhHhj9RVfldO4+qTBNkvxxuu1Li6DeRg1VVHhtU5gns/4ftfChxPLwvpll2393aNMGX2NpGAnr0K
Emz1Dg4eJlq4Nq8MH9m8KtZYW6CGdJcbUkPSrCAQkUlKOthFAxnW/nbx+Q9QjbBNd9FbRy8RDHFS
0+SZwGdQj99OYU4CnCVPiRhJTcx/AtUzFPgE/VeNsguuQPuLbEIFaGIC2gNhKCgh4HuVIlBtTGnq
bf6Tmw4YNQyGEUVJX7w0AckB21Vrh/rMWnUWP39o68e+QMC5mPPCuOBeG1V98osE5C9BRFS9T119
CiROupfzjjKEXyjdCPg+r6fHjQIDSCkCeLjPSE2FJfn8JvEbTxHz1f5qwcISuDjfByg25HXUaOQG
a56Fybbg2GX1dPb+/c31SAK6aTjxNI/ejJStQH7VbrPKiz9Tv5Brqy9QSCvgIRJ+rGf0ZnDIdEgN
M+rZTr4o+1nUDW+MtXYPGmwyHzUgQFHMYBNS16kbUAX2LbFi0OsIzGmgU5dQVb1t4m26TUdjPhce
uSjiZHGBOkjS+D4m0mn5uJJQpaR0qSbpc3MsMYh56xnLw/A/zIvbEqbsSJm5Bd0156TwdJ5TQMsa
2Y0M6fTDjn+J7fuhR6OlDeknAWzTtFsDIK8a4UkhFcn0zCEUyagJoW1qmzMlUFkRmOv1WzlQ9wtL
ajuHofHfkKF6NmXz5yqGgyZnRQp8S3AaFFcprTOB2k9RHLrkaVmcuXvkZic50rF6UesFOjLPLI73
K6wrk57dTn9Kvur3P88drTwZYiLN7xK1+a0qa0AMf6J2Bx+2RZI/ZqST3vfjiImzP524iRvKj3Bw
qOqxfw/RfKVHoQP/3DnFBSf0mmOUnQuQJ7NKAZlMZYeWtB6upAVazU1kBwCpqhUARfx2AgPVXpIM
a/ux7R5tRiGVTzfOALbm+3NPNV5oblwdONcZ7XY5rrP1TVdhaYnBMTcjtiuRIyTT21HcoZm5KWC0
RmgllwgA7gu13M/t0zuM0L1f1aDw23NtsRmnkMnzvRTuWm5pf0MLfyrvKxs2NCuNEOXt0KjpYFzc
zkUJygSeXpqr1J05lKTy8RQtH5WI2GfnrzoWZE566ZZ3zJVi9LNzfW6I1605htYhhexlHOgtA3qN
IeNYM4hKUREC6e6fYC+D7iW47kSrVdolEE/80CNXdKeqMsWBFhVlMxkEzSFSKBJdIGScv/qdtpO9
S36CYLlB2rsVZU6mKh2BdBAQ9r6FCnxEWVO+vlxo6nTPoP3/f9HgNLuG8Wq8+klmoQ5zCcc0op+G
wIOo1nbYuA5yC5HNfpi/oHDhZ99UJadQvblszdxyOwOTuyyKnMgnzEZlUha93Fo0nsyK0JhF/Kpz
mIcHwMq0gbjv0teabf8ERSJYoA4e74fo0Vpv5IGihvayrti7xiK0LweA+yl1toMllnuqFR3zABNN
02q9BQYakMifG2HAiOceBif8+y0UqYFbIo7KuAg/CWfNmcnbt37BbcGDuWTf5v1uy+zWgeI862Jg
U5Y/TkM+tPXiBbFJFTTGOTz5/3AKBCRKyzpG1tDrB/8T0nICfFQrgYbbhVmmUeT+jl5YFMjKWn/w
cKn8AgLaCXTburLWDcRwvFdbT5ajupLD0vop730iac+pasVfv2lIMSnlw3B3+ZKxoBtkCudvHaY6
UTuA0R+AUFJ/SW2KP6jLWHVCEbtbqoqQCNujOjJvLhmrZ2TaFdXKqDlbOnltdMh4udsAz8DJQZv2
3VzEpPOguNJSTmoZg0TU82aFkkWFPdyETxX8FQXxd2CBXaMsN+DWSs7d7vnnGXTSn+/DOZvS4qYq
pKL59fjdbKaXep+vyuCVN0IJ18+SHTWV2YQE6AwdlGYVhRZnvATvW+bhZL6SlaE9H5HxpkIOg+Ge
ZfW0pVN0uW7BALG/Ddi6XNdcN14whoJXFancciiJGX7DemnApH5a4FZ1GW8YldKp/NU2u8c06Y4k
krANBWMBb42qO/u6B6Ht5sFXkWU9AWYxyx7gjQwKR4B+r80yoDPrpqGch9cVPADzVjQJhm1HpJFY
sCdgtevlyL1fJdZhXFIEknLrKboXVIeWqv6DGqVZhg8vKeN3L7DykRaAeMLxn471rV8lhqU1XDBR
Yyo1AZk8rsainIVspB7WimLiC2/w/kZKwclYukla6UJbGKJefKtQD4COv9nk0QEDRtLnijtpJLkY
wLma1t3o6i7eAtVQRVTYxicC99hkv9ToJuhHSXzAjAusRvOcWtZJhMMUplSt0Lu5VFxkEx2dMc0C
seIBzCyTu2ZjBgivlly8XIWUhwg6+Y1yYnJSByP+hoVZlo0PUFgcMpgRcc7nKHsfxgObTkOMxZGD
sjpRXH90gYJvc9kX4B94hzfxQjHvtF5PaOO6touEYPXqwHUSq1uyu+jN30X1ak2156lI8iW7yjKH
Z3M1O0clhzXZMb44VaFbPv1mpp6KWVaGPWW/oF4wttqUcLWtuQ+Vemph3W9W0xcPRlsxREyl//ie
st7mfQujOupR4vG8i70TK7Bvw7Amy1oCdl0HhlgcojUkvwg8//YT6Si030+zB8O4metBV/2/mGwb
J8mBcPA/tKz5hxPjE3oUe9eV5okjDe8zcJByTRXOKaMXrLS6+jSITYkHI7uVEYqV3HpwAc9a0MCP
Vo9h5wQ4nWQe9j/Qr2fSAB7lyNnmqMlbc+0ZkNTYPTat1ZByswNcj9NyeCq3hz05x7XSxYSvx8Lv
bMXFR7LRGJUJ1OQjeVQnYBTY7kOr4G0B91Vw4fjZQZhC92q0c4R+RtXOM+delWv6N+DUJjNmAXAc
1h+l5Xxx7jtym9AsXwBfKr+5ABroRO4KyJqpoY0a1cQ4J2q3B+BWLZESThL4uWebWs6F/UimB4G/
TWhumYw+w5IvsRW7yJFb7UzI0Omju56f8BftS1+uup/kUO6mF3NoTeOTARxDVNZrgYNNu8BYxYZh
1V1vYqOX2HSAaqFeW+LHMS/2GoiWtGWW+21lbcJgKUP3AFRM5joHU7x5Xp7dxr9CWxGqrnOJr8Ww
1uC0LPBCtqRDLiHPC8hyNoIr5UPz/u1v7RT6VNUi/cDS6tcX4sSepxfqB1fYpM6kqHAWfYOuglFh
tOWxLysObLGol/NyLgolnJHxo2N+fKbFab8JkDUEBIX2a+GQI3BneGHgGTOSWcLqa6CnnFggJ/Dw
P0eeTOO0VjeG61fciYLDAhCb16wOgUQKa9Wnk8lByD0tEawxjiCIJ/EDEkHxMTVn1DdcZdZEp8D3
q6KTdEVBxvJKr2HGbyTNlYj07vocheDGEIlxz6elI8gfpnwGLZ+xmTNU56RzG+bw+G0C04jj0C+q
+4OGm321KDI8it+KYBTbuPB3I+nFJ3GSBsuYXQ2qNGJ1lIHGXt67UBTedefvFDY2IdHiqHNdkP1k
G7E3U0OtrRTs28FSTW0zlA74qGFoIB++Z+rGgWfvl/hRC+ky/Ms85CIpy73khGVpYwPS5zItvBGN
uZc0/jDxYtnLpbYujYe98xJqtyj0vIG8i0Sy1WWHIA5CCYwJobiaSDoIaLjjBLvRgNb/TmY9nPVr
W0dCUcvYtFh+GyXQqR/GANmNTeOXvFcYX0iXDiGTkSmgkQW6bnbxHLFmcze3dCSdCltw5AsyYwV4
ez7mQgU1Jl08LW8aLJmju8gz8GDsE0i4qtDrBIhvgAajt0lstDSo216F6emGIlZM4bVAUY8nXFZV
8Zv+N5pulHpNOzBVabSvmCO+hRxMJl48gC1aS3aZGm/6Gb9/0l5Cuiloo0nizM5+Mq/4EgoTykOS
UA/LTnEYe4ErWLqfGXcAL0yZ4VaiHHsz6/ZMARA/cRZzOwupwpeW8EvtsntIdPQotvlG6xjz6hSG
718Pl9WBD13xZHCAwAzjG3GBEeGoTpMaWaahf35gIa7q93LVzLs8QL+wHa8j/M7nC3ukKabcq3/0
ivQkIRtB1xV9VWXZ2xC2yUMrZBR6wl2RpVpSRFIKIOeclqaNjfy3d3ZDy/sJlwhdnJv1jgU6mY/8
oj9ANmuBHKULf87zdsvkUP0dIbUniqus3lmgrXqiKVTs5zm87BUWZEgz2hIDFiiwAVbEEvAZlott
8I8mzHtHTAIIP9GfrJ52J0KZy6T9MJzV/T9vaGdf9KQLoec3LrUPog390/aj/Tc3OAzUywlQKAaW
SbmBQTkFi2of52jd67cFEsFuSlNhX9I/QA9GtSjVd/g/VfZhEtSVZaRCenZKLYdUrTSn864h60NS
5O0gQN48O9x8E+JZwAcgtsnqzMM+FqMwVvtTsruOTD7Rn4dwgn8C6NbiULjnpKrqt4mzPcVSeI8s
g95JYMqbGTse4AXBFGMn1Sd1VyUOBno/+zXWObAyHIj786+vXRoUGVHDzOl/dsbwKHScCJyHBs0s
LHCBg6w/OvySc6B5XfKRH1Fw8vtjVBykfKDgVVMq+WTD7ZQI/1OFTS5O+2v/gyR+vDVlRgVlmZ7p
crz1eTJN1WyWuKGGcINe0K51y2RankVKWIkDda4pwYf0+0t8IcCAIGHElGuIAcwQHvYGubkFJvDa
XTqqmCZ0hj5Awv/95aPofEJ4JUKA9SIENqECETMJPILu27cTOwhBvE2n57UPNX7eNpADkbvcEjjT
LYlnLe1UKI6vRVVGevgEvzlALTzQ61CjCxUTvCYW6UXog9id6JkCmoti9Evc1eGoBSeJDm6SpBNN
R/UZuyPj7PUUwIGF5b7llFyOXEMNb72knnD129CdjttXFnpQMaVeuQ5MnyvwGhGPyIQxDABkMt/F
1VdGiuokcDlt5ri4hk11nYtcoqMhoxw+EPLSKyWpZdVaZ03j+nlWJLdAIALGj2n96+2geT1XRPGX
8QJyNs8BEGeSYAXtnTgfbcJwIO+E/dZfu3w5Fh8N1NloqexL6vko/i1lhg7+G7VpO5wUpp9JoUoP
xBay+Z2xgFR4pjfOw1S2IOtoP6DloL7kHtp+LNa0C5A4RQudz9xErj3bMmlZ2lB1UmiTTtMp4gtX
ZaM2S+NqIBhvR4jdl2e39gJVn/NJ2nzX6CXegNNDtihHg+Zf4Qe932W19sczSVwpv02iriFoD5Yp
gKHa9fUWLZt7pMc/TZIMKgTO7VQeRFJxYHgUhgGQ+ZdJ0FbpAY9D3dVQqoTqQiMUkDsniFVgqXxA
CXUgs4RYNnhuPY/W2mdetc5VHxaN1jjQTP7reauU5uyGyOR7kHbgB3maMKFZ0tLenyC73f2i5vE5
EDBrUlBN4+rdix+hQJtKKzxG1jvYxkdAJ7qmkCloLbYEjPQmtPtG/prfCDZ/Wx2p1tMU1CyUfmwn
rIH5Ms8csZTeO/qigl6wkojZvD2NnAZq/m39n2JQEApKXLmEemgx4DRgsfdSrHiGGco6nZrJq8YF
XTjAdwXDWude8QemYDKXoVd7lQWaGCFA24guMOQsckm1rxtsEN9jeJyCy1nyD8mXCieZ09iiyL+N
kLkwPU7TaZlu8ZG4hDoOVwXzzNSMkCJZvFfo34SWx6MN3W4KjnN/WGFnWONHnMbdJYE3mD+wecUN
JZWR7NDHhuEcWulFQSs0bZFO7NMYwAk1YvGqO2YCg668fms3ZtYf7jwFXl0a8a0Y7fcavCrIgU7k
BLExvvy7X26WdiHSRYLiPM0enm/5SGntejRzozrY13phuH5uXW3xN9ytS6Nu1izmFjZZWIcjEnxs
TWG1+Yw2NA9ivCkBJv1e+MDhC1uLlYqEEVr/qtStgyfJn1GxcLWMSLmvHXC0opWqlDZCa47IY7Ch
o7okc+h7qX8xxxGm2rb5IlCxxfzd9ULYGzbY2OjkBifxA+JDZVWVVdVQqc0qtZq6FgHueFjmY5Aq
LHbc9gYOy0iyfrMcScqbMNOo60IFme2Y/ud+Dqz8V/DjmL+H8SoqzDErt7RpKsMrQ+oud3JanU9J
cMgilMBLBd6gPPrXAu1l6+MjWM8w/m2icBfaXORJ9FhPITIdd5kogwrlPE0B55R7uQUG8KD509HY
C4YGaDoHVOQnlRDeFf60ciBk/GWaIzo0nKwIhj86Lsd+ysDYLXPK06ufGl2JvEdR9O0287ldWK5g
jN1ZqEFzJUcbU9xvH89GmsV2G9k+bvYylSnwNiQpTtAdySOPSbxcC1qkFUh97Js91tavMWt9KV9G
ibwlUpabiw6fVVChYw1wD9CEyJNRC5Mgn5ZjHhRBIwjt1a6mkXxuitCkgEIEmiSuJXx0/yN6Gx5X
iUzNnY5+n/XNljr1on4AVtUzfQY/Y+RpfXYcKksK5N/Uk9qmZZQmRCwaLNdMXhJrKeeX2TwFGl7u
ceFnMRLvr5oYfn/uqi3+Qq0be9VySYFiOQmUOr18UJIC+GwF0whbDIQFIjc+ORWFE9k4RmwtJemw
IIkRjHhXJqes1QFMbp55nGq1KuwL4bxvc7jaCKIwRDlKwDeki6+iBem/pqGAgTHx4Gm6cLXpN61l
XOwiCMBHw9UIb1VC/GNBhGDmxlkfltV/yPEms/N8znQllGUD21YBzu4tw88rOJbHXyGFNt5n19b4
A+tiUPVi9UXKlDjbij+ndhZO/K50noq1e6pE9RLVjxbthm13ZrNkqLU9ScItgpGrWEsS1CcsTicP
zY26JoN9clOzfB4/n5zZkQLfYJdpPfrADj/hNI9X8BNh8WRqjWEmJ6huUuNQwNoeW4r/WHtJJC7K
yRm6tXBdKrQrEgFix5n9oxzVjXcv6+WQMk7UM5b9uSsC0g1zevu7nJaFpO8PI+UTIKJVqqF6oa8N
BWpsazdU6s5F7wyGlZsiFLvi4ffwiNygjL2mthzDtUBtvdyx+FGlY/hMulMPEA3OJ0LCe4VQHmns
rmPSI1VtUuJZFs0f3RUtTiI7eL1dumuJOeHvIjd+CYfZrYjFuhnTdlmIMe7/952pQpo4o4qMRQi5
fq7e0GqQ7RaIoCNqcfTFBPpBpmgO9Hnyp0mKNk0iM8QZwh4+EN+xuIGW6AW06g22P07C8t2soWyA
lgDXof13VhVqsW5Alc4f3KnR55DtcHavbDfEeHhKLa2HZdGocdT9CWHek78f5b88CdgD8vITj+GA
gPBGz4eW8o/ODUGkSbAX5ZBaqeOx/Ie1PVwgOMNFCvgWi2TyxL33EhDknbzpoV/Liz1bn9RCEbtl
NLsX4iv10QBroyucGw3C2sArkMTPQmX6lXwkRy07kcXr8FV8LMFkQTfKJe7vfRp0D36mavqrcGgo
2DXgchoCmyYtcPbicnRXW2vDofX/znlEmA4/xsrlqMG4iHAR4O8Oiodk/qVvBoXo7Msq3WbmhqI3
0U4eTpkrg6yD52E3UArP5rQyYo4QlDyVYwqo6o033UIF4UjVaP1pjrN7uJmfTUPq/WKfz2nb8fs3
YeR/xuh9L9kZniHMKDLleEFgivBpdTQ9ARQAxBCJe+5n5cJeP1NsceCVDxceDNMc6rLuKZ6X+YUl
Ky14NVUqgGdM1LEeA9PyhHQ856shbypBJ2GIMIFeXB5Ihu00YL/6qMtraAZO3At5Tq0sA5RAXgMR
h1gH0lsNE5vod9gfOjn6+k8iJtLntfsLhSjJj1dRZZH4P/eLvAXeMqYNNpSctAggnCbPHZQYi8WY
3DtRDCmksnD2u7cIRW9SiBUbk7rX9Z4q14hxQcBUVlPfhBdC/Zw3+dY6RvG+FD+KSphQFO2Q9TDn
tdTvv8h6hC+WUx2q87qzQYG0WQhEQO0FqA/5fes6IbUBZmx8hCKa6v/fTJdWi88vrFEhlhSJ+yTS
C22cPNwCH058WTb8F4gjZ15ye7Gsd5/n5TYHKlpwQ2UJAeOSdQ1xUnE0DDoII1u5hZCJ+SKv7AWJ
AtcsXFFmv3fGka7pfmmyUIxZ3eL7AlkM9y6aUa4nLzLoRYyue5SYDbT0aJKgBPUsBsXOvZeNvz+5
IOlYuM/VH0WKJuvaFrpyNzUfK4/vuJ56Sabxyw9GZ2L4xTgv3aTRBxUYk0+fvsaAddE1vFoQ/oCc
gIpxEzvUik/evLOPFV8uKt//obsE87VkeimOV95q6STF1kE4ZbNf7kSOUJ5N/moiOGXKkjM6hPAl
5BoQ6F7bgCDoFd8U0vVuoJD5QRLWcugcyi2oMUaWb+NrFZ1ivdWW277u/uhzAfY0Xnm006rvUW9p
KbwizkXKrtUNz2hL7AaBiw49B+LRcdyaLeOHAt2KHHBNoMB+YE3teqPNo4FZluBEb3NcPTKgasd+
3+rbK4Woor/xyezx3b354EUOrCYK9Ii4yYph5sZZPPUQnVNVqk1Hv+rHfwDvj4xnE1IQHnZ2TLiG
otfmWjFeFlMFSKpjLYAv8/A7vI1H/2Wfe+uhps3ys3b9gNR3+l/MXmQ8V2d0qOy89WFBxIP5IgnI
muCF8vkEPM1rHP1RbQRfv9LQYIOkWeFFC4sQnqiG3kDDnPP0f2xpXpYBG7mavE/mj/3AV3P5M2cp
lA+KlnbClktSoHxyeXwvPMsy1ZMatO4RselHT/V8MwzPBQsRiuS9/tLBDP8KW3JgFCD//3HCrMyu
VNwlIZbWADTqlNiE1fabrPeI+U8ZztfAGPm73Y20AxlojMJiilJSDCESyZ7+NwFPvoKKsFuM49Ln
DByKipJA+tHV4vS22AbGNUVJJuZx4kHbX+sewXWlLkCuzyIFoMHllz1iItLAJ1gfOcJyox06HOOk
lnALbhPPSNfZMwf9YSvRmaFTSEsXM3rM8+OphsGAqae6QAGDzMIrO+IxamljCqX2olqj3QT0kZT0
oicZcuDhu1ndFFcXRMjF7ztbngbJsPWBt5zlgoy/HGpR6fv6+u/KpPqOhyGs8oBMhyz4eKsQTqO0
+Xnm+NzgYTmxElcWloN+WcyeaSRSl7U8CzAUNGvcoGuQYYy1ebGH7mDZewqqdVLWusJI+1hXkhsp
9YOVAR+fKQqppppofTT/6Hlmq3l/C17FWToHrLXfAKLl9YcbVHCsQRnDG8zdaN9L7egjbjn36tIj
3Y5XxUVLLnCpgiScnlez3M79Am5fyDwU637YIiU9z/JIgtM1jGCB8Ozi5czLSVkmIY2rfN1Jub2M
BSmWjhkp0TLBlTP4z41S4Xfr7tZiVzSTH9KMV7c5aHJSB/lDDxAyugQW3NuZ0ZRlx7uNHpwO2R1G
CJ9Tcf5UQWpa3BLjwVKNp8WhhcAEPbfsBkmhPxs9uEuV4yUdrbDh3w7zqYyxkM/+mxk8KbXwMnyk
qY6BCV1gh2eTUX2J30jE2lGndv6cq7clnYT39pTU+Pa7ZUxqynoKq1DnaugAohglfBcVx+gnhbaN
v4bu2t6MDVzSCV7evaqA9AgRGanlVpxkXSVfmeMbHC0IZ9nZXAOVtugZk44ImNKlCNXvgieXi/Ox
k7pIXhVq9LfPd6Zb2Z3zWlNVUoME8EXT1C/TPpANONz93o7Kg6soayl1CjOuCZ7PgrXyDmd0BaFS
99QkKhLtz1/GqZGcg8UZUa+VGEc2ZA7eHNWxrcB1QXRbZJkCJDNceLyLneeBdjgg4gs5I+yFjnQp
sHZJX93dWZkpihp7BoWdQt3yqKo2NUrxdw9Ter7N2Pz0g9hkMHSEfgbIUFX9RYQPgIpGv0zwoGGP
dZn63WCWzHmdgYThYzaChUSJpFjOYK9d/+SwpRMdsEQZ4vu7Ctlt6vrOYnCuFiPEANqkH0lRQgKU
VtiCbWxHxLCj+mZJIZuCpD6zu9ThfFUj2Wlkhq+3qjbTtyXVqU3/47SuA+X/1maR1Y394JWnVEKQ
C14ec592qJD8d1BBQvcScZwLxWCqJ+O936XVFP2blULcI/RxvnyULPrANmlP1txYr2Ml2DucU8Je
vr3XAtEOaD7ySnz3aHqKeITLfn7tEftAWAHVniaa4beSO0LFAHWGrnAfLI/iLdt+zDKX73U6R8op
oh1cZdq09Dr4IUPLV8iHCW5cMk0ICZlbJFcbcVIvWvIXHsaI4WcXLn5Y+SdaPI9ldQ5RJ87bmjdb
fqKOJSMLcHwvHYCrcUY58QyYtT5qKqHppu1qI9XEo4Lmvh5dt8Pdunpmitu5LFIspSFHH8wnHG5h
c5HFhqDsm1VDHQhrpXqJT0Y9H/E/5L51Ugw/hsu36Id+wkV81ob8LrBLXMy+pqb2JHecdlOb2vJA
/JdpoyQBUXoYmMawL6UOFq7DrLiV1fY0GkbIEmg1J+vHGKTaPGuhcTAKZas3xioeGkXHfdWahMS3
3uSssks0h/fIONZStBmnTI7+bDUdMN4Ntrvh/t6r6VgCX0VqqEQ2tPAIe/YE5tQStULM+MAHk6D+
ZzzLsFOV4F+2cgRKUCJwAm3TDVhaNOdcy6IgmFTT8mfiDxgaC0Wb4AMy6T+axhf/wQXvsp52vS0I
qS74/6xRz3Qu/hDd0dGGlRtbFImdNaXMMRkz+kOShXKcD81SWoW5vgLZ9iUhSRArgBr90dWQtlCM
Vr/sXMXmT0nn5wQ0tlkske2oB+c/ia1Fj3Ycv8oKQSvPaXZCZow3c6TbT4VieVPfnQ7/x4/E/4c9
JH5SYW9SXOwKIfZzBQdjr8h3gD/rCgwXQOC+ZfsvgKV/h6HSSNQWLmhP4sEETkGxu56HH4RQvAHb
svOyztFW35a+bJK9ceyx6emXHSmRcB6X011gxnOOgXpNpRydTMpYT91Gh+37pAD0MtYTmkdH0icC
ytwYPR6sRlaxq4sWYRgJOh+AHzpEzgL/3xlne0KRmTZyCMblFBmMgc7X5S6w9kq7wZJ0q0u00aHz
WqedPd9URtIRI5CPXqvvGywMJ8WGrLfIAVgvu+6p9AG4N1NmVmelQN5RUyjhyFrdTtYYwXvU3gRx
inJ0LA0+/peJyGOqkgoi+vAWD84/6vuuvXuZrAruPAJxzE5BxLCGZ3szlmvsU5FADrnWE94kwuxr
JyM88F/BBRxibjieh6ETIgLpWnvythDBBKYJG7nzEHI7fR2tEBUDaG682n7OcrFqNF9gRSoU57Df
JVs4pF+0qYgucbv+dJMT4IcOGqnl45uI74q4Qg82lRJWIA5/q8j5pjUsNv66gIqY4P/VElc+Zhdc
N9BtIpFLM118gGxnTxab2xfhZoWMVFvX1g7lk/U6Tu2qu7/7qdwfgBLEoffPYIsPaUpK6YxH7Px5
nywVVSuCPi0ccJd+zqRUQ6hPA02CQq2PHHKU1ZUddIZclvrmmGCvjboVr1psLW4YoKaXvQpLA2sj
AExSKVqJb1oWaiNGnN8zk02d+l6a5yAtO0SMi1HZcjCgOj95GVH0W1i1POz9JI06DGXhoTXwbp6H
RLv9LaVMnKUsryF0i33mcVUuPIbROM3fQjQ7KFS0Bhu6OPJNT9m1Lrq55U8P9WAQGy7kJVlz+wDq
kfeKMh7Z3YDqhCBDolwJrjuZuY1/PxFcId+UKcZbUGy4UBs40wFXUxJv+xfxH4ICaqKr2E80QHaB
NK9Snq3DMjkoOyGgH82VIMAQz0LPrQMNmhGFLWHo2pF1qzy9eRKf0hwO8F38s2R8KinaooNyFiXa
AV8XMgoS/8ioh+kNLD00vrTrc4cGXVFe4i3adyAKEpLlZK5vLITHYUOH8leNUWtaAl39iXK2uUAU
1VjV34jH7wZPuqQ5Oeml4DQT/neOzIYaodLkwRKdiEvzdGmPmV3G0rVaCPcFHErhVSto2HEOt0w/
w3/KhbXHVdxzNn9qY5NUnB5HARlbAG1pV1yFRIeJGw3OEuZuxoDpnZQ4FbtftQTjulKz2wH4dJ5r
2LMZLNhesAMGFsLiKpbbK/F7Iyu5iq9W5wjUFUQzVvRkkZuAtVJb+88kn4Oy8Y2C5s7Ri3KN/DTP
AKp+lITKk4P9EAE53rSyZZExQ//hVMPLNoiwe8+rG9RKDiDtUaUjE+lvMLojMJzWqI8Z8SV3dgTL
Flm7F+z5aq05WKQVAroSs3Lgk37eSKCPPFPz/5uNOFQ64QAuuNbIrdPdZv8lEcjcqaBe8gyV46zb
2ahV/GC8u9d7q+xDqnTEwlwwov0AhzIh92+X+GxYo73S6LXIISZvKyUKjX7i72r70nDcJOQnZZdB
jYcfFsrW8cSY2IM9hvAW/V5gC6/TfyjbsvPHfMt4rzq17QQWmr5gixiRJ4UlqsoMluWWVec/USqL
8Wo6AQCzrUaalsq+LnKaHGp8l5XdJfu/7SpWMH5GxQWDHXEv1lJSpKFsumuCMgB39V0zCN5vSeU6
gfIf0gHkJUYbzF5w0pLL87ftJhfSY/Ka2BfVphfKT13iJgUt+J1+yCc/rYB5ZTy5DIV0hKksKdBk
ltY/aHYdN9pjjSyQT9Yiu8r/uFN8Y/Jljoy5IBQuQW0l+WeQfVcZU3bwt33UX3qucVbB6Cnja6JC
oX+/50QotTu0ve9lPfAcBOtbRZbRbVFEl6l5d9cIH5FJdc+U99YJRTbTTN/XCWa2bKCvIUTy9V3f
upaamI7cd+LjslrxPY/58zHMSfCkamw1wd8lsW8b1zTO3wXoW20jw4RVngRdVc9ckJRvDVOmb5QL
UZSy1jW7IH7c+NwZRRMtfULWGnayJQknI3BjP5jqEwEAZmqSwO8Hrp6rom0jMJCLIOithFP3pGoL
FGrxBQlTrL2u0idfSerJvs6dQPDTz6/5PNT+nEkM7FBQhsivwF8EAQrnQ36s8+OpHJwGQMST2dzV
ndb4y/5QckBzpC24ZJPG5UyUhwkD9cUrIbxgbFv3hvCGFZ2ageCX+6SZeFPpWBePkeh5a2E7v5Px
FTOuIEYGp8xFBXYLvmPjj3y33ruKy9RRzrYwy4wwLeiTA/5SQtHWDMfc/G7DM/8k0sGn0eLMO4DZ
acYAHw/d/VgpGo+6NQB6ilv81DWpklRSat+OX+eDrKQZeb6QZZqXRprpaTAgIaFznmaNZuKQ2K4u
Yfr4vxSPlp8OszYMxN2dN6623Idy26xYBwYLgblQwZ8BETQR0va0N6preC8Ue33prmhav4sRdqrp
REp4IzGCk24FOEObLXFAnhl7EfG7MlGVa3jl68Lbh8dKGt3ZUx2RgKkMjhZJTqk6ilW3ksiyxt7+
ain5+qCUCSaA1TYYBFKbLxg3zpOz3ev5fd0rOTnz4jLMde2FzgL2n+vCCTfew8z/K+o+jzdEzMci
U1P20ziqzN0lJrx5LAC/p54G6ztIFfL7z1Fls6hs7rvdmhpCb5BPHbhfRYLErSLMtquRcaXopoEo
ffzc7Mr8ImqWd1UykpyGQOHBdOUbuUP42iowtiw4Eu6HBaosFNqdNEHYf1UI3Mzhg9JoT+CDy4hv
1A+n3uTDN3OX2d0NcAeclHirE5/96Bgqc0I1rF9BApGaAjWlflcU5xRVaI9goYpYfajcHUxrQBFR
etE3zqap9prYXULbbsCL9ODmSZ8/+DJshzzVuLTlZ8jr0lkTjAhy3VH4JSjGLF4q1fy1OdMmu2j9
lI7Z+cnS6ksITVxtGEJ/oJ9Kn9vRkyK6V//TDnaIfruCGKnNTjSJ2ZKVO9rz6ug7/VIPoLprMj+x
mE+KqGAmRIGiqIGUWNaj98gCuK3j7gZdA7heI2HjRV9AXznQDmRwOZQ/+rh7RqQKuTSu+XtTRDNQ
McudRtOKhteR8UDDOAurBQLwiIdzyHgTq8h5cZWxTO8Oaqh2ROyjfopTeq8Dj5eMYVBf3Rk/06s3
pA4gaJZojWRM0kXe+d4M3Ca7OYdAGPw8fHhUEa0rs2e8EZSOVmZvYLjPfErw2ooJ7JZwx/MGOC0L
e6/ZEV/eMhN4hwhklb50tGQzaWNZy2d8LBK2Nfca1EeK2/v9vwqG/8icBWV+qiBpNf9rAgwQkANJ
dxj3CHfCqJZ7gZJ6UEj+TE1EHSIVd8ckZM3+899NXtCAOngsABCGg5NMwGMu9kLJknwutb/izUTJ
Kz5woy39tUW9nhrB8LoR5fnn7DaSS5RNqQRvtkC94gxU99s+ZorxXBDWqklPj3Vs7tr7VuDDX4tJ
1+iyknS/i+zgrPtgDbSO/rZ5QsqPIR0mRHfTOHN5E0dRZ/BqLWETLlzTmLLplDyUHRmlkC4tqTZ1
CpMrP19qhIGz1dhzcMpYL3T3gRnYH4RhtO5UtZ0iQTbzyeRbzZJ20KYQlxGRqs+hel+izRo7FUKA
TlRJp2DK9i0b2KRB7LlPcFwd2+0aa8gnwRam+ZNJMee8q7sWO+jycVh+Ob1BsD5cZz9u70tW7h8d
1UjVoG1XS5VmtqjbQdKHEewc7EdNQu+ZBpsA0cgJps+ASDnAfg+LSRe3NlqqTtLFDgrf4Qw+32Ra
Ob9KVJ+XY8OrEv6nattYET7yXhH8uK7K9a9EvcQh37249h8vMl6YNM7K2RaT8UMVRIOdc+mHtPfS
+v/kYgARhiNwaBozTFd6k5+By8S5tLkbQoLTNapQ/sr/T7Wg2aw2rZCykrXrqkqY0cPuzF73Aft8
y0hySkU8N/sDw/41Ioav9BRgOIwpUjb7bWlzuMJ0vug87CzEetQLA2Nt1m/dnmWvX98/89XQf0hB
WyNO1BfF+Y4sTkUlmx03aDqJcmDMLUDSYpSCHU3XbtVxLHhEz39o2+iN+GakWv1YVHb1mzl9Jrq2
GvSZ8/T3Ww/kH6ENj2QZ26REI74kacAOmkMctPbzqmBI7PMIuPHM/SlgZozCl7MuIp8DMdeQ5FPw
CA36Rvp4yVGFCA5WnFe9ABkuP53N2FQBBM/ujHgotV755R/P5UeEEElNWEqZSKvV9+A2eCkShCG/
H6PzAvK+6y4MOfdeFaZsxlfFND+DP00h6mOzMiCLsj+qCEiBnnAf+KsEsGv7M96RpiB0zOFo0l7v
8el32CwXM0J9cx7d2liLJxySBRgIOm6qsBpWLxWnSfboKBICS5HdzzI1rayVoDj4wMb29YD02075
Fqxq/qXlG7ehrplsf+0flCwe621GzeZrn4KS4rgc2quWu2hbwfsh/3ikGoTbL1oz7JuZBiAnNSGy
VpKDXYHhbsddjy4W1YSwXBD1rMeVm7glxDWmnsM2X0Xl0L2Cf5fa3DyHjk2qtjTjwK3k2cvRrc1F
H6mTV1DH0UUes0HEa/SccV/obqo+hDFwrJcKFkvKP6OtwHB6PfmuvTkEUwmNoaQXo7V3TblvCOBg
eLdCH9I4HSgMG0429/eak6eDkezEmeUFkJ6CIer3WsMGo90lrYzTTf1PlJgExDC0ZFgB03t4jC+x
k+pVOUfDRMKNN1OvmWIt8wFYE8jvCM6ZATvfRzv5QBsSapj46CbQbNDC2p+VWcLBf0fVd/wQ1tj/
41C+PfIEUZWlCfu/yBVmcMZjjh0FQBAXDFzg3OEPBZl42r4GCmSE02mMIwqBR8J5H3xfGa0DJtvh
KlSRluhlhzErHrhbxVR27/Qg7UzBkbknAJWDw8mf7Pgvprmmp6UsFVz7vaEpGYf2n2hSBVT8C/Rh
RTU7j2C6YcGpot0j0W6jSAmykb4QSXDISYOS44zyr7OhlOeevCy4JvEdNeYWHl7FRzqvA3tEF91/
iPp1GP2uHknz4VjHcu6m1eUud58QtBJncMfUreEpnrywFcqQBNNPEsFw+0NBy5J6SNSS+3heaxL5
Ja4hLZbWv24IfmEh8TZfblwUdLdHbMsXXGZbo+alyvE4rO0fToWmWuiRttJaEbp+QZb6zp4IB2Sy
qaBjmD7TddDckQ0MT0tipwxK2sAJF+qQ7fBWN7wCQiX+Kxcl1q/IGVsh6rQAAb1xwH6HMNua1Qrl
NHDfjKP88saMiH6UTaDYe42TFoXrZUjd2I96h/G55A51OpX5w6W+eEQR2Qji/BA5de/oKI86h9zc
wiIXRKGUv4Gh95yGRh3itOmcNjkcBeZMJAnuK8UovUAuXuPMQq9Yz1nf+rbwnt82H5XrmWBiTdn1
eY0CtP5ADhZzNg7KCTWro5KKORj4XAWYWE37RX1hqDyGovU3gVlv/uRpACE60xqo1CaHcCahCSWy
Erb8YVy/BU21vEqgdHPRwExqr24S1Eqo5UGFzjWYgF2gZyQ/JvmV//yapQmAleS3/JztedbBBrxM
m6BudhSCDQuntqDGT+Z3gva+Q2OsZ0qvJeQoBqXU13mfYy0fVpJAtK6LL6ns6eLd7vXtfwLhTu4d
qSfdhyvJy7rcaSa+9rzQs4FzkN+qEqoh12nA+Es5qjG3OCbMZ0TBTFm5rlYgEUPO/DKN+RSARwIb
rxbvJT6mUT05UiZmPzlYb7LYFKmdatI/vHPt12vRjcnLvq8sDrTKcWg/jmi8ZKhpK5AUPwPH28Tc
XlrnVsBlj/JZnHpIZMkN7azXMVs9Ku+fL/SiFRuPDZNQ8oSzIWz3m429Ic75yL+qqvqdTaLjPX29
U7mChNk8wl+R9T8I5T6lI6Ssugvwsff4wOkoBZGOSI5qY0Rhj/DsJE1BKRz4P3e0p0zPkzi1RBp0
tDMUK5n5GV1IEOkiCir4h8l/IKKz7e6nSQavAOW6qc1TFtoS3UDqcxCL+zIbatfoAHgmueFh8RSH
UPUzDR+H3BsHvZkLX27QeVaZl7UBsfZLKtkskPA++IEzSWQZ4g+wOUUktOswArHnL+sbzerslxzZ
ENm+dYdZ76M/XYEhdfLscbpa2PQ5Y0pYANJmtuMh1NGw/hKvfGXNbxMVTI5lufd8gdSYdKnUpxIZ
zKrr4kS0UpRuGtRhCFrApvOtXoECPPx8KGzkDlZyONCfDn1/f/6ihtnksFIDv1SCRfce1C6pgxRt
3TBIWGKTBiKM05LuXhaK3Uz4+zplHCkxk9xUQr5Eqoeth6XVLwKf+cL9wLh2b5y/y5dKvo6nTlSJ
5zMua7fwqL0KW2JVbMmxfTZOT940znMaFHFfDvPFoe3I70aSS1i4j6m6dDn7B9E8pJcKBdjpfEFr
KHHJ26IE8JNuBsdm1fzFOBwP0zFlD/TTahxKiNfY9ehHF6Kz9vz7RbQ2oRywbPwT5XfYjs4pLMGD
mLdOxxmdFC0J3339SKP8wtEHtnzl0TEllAN9MTlcRm20RWkkKnMOxB0g/iig5FyNL3BxrmGhk4r0
mKglRhPozznKnDtG9/3DATAWBcIdIlYN7m728pTWTsDv9PbfLQxpkZFXtU9nJ5g1bc0ND5XgCmuI
MOypo61tu3Uufr8Ul6m3huTMpyrsvH8P5sNjgGCNF/KWvzyJZ2Qdyl9sP6X9B1fFk7EbO+nYm/Ty
wc8n4kgk7Rubtc4Q840sVWRhDcTbq5e484q7O2+ObzdRCUMlPUhNktI4DkHfpuawPjw1cx3wVKRp
hlalES0h3FAjkZiRydaGmJAAVEurRh/IzRuRBVMZzyequPi6BG5pt3EqDh1slMXEUSmzJh6YKY51
N0uNNz3qvqtEv39dCa7FNCH8nLrM6k+t6J7H6bb6XcdUknnWU7XUWVczQVBtWUqcD47T+0zLmPmR
z/xuwD2nobndqsF9TgArBL6QHOMJfKARZpAO0eAQ/s4rv7j+YXbXbymqejPIGecMnEtY44+qCvID
yQM9N1qU0s6L/UtPt293hNAVm5WFKoESoyuPRDjmgBlwER0YhQPiVhda701Ma5aUCcb1ALamNPo1
TevQ8MVljnG7swm6SYL0748DdPv1I8mRiJIHqY3pXtgdIVF2zIJrCJhjom1cwjWL+qPooObKT/3F
c10hblUUtyMlo6mTAnz1DSfCaPt5b06g2Xav6YltisuDEzsvDAneuEjvtFZ8PSPLs/qGxPUtHSX0
4m3eTPmjEMppBMPxZ+ZlX7d6aY/5mT3UinRcEgwnWw4qqlXfD/Tgajf2DpD9J5NJAcSN+Lgz5KPx
lhztakzyXM/sdy3pfGy8+BeWzHslhu+hIi0xgRCiuw2ju6LlqOdXAgAYA+Z3q3kr1KKcYSj3a7Zb
zrInJRd55IkvXsPcy2n7AQCclk0PCnBEuKSEiKHDEQBA2mVOYb6pTejmB6mbKmURp7n6PZs3+Z4E
RH5bLF/TtDc5oB55Me7y+i+tn0zE0yoPrxUHbZf3UT3hcCcqn4aa4vYsThCbJ+iz5P3zyOM3UBrj
hrwVD8gYEvGh/fzKLJL7gDpBIJvrKmIZXDzaO70zg+ZHnHgODpNSlZh3oOX7GEA6Z8aEhULTOhLa
wjUAOTW5jcQZYTQt0IV+mW9XYoI13d6RYln6d+WP6VZmQslPrs3reKXq3fmKWFX8ICf1NSI1907a
rjvu6xcNOxO2CM5DRiHaQBgrT7o9GYk7LMll5P901KA+gaVfyIs=
`pragma protect end_protected
