��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�a�ȝ��j��^5O�w?�cF�9�X�>J�l�^#N�c����~�gZx��A�->(��� 0�Cx�M���d=�xK[�>��R�r	�7�0�iMw��%
P�/��< G����ő�O�Q���WDp@cU�Tdԇ�b�>���nR1�n�)gA��Q��Nr��9+Ȏ/���i���݂b�A��碎G4�[����C۪�����v��T4w�5�.<��W�~�iDۆt��<��sK��d�hI���"⃣�+�E���K?�r�˘%S	��sK!��m�>�t�!\��.�p�E.�#���P�?cYs����2�N��ڵ��]�\a��'6$�u1�c|ʵ�p�.(��hF�ti�>�Q���whR^�m
=��g|�������Q�,��\؊��`��J�Y���4�@��D���瓃�H�˳2O1���"��ĳ�z')V����eđS��__����5В���>���@[��t�]�{�[l���N�U'�JTrʇ��n�x�19��j|��|�6�<���~Z���d��x�U�5JQ���]:SM�/�4+m�n�d�� ���VD�Dn�/���;�Ė�'���D��s��J8{��,��#J�S��@���<^�_aM����6>�G�\��-\�*��
�dC7N�X.�Z�qXX���F��
�WÆ�/��I��sيA7����D��?��,3��KRH_'����2��}�C��}~/g�"�V�����m�uo�BJ�f���1�_M�B�h��'�{�ӦB��E���I�h[;.9V�%Ţ*�f2bu@ Xޚ�@&"�'�[��gǢ�&���⎜_'+��=� \��y�*O���w���uzf ��2�U��׫��f&��(j��zX����G�>N'
���W}�ӯ��=s�I�Q$�$�����)S���:,1s�f�Ţ+%�,�O��"�]��Y�8&'������^��V+��j�]�)�{=��$�m���|Ŭ�+��,ɄWk�X�Rwm�����[�eQg�D�ܩw���nb���<Β���bx.���h�D�}d�"�����Gp/65�('T­j�0���P2�?j������=�����.)�X�	y�Ff��c�/��������� 7Dk0�=M��&�;�AF��r�N�.ɛ��`��(�쬌6wZ��1�Ӑ+3d���	�O��c��|clq��{�gU�PP�@Z�5`����U.U�s�1@�N�ZE?�/a�!�R$���݁klt��~nm�4�M1��7}��BZ7W)?�qP��hv��S�BFi�������]5�a�N-:'��F>������}��VS��4����Y�»��kX�1�[�{E�*	��Xos������[�����@������Al����5��F浛���U/��"Y�j�C��W4�Ɯ�����E�{"�fCt)�3.��S�}%��5l���>���'<:���ڈYv��*{�Rmޞ���9u>�~���vz�����a<����k���g�����V�Uq�G����;�VsӦԇ�"��kO$"�e��;���Od?Sz;��c�𮅺&^��3i)ڑ�*�u���(�`��U�W�dTB�C����`�.]?xG�CA!�Nhl��:��Q,/#$��� v�jD�d_��R�\lxm�}^|68h/�i]�k\�h�l�2��o��I.�Im�EG9xk��ѽd�8ެ�U�@=��t��f��S}��@\��6}������ s�B���ɜ{�F�&g�
�FI0�Ǳ"��H�zH�j�l��=Hq[�+��㿲��ċۨ�\�C���xƕ�h�* g��b9~C�ޘ�Y�����Q�|>���R�FUY�kyŗk'%b�Vn�y�?�_����x�Z%M�S��Aj"�2i's��g��5�|�_A�ظY�S9IL�r�����j��C�"Y���n����d蕖�,�������Cp�Me�mi:��4ʽ	��7�^2i�W�7R';)�p�6�--�Ʌ�"���h�v2ѵH�i�}��Nki�����Ys_+B@ɟ�Y���� �nv����.u�8�}��}9�T�q�߫��*��zx'���2�ޤj������?�7����-Ic��MH�u:�JL�hV<��S,1�bSܗo���D����
:� _��!�;��q=�.�;x���[�[�$^�O>�y�.�U���+3u�`��D���ǉ�>#�+W�wC;��1���+��Jz�u���T�s&}n)[*�9�>�ِ���X���:W�P,Y�A��������i�⇄{T�i����R�ճ���Y`j@�@"� �_��Gl�G�	��Y���84MkS������R	#�����C�1إ��9`�T�خ�v�B��ʥ�����乵<[��"��b�#D���K���W�2}W��>Yp���6��X?<t9|�]8�u�kĕ*ܳ���'.O6���n�>1�F�f�z��i�_��2VSÜ�ޔV�:��gm���j�������غ>���H����!Ύ9[䜢Qc�E��e����yXF��v��3�>m��/��_�m����碀W6<�Og�����G�#�0;l�Y@�:ue�U�̚9��x�Q���tsT��,2g�w�(����V$��{0�3I�R7̛�_��DH"��b�Wه ��ؚ|su�z�;�C�wͤ��Fue{�hV��/ ��x�~C���~���$3����DR�>K�dF���: eOt�o�3�Eew���\�sȻͥ�w�"K�Z���jp6���/T�vPHrh
�G�Xe��φ���J�A�ɶ���o�y��}i�$��_{����U�>To�]Ri�\��]Ey�ٹ�b@Mߝ����@��l��gE���`����O{�qҚm��Nw��|���Z�KJ���Z'�]ܻ��$k�]����D3�$�f����\_�+?�)�����5:�!��9K���M�Ӗ)��<�S��N������V~����iT�-舓P�l%����Grj�ĸ⣊��oP�<��}�,~C.�+M�M��\���.R��^+h�9��-9J�b5�Tڹ�/�5jMj��:��D���!�Lx��3���t]�H�)z ��
76��NaR�֬%ʙ��Ȓ��>0u������;(=oMќ{�����������*P�����F4H` ���/���c��:�I-�v�����2�o�G�,?[<dJ	��n4ǾP��081G��*��n�����iԹ�!8e���H侘�V��G��7f��v��{�S�������
��r`(r��8A���{� }�v���+E1�jϢid$V��Q p�Ɂ���H3�#h%��M׿���˗�1*���
_�1	z� ı�lG��&u�:]�x3�'t^1��̓֋�g>�i����M?3�����E����%�S��]��)��j��zGcT8����{��~07`C���E(���E(y���)D�P�J��W+YC��U\�e�V�*�@ݐ�smp��3���f������G?0�	-V������H�5�~���+1�w�Q�N�
��	� �-���⹅�7W��N�-ȕ�Z����;d���C{E��e�����>��"�v0���Ɏ^����ᗝ���~�ʫݏ\�E��x���Fq�+�䝂�ei�A�겛�r�x�7�=���zQ�<��&�� �GA���dyC�+��;���[hwv9ڕ�����'�%�a;?2y�9���TGC��{��	͂rEiF]�+��r�����;���d���SJ_��Ľk��G�mpB��1+3�%WF�tN&��3NmQ�n�����h���z��]̷ $k��̬JE��?����'4+.�R�i`r�9D�-N�z!�ۗ�`�n�u2�0�9&�����ץ�l�iǉ���'ى#��6��F?�p$D�{DQ�s�~zC�]��/��7�Y2�h���*�;�b@�up�3���/E��*���ԧ >���*�#3�����T8�9��</Y����ݜo���w�d�`~ �}Xx�ۈ��OH,��9k��&���}Ӝz�WuW�t
I����$�I��u�X��i(s��\��U;.��$��Qq��l'���AlkL"Ʀ�-�g�pvc���L}@�9h>���(	�v��\J#^|\<AЧVx���a	AЕ�<�zѦ��~>����5��~2V�-l'o0��!'5�Uz��-]q�ܖ�h�}�SFx�����A�i�m�-�I�-=p�J��?������&T.y}�o�b"�������qkc�M�$3\�K���;�&�U8�6��َ�ޫ�[F���ªn�N8�:PG����u$����v�3��y�?.�ywC��� �g;�*+���AN�[k�ߨ>�KL?+�g{�Ō��K^�
 K�]mb��.���-�2�ȔG�����}Kn�����I����VJ�k=�Ռ�J�{Y0����Ƙ��G�>�@�jTѢ�U���H"��,&W���,��y/۞�Ր�wH����!��z1����ý���I��bj�����
��D%J��P��s�!��L�V�P�f���C�|��)������oZ�}R�EGrM��P�+���1M��\�V�蟄q���'n��?��4͏͚��JU�l��l3d��^]~j0�4�ii�\�R3=�kX���pi��$~����x�镮w��DpDA�#��g�ͦ�7�0G�F�y������F��%����p�u$�H!�S8����4�\:t�4w�A���\f!�'�{�E(χ��_���� �Ux�-��Ӏ43^��6��vָ�-���C�5ܰ���JP�%��%�1m�.��^�+���y���I��i�{��K�};��撱j�oB{ǴPZ�xV9��3\U��6(���?�6>Ϥj0ԗ1C���O.�X����D�2�9���Z��엁�!�ܘd��H%��p�������y�W�n9��Ε�� �Jg>���-�?YC�H�IHtaY�"�&�l;9��p��:���O��"s���]��L�͵0�� ��lF�����s�E4(Ǥ�?i=6�y�x�.���U�R/<�
ܯ�.ѽ�� i�1��9DS�����G}#(��);7R���d��9RK?��R�]�o1s�h�SdD
@�A�Oz<xrnKxD�%�AX
�����!�Ơ��[2c�t�y��@~���2����Ti;��ǚHf�����>',a�+�<r~ıڴ��4ͽ���Ъ���w�U�1;Q+�-�|����$���ܿ45����g)�7���Q��Eg$��.ʐ<Y�[�ƝQ���T6����J�PO^'�%��;��2��"v7���i�D���3��2T�&W]�Í֍��X3��^���������?�5Lc����Ih(�y����t�}�C(��Oע�w�J%���� �t�|v���j�/��j�3y��iSZ���s���M���3�6�I���[O{Jf>֞Գ�S�5�	�0wdZZ���Bp��SY��e���bfr���2�e:ֶ�x�պ&){�I	����O�c�~~>��$���s)�e�q'��7�ZЄ����9�%g���vJv�Me�?���Iݝ<��7�r��� l��b�M�뾛��*�\7;�����2�Ĉ_��s�����v�]����^µ-�,�F�~ܭ7�գk��,��8�Iږ v�sMJ�I��}���+=g.4�<�د:�yX뚝�p���[�D�/ޣY�Y�d7Xf��Y��<q�owd��X]?~�������Y)���bVKn��I$��aq��|�i�s�EP�������"�ȶ��/O���䭋���wZ"UH�H(Z�6I}~��Y#�3v'ʎFu�' Y4�F}r����c�&L�?^!DN���]�vKj����s><'I��5၎t�95U��V�W�QeY"Vfz1ɱQH��f��˟0��X��1'Ǩ��j(�A�+%՜�HN��us���0��[Q����f�Y���X���8��ހ��`�w�q���p�8��J���[}�������}�Ȅ�m���S؆:�l�İ��@G�0f�t�(�����bX�IM/�2>�|�O�k�/�r�N��#ey���`}����G�r��[X�?��ߌc�j<d�}��Bb������#�f	9_�Jlrի:�	�Q&�W���%�	���10������jc�+�^p�~ ۨ��ن�����MϏ�0��њ�&b����5�3�ut��8�1_HR��â��/n����*�`r�W/������	W�5�2�q.k �8et`ŵ"�n��	��S�Xn��*�V`��Gm�n-�ʝ/��m�;)������K�u���&��Ŀd7���6��>�$��1��(��y�n,�v��+	��|5>zXY_�)�v�9s�N<�=���RI���� ���5�����D ;C�pZi�J(�] ���m~���8��`j@�T��]��"�f�� #'N�¦�$�l36�^m��2�f�|�<A���~�3�B�:h�޹l�!�ʍ���xdVv�������������>ݍ�k�ǿ팼C���S �X�
���r.G�A	^{�<5zB:�ظU?:@����>T7�3��E�Nc�o���fGKUT��F)l������[^�0�u.?+ެ_�ϼށ�����>S����X|^%�`��Z�l�C�{ v���H�������e/�l��1'��8�金�y�U��c�|I�hTшl=�ȴ����>N�+�X?����:��� _@��w�g�٦A]�79���}��t�L��Y�����-�R�|��&MF�z3"g���D�w�c�FvC*�
w�ӆ]�2����^�D��Su�TꟂ�	��B*��1�v�\�j���������|%B���2��:�R����R�ޒB��l�Q_w��d�$6��
�<�wU�q���o��T����� T�0���x����*Nn��)*�B̤��s�ċP$)�j��캩��9�|�ݬ).��:�I�����+m�K�&�jЬQT�1�12��8�<D��zc$�+�A5��ᴄ˿\w?'ؾ˃�+\D� �V�A�pW��Zd�Cs�_!���I�A9�&�wu?�`��W<��z�18�n&��raA�WF�%��ҭB��lԉ-�B�� ����8���9j1��R��jjR�k/�3YT4lI�p��Y���C_�㢊\M���2�Z^7aNC�+��6���F"~2?�c� �xٺ�-À�5��T_�R=|�j���z��t����D/�en�����h�Y�B]V���m�8���H�\aO�M*�5N鎳��i�t�\��^�­IA��P"���{Y��N�v��m5�=��}���<E�J��zE0�r�t�W�!i|��KF�A]2���4^aE�"�k��#�Ӯچ�[�W�<�:�ܞ����<ch��tQ	���p�%�r��ݙC��y�������;\�k��^ �6ѧH`���M�h2X蓐7Q��C�!�w
~��W����T�.�4����^�襧�Ŀ�um�^�g�J0�b�o��ӻ^c9�9G�#��CT������o[�y���US3m;\n�K��>)�"U�2�j �
�8O�㝌m��^Ch./=�k%�*u��&�$5j�1KrAfŇKm�܋�k�QJ)}���H���j�m�G�e=�d�}ǽ��G�M�NLCw����J��k2A\t�5���3Ɓ��j����:'S���p[�#
���u�I6�Ф�WP��H/�����9���,�P��+5�JaiȮW�xu��(M~�)s��L@"\t
	!�-�a�'�a�!]��F\k#�44{M��
�;�����2��<�zf���$0S"E�aRQ���� !!�ίM,/�p~o}�O�����^�%n��vΰ9R�/���>���A)Y���C#@z@�����e�&bsZ��uP�3�YnA� �@p�J��.�г���>N��Ԑ��<9d]����Ј�M���p������6�Q忟5�{!;��bj2FUݱ��!�hB����R�*y���}���N$Ƃ�u�M���u����zN:�MH4~�)B�%�y<��Ae 6
�jpwFC�\G�	�7;E�R�-�k��K�⏭��])�\�T�P+ R���93s�7|�B���¬�>f��p
x8�P���bj��]<�Pf>�+�|��QG�)pW8%�~����y�@��W���b�x6�כ��]{`� �N_�q����H>Bo;i("�0ܣ
 "��u!�.��JI~�ƼL�Q�q�!w�U��u[7f\k����X�&�n}(��-Y�X2���|��Fn�[��a{97	ߘ�s���L���7�o��d�c��&y�0�3�I��v���;�] ъJ�}�?^S(:[X�*�!�s����S�(:$G�_�:}��nI�"j���*m��!u֫����d�����{�}��F�[ը�1�Y��@�n�ۗ�`!oi�i�υ��ǐ�k�_)&v�@h~����P�4���p�j��.Vb���S��j�Y���M�R3��}@D�Z��\�s�@L��M�{�1W�� ԟ�G��	�E�z`+��ØOr2=�l��/!�Ӝ��[Ԗ��#������(�k�i�ڂr�I�23�):�sɋ���_ ��F�(m#�<��VZ([��t���ӳ�-nOۯ�[��FyS"����{�o3��Z$�'���!�l5;A�	�S2u��`���T����_K}����C�ӝp��>hi�;nt[��q�e���t~G�Ib
̨��B�S0���"�c�S˧M)�ks���bn�5T��5=6��!'̊h� A����;��[��d8u�<�����#!��o	�����E����̎L�&%��m(�������r+.�����.F�f-��$�$ g}�QE��k�v�z�PER���n�����BW�̶k:
Xk�B<�f{�&lE�̋SM|RΪ��~aǇq�c9�
K�W�[R=�/������9Do�'����p9��z��,�"���E�6ɖ 4������W�fiJ��Iu(
��"�½E�O|G�S.�#��x�ugr��8l3�+Q��8�$�m��ى	vDQ9������+d�Rg�g�
O�f��I�G��J�!��PE���H`.�����~z"�iv�����|W[���sH�����sk�g����g��� +ݸv��i?��>,���u��Z���_�S����(���''���٬k�ӂg떭��qV��w�ns>�o	�z�ѩ�v�.�"�34��7Y\�2��T�զ���yl]�Z�eƽ��2!��� ;����88��1Y�cx@����_i����R-�
޹��.��#�V�U?����۰	�`�U_O5e}���fS��+1�N�[&-���܈����83٢�yR=o)&�c��0��Qނg%2�{$�:��1��������Mf�)���A�L�}aIe�n�g!�*	���9��8$ԁ�k�F����%��Ǩ�댛�ٺgL�}�)j���֞�;x�H`T
<ף�n�$�֍�!� ^``��$n)�,����S���FO[jt��1U�5W��R��z�*$��q�j�;^���"0�O�U���^ �@�27��75��Uٕn�@B�^�Yժ2����{�&}�K%��0F��aE�=FĵLJ	%ʝ�|#T*��F_����+7h0���RY�o��yR�츎5�M��N��76��E\I�_�B�D$C_���G�h���n�d=�]DΤ�!�d�Xȡ���C4Y�����/�&Ku���;������J(��ׯ���(
�ϧ�'��a��HD�B��ՓJv��v�\��v�<tZ���wap���|�W�*�*^���:�ݖUl���?��Z�|**-�d>?�Bo#� '��gO�>xDW�l�	^T�%���~�f�GƩ��ʅ�		^�O*�|��XA���� ���u�b�TS��:pʌ�d�n�� G��qY��Z��_@ں/�]��|��͘W<q���M�\)3��L�1
�f~k��^՘8P�@�<ߏt�\�v /������F?b�	��\�D%Juk�N!ADtoM>{ir�=��E蹖1&U��فsG���\�:^f�,r����q�֫�>*�A�%-���Q���o�|��M!�pz�Î�@�E;WÂ�B�k�/���*c���βh?�ث����'���E�c&�m�Ib�j�y}�8E9S��xa�u��А�
FW�|�%��wa���pƼV�(95ª��jt���(`��º��YUnΫ�f��>��V�qΥI�J�����]Z�d��_���	�P��a�)����2�h����	��p
��u�G5�̔��%��~_9��C�!}`1h/�o*�j�O���G�|� �u�FP%Gz�;N{H���ߌ\(��&�A��`\/��1���bUs�Ȇm="�ގ�X�3���Ӆ�A��:t���C��p�"�
�8�p�f'Q @ٕ�kt�~�\���$(���S�DR���!�զo��F�m��`�'�2[��O��"�,��.zF���ܩ�#WSY��Q9l� Y(�,��_]��U�R�_v ��L�^��_b�*O��S�i�:��+~����po���Q�cQ+����"j�� �� ��/���]�:S���v#:[�o���m����J)��	0'U<a�-�,ym�� Rq��rB >`����9b'(���ѡ��93vUW����R-i�G�[6,�3�`i�A�[� �5Ə��m}�q�%ٙ�d�<vIQnc%�g^�9�_}��A)���������'��6#�F4K�Ĳcd�`�&mx?Y��>'��-
a��Q/�d��JC���k��(W4���8B�阎��q�P�D>�Mޒ��BSo	Am�v������E.��	���a,���:�v�r|�U��s��ޕMn����e֜3g����xs8��=��g�O�Y�l�#AV��%x��.}2:R6v3E�k��5�䬎��.��!d�(�t�:��(��)���,Ke��Uv�sqA~�������h�¢�_�A>5�2�TԲZ�0R��/y�m��5B�O��U ����]��D��Je/T����4��呣���O��Q�_A��x�a�i�d����*��4|˲3=ݛ�	��6��~�+���^oF��̽W����~��������z'g�JU�ihˣ�;�3�`v=��I��=V��k�=��}-�8�D�m�:�- )]�>�Tw����G�l�}��=�+d�/���!��a��YP~N�3�XdO#J3�FʇOR(>�G���o��Q0�p����4��.N��A��?)�-WP�;����n�WV�+�n5ި�Ǖ<C�\�Â�ҷ�m�JBκ�J}Y�O�\�HɅhx۹�d�����uבd��U��u澄�~Jn�+�ۉ�(��r�����[�����NξQ	�5�`B�}�:�$�"	*~�Z1�5� e&R�{PjZ��k�^z�A�4-�$��3�+!(�������/�.��B���2Q&�q+�fi��%�4�E�����$C�$e��������Z��B>�B�c�ѵa���~��� a��mmY�	���������؄k��t��|��O[j/�fl�(�4�"�4���A���J[X���!�y^�gP�`ce��H�tD��4�.p��"(�Ǡp�$k�<��H��Q�[o�W�J2����%�/~|$T�y���$f��|�;�B�@��!�D5�群�1�__��0/��0*	�vSt�<��{"������N˴/8��!%%�.�X�W,O���&�P�����}b���Mk��a ��t���Iߒ�%mnUaL8+�|:�}=�������>Y�{R�#��ʥbXٰ���� c���_�K"�\��7�U�����!�Z����d:�'9����g�1�B&�̫uYW�������V0Y�^���A��'�C.�&�x���@���i������Xo�Ul��Ǌ@�1�2)&�3�����H7�?��I��0�´k$*É������Ǟ��?�7.��y�\=:�����F������������h��N.i����xڟ�T�ĄkATp�'K�zf���
��d.םiw�0 ���Yl���@��`�7�9�C�Ut�x�OƑ+�;f��� c�eUA_��%��P��2�j�E�TM�:�H<�yK���l����H/�y�<�ȳ�}4�a��ݜF�!7��*W�D4=��&�	�R�ȵh5z���B�l�X��F�]�G�e�K�R�a`}��`��	��t�5�-�g\f� ��f��z��d�>���	�e��y�պ(�r.2w"_a����z2Glj�<$?h�e�vM=I/�k��Knz���k+��1ݑkW3��i-�A�I:G���y��<>�H�yI���`�`;���n�RT����'���/?�X}�s!>_5 N�I��ӮYS��;>�(wp
���*G9R~��p��w��d�|���5����W����������!���c��1���lXUth)f��  �r=�)��.��b;��U�'�����.=D�O�y�r�/��)`����豏)"�˸�cJ"�&��O�Q�*�į�[�v�� ډ�N͏gP�0�CnnG���D+a��h`8��~|!����c>%�uz�o���j��`��~�nlD�����t%�3�a@}Z#ɻ/u�&qѝ㱽\m�(�Ld�����vdE���9��UɆY25�z�P�'R�7�F��4�%��b�t��<�ia:�*�����x����z"�Ÿ9���T�����o;��������y;��g9��RX��g���p"���ط���髚�7��G9���U":��b�M�x7Qba�S*
 ����9��|��QG�N���ѥ��F:�h����$�
�u�3��u�P�m�R���m��H����S?��<�;��p�K̩�����^�&�A9�Uh���(�C�*��.��ؖ�o��J�f�#�"���U��P0��5 �TU�K�#�ޓ�@�½,�NV�D�Fݥ�k� �m�>���j�ӝ�����H�[�sӳ��wq]�C-�P^�z����:_�-rU'U����+�v�aQpj{���G�9Aq+��$\�mϷ��Dv�l4`n:	�Dط��bZzlUJ.��耙�������%!����=�*������(���8��������q��s��Y+�~����/�}}j-���DDbo�N.��4Q1䴂'��=�i�i���M5$_#�,��ty�ظQ<���[�mx!Q��ao8F�$��@�E���و�k��͹:�vr����Fq�L� ���m�u��WM\�.���j?;�, 7���x�#� >���u�C���B8��Xʜ�>⁭��1(�)�厙D�?��~vh�l��~���g�aS}�m+V6�3差g;V{b���W/�,�d����dW�7��}�@bBtV����I�kQ9��sR�]�Y�9@+Z5��$�j��t�
�)�����Œ�y�fE��ng����h�7���d��Q8�g�a�ӭ�ۦJ���{�{݀�!��acj��yP_�jBq�k��&��J�8�h���&mr�e���}eC�	�e�M���B�s���M��{�W�M4�n�;�m�|������ĉoPya�y��%��	Ԥ&��"�v8�0f����Zh������Jg�6[O��'��L1g��#H�A��!gY�Q"�����\��x������{������~�<�(O�����r�N��
���_�$�RG�#�%�p@��A�(�,�	{d�3v�a�{��ާ)]����<�����5�fI+�/��2�/��/�sqA�M���,G�
��&�aLo'- �.nX �Y�O���Y����"��n��|-]�O��dr�G���)�C삒�������:�	f`�	X�9zIm�7���94���E���۫�]�)9�eM���>#�9�e���Ó��K���c�g-cs���R�jӱ��+�)C#t�w��z�� ��>�Yn�G*{�ܷ��?���[
Sc>i��L�`%�x�,�
v��n7�_�	�f�	V���&; ��L�ʷ�Ml#R�$(����`���Q��W��լe��L�x�m]4˵s��Y��^3��.[k��6�
n���|��g��D/Ͼ��l²h&����(̜rjbE�Arl~�p�7+Na�|��N�Ҝ���� ��R��_�v�`�Q�+`��a���&��t9B����O@��,9�lb�ڗ>{N��yx�i\���%	�*��ۯW\a�6@;{���X��C'i��_�C6��$ϖ�t]>:(��<0.��^�QW�:`�ag��e���}��k�(����c���O6�U4x��[��k�l
*�3�X,���i$k3p� �&�Gf�hV�h%#�F��9����?�.S ���T��(1)wTi4���eB���-K��((�)�����lJ��wo�Y��
�B�g-��Nߟ���W�(�`c�\ZHf�q��d���{=G{����5�����U�D�oyI���� nC;M�{2#A7?�TB�:�uPv�J'���^9#���B���~�Aޓb��x��EpPL=6co)�w�\���8�%+�
2��x�����=:�Ϛv�A���v�> C"��4\�<��(��0�7b���'�x���3箟��fK%�k�+j}V��۔o�p�@��u�U ��-�ar��ßN�}����Yx��½;vB�alՋ�@�/�3$uo�ɫCު�U0S���F�,Z�O�Kb��
�vͪ���Tw��p��jN���8*S}[N��~�8�C�)}�,��1�>�]�����lTsxϙ4Y���L������Р!hf�%�B-����&�hx�&L���,jD��N�����9[����U�9�1�*L�j ��Ǒ�
m������+�W�����B.�%?��+��I�d�|�F~�b�>���5_
, �l9�`�}��x��7��2�:	�e҃�p���w�rZ)�5Q�	�J0)�~��8���(�������i�L�/�?�F��+L�đ�O�l�E `��
L��3���[o��Հ��vB����R��;>�J��O�cc+?c�Ȉqz�O���^A��|U�����<���`��뺋:��&����R�F��FN��'S���[�
ftDrm;˾�I�C�P:n��7ۊ�7r1.W���nl߅Ə���7��%lN\��o�g��K,��b	u�Ce�ϙ	�/�㦗øfm�����9��T>�i�t�� �K�L���[u�$!���_T���\�_.��\QE��.JY�e���T�C�7B6��"���8<�Kس����Pt���8�ף1Ǭ�Ai��q˖�l�S������;Q^@Z?�P���xE�#P��,�L7�N�uh���f��ab�鷟ȿ�k`d�%߽6k.R��䥎1��O�oU
��A�0�#(5J����w6��uH�Q�A��,Z�]e�c3C����0��[�P8x��2�W6�����T�\�~�X_g�[�WUE�l:#��g. n�`h	r���e��~�dp?{+#R�q㎖1W:^�C����� #ބ���c �g�T[�a��9�1�2��|�LK]۪�N�/�d)44Xb�b&xV���X������.Am7���������4�Yh�R��_�MP;�f	L��'�|���h�ql\U��ڎ�>A��2�&�����~��o��k����Jy����C�!Q|c�H�����i���"�ﮮ9��Xs�a1 �4�ɱ56Je �p�9N��?�m��`�c�2�"�A�
�tʃ�Q���4�f����a-Q�̹qO_%g�����F"���������jV�ȣf���n�J�<�:9S+o�*� `�xބm8�66�����.�,7���U������y3V�B9Py8�,��|}u���
���;΢�3�ECh�{��7-��a���#����7>S�j�S�\�n@� j���� �`I�J��%I]-�����R��U��ݠ�>0>�;�_�uow}��JA�)-3�tb�&��/�=���E�T��w�`��p�7��-� !K���d�dM���n�R0����\�����ь�-VT_������&��g%M��1��	hA~��勢�<���V��5i��p��@^�P����Y�[k������� �\��M7�H'�R�s��X�>h{��?p<�O?v��Z�y�����G�ش�M�s9�{փH���<��z��:%�H��
Uc.k󞈯'ҡb��''xg���=�Q��?��5Y�F�)Р1���y����t��Q�ʂ�DSJ���Nϭ����h��|^��q���Tu,
���=ݪ��I5�*�̝C�ev��v�/8m�&e��RݦY<8�w�qx�5n21 ��`Ղ)����^_�jo���~Y��N�������q���㸷��m��J��T��0@5�#�w-��o��C���y�0�]|]J�ς�$$����lԙ�y�������	��Sy��f��E;4&�"���W�Q� �v42k��A~[���@w
缴�����O�Șq��3S�����k؞kM#�d�؆&+p���U�3S�	J�`�/d�7�i8��4jx��R�d��x�@�e�ae;��[��7�����C���mҴ��΢�2Ua˜�St���咞9��0�K��r����Z�B���9�M���W^I�h�-Vh��H��)�O[���3�$�Z��ň�:��JyZ��-^C���5s�]��`6�����Ȑ���8�Ϫ*�nD��ORk�ܵ�xmD�Q�V؊R�
AD��EXG{"�i�4g|��pLL�n���آ˙z�Qg��$o�M¯�4Ć����иN�[�#��gD2���C7�V9K�;����%2�5M$��i�N޳<\Y�zlN|���8]��}�.���)��k*�8�i�����F�uR�EZ;i��݆J�[�I}-O��Cm�(Y��i�<����!	mku�u|Ҙj�����U,����\S$.x y0��⶛�'?oԒ]�rY ��u�,�X�pɍ����)��G�3NqvcpRٲD�a���O�o;;*谪����'�<ڏ�S�o���P��<�F)�f�]Xy--� �"A>���*���ˢϴ��Z�_����˖q�sI7
��������8��T���e��A��e�����N�����e#���I�9�9��/,�[s|�q�;�ӻ�Bw��+H�.N�hd�� gr
��;�L�������QϦ%��G��?�x �l;4g��+�T�7���a�5���Y������HP!ym��ܗ�uN*�f�8�8T4�Ft�䊞���~��}�)
�!�C�5	��v�/=�����k��ނF����%>���2L9�}CmO���N�_�|[�q;�X������T;��r��Y�11J���b���]������\&�?�#��@�(-!2�YFF2s����b�������v��ް�-�N���9C�U��N��|qXf�m�r�
Y��BsN��.K�_@�5�� ��כ�RCc.��E���8볿�r�.߇jӄ���ʐ�d����X��
-�����PK��K�Q >Tr9x��{GR��_wQ�m�s����-��a�t��A�U�xw�����S�~��� %G���:��x���p�qJ��)�
��U8q�,��[.���O��O��ih����J/\,��d�|;^c#$4�Z��,O�" yΜ#hP�Y���L���鴑L��g-��J1#p{PW7<��M?���hL�,���3b�@7���#�"��w'lån<�i� D;�Pɘ�T:t��T.�Uu&������5��`�6�^�٢��;����c�¶��#o��J�F/�G�^����9�ek�H�yt��5� ��9 �ܯ�߯b���b�SΛV�'h�j�+A9"��k��	s��&d�ȐR�&��T�c���Y�Y8T����m��Re�b9=g�)�;SA��S�.N��4�Wٓ��~ˣR�W�
���6��;�������7gþ%���R��o�������yƃ���_`�}��o�QpH�{1�:_�-�q��g�]��\�N�1��2�����=`�w���v�����w<�L࡫�;㸑W=�aD��a1L�N��BH��\_;,}k�4�T����Z������K4/�&1w���׫&�?�~z���s=�][���<���>@.� r�i��i][�S[���-���>���+�������d71�A�OH{Pq(�ea��50a��^����y�l�j�e�:�賜��wg}iD�.&{jj���t�G�Ԃ��v�/"�]Gm�]�t��`�offS�^<��r��G)璥���W�U��7r'7����oD? ��8A�q~��=�*��B����t'��%ko	����~��1W1��oE�;[���ă�6�v�y�g�������M){�x�lfΐYڤ�����t8��G#6])0��S-ք ���~��<�j����~��%�AL��kk���:�)�V�4}�C�W�\��:eb�������1͹�����_g+���A�GT��נM�MtZ����ӷ.��U��V�RY������-7����v|���[��8�}�s�
ba��eQ�zg��<�j�NB�3����8?�|G�DO,bc�j����k��n��٬�q=aG�q�p�}ҁ���Y-��zPS��<}k����h:��Y��`sY�����!I�l�{���A<O���8H{�V�����:M}0p�<ϑN-\F��^�H0(�K�6��l���ݎ�J��T�V��nnt��q�GL`g���E��c\!w�s�D��0�\@�
1��"�0�}Jd�h=����~�Y���G#��Л�Q���DEƿ�9����q=�`��\T�p)сdЧ3�<�����d�f຀��E�Y=�)@/A�O���NE�a��L�%.�SF���8�{��o���[�>82�^!�2��|*O��PL2�W�;@e2�j�Q�����'�������H��z�|�($���rY��M�[�3�w�L��U]�l4+v�.d���/�bpxN?ckˢ����<�W�n[�kM��b��?tLCs* %y�?�a��5�!��U�lFD�4jn�x7v��ci'd���OLz~mSW`P�(���տx�ʄq�8�Bn���D�۬���c#Ǣ5�yJ`V*�O���)[s՚� �6y��νY�C���S/�3�:v/~-�֏
0&
,�s��&N�7��rsg��|�U����Jkݑ����d�ڗ\Q����ΜR� f�ģ��9��Uee?���A�,T���5ڝ#{���D�3;��-z_�����K��2�F0HrzMB�5ӚW�=���=��U��E$�sv����� *tki��/��ݠ��E�Qy�PL�lY�j�Ϟ&��\(m�N��*��;C����J�f�K�!�#�@3{��+3?aW<�	�� �y�>u��I1B:�P�tS�B�I�I9��? 2y ��t.��<A���þX^��G3s�h��t��4��xٶ�F �V�E&|��q�8V�l�
����~���qN*�jkz4�d�⮉y�7x��M*������(oH�c�D�f�s���g��+qD_����']?2M�t��B�V؅���Gl,*TƬ#8 ��Ti;[:k��J��Qy����Ww�㷲��3F�OA�Il}�����T3��������*P?�1��^(�����O$'�zrx���e�j
IS�&�Oo`��6�FbEj���v��k��c"���1����0r���Z]鎫�7	���gc����h3r��|)2�K{�;�\�����E�B-k'��t��ˌ������\����*)�������0�X��B�_�LHM;Q�f����3�o����T��Y|(�*ҕ>u�}6tѩg ԭ�8��FFz�fDm�[8yt�����?�
�2��H���<�ieͻ�j����]�kSm� .�z����u��&��܎f-W??�I#�z�FxU!�ISa�:#���z�P���)Ώ�V!�θ	4C�0��x�6_[$�K�3
����F������@憾���k�)��0���qUx��Y|�͗�G�_%�0%�I��CY��Χe�8�m��;7Oۯ�%�����j薶S?y���S��(�8�7&��:����+��M�Fd-j;�a,�q��#��:a�@�����;����-�0~�$
�ؒ%g��I����;�CBxT���(�"�b$G�rq�-U"�Nf�s Ao����}�	��:�b�(����G�q�ӈd�M,P�]��5iH|Bƛ\^:;G��#�;:nu2�흂�Β ���O�x�7Տ����������<��}��yu{� �*��j�`E��i�a�\����\fj�w$��H>(����iLk��:�#Ӯ�"��?�;v��=��ۊI�z�m~�X���{&Kt���F/O)ǫ�Æ�0#�ÙՓ{���j�ah��mC��2�K��Y2;�$r�^J..<E��γ�� y��l��0o�C+���Py|X��&����Pײ�xLX�ߦ(�#s#q�[�[v�RW*>���N�������q�zb��)b�Ch����O�y6��{1������hR�s
R����y�`�#�Qh^����S>�����U,�~0��<�g⾧��HJL�]�esq��\��,.��P/�,�gV��G�'��Ѡ8�R���z#��(�����3�!�*o�~���˶���m�Do�?W~8qb�=
&ލ���:�-����� ��a��$�Ro.6���:���O5�Sj��)X2��ӧ����"��O�+c@8��)@��"_�L��q�v�i��c�u����[_M�$GmY�Y������9x���N��K�Ŏ��}['v��w���'t"�����4QJoG-�m��L4,���[�������9l0mޅ�d��a����M���{�>^-	�D�;���Ĕb~�"��~�0� �<��j���~ĕq��&Sc,Z�)/Yy�-
��KW�U���l@�j��PsSP�#s`чܶ� �I��h����Ey�����#{B��*́T��K�)X�ވ+��������m��E�;qW��m��T�٪|��f��3H�w �ͼ����?Dm����a�jB6�ySM� �E�>뾬��2�������*�q���f��S�i��,���G͇̒YK��O�'���q�;>
��!��h�]��D���� �KbYQ�fR��V7�m-F�-\�0DG�.�=�Ts����ۂ��φ����-�׶�󼐱�Pg'�5�&�ф�<�:rc������s ����d�� (��M�g=�i��-j��=7����y����1�扉'w?R�"����F \�צ�!�od�b �һ�r2���6D��?����$N�q�o����F�F�k��if^z^g�e�:2��Y��]��8���xD�)�xwB�;�I�%~��n� ����2r���a+�����0)�55�u��u}�'�@�8"�0�V^.b=5|��؄��FJ=��S�յH���m�����\�Z��3� n��uqQ�C�� Q��˧�~�a�U�� �d�y ��|N��jԏP�V��@vB�p����K�Kb!�.�o�-�R����E���\=���!\X�=ޙG�����^qO�� f�sRYU�+d�U W��"=��_v�Rla��_�Q��4�W
�un S0��͙P�[�3�b��I?y���}j�ү��0�$E.Aٷ����^�siJg͉p�����j�y���>W�%�LW�2�l��h����"���| ���u��7=���O. ����X�"A�HSF ���e�ÆW�bM�GnU�:��d��o �K�e��B1���v�u:X9�[�ھb��Co���ogq��/�i�ڛؿ�(4G�P(Ͳ:�r�"NV�NF�Ӄ�)7�Fc�C���79�ߥ��A ���N	�J�)�ߵ��Z�eK��-�<�� ��1�)9
+V�fy@��<t VI�cIZql�4��K��K��-2��Ř�d]46�E����Þ��iS�
 �ʩ�{d�2|8�ζ��WݍD 7�ex�
�����R�5����t&��e,��e��ʖ����㨹=�I� �;��Cn��8gv��Җ�b��Ȗt��`rj�V�Ƥ�������2�~�ȹ(�����]��8$_E�w�����=�ɏ)�Ru��<hf�p!u��Q�r�]����s�h|�k���5��8�����S�Δ'*�N#l�/[F\4�~_�#���x��C���0��k�n�v�jۈU3N��� }b���)v��?�F�CuDu55��vv�&��H[�|_%���eֹ�zŘm�)� n1�a�!�UoU���/��h�G�[��x���{��E�u����\x]$\;}�٢����*Ǆ����=8R��l�FZ���j+L0��13]9�"{�~���%8;����Si|�z8�=��Q�n����F����?�w�rzqF"�����:�~���lЪq��q��L�V�o�WC�KW) �x9
_��j(|���r&9�"���7_�稞S�Ъ8p0����Ȍ'??JyE�S�?r�]�)�N@go֠}q������ʵ�B~�c�Q�e�ǵ�a�c�̺�Yk+�H��xb���L�x����l/
��֋����T�0<�.��ΒKN�ڙ�mk��1�������fL��_G������'�lB4�EY��+����%�FZGP�o���2�յ�Ǖ!��ᑶe�f1�&N�dIi�뭔�r���Ty��8S*B�����3�ed8�`�p̢@�?���S'��L�(g���Z�����A�	[x��&oHl��O���9�������0{�8��ƿej׸�npm����\�i�
��Uc��Y��
���7H�F��ٚUe�C�G�g�:dl�*I�Y-+GBȇ� x�ϧ6g93|0�p��ƕ�xT���~���� rW�=΍�,��KR��#z�8���h{![��YAƭZd��-�D�W�/=f��0s�m�� Q`�0r�T�z|ݦ��	{j�Y��r,��%d�`nf\g*d`��ڪ�I�,<�'���f�DY�����֓����R N��J6}�q�Q���i
�ߧ[�%9�xg�U�l��H`�U J��ݺG�H@�Wf����/�n��uel FuHd�c|�=	\I%Z�ڃJ��׊��7ϯ	�fiͭ��yn�h��@U��w�dZ#"���I��y�?�%��h�����9�/qK����B1���1h�����Em����T&���a�s�j>��;Fn��R���"O��nY}?X�7���V���
�w�6J��m�����|=���x�x�(��:E>:��U�l�E,��GDM���Fx�5'Y|������=��LT���8f�L0ֹ��⭜���Cks�t�>(6��,�ǥMypt���0	�ߕ�Y��j횂f�؆R�~���'�:�>$b��	�\y}��D=��A4�[A�������P8���4��8cQ�杖�:%/��/Oy�ލs�S.��)Eb`�(�RR�Iַ�<�x+&��n3?��&^������9�]tΠR� �hr����Қ�e؎~����:M��}�J��w3����h��џ09��I��X\�`���K ����/�r�����B�t�����^���<���� �i�V ���|&p�2����*�1���tp;i䔁uM���ȸ�0�ٚq]�����X� �,��rR��s�d���>3�<�#�����p~tJ[��dWAbI>�I=�??�]�%����{�L̝�Y���b>�e��%��D�i^/d>��Û�e�c�u��슍��p�T����ԩ&��T���E���+�+�J42g�E�U�ҭw����u�&Bb���nBȘG�X�tui�T�]��QE��"eԪ�K{�Y��쩁���cOuG�@��>��_1��lm O�Я���Yz/lO��07S����!�W>@�h��Uh�i��v9کS�Q�B���HR� �g��<�Z���p'��^�21R�	��AB��r�u��qBf�ɩ1ZC�V_W\ں����a�h��z(���f'~:�"���~�r6]��J}�4a�F{�Z�x�&�nЙ�B��z�y)`A~~��&�N�m�k�vs�=4��@��S��?U�o �ײ�Wh�Tu{��Q�v�pA�����Lv�x`X>[�(~SE��X��[-�(�̜�ktd]��/��Ҩ��Pr�)���(I�L�������4p6g�qq�ۚ{VQwmՕ�_)��VĈs�pcn�׷L�힑9�/؀��ښ�'$�d�~����\���=��=L�SU��?� ����"48�������c�B�X�&wԜ���C`օ��]K�m^o�*��];�	�
�����!w�W"�����j�F�沋�i�>X���*�8a<����v�4I�Kd?�_���9�#��E�����fb�U���ɲ����"z�Q��N���*	�)���τ]��LH��_�L��D�.x�䪦�.!<�$���9ƒف��v�����p�pe%pg�v#��Y	�%,(,�7$��ʋ�̪�s1�	�El��`��?u�w�bc���L�s!l;:	qW�ڣ����N5?FW�]#��y����X�6������&�%��tnA냔{��4h�X��&��N���d����_����N���$��{�#�G��\���"���xHF>��`�|�n�o�,�{%c\,^�ޤ��$h�-  0�Ź��..w�7כ��?��բU�K�Y��In[ϖLJq0������J�1�L��A�/��F�s�ԛ�^w�{St� �wN�Qg�����ҥ$;.
2kxN�т�~�'�K?�����D�0�����ZB%�:����C�N�	"�eW�s������Z{�6�>���y��a���/��ƈE�=5;2:	���z5%���L��1��٧\���k��I�Ҕr���
s���b�8�:^��!T��6_�#[�C.���C����\��kտ�!�b^�3>��Ǿ�tt��elݑ!#y,� h&����=sh̳n|M���+(d�!�ǻ*%!�]�h֨ڌ�	dB�{U��_�pD��~-����u�ZX��k�%�n���>Ē�i��OWZ۩�/ϤWզy\!�!2�ͨ}�<9�m�5*����a��"�n���Hý!�7Uб�k4�k��\�}�>&�L���:�*��ȅ���Tm�4%��H��]�|�	b��Z �,O�Za{^ԯ�x?��fO�5a�^:�f�"�L�ص�C�����v��Ѡk8�5�pU	?@.v�+W~��s���56�?Y�+������"���̰��KٷI���%����\ tXk�����G������B5̻P����>,}��/�i(����&��w&7��y�»�%|�;�!;z��0s�PŸ��$�]h�9R�%�]9U0�n�3��+�HM�%�Rv&3Ǖ.�ZtQHqCv�9J�Qkf$�i)���W�|.�X�[�"6����ժ�z��8,��x��Ȯ�EZ�����+��@v�V��G��Z?�d_|��[fUyFcbS���1�3\�`o|�`�9�QD/�qU�~�ݨY��)�#w鋾v��#���1MF�X�*?��8�h+�{�#�Muy�Y!��(�-�m���l\�B��Pay�N��k%pk���.��g�/�����n;�/I揖 �h�ȋ������N&��v���>��Z-sǶlh�.�NӨ�p��|4)��y�'_Y��|څ���ȍj܄����P��[T!$$2zB{���}e�����
�6�-�����۽�0��)0!�~E���_ҧ&#���
����ֈ%̰,(����H�ο�"m#���:Exva��bx����W�=Wj-i��k�.@.ɧƎ+qcn��zd��m �q0�]7�˜x�Y�����
���x��Ȋ2�;��&����3��v5�c-��BB����>��h9DBa�k��)�#�r��N��N"�ȓ���EE�l��U}��5Ae�}K�:�V|�ۥ�8��f,f��|����m୬��dSJ�>1���6�5ӹ+�:�pqF��I�0"퀢a�'1��Za<��]��S�KI�8(��>͎�I�ٱ�3H��o���X��1�l���S��ȴ�`��2�Nnc>D��z�sٺ�j&8k���aэ�~Xx��M�5�~�o���z�J�δm1�uy9�K��u�Ñ�$���XKҺ�w���^���~:|����@��B�E
��G�"�gQT+�6��<Vx/�������%�=M�4	(]���)�L�g]}�Uu��U��K���([H&C�Ā�������^[\��>'��La�9-5���p�l�D��N!Z���i@���@�eGs���j{�Fg�4FY��W`�0�n����w�Kk���=P�p�����f�6����?a�/Z�W+����0K�YҨRv�c�����iթClPs�j�^���}9cP������̃l�D�ECυ~��zw	ǟ�=�8�Q��,a��]�[7 �����'���o����5l�z߷�3co�<k�7P��95�_��J�a=J!�3���C4�@ܑ{mL���:ȏ쉆>�c ��҈����oZc@N\�{�R��C���X���^LN����s3�hlc�,U�|*%��������+ �k����'h�r��}��Wb�aͿ���aX�oƸ�hj�߮�]�LZU�� ��~a`[x���<� P����$��<�@M�]�3)^��# }���A\-TA�@ע��67�U�Hu�\�nw�4�mh�s��щD�?���i��|M�_D>f"ga�<p��2��G}�xf����
w�݌Ej��yN�L�b%Y�31�+W�<�%k�А�z3<��W�K����T����\V�oۿ�3��u>�T��j�w�8�q����%U
T@�/�%zr���U��/8x;2��F-{����e�\4���pj[��
b�!i�7"k�[���6��3 ��gf8�!<�m8ӄZ��3oJ��7<���Wt��kOX?P�D���f�a>+3ڸ�m�����d���D��'2�3�k�{��^��e�R+���C�DH"�#R��}�������F"t"�/���?�o�����D OP�u�)�K.yw��C.�z \�YN�e�?൝�fB�ZӒ����Xz�9�꣄�����\�V�c��St�X%�뛓|��k���LI��O�Ra���K�VY����{���Eÿ@ ᘤ��� �h�7O%�Ȯ��X?>�>��w�(G�M�>W��w!uJ��c#ɏ}�߶抴u���13lq��a�	�z|�e��4�:xI���o.Z +i��?�H��݊��V��8�
��?���妈���G.�Bێ�B
��ō^ٽtf�>8-�	��;|t�K�s����E�Dܣ�����7�cm&�<S�-%��U�KX��y��ʁ�^h��N,�3O�q7]�����	V�&��r;�L�%���i�ɋD�R�8������������'��H��R
�H/!��3/�B�?�����S���#������^! E�������@}��EG��5(�kR2ٓr�L�$�2!��;�E��V��ݑ�NM���b.pI��u�(�*a�U�S��D����V��I���U)�C���|Lb>���`SA��j����j#q��<	kVZ2.�+}���je���Z�
� �Mn��*�8y��좋~q`���>�T�<D��H�hKy-0�,���o��M�,�8�E�0z�TЁ���ca�3b�L�IG顆��H�l� X���T���[�����d��jM�/<�bw��ƕ}B J���hI,^Jc��o�&egִ�e�Fi##�s��и�Ƞ��?J������7O퀬���=n��_q��ˮ�Y�Q���ѩI�RHɠ��c4�p����6�{	8~4US��r|�Ƈ>p�h�=�����{��4�/`øM��]�=]��Z��HW,�A\��YQf�$�I�B���,`c�g�5���Vr<O>A��w�Nk�4���>H��θ��7
��z�Ș����A�% ��i�u�����?t6°�y�"��eb� ��NY�����"u
4�4�eʳ�ig���
Dp�Mg�1�˦�	�AA;w���2AL ��*�go�N��
��ءQ�P�cG�ך�Q ��;�b�Vճ�'�؇���+p�o)�;ƼKH�v��@�A������6Պ�z:�۝�0W�(�s*[��6��㛽�)�u��}\����$ �����dZM''g��ct�l$��θ��ϡ�	�oN0@��-V�Q�����g��-�pb~���x1��-bK�Ž��J�	\��T��2��!�����86;ј�A�I�L������|ZJ �q�R���1��i.����Pa�j�����r9�5w��4��vym�Y�����XT�A4�����8d���Z��a��b�S(��ķ�	� ��ы-q��&j_����ER��^m� V�:p1:��l'�W�Tf̖3�<��1��@���������L\!���S''��녙8s��<�^�-��R%���W��Q����D]=��1��+�3(��d�;� 2m����ưW�<1��3��v���w��)r�%%^P�
�WG����;A��@����AjPn^BI��A����n����%rb��mHָ�l`�7G;��/��0��%��\�B��Ҋ�Q��=�m֍iD�f�W��X��gk��?7�a���͕I�BW�����|/�r�;ƙ*D���fԬ�ᐲ�&�䉉�{a���Sz��w ta�XB��K�n)���t�Ҕ�E򺠯O���zF%&��֠y������E��b�7G��%��`D����3�%%s���@C$$(�IF�7$�+�"3.�6��}�#��
�X7���J_k�o�e�3�;� ��@ש�S�������C�sǼ���+<�칯�;�����y�ȴ���$�q8����.�o��\Оύ�iV��{,tp, ~Gԍe��U�����z������3]���������M���ǤH������9���ޤ�E�l^)��������YM�N�k� 5�+o���%����>�EM�K����(_�Ƿ�]��K/���4a\�3�_y�������FOGy�։�9P&/~0��zds�P�s� X���U��;�>� �[�Q+xJ�u�O\��ž۝.9l|Z)�O�|j�8Ht ��+�\jL't�2/�f*#����>��������C t�߹F�,�s�_.�c�"Q�!�C���17U=lg���G��ض� �6ܵv���Pr�d��,����" � a�X4>7X����m�x���o��� ����<mNel\Jbk �;i�����O�BCU�J����t�Ϥ���
;�p�J������ �,L���V�:������K�yXk��1?�;�eeCf<�����ٛ٠�=p�,Uv���ئ�&*�M�Z���f]���y�ĵ����=֟�/$�$�L�b���f�ֻ�˕'-ɕk�'�(3�"�Ͽ�}sW���Ъ�d��w����n�^G����_�װ`�_�*�α�	bHb��T1Z��a���Թ������!���1�&��p�5�m���5��Ҏ�[�\�IR���z��r���Nb�������D�gdaU�i�MEǼ����/�6X�����K`M^L+��zc�8E*�~��_�8!��Yx���>��5�?EM�����_\�?�����Eޖ0��c~�vd8��ď�Z^R�m��u�t���ǻ�O������$���`��O*^�)tjK�q
�x�8�m�K	&�8�Zu�͸
d���U`B�@�\��!Hv�\B���6����ơ��G�*�ݰ�}e!�!�@h׭�1��
�U�Gᘭ(LW����5���� h�73_W"��Z*����/ތYG�������!U
�-�[�,�������!3E�hiu(t����(~�=�C3���̍��5�6�W%ؿs�;�.9+o�$���i����!*=`?�-�a�Jf�r�G�ncGu���c^��Qr��E��#B�ז��`;�/�nwe;��cM��:���^�5WdE"i�.��`BQ,�QYX�%�.��O��z
�Ӭd	e�j=wN����5i�5��?4o8F�k�A���+�'�]X���q2=��Q��a��U���a��>+��_��F�o�K��LL]��gp{��@�𚊆�Y=^nۢ��p9��!a��DN2W���d�ݴ���76�����Z�����e11��ݬ�ecܣ�������V��}�S`��=��`�p¯a�V�)��w�p2��WxO���K`���onԵ_O�JVrX�6x)�#��*XWQ�s�B���˒�J5�X=����R}��Z�嚻�mw#� �\�D��A���5��'�Ѽp@��\r��T>�@ݥNb�~L����{Vjn�±Ov��&r��f��D�YR����݈�S�o����i�:,�����Y��N'կ��Q��]������?Qz�2�	�)�&F�N[eQt�$̪�?aۖ�nR�m@}��y�HY��\�����(� �L�'b���b ��^{��ˮ[�>��;Q�$��E6cՌ����|�7$CZ�V�	�blY2�M�֜��y�x�*ؓR�@J�!��6�g-� �<p�z�������Ϝ��Mkx�� @4v�{�l/~
I�}���'�9Lik����ϓ0��Q�	��L[��SU|%7
��pH��фO�R��eғ� ���>��/�I���qD��=�D&㜅��[��u���pM�¹�O�j\̢;M�`���<�f���|a0��ReJ���8?'.zXn��.�F����) i�r	�Fq�����4��(�i�vQ�[o�r>&S�|X�6�/������&,���8�)�\l��n)��\mt|H����07X�ۂ��b��ˀ��4���b�H�Oo� Jdl>.d�]���Q������aKE�	��
O�ۿ&�y�Ӓ�I"V]�O����F���s��&G�K�2bL��o����<?��i�9��F���?���E`d����G��*����9��:HG�~Z�(�K	�Oۧ#io� ��m9��rq�����*�ʸ�ԫ��apsqsk���>"�D�ve���T���y+?G&
��ϥ0�:Ԁy�s�g�f��3����Ǝ�b�f��-z����;G��ܟL���߽�~A�93z��Hs �4n@-W���I3#�K)�ۑ�V�z$I��S����^҂X�y��4}SWFDK��D�̱���g,����BΟ�D�I�A*�J�,��q��AJҙ�X�_���B�M��	��U�']�M8娛��!�ٲN�h�]�r捔M�Zl�Z���^���X����z�ϴꝡ=QQό�j�Z��~��A����\�� �k��ӁG���f�{���\��A��n����++ix鯬�;��6Y�$�{��r���zxTX���W����\�+�l�X����b�;�C�WkF�N�sh�,�D��`��"4o�T�n�OQ+�i��B� �"[�E�	2�	�_�Y[��7�Y�����"J5���0��!˘Xz���^X�2ދ�܍�I���ۋ��m_��m�l�Ll�gIu��ާ��ܕ����ntĻT�DQ"�D����L��&s���s)�1��13���܇��|8aǹc)��5���&�8k��&8X�8�k`��^��YB�Pn�����$��jnm��P �H���A�鷵���������?�4��̎���؏����E1�:M�2��{�ΑA�5�k����}���8p@#S���i�Q5ᒝ)�#P�Gd�M��{���D���o[�r	��IU]��7����� �XD�l�2�'�G���v�jj���n@ؠ�2#�OrxSm��M�| 0Ǹ;1�f�����0p��U�Fv"CzG?��aN�Gp��6P�e3�)��*z�u�{t2�n��f����?�P�X�?�Ӆ��\�I�p[���7v�g�#�����s	r�������H0�A�dRf�[�dڰiCG61��0	�M���burVtIm�0kCGt(߱&�k�5��K@9!�/�6=���/zZ�*����+4��2|�bL�U����	u��Ɵ�l���,�z�t8Pc�C?'CIEM�ǖr@wleA,��(���?�!�%{m� a����'=��q0�.�D�鬰����TS4�.����
��[�Z���1�s�`:)������Oډq�U��� �iM�j��SC}����'S�JSrʴ�H}�$��&#�m���PW�#-Xˉ�\a�ii�3�/d�j�k\�]r�	+�����~�xk���~0r����o$���Ĭ8�|��U<y�ωɔ��kNfR����}V_�X���tW��y)S�s��[�0�i�a�[y�J⧛��_(>�1Xj�YP�,��b���*��X�O �5J�>�ʻ�f�mxZ����!>."w��2,��u;~%s����\ H�7�/�a_�)�����u6������0>��!�Nv�}l��W��f���:,��2���k��� �>�#~l�ݩ@ʐ|�Zs��Tj�/�?���*��!�)�r��2�������4dc�I~��V�B�f�J����AsĆhJ q�l$�0���-��A�m-�������z�7u�������\ނ��k�����T�B�W�6]�<d0�7�gd����'�"�s��A�Hy)c�!I��Rć����cwDPu�ۓ-a<����Z�?�n�{�����M��Ȗ�Hs�H4L��0rM@C*=�Vqfj�&7��ξ`�$�	���=`S0���ܗD��*`SHlӍ�?F/�Z��F%XnhrZUc�nڭ� g�)�bk�z%�B�`00�L\R�W�է)�Q(";4~k��j��J��V��n{���Fb��cgAW�#�&�����%�7�c���J��s�Eg�����H���������5�E-���+�_��9L>�a�}`*��m�T�`*IG	�#���i���چ'1z��U+���>��cF?�����BR�x�>����D４w&"��h��.�,��ߧ�l���gwz�Ll�L�ɣv!���Hkmu�.�/��'!{N��&�K�(��^�:�r�2�W���@Պ�d�G��?M�t��)�W��0��ekc��:�Z�#b�e����[4��ꮚـ@�`��� �+ꐁù�f��ۭ`���1b}����n��h~F�e`3���U�9oB�䤜�j�>�g���'�`I*��t�>���VS�'`�wR4xr�*�