// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
/wGAjMTxMU7yhhE/Wtwwc7TL2It00X2RRvSgDhFJnvKvVMYg2C1k8i+NbRO9EDbe
2EUcqgMyWZXqzNgkWvBCCmhE2YUUXfI3xdl3ga15tef0zrhXF8JhAmNuPeCO5tGW
ldUJ086XB8iy3R4w4XoBtgAF8DZDaArW8jmy/U3lrqUCgJDlxv4Ysg==
//pragma protect end_key_block
//pragma protect digest_block
KR/Tkk8rWYfiXrTQnBlhkij8Alw=
//pragma protect end_digest_block
//pragma protect data_block
UADNUwd3hpTQ64sDRVPdb2/ZTJGTRDgIBnll0I68VuCRYuB7sYatrLNw0Ucz9F61
/wpS2MfrlOUXrAMEcOk37tFMNRwr1AXeTnD2dyV99j+bLdy346sru564MWL2mn1O
XODjYg/kiuwCv1DwgTsi96BSvZ/mUnmxGCZPCMHc8sZkIqwHIiaUYdyQ4BRvVpHk
1fBR6cjsjRb/uIbydCUPijbbF+lhZWLe1Vje7qmx9In12bHclDR3H2wmuu6DWFm4
uBcaqq0STECqFCaMaa91F+b5oQ4sEMD7z6k8iaiFOosVhKAugbOGS7XvZ23Isqrs
0r5BqoQpeZBl1nLNtD6+P9MNHD1puO9MrNNik5r2S9PrG59RsLNJaau7eEGTGRV8
y23HTnF/jiJ2/8J76S4OL31KwVPCzSc6VEAjJQO9WhRPzOAV9fEs6IFgM+0wKxB8
ybaQ8RR9y2zJ38Ts4w1Pi9X38ZSmXiozrjQHRVUn7Gc0GYaFgW82x91LxTaq6G82
ufDq2IfGUaGFIxcVJyBY19WiDopbWYUkfF2rmGNH2WizQYnvsywZsb/kJEfV8cHf
JH9+HlTwdv2XsekeCjMub9MSY5URMwRM14W7wWEmZ0pv7QJC66eRmBXkUY7csexz
WRESflujHVf2uqxiCRjlLGV+sMegq85ME4vW9gypcCLMoafx+dEgK+48iO8FDX7X
uhSFa1Ocuo+C5BTrBTn9NX8gqxEq/sJYABnd7vS3o4PtH7M1lQci7/qm+DAE/vol
wq2ix+BIo3Sb7hPDk0yN9gvbm3oHFDUGLJdQw1dQFv2JCRsNXe4AyR+kc0KK36A7
rOWEyJmEKu5gTR5bzlTE4cFSbxTi/c8jM4knLPez6f69TiVdwjVk+lVJ+Jf8vTh0
UmRs4yxYtAXtL+jvpCxeb+2pjvTOsj3QvLNKK8JzZrmUs00ZE/4mc5zzKRnzn/5p
lpdmJMGZnI9CCS+U3sUxz3KqPuUV+49Z4k4JiKepv8E3Gu9KlWZAKlYQqRtf9wtN
tlvkIh3W9wViRZR/57dqk0Y8Q+9R0bZARWpaNSWgNMKQyiL6roY720/nVJakwuZv
x1KtZ3dyPsbIjoL/4zzPdVAZA8qeNiu8zcQaHgR7z6L+2WSHoDxzN7TjNefYj3ue
5J/HaElywlqANhOegWEn8R9iIUa40s47GICLPpPSapHmGEQx4T9DKZeqNuq/G3OM
PmCsocOHrUqB4R7v4urkIDvgU5c1395DdnGRO23eiQsUUhKv16yqBOjqSvSE9YRC
l9qe17P295VC3pcCUN/K2oFq/gzYpLg4tCA7O85rk93Xns+3j6dIsmgQ9kudChfd
aYUq7hqsb9gIt36h1L15o1CHEejWcPhsCEMNd3AqoQUAJsoQgBAPvd6SnwmmeexQ
A8JgJ5JpvdkqyGpaqLQRj5wQ2qkRuf3rdfPjaMUUtn+RP/Tv11TyQR2pxm8sREpV
wPiZ6cc1MwZSdy6zYHUK416NF2kExhJr+LRQXf6xL++GsSAuZH5j+2vrYMKrRPS4
FP46k4DKnlZd8MlW95s/sHQQdHvz3WIDll3RM2ABgauJ8y/91Ufv4CFWK8zdHNGZ
rtPveesQ+xwd1dgtEKk95wkuBZ4JjH4073PwkZZ+YWuQiobsTEkRBEfVXJl/f/nW
0BFGMMQBYinQbPQT6AHqQvDLXldNda+7ZFkjjHbDHVu0y5g/jenXGo4mL5ybNB1Z
1fP6qPU+zePxJSi/gd32aIrKubd0Bf8fR8z71dNXLWL3MNccdipLbqzcVPa9iqY+
kHCnB5ZultPZTKxViM4FGq3YlpXir67LPACqVG94muPdrSrKNRlNjTHL+gGS9qwY
nmtQiWLFkBLf/ZKbdLu1UYCqMY4oINjrfx0P5XwAm2ele/OmSAFz53CA2myMbI9X
Ns1+TAV4QrDr2C9r2mvpqtx/s/Xy8cP7HhOX/vABQrZnn51D8LQATzv6fHCBANQw
rcbu6qLqHTboN17fEZaqgDD0WS+adV1PuSHM6EovN0i9GcBX7IPxrxP/OxWn4JrH
jEl8j0dHOHgCnKrH5umUmfMRspbDA6s8FTZ4HrsmK/BZNCQBPthY9z4Gr6DJml2x
rM0+d/5BhgenzTEtsPiMuCM3uMhN3TrY75LOj59mItzZbwKXT22djr64mEmQsLDP
A/9rqt2Z231bRgc3xH+s0KmsejFQRv5W23r4KHVnyoVlVmsO0BYA0YFWB1yi+AWL
cRWpmXhJFkfjWhu7O8av6uoVTrvNysQUahp5VpJV9STpnikWxHvGwgZO5BKgJ2iZ
m0SwUdcl31cac9cxkN6gBRgUjU8bG4vLk8vvUbHprxrX/TFF3puracweLPxEu3mX
g5UnWHJgyo/r7uMIs4uPbrsqirdkOCqJCcDFypHMEqvhRtIreioi0OPp3BIJWR/7
bKEXL5kCqsBuqAGR+FV1m8GTiqeR5AJQ8iF4fBqN7BAWExiGlCF5ZJlVtLKEKRyi
wNAAPmP4snkL11LSvvdaydJx+19cmhlzZNrYfzOez1t7yWP5PosHt0TlThjDJ99b
nVAwWygg5ZnPH+fkh3J6RlUazqvY2Ymu09SIGke2l7di+2gnKDsQv/hbanF7U6n/
PXELtFrtzoUVVH2YSaWytZdn0e/+8cM95swA/H+bfNkBtCKORYFL0L6yVmSuI/p4
P8q1Y8Yoy8sr6j6l8vI2pH4Mud2D+odNpfTi4rVBUUXDHgh1SfaRAx9lSLODdOMd
/VfKmK4w/90NoB5stg3fg19FAWIOJVyQ8u1gcWgtgdnSPI0h3A8j+cUqrExEHcXk
EUL9cj6niTnBed9M6llYilVfJettXYQ7sY1bjpruUYr+skI34FDAXmKTcuY7QSqL
ebadGbOfmp633ndwNflUmOJExIClurKfeYN4uBprFCPYxhbwxvOmQECW7N28zO8f
RsLQNhfvsqsHDuuDWWDwkwBEs4in/mDtB7Uz7e7QD0U5LysxWcFPTtBBAsEcsqdX
VVGEBf8YGJBTxoQpO8hs67MzmXWdCJWBS2dTUGDzjPmn8heLBq5+vMJT/q+pUzKZ
zNHlWaYQQpWKPnxb8mT33X4mEvtoRvSuL4qWhChNXzP8DFaiyKMQOOVuOfmcBelZ
Fq90j6//rL62KUs1U4LU9XjSfhx2cuAHWCtXW0h3CVqy0lBpDgqZJ/pkqKd/5dL/
m6Dkog60FfRVMEq5fa663NZURaySfCBDi7ggQXNNXlS3tuIx2zcu+QMwrhS3dw8F
xLO+mA9GiwYB3qrWqbtLYxHB0p+obgr6qShfJD8kJzwdg0+3WSOqrFiRl7aktIZw
TKa3kT9DtAUhWtuUv7NFlscUmSDg0Mu3rBPQ5vow7tUFcJ1goFvzDgN1RFVtrtNQ
VDYp04powGoh/qrDsnmgHHl8enL87tizFx5eA96llI/yDK4xATaKEl8BjeCq0SPw
vZgFrWm3oHNHBAezqNGU+8+SYjZvmvMDTI/LAnLobQhzjoJIGj4EH4lyANsQKhwq
ktbSd2vKcFqFVgTG+CGTc585vWWAfhVrxG8ysoLj0ruwBtZP2unWd9css5yqjZOG
GOk/jcUBLqZSHranetk7uCjccdeGZXG9la6uqQ6PHvYr5m41b8DUDpYxvUsOWd5M
lsIntGonuTBsf+//T2PiRRTLNuWxN494bUo194ok2T4iUTjdW8TU/ASaHx7jCgtq
RZq5RcF4nktrcyc2XK8K/YRfOEZOd0bYcE5bGYRtjlLGxTnMc4JwG/A2/BR+qUEn
dVc54EqDTQlUaOZ2U4c0ryaUSzjjzzF3fZcDMq8xjfsJjXleBugaWDQHIqzVdNth
bpeXSjHI9C/sQrVtV6XFLWWgM69m374dbMCjtRGyv70uFeo++oNpFqfhwrIPiWz+
VY9auFXcVOW3M7RtOs0KP50zj/2Ff2eeCrC0I1HHZziZatGmqoKif7OJcyAJJlrR
9iQm1tnwN4QIUDKWm6RfnZdGO56ea56uPMpHf3qBcAFW1neBp5wAgmKTLVrkQZeL
pvVhZmRcgckSU+Vxw4TZ5t1MJ8HacVo5LRjL0liivy41+4zPrf702XtcqpTN/tF2
3hGCj7dsb7NBYQlNeQwChGJ/k6RNfIIC27gA0zn83dGwXMaAQju6liY8v9X56+ZN
CxEJYinekTGCpC4AWV7/QcjgCWlnqajnLqDRNNW4H2A9JY8yMsau0eqAN7rqbVQM
nz5Cvo3I9pNnrggyGaB3HCkeze1ldDDDHuzJ4fMSrUQPC8jGbTOJ0ic3u0YEahYK
gyMlW/OrqppuXYmuz33w6Lb4S/kIawYvTMK7vlDe4S34/0NUBMgptx97kp0e+VSs
L6qb2NlvbizhB0SYWo7JFAkFGFTjYde/7IjtE9Zgq/ZCQcksckIxxR86TLDrCKZl
leQNBkMayyXp6TJpDc+7lt+Jq/VNviBUySSJjd+8gGdE+4WPJFWPbAjKH5QQG6Pu
0WYI7vk9ls+OFrJLllJgVt0iG5oqbayhJh9hynjGtWKBuxqCLVGDbeM2YUEX5CPy
/sZaXk35E93/8LycGicEc8ev4qQFLXWBlM+lrbbuuaEmIDIzgr+DFPit17erM0iB
f1yfYmHIXTFIqmLidaQKN8Is2abkEdGkNNulaMr9lwvfbVUbREn5rENzXab9hfkr
62UrL76Sw53KzjXyc7cP2fqxF0tjKe3ifEL9FTY2i4lH6kswWetuCtDAqXfAaA3q
zd9vF67VZX8oEt21h3wAXRr2n3+Nyj65wT4vhWNflj5OWTLzD+voPxLq7c1P+YAY
h0M5BfFr2kqPfJ4vY9AmzTPPf3DYwx7dyUhn+qttHgW013GRtwNKiwKRdJEzN4E9
Ge9SI7keze3rgbQfADNDEupURJnKmperL2kkL5xLzHFivM9MtxwL6tqass6lsSb/
kW18RS8fndu67v2qzlrJZcyDGkGxlgGTewetEZgCpSYm6mpNAhXcs9BgMj35s4gh
G804w/7w/NBls5nLB1W6I08xVFaCx9jBKNYuZA3AHmrNGLlIBh+POBglAeJ4iCCK
7Ksz9jyNKVC33vdlyZetoD//xp4+IiSEneNLA1g/aAnZBr6OT7vonu7vpC7jvy1P
SpMkQC3+uJdUg8+RmbTaBZqtxC3eUmhi4oPFWtEJgCj6eB1oJk1Tk+TDHaLd4wM1
Tre8tj0a7vTkOlTXR69GSZdbC+3yBfcqD0TNYhD9z/NlL3Bp46I7mxMHdONGGSd0
1uOySOjCtccBPHbbESAzCeBiJh08pM0QX+Bwph9C+ggllbm1YJMiPp6JeNyFIWJo
k/42t0ycly/BPywR9eRkPhSHNjN+ia7JCw6i395i1XJx81N77fqhQFfGzlrViz/4
R+v0UHJTOgnQKUk7KC9tKiGVqhd8AG1Mjr1bku+yV3t5txQvxaL/beLpTJwdTpCg
05hxfL3PKkJdPfcSElVKEoBSe1gMqeqetEPtjAne0grw+zvEK32WIIqo3mxmeYNR
oNHp1odiM4ajzb9Xo1uxfp36D8tVQ80wwg2+a4WjTtEEOv6dnIoPas0ekE+LcfOm
lXkPAJie/ETpOfA5mFoAZpTu/xcoyAPCe++m0KRoLAnw6vNSIah/zIToVeJQhmB4
OmnsUBNZg6VMGkMktRfVOTqYM4U2N9JAuFOIyQ6HmWIicYOwyqg2R6LN0uqE0V8N
ozMQXx4jwSxR+eyxUkhdRDGFcgnylC/RAKbm8Zq1ZyjMaX93RzjZpE0F3L9R+umO
yIRRXad6AtS7mnxhV1+ApcGp3ZdT1Dc7Z6s6wBl/rt4uF+yNKiqucpDoJ4W6kVke
fMuJHqJlzyWXCzR8l4jbDvzDQ/fK0iiDeGlarVun5l5Rlrdc5TvTZ/espVcS8eKc
vOBxSECkdjQmkm8cijZ2qOexCHc6CIbrLnf6LRKqG0srMiidyt49zI6juEvH6y8s
EEN0K7NV4veI5ZwINYGfKKTouK3+lEqDTGRqO7D1bsBDdfGw1JdUA8sKyD28J7BP
D2MoUScdTPHZGvsVq2rChNuZ6ZVheYJKL14364IU4pm3dQt7ucM/SSRR6n+F5ay5
22uHSVtr9OA9jH67/BOkj4WuNkV/Px3uusNVHBZOp3a2eysfoRU2ZIvLTRdlGUAo
XM5atxRmyEGcA3GLdduSd3mM91T/hJR+YfRhZDr0aIKINxrrcxSs7N5NoK1xRkQ3
qJVLCO9hNCqWGHd9ilLIYIQD/m6i6pwU31aNMDMCn2botAdoEcQOh7GH/Ik9zOvY
5OWYrUQAVxq0DBqTHXneBGIETeQMPR185/3VV9347i4LL9A5uZTME3ai+kXJMjKm
oEtPvZmqUlwh2TAwpuMH66HrVtrGXb/KABGZl6Yov2ndFepeSCDufzVER6dkT7WB
43NA92tFRkH97J/2V8NyLYCtm1OmtLB549YWyh5SlUiHCV87cEpvbxN1CiNraXEg
mlWZ2hf8jkFpjeGHOpssAx4Mcc3ZHWZKA1VfAsWVZgS95J63RBUhlLJw3ZEFRcJ5
kx6zxEOJloN8ABMB2F8uk5xvEWdrY6U7NLK71nuLIqYww1sxWEYU4RMjDDhZw58K
26QLzgHjcqo1AXPqXf3jYxRk4RwnWT4IU2ED661vQEqOQgbM63Mh6pE1BJrfl/L3
uAAFiSptxsslbEZUbqEKFdzulgT+HlMtE9PCP+vhEsMj9QXNG04Lu7NxiKHJnLrG
8KoaVyV8wMGZ8B+b6fjm8s3w7T0JQp5wcrPad9n3iLU9w0AfDDbZhUUGKgfqR9S0
gRtAaNvVSUT19Q+APYvWriuW1vcDGX4OBqlevLkeLpfeT2d/vGe5otcjhAbYov4+
rmOeheC4qbab9VjEhfoYe7mcWUKSJtzeRndi3mpxV2BGeLDig2soNIczY3VopHDF
YHIp0j8mlTA11louBI1uT2ZWmYLsI9AvmRapy61wnODuw5jR3qTRQKHt7BqJZpb0
6CyZSSfcTLQ+KdTXyNeslZ95Y12OGBm7hpWLnq4KvzpZXObH8HrDobLC0zoqjh+H
AgLJDgeooKlJBbR1GYau0L0eXOSGhRaS3pmHIutn1d4bMCHpqoQ79n/xpZTGxHzp
lN9LhadyAgAicTPOw3niFab9z7G3Bvr8bTTMeMc8GeFl+npmtNqlXoqhvBzhNLLz
Nxvaypuu7mrqO0wGCUWsYPrJV2jTLvUQ4gk9eSJQq8p7Amwny1Fs+4Vi0fBACxNk
TvqibPajdf4MeW/0/Yl4e/R9/kch2aNftvH3D94DtICy86BSJguy7qf0lYj1TIUO
CchT7yI+7YJjJ2uUK4jeqoO60Wg9nguWky4FctD29E85ISzdZo+/Bxn7A5x70fu4
gvNx6IKtcWVZP5TYYp2PCn32oQK7BV9XLLVU6ZCBk/qUuCTsvAUyBBozoNm51A0Q
rTaIcd6/zDb9OPVduDl0IHjUE5FuQZ99ZINgTBFrmZqfks42dc1ZO3euFOIF4/N3
UbrVKB1ftJkLd3VtWtbJe0Hkb8HF0uekVDYIonbU9OBT/ZaU2U1s3dOlJtoOhyvR
KnLnI9WLfhk+I7wT73/4POlEwIXtM4n8SzO10MdkgZOOmjCapfEqh3SHv4f3ETLc
+keFUQbTNtPN/UbejINfV/EhOpC/iSopKuR1GfeF8IkF36jis2lX/BNpmMFpSxp9
v8gvpY3qpk3OgfXpG9xR1zzk5W4o88lnrSaMOQafkzfmyuqBBcNHh1gus7zIWViW
DF94cxeCsJbb/m0uqupTXyg9f12FLmP1OZD44Z6UjWCfU44bOPNr1u0yvZn1+dE0
Yvjx8k95f/AcvBeKjOTsJMbImNIXX+yPN8kBlvz9dazM0rjbCfaz5+fs2QGbXImz
cO+MfMkms66Xdg7pVEcBzIqaKgYOylM+kbfxLiOjvmv1BeiyIxU+/IjQVCex92I2
+CzK/xMbLEjAD5ulCcQqLjsayGjMHS6U8yoGQTB4B6Rdoa4bti/z/cWmdzeHZOqY
hKM1vjXNU6zlJSm5gEdAsBkGexMGhFQtY5tCAJw1bboR2H71chjYn9HXqMCjApSP
AzhX3dOGVbkoXi5ziHbDhmB9AMPwamHrAY2biDGafhoyTW7QbikBnQOVs6nbFiPu
YcjgH9CgFDuOHP0S1rzYWZ6ZW7zM0JxwhOhcI7wSFnXQL1+i7+MBzLo3DFzHtdF8
enIzSIwG8Q6c/tlkbwd41Vv+xS6pDbZEiUojCeWOczrYTohB2D4FO6Yyw0BEP56R
5mqCZjcEVhe9kOof3msHKDzpB7Tk0zcwvJcyDZvPYFVw6OImBycQthyfI9Qz/xuo
RXm21FMZBQKy9CujLFV5asTqJjOnI31PdtUu2lBELDk11/OvwRWfOOcB7OjT5na1
UgCiBASfhb7ub8k50Un8ROjm0C6uebrqHNZdTKPGifyRpYzYJrf8EIY0ArXirRHN
DYv2r57lqhw79v28WyKwCkYw5wNG84/u2rymGBS0FljWKt3BvBbUHF7zxtPHaNiy
TthGICpjsilUGO/8FnaPJHUdTyEyVSsu7gJtdZ9ino5fArtwycwaXgEqlVS7CQvZ
pz6+0cdIkhRebIYE1R17JRyos69+2VlLu0dAGDSXCPWSLElQxR/UgRdrgMjyWUEI
YHWZ8bVF1JlscnhbZFdc0JmfdifKl0khqfQPk3MO8b+9cQn6AjV0sOp/5PG6aeE3
RNEhROwBH6JVJ4MhCRRk2P7B0ZsFxV7cUyZT2i1kE2C1l4WnSdkQV3xHPTWhesLB
g+7bGBOElS3gd4Sjd+RTRNaQQy6P/4puEEr/ny3c942AHjox1gZMcan3FC7Tzb0C
p1lmxFhxg/rsITrDgOcL7ud75ZZfimhiys1keOnJ1bL9uewoS7mffZ9jXHGwVsAz
77VGPb9oIHwAZCI3k8eYbP7KsPq6gAeCvI72w6oZEYldLp2t+cKUsKBs6NCaq4do
QPXbjL86Ln+7zswzQVTmdF8dfGoYoQifH7FbOfv3nYQi66+JizwqhKRG0qHxa1fl
HvSwAauDowQgSOSjRVNN3bT6du41MDdjPgiRHv6zG+MgbmpAQ4GXJv2Iu3hNyncJ
8Qyrf94JJNMSg72I/EI9YhdRX6s4VtTjozCleWVtK1Sm5ZvY2WPA9qcC9PMgXYJu
rO66/7RBs4tT0PGNB/Fto1k1NbnK382xdbrEsTsY8OYO/DKzwb8Ja2O5OLAc2bRN
pZFT8UgHPFeLzD/61zZMKWq+6GBq3qhUAUC4RWCrKNvrk6O9GsGC0DCjE0Gw3awZ
kStr3oAXU/aMs5Lj4IjsNA4BGvGWkdUI8wBxYb3o1dZLZphhAfY5HF3aEwkhFMrW
tLDRR6Qf2ai5+rdtX7eNyTzq2fdN3UHJLzYKCZlyhR+hc+VpPUMcBnn0BSjeRWZ0
GSm4zA0dz/pjS4Qm7EPAeTrebolO+cRn1x9KcJ6QLKTOrqBqpXL6RZoLRHIimUhl

//pragma protect end_data_block
//pragma protect digest_block
pkMB9NpW5OUEVT1q+v5IMRGyfEM=
//pragma protect end_digest_block
//pragma protect end_protected
