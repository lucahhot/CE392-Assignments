// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
O4bYaCfhjuZtKCH8qVskd+vCNcC6GHCCE0mbr2JQWVRYcE18Jk408zlThc1DR2AF
S0Ao7oUf/9/qaqx+EoSE7vU9g9vRVjGGc1clv9ahGePavN+/093rWQQK57sLhGi+
e6vUy7fjbIekKBQGq6dbYn5x/Cs6u9K4/lkG0A9tr5Y=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 21808 )
`pragma protect data_block
A5km+l7jElW2D2ECrCf84Yf56UfZzeKMgk7OxXjG6DTeo0dhaNIb1EAAq+SZg1x0
J8weFJM8Ri0uSy8UTWr07cuEcXM3FHf700EzlsJ7H91niLOt4Wc/JN7ftDbsDIsT
iAxv8LlP8HI1GT7H7pa2xHyqV9femcaLEurmc6rn+LN1U6a+C0y1kdml+8kbk9Qh
m4dqRR549Y0s79G5spngDEZMq8T5jm5Y5ygLc402rprwzKsWpb5985HRtXDyF3tw
A1nb4TRudJf6L5A8+u1fgiqlmqf4IdGiKdjNtcqpsVpzTJoKboNh1ecdBq0kIURB
nR7P593phHgnlFaUxbAN5OHyqs+l0R4BQO680bDvfafAzTm2GyukRkCAWAX+hji3
NEeBmeRxPz2AuTVo587LEe16o/yRGU1XuHeUfTRe1xtyH22R4P6yHH1DO+t0MPZn
HWur1VyLlGj7CgfdXmMzqjDjnep+JhvhM7qoPJB8KavKhxdkDJ452+vKIrQi82aj
9MYoBI8QD0y+E5Oxb9OuLHSy/wrEObYKhAsKlBO0brChhd0jikyp6RUhKIz7ZF7a
8C0jHVVkQu/ckcS8P07xN5GeoH46ZNyymmmGyr8QuDx92keGLGsgBpxiuWf5ypDt
HPvQkYfjTDIhKAovbU8iHaEI++oC+bFPlzcwDuM9/hadOtWrnG+VHdcoYxh4Q0qg
fydht2VJhv+KpVw9fHQN+m7z1IpYoyHVyiMRbElFqDUebwI6QPt59gaATnAFjSpZ
Tkl3T9ilT1NoSUqW/VxnwrZGrRtW5RvLMfO6xTgXGQqybMFQKyk/Gi3JWbloyh8L
sK7V/35+Buwq0PnrMdjC0EyMfshKg06Yrdx/OgLCCBxLi/7Ai9YUYYhFpOPt7X5T
5DFwHtRhJyW/v9SkThRUnhryadSYbaeIcXapCKUQYzDVWbF14TvrSPPl610Fm0F3
45K3ETJ0/K1vW2uZmRQzc6IwQwkDwMjRgH2oGb/zNixNQussq6EuzeewoFfM5gtT
C3vAC6eGg9F0QglqKyYrDh9isi1qcKQfvhWsbkmF0wn1Y0kd1jqoQYD0Abk7Lca/
dszAvsJacYY53u6Fbv1ARa8s2IPP3MhJDtrVe1Ok6f2YFClx++39fiE0xoei2X/Y
yHJKpspR1oNyuMUFa/fDZT+tfQpg8jDNiYsO/+kMHEI8VuwcCe76BDa3tyeqpkJ0
4GXuQ5OgyzE5q78YCMCCqBVQKOEsy53mL5XN4hzCuHrSpQtA842Tek5wB+64q7Qc
CKQxo5Cf78P40zC9l9g0cd6crC7/Kch8bazOkJZXDNM5mqWkbSm94D+R4Ak7LH5F
rmGxBjDQ892VGSww+72r9V2C53YnqJlsO+XWHv8Fe3XAAIT7o7O10vQqLgAWsWxC
h3PoU32qw6CtgbWH29ialeEcgMo6zDni9HLXQEm2Ll8k60ZCuZUi6iw0QpbH5oL3
SG8j733PwMJzxquvZWCMlZTPSSWhszLK36QJX8G/WeVH9OxjX8imqgiGrrvAihrW
nSmWklx9y8C0xt5+O8Yl2ScqQ8W2o8DP2Da5HCZaSwMhp924WpFiE7es3C7lb4bo
E2/iWv4HfSx/CPSBSaZFe17ttKWUAtJRZp5hXF/0ReejbD3fB+SHUq7qWB3+osqp
n83VCJGB4vrVTGlPuJRmOK3wNlrpqVwP78QkgOfRi02liijg0tQqcG0cfXWBd9v/
zXSC6GTiCm0gyemPERW1TiSzl+sNU0zgkIhOEGa1i8kDMoBtstNgqBHc+YmD4IjI
fXJcpSzBdOCRL6O/de2JBcgxW7hvEA9vwPIyj1te0gGJ5uO/FFEixmdY6HYGkY4H
U7gXE+wCbJU9CUOqnq13+k9k+drA8ouUuviNallz9wiV3eb6qw1L6dd4z2iY8zhN
frZK7yWbKF6kHF07Pc5ec2id9KKtju5oXQsVDYlf9VI2W9Vi/I71aoO+gtMno4hM
8+5opjmY8rezpRQXLZ8TuE5Sab8o7DFnZyNVetEIbtNQl/VIW5Iu1fE6M6SPPA17
w6NfU7iQFaNioHYPcYdz3zGBe8WPPWZ4Hb8sp9glwElsXMc3h0981H1MWBPiTmrv
llOgWVTM2zASMheVntTX45sbyMaz65bqO5rfymSCqp3YBSU5oqW8MVXhpZP/6VyM
BVf0RxuhHVP+4CWfOLldSdJ04Uhq5acBb5S3sxAzU0wc/GazASAf3+xEI6z9s9YH
v2k+ZgjpfvTFqS4aa6Sa2dOueSUFtuSMCu0iKTrEfwfBXrRyMtgIwaKJVPHFs7y+
rOJVI3kc7lF+9tiqOO0xuYUhU7c78vqjHfFh8jJ4CAR6zAb7e5qQ7VjZEo0PK6Db
GkNSccUKAfK8IDlgvFMl9BUKk8fmugxINIKYnRXUMg1lkEksirxFGayQRusktm5s
QL+Bq6UHeyvnvifktuu57nZbPS3NRpVz+mZcAzPRgubJpI+iu/xdsoPaOohioiAx
OMf7J9DmDUzf5/9GGNThVd6mYwd0WbPktEGqmbjz0kN9eu7lHTtx5W3esp5C6qcr
beZyS9jaxCnj2KB/03nBWs6IufGrzMAXwSxXTGhR9slI9nxh9uiFQr7Fhc1hSjMX
G3Aiyi9dohAB1+1BMkmcXXswI5FS1s1Csg5j8sQaDSzoQSZBJEx2Hek+96FZhWoX
JTm7ZP+PMyshA/jOAiH0xusX1oNkWDBvnYtl6ERJu7Le7XAfkv3G6kbOt3d1wy0k
vk8Gk/tkCjflnJdSkK/303S17PsawDRD3/cmNZ4IufMIpFOPlaWJ9KZEfpYJ0mVO
BMnAF2V49iosvBcPAK3qiG9znaZsAWSkm7eNjYSyCutQue536mG+7W9Vr1v34k23
2Z11ioeWT51/50yZDlPpuYUToD8gc6tkY5MPYJOoBHm/1xAn/aqcO8jm/ZmyrDHS
heHtoAUQqQCPm8+xn1uTTo5t60pKASHkegoYv34VALGbhkUToH3JYLEyqXJsxhuj
VbckwzvO1kJAraP7mPnMy2o+BEBU8YJqrk0j5LVpfINLUVGSA7GTQqKq3zps6VP4
TWjtyHa/OFOC7xM0/yxDd2Dbu8DKGbG5fvUoUEuW67QvEhLp1Kh7uJgBTLntcz+m
Nt/h45lBnRX69B2jB/erpQpF5KPQ0vjCY313/oBc28L4xn8y5naRfx4/yvma1Ufl
LHDn8GzD04/mjQ1mDpNjLSgJFYzM1Ua5MGBRykdFMUXW9L89mFShAUYEYVAxVYpe
4nx6FNcH6ZxcfEzzwhte9X1Hi914FXok6X1WERQFcnwhCIQnYlgjJdHCnN82TFPi
NFimGf0HRFURwUsGsvADRpjwS+D8k04tvr8CIqiAk/zl0sqbE90d7PecoXdDh+Ja
MOTBV+HQG6YAmhmF2TCuhILN81SnlUy6RyTaeHKHKhK3crp9aRrRxdBmc8wSjDxp
kVKO037XwFtz/7+mJANZSjK3n6j6BeEjEcgiMbcNh6fHhsKlkJ2HQN4SQgMlREhp
HnUjX/hFEclHPe1Hr2DMboODqxhwAZQHiUTGztG3gQKiJ2OSNEA4DZka+Z9MEL4L
o7I44YJJMQpsHRwVraoxCZjHcHwFZ/fclJtdC9jgv5tl6EMQkEaw3cNluvmIi+0W
qnI9enEMn6w2eO4TpBwoQv7LA1w6ojNIwqMC4EgISI1ue505Lk9fHg4H8UiCP2Nr
Hv7mlOenXVfnccQDy5JqQ7DDdfHko4dJ8R4CD+H8Nvm7KWYS5WAAXc5IES31EM92
k36ScYxfSf8IldMZuGzXvlJ1lRVdJbmdGgIXd/y4BmZTrPIPguENcxuiOGyaHXGX
3NPZtz2E3sNmV1OuemPRCunhRBv7DrEbF/j2d+c004gpbEzromThpFAAZW6mQrTn
1o8niji+oIbOEmW9XRSYDj9k8X8YikRA43ZeULuKSeaTsAz84j2lNmZOMdwoo6k0
knmEWxlUtvPKFjEPELPWU1pl7uEnlGMmxZ2GHr9azMwZVhtkognok2Hxq6q5Z4bB
0uxbUUmWfo+GjPHQl4tgzI66YywbBLDNPmmww0DZHrqUx3tI7UL1otnRPsind+vY
MgAe5NYh8KEWOiOPJltqOQ8pzXjHDj9W+dYy9IWcuHbcVoYNTEJIkOOU5947GQVL
13oy3bMjyCf3WPvEpU6GohiDFMQfojpsTpvykGytSWqnMlqcR/aPXzj8apK44QI4
kBfZ76v+ZuI1LtkYtr24ihxKM4a6/eLy2Zrt5X+6eeT+dXHtIWIvYRC/tluwsO+8
Rxu7qizPqqGgDkrHVbm726/2p8d6ky2eVJLREZsJmCxh1GqCWndDvpluek3+0/wq
u4S0C54+sglZvk+J+sSBomBsioxvA8UZTSDHddLV6DpsqsxeBgzrYUr63A6IuUEk
Y0LNgKf/hQrtzVCxuz2oqith4OzjSmBkL1t+ITZ4TDXiqMn+am0jhErhejSYsRd0
2bZ6cZuPW1h/HGHSwOGlaA1xPVTkfskmrO4x/E4knqLBTvpZECDku/TSoWEacA1d
zpglWn1hwyrdonbjPPbvtSsVtPi5xZsDhM4Tl588Gsb5ZT9JOAoByQRIz+fnFTgz
liLw1RfpsYF4ALTZ73AJn3WJSxNhiJjKXIW68LR5MQyZefmpG8fspyPLfjR3RP06
TOYqRGBhL6kS7bDyyDgjTphUYfo/thfODGpj9Izkd9+YjsdqRqKy+qDErQOBBwBG
QHHSNIsM7+e5KNwiewhcej1BlWogvd01iqKedjvoTFAvsYdEbVLuI6qNNXHmt/+W
voNu2J3hQQhTnMyxWV8feWc72MfFTty0fupOVFwjTLEvl9S8dpYdko/R/+coVCI6
dDS+ESdDngDp5OniAwMHeb6mFBvckjOZ7QXXjyL3n0XoyWXnko0khDzMHcG1hfak
6GFNSJvcXrb2tSrv2D121EoKzyg9EZZYpenvnI2edEHVjgCDENLVU7oR0UnaKBTl
Q+tX84acmfrmHkI9EPZG0Ibc/bbkApQHDsAQTgDx7zvttu6UhpRb5dpjUmKsDTtw
sEhOzpHNzT4Ss0NcxJo3AUpCjz4O9htbeotIbSECvRPVKKwPswj+HMySeci86GmR
3bX/J5g1j0ayHeOifKRII4/YJJHagcXqzdSu/+CMk39T6JGNgWKaO+7KGP136J+T
X7snKjWB1nbqUGN9Doeh6WePrzsIroO2exacsp1EOI804h1XYNdilum8IPeG7koC
6q+Ndp6s+yG/wfR0GKCJ5S/x3T9P/dWVN3eWwYsNe6MsAf3m+J35U+lBMT94D2ai
eRqq0j6apsDtA/w4mGhAGfDZwSgY3sx+uDI7HeXV3Iwp84PA/N2xLYPKUNbCeW/E
UG1Bbv4KIsr0QcpYbVtGJq1ff98itBtMiXXDRlwWV4VzCdapZ+imso3JXrTTQdo5
b9fFCgZ3C37toORBbvuTGuFp1VsxqFsfj1e6/wwGBNHaiP1S1WtmhmcM38nhO1iu
fiXiU0PBTbGv79vKfV7AfI/joSWdVEav+z1P3nAaTHpGfeHcVcBG3yY3IuIZJA2V
hYOZtvqCfMvVNfFbSZ7t59O0Z2C3RBWbe+pVY9kBZP2xI659Ljw6okOgaOappN4k
7GSmH7OMbGc4MdmhJdUNm4qwt3pTrCr3ZPS2CMu5/QJrevLyhLQeeUDwmsjZhy8B
Rsh9z5FwuHUSmlIG9TXYSxZq/aHZL1om/cVZIwahYsrFr5KLmjxJ6rTO7uQwuEKw
Ia8+x8PZl7apJUsXX06mRAQsZj2B3IiZDR2QKXDLRYoLD/x0u5TrsrpYQznuQ0mv
0VMcuwPZd3pmwUVttNLxakN7Uh+W0bawzDkWjFGzrcNCVIGbqsUh1P6MzXsp154B
5Edgf8XqJsprSTHTCi3tbkFgfLw5Brx1kjDb2TggSWyscidmb5maWHHDH+acrYMZ
ANK0PKvgYKHaEmk+VTPkJP/6uNc/fPPeF8yH1BNyG4qKZLIZVqG1e6xn2nsUtTIy
CpXwhy49DeAuXzBkSLOaZWgIQSFMPd4MLw+9Daq4Y0sy7Msn6mYxuln5Qe0cX6Sp
NY3TND1FAm88zO5RE9vV3Y1nC5z79xlt8QFLkImycO0ajAQ6j3UgAZTM/eGeontc
iFEY844WJ6VfsqPjA8A2jyU4H4A7zR7VP8HimIti3wmu9j53+OzmsBvp6TYFisCg
HWLngDYBtjYO9UiC1aYSGjNWCY529eMOsjwiroBGAf82GAQfLqger9ru6SNWak4P
QHxD71O4udhhAABUZpDqGSJ4K+mOugdQ/vqmoB82eNNlvkJgvfB/EVAv0nNEuKTK
jpAx3Q1JAXfue07GNVxu4/n/qli6zHFOBuzLcqp95CeldBuogGfpQUuAentgzABg
gZnWcUBMYm50vKhG/44Qp4xyT2tENOvmsk6AwX4DSFuQoLVTgUT/uE7OBSXXo6rP
5djaHI+5yO8KBrbe3Adv7fO8N6vGxoHPqZptkmeXUqo4leXvMpT1HoBmGW1AZ8E7
1Dp1eE0KubILpJyGQFsHtPAmf8HwkueMzEtFwOdSy7tqt1KYHTDaLQionNhVE0uq
MMD0MBwLJepNtwgk0SsukchrOREP31ovLAGtPPTBF9KEwkEGrLAx751nDIEs5dNZ
ieeb7efhurmR/3TAPOXxogNO0oArzBpPuiMTW2lkD4ra0zAFxZhIspUCXJRSzspG
oMaKI7dmcHt1HhTNCg6M/vuUZPZK2N2CmM2rmKqyiDz3eo900kyG4Zat6RGG7zI3
/PbzfXUbIxz/0IznD5+onIbJvBsF+C6W8qh0gqWeoGic11UXv++ATlMd5gmLZec9
1cN+ILwmE9OQdpXHMsbQXDQDmi7akJq0LVWoxx55jDFt/9rGHKk8QHw3ydSr0pYq
tkIZQskeTzL0MJzzenQt4En0l0ZyLC3ZS3i7kUfg4Z9XTeB6eSghdaG3HS64HODi
cDTLbo4+pevoBxf9qM9cJlaQV2zV6MVS/523sB4uwWxR/HttSiYLjKQxUdlJW4b5
XGL2+s81ppv5YRa7r8yNu3qOlIerHAfY+wh6xN0XyK8eO9S2VdHJAiNlZ9kvy/bt
xfoUGho7DbaqhyroRDh6j/i5DmjZxSJKkBq0ZCwBv7U2kDVBaEaJPq3EohnCw8Bn
GR+bxWWnFQmFOkHWNzQWqNiHVREe18ezMdAupQFflIU1mAkbxueAt9fLkGrgu4q8
jF1F8REbBBGf6E8t4SUqXPF0wxSybDr51mVQsT9ZSVdGDfJrPZ25bCNEgjVu655J
/g7Tq4ofK/U6VpSUD/SF8PQrpBZnnQx7p4hgbGcHWxjB+MIEufFV0zh8qCT6OVw0
0q9dWgHIrCDZ5+2NpcYFqgHeeayl9N7+i9ajE/skITrQRlT6GPy02uk9Hl3gE09y
C1HiuXy2mG6P7KiFfajNs82mL8ynouJCjieOSKqoonAMhsQbKd2VR+JaafwQq2i9
VC26eFVPVNHZERjBNZ+igd2Od1H3kwM8W7YtohHfxovy0/WQeCnKc6gKqkHCL/fn
+x83YMwStgviOUR2HpHgaAQ4D7TXV5b//HyNOo5KP9UUufkRGIGQaOycq8fO2OSo
DxBPjOlKJBpmeePOAzUSYIMVp99cFlqrJuTNq/CkbR3ESl0jgLO0zsukWkOPSAr6
ogPBDNsN02AveSTqV8TVzDU2h3wT618WkuTQyuHRvmXm80e1LSSnYw5yos1f8AdJ
06HS++Pqs3WdxT/a1K6zrDdTn5bJf+dxKE0XvxmM4H0mq3D3o/BieWPlOziwO8oO
KWESyG0RKqpY3vvDBkDW2Y0nfWekMa5I5LJn/NzRHZhVQ7j8fn4pCQRGDabwZVdC
yMRjYBO189yiZrtNn9d/xcNvE6MuYyfOQOtllwf3pSjXP97LyIrfKtGqrxnOS1MG
PBF7g0KZJzEP6e0K6Ia94cfdRwyltOG/KxQl3WCeq3xnh4LTPgVEiT6saVw9ltZY
5+3vaIvW6ZtgQi1f4nhGAiayQg6zCvl1BlXU9xvV6wMTkY8W+onKEsvXJvbwxZtq
yqa6dU+Unryh2mAE1krMwNEEMh5IKp80P5g0wNa+Rr36I2hmhGa8wPCnStIJjws0
gmx9J/hFQte9epCQ3aUQSyZX/L+zN4qeM3/nYCS+p3lnLuIYD3wZjfW3DVLJso+C
x6SMHPPC+Lmf2HMKafHcAcBc1z/53IYBnFClpXPnTqKwAzsYErW58pVzy8AYI7ev
KhP7MQ1JpysXBTLZa1ONIQ4SAP1RapJI+1kU8MXHK++yMEBJ8JwwSNd1p7Avqb3k
UJOK4qYmGBgs6tyrvML8gNuNIeVXMY6I+H2EEFaI72Oi9b8Co6EtgO9TXGPfo9AW
0WE0NeQbnCLj2iiJjHOAYvV6y6ve7tGTZ6qasD8/ZnleSzOVoBK9CJMQqoNXukZZ
kAnyxhW++qxYPbMZGccQ78UcuTHtxlGPoxl7PImwG2ccCVdkLPPfPV2CzXd/+4H8
mzMHO+4p4ANPQyhxdeTRr/y/IHyVYt5A9CT6dOOfDUWXMmfnt+uTldhNoyrXKhFU
cXgikmQnW3MaTvZZpIrksCaGaXaZ2BIpRZMHVWbho6jgZCX5VOLB6HOt7ZAo/+bw
CnNSo8zHYHtdOVqxGXJklq01MzIcaecO9DGL3S71LaRhQponTBKexG7CV3s3dNeS
jYn+0rF6X6KgMm79vQ/kcaLvNsP1IpOvm/5UAtNkNm0yaBGSzMhI+CkUdGhfB56F
/m5pZvPAQjF0dKEqZJQ8OBfj4UUD7a1AfB/ZIVHN+kBI/mkmBhP9E9hv5B09T8+/
OyLAK6l3nrS/6fMOFsYodOawBQq8+hpZJ648DFekUFbAeeR5sca60+obbAAeC+U6
zxcQhHJZtqOFhM6m/9GZ3ES+IvD3uMhcd1Cpo6f2x3hSPp8s528c1T3gNyOT0yWE
OiggwNzPIabv3ehaAD0dfj6f8pY27ks/M+oKzqj9CwwK+HGXTLPNZASNNOSd0rDx
6VmxABQzBaUO1YY3wmWokTKO4c3iTfUbuIJTm6qI9Ut9AFrB7xz39SuCBEWerHoU
rjIVHBWu3E/WAwQeeD9Id0qaB4NEdTwYi8VVM2WXdQMlm2eTKEWlp05F7binG/8v
b7p79TE4/rKKGGXT4eT4BUlnTmuAlfMRewD304ddgL1yMOnRou1k5bldobspVwAZ
AMRyi+NRKxPJmaR6A3xpNw8x+h4o4++zoTJEfeQS6/oore43HOpq2j58JQE7tAyd
07YT2AkL0QPHnvdvv5CwNyj5K+ivrD4xip0fmzTcttfoPwsgsByfotzuztegvWxZ
hGTbUiVbVtchlpROd9QnZWy4Vib0IRNB1VPORh+qNZjRas8jYv6C1zhrDLf++WO+
HXUNSI2Y3b5lHJB409GdKZWYbRkdqjQc9VnYDVtbm8Izaf9A1wnnGxZ0GcFCT/6M
YnYSWO4CdIx/0kYDERBpJj4BX1lWJNnjvfd/iMGg1+lmiA4UGTQxueLaOH5FNY1A
U68IPOq3vtC1OMcSCYDxUOOfjf5BXtNBGrznG4Bd75j3WJP/iIQZ/O73YujXCp9h
0PfXax4Uyc6YmrqR08DyMU28ww9UN5zBSjrUw30vyJq6qjq93dKXDOKw8MkKlyQm
8QVwPnZtulL2peqoY1pHCpRLWxuP70NNP34X4Vr5FWHlsG3KTFcOHh5X+TGqcUZz
gjiNskH+4y81IJ6sHR4j9ineQWPC/6qDOoMUnBv7Yjk1Bwd32GGF1bnafOnCBGys
eerwBm5cUKyEbpHQFVqoA2hMk10YgXdtiOmC2SwlOyDxdn/eLlr5osQ6EGy51VYb
m8Je2GXpvyqQmBOcc5tUiL37Mhhlv9ZzGjy8nR5FoRVInR89D8RlLmbxl6HRhyHK
gwhH3kCq6o+OZyIYMEVRm9iiQGa4zCkCyp/cg3CHW+WbqOB0U5T4atDaNRpuh6rn
0ooPK4omqK/fHpCcO0uaBM4IoVQQVyy9oDslVdyQwNU4o7EHvoIKyDGwo8RjKFSI
9u2WQQxkOt/gDroHVn1KVqtM8yZc8p7ZeaBmlZW4wWqsMfBdtmtO3N0+fxgdRUSM
zkGbgFcQ7I//R7Z/jUcH7eqxFjicVjWq3aSn6U+Rh+WxSUuqednoEILezlymZMzp
cts0o8SVTaXZN1ZRDCfMPG+zmFvNmAFh31Yat5j/VNffz/sHzqf6kGeIeFPdjmcW
8js8zPV0Qu3fZjLum+EOs6liwmGV9C04kX2vvkcOv2K671CiVAEutQqNKRHXwPA/
KfoWBNyHmbqu0W7hiuy0E+BoIVxgu0Fjgi1oyRsFRod+1EpqqR+3W9PRhzY0dMhk
28LDe5dd5qNh1s0boxra8Ylg2vO/QLJbvejSpmXEUONBHRlrBNstU/pm++y1pVm0
GIXl0RzaKYpGIDuroXqqe9Z3+QP65Ohqxm6B8VJdGemOsl1pgYpDXiQ12Og3psgf
cAVQRMKY/98mTyZE36E8lfGIz0KF+qJMitT9eZiTp5FsyL8MvMVGW6oL042u3nJj
s0Tg+spPFuv7v/Ahlc+4pdNfgwc+ECrRds9GOfMCeSxMpyWp2/Sw0fs89fsAD4GN
Rqb1ki4iJVevdqOR/U0bdKIhRWpiK+6NbOS4xq1u6kHo0toYUIE4nhOF4INM/qDE
MNtS3uj4xEx4VQ62ZW5I6YvaFoX9yS+6tM1tY3X0qfVd94YmjzQF5th9PGRbb7n6
YAEcE9h5gF7kov3mj7vHiqCM76d2UVgEbA+WwHirOFsmUGaCVR0j0/H3PDdqjpPy
FEicAnr3iW7Rq2D6rWbb8SY7qUJa2w0O4tElFnheHAQChsrVc2sj04RuC7hX1h60
tSvMEg83ZqVPn2QEagaW3lCDVz5T8mZQ3dKKhFndddXvaMirXDHKaKVP2w6RL+rH
ojE65UiaL1cq3TKlPk68P3W2M//B52rULzw4JYhdjpcCzmFGtJ3olYzRxwyMXaD0
PI4XMik1eDfrBzNoW3xHB3K1RTxePFjMmJ/iuamcSEKBKYrUOal0ICYQIt9UdFqJ
Q28nvl74YJRzYeL8dvcGnj322bfGGNGFcaYrX1eOO95sR9qrVhOefOcKu38FCIxh
Yu2Kkg1Cxi8SdQWtb19neJ862Of69d9KeyCEmv2q7uZFyoQUueftKzNSk+mu77DR
dfiIJ8VWD/WAE239Q8IuL1K6ZEdeySqdO/UoyBHGER2IAWm1c9VDYQTnz2Gk+4+N
XDVtrMPZa1NQvWCSpU4oV9PZQw00NqKsRyvw4EOTdSyJECyzbanhDIJVDcZFeUxd
nd5El17Xue0MxGStr9tQqyggC5fAjzr1cLLXMGNo65x6QUpGRjBwq5QrwCtOB0BE
MTLaRQbSMe5HICcYcSWlKuN8Ha4ByTa6nONe/BsOw0HmpYI1APEh1Mu8tz3nsfdR
mKZu7/yQODRfENiYGfocmpvi554reHmRghs9Ji7JHrGyonPjEomkSjQc9JaxZXoO
LRz+4xqGnakOmFsFN6+JcKYzBZ1jREoCSR5Pf+C9R7Vwqxmg20RQPMVdubr9bYDS
2fB9TUsQLrc5g/LezGwmn65JjKcPE6GsvbE5Kt7ECiEItpXrXpxgeGr7is1uYlWN
FCmMLH6/mmSa9M/rj032l4pPhVCtA1WRDHKEbHe9oiDas0h4rx8CWxj51pqis7CF
AQ+tacVhZAxxXxX5Use58+ZIGG/t+4LkzKIOFx/5/7En8rfdpsLmj5FqTJa3/uB/
/7NB3HUOpY7VfkRLVP0tjB3yS3mf3c4tOmWML4qjMtboiTl4Li/llA7O3uBSTdOJ
Dvg86I9TjX+dq87CEDGVug3SFZ/78BI5ycepTycMn4Lcuwj2Z9I9ERGwf1MJoJ27
l2G0JdeCQb1sIrJOo4/ZIqLeUIYRgl+ydFW6b6kFqQRsvKJtVmdDA5xp0hqk1qz2
SyUyI/hPzeAL9F9JuX2VFgQWj546QkKrBauombscgpw0sUyCxutKi6nrM6u2zls7
Cc9Ns+r+6wnHXiS1Ukd9O5wA/MN5oxdstetYIXLBCv569MKxfSNOD1VEUqXXedtf
BYkQAoTIbIzJ10zpukIeACcJMhwFB7kg8BdN3rlvPL07v3ahJPumJu0wQzPYXlCT
Oo77vtN088cJOoiMvBTpZ4dtyJ2hqBdSgEIPMlqwuL7WiuhLwUQuANXtE9bbe5yQ
oMWzj4WeRXHTSvhvJzk0NKPZ5j+IQarRrYSr6/0bVd6lzDtK/jVIQ7nQC4ohFI9P
M/h5iwPriXGqV7VC8RbvxIpkTzOWTp0RuWO/agW4MsnzGrN3mTtkQwmcdMuUJmac
4535HfNQILXnbtZXldo9vUL/85Oqzqc91uw2ZGn+Sbysl2A9ev1w8ho7sGw8SjT4
fZdtCBZg5WQ7VMaIQMoBtEejIGVXXN7y/pmbv3KR6bTxQ8X1vuz9mEzvFk6vntaO
cn+2vVUFyty/fCOa70MauHLBwc5rBT8QJ05dLeC5teec/DiKvHADdsp7TrBdTr7e
Xl97eTSNSHQd+1J4wHMcZgHRnLZXOnm4D9wzkZAOjiOii1VhOdhqqdzny2PxWpvD
k9rWKnG7LPvdGzlTqYXg+8u37q6txHITC5+tA8yH1Szq+tc7E81u9eUXvOodLpsX
zgQhaI0mwywvGqG0sVyNdJ2lxvn/kbpgISh9hUfOdkxX/gtB6U9SuqR327fmFPuw
SeAdB56UF8pJaollRioQ90Bz+6oiaducxtdCAe5aJKlhmH7JILg/tsgyymz+HFqe
J3wR9yYseZAZrKzc+vSeIBDRaWLFR2amPcZMt/pqNYLRKrKjtJyZk/giZavRRdWF
8zt8S6FvIo346lmCdI0u4jEeZkb6is+5mLb41D5jc+IHrdszhx72cz369mhRCllc
VNWlqMBG62iuJJmes2aSjsqkrG6LIdHks3bZMDBxVUohMWn20dvTzXMCg6x8/ANr
zFqu2erkvp+3If5cFYXSjvGWTRZMYmnMpnCKk7jr4XioGFrUb+ZYdZrxwijvfSCp
jUkECV2r59HA36TdVMO1CMWitCKlDc0iotLEHf9+yg1ivBndp8CGwUBtCbuRkT8x
jPGWT5EiaOA7Se2G3YnyfNmCckjg8zEhyLASkKwj962eDTrrrxtgM19zrFuet4E2
z4dUMqHMPzK/irnXevRyQDE03eFJXYQMBefGlZ3POJzR7mcEBRbjqqTIPTBmahYn
Af2suuWFlCZAxQpIJc0HnUxDjJXKRtUfFnR5ztQx6Bthj+H8Wa2R1ra+gtVYA4rO
vTU7XDadn986FOSkIJk4bYUfVkR68Mq/2YzsoUu6zE40yB6dvPYZnLRYJ6/aCUM3
pa4mMpteq3u3El50SlNMMI4WU2GEl1JpdnOGnMeUFtLc8ZfRSFFqwUXFsx9PT0ow
0jayJCs00ve1P9A+gf5A/S7Bgm+DESjWqE3V3zV9HlfmEXzBnf97I9duaHECHixt
2h5vAwEqolUwHXMM1GX2kgWOJWxZSABaIPf+8Li+R5tmhelEmd0wEt8BeftjsZlC
sie6Cas/Tg7CKLcCdKOHoIxvgtxz8NnuTdV9svuf0k4XJu5eISKsle+Y3nBYfDbk
LLon1+zWIucqcDCCtR4shUoOKLn71gbwZwHglbvUuuP0ixgZru3m+UtXgmOWVGui
NkrRFmdgo+/tlO7MSW4gjHXWQFAkRIzsHTIEkYsH5DFaGItsUPUWyprr9at1MOcj
tMxGPgNxIX/eJ7Tm/DPfQ/igCcm3f626qIkKF5um7gzTNtYVN8QDKKcgUPTdgt0V
aAsAcqdJLPJGflNNVZqtZ8tUPqe5Q2BblRDlxkrUxQ1wYrFaFkD20bs97Y+OvfQN
LBPVPUg+8j405qD+6cFVgFGFuIXxo5iqBMQdMCpdoIflLqQ5T1qeU5R+Zonx/R9I
WzPx0naCavQFXqFpqcnkejuX16yfQTqCxz5xs6TiE96mQcdX/ckVYbSRjOPWk7Tk
YDkczNcob8Hbzy5ho1JJaaW+2+mnU18QxUi+YQ+awKgE/UYcAYZJXgqUgsGPAUYD
l1FtzytXJLq0MZJGdwA9FmfYB7AnBn+f1JLlyuQCycCzC67XAmtEM4dGCSlJhPg8
1nPdL/vXidQvecdlk58chcap687l52Jj/7npmJb+ruJYIUgqbyZgg14rMdazD7CL
OCtHTI5OnK9p0LYwR/HXdt0UHYqAw0TYF2V5QY62iI00uByafYNmqhpGBN4ml4gP
ISu3UMyyF/bX0FqfKK2W3QVQsjz0i00r0vrn8y9z2VslDOUAsUu9yRiOHk08hdK3
D/PJUbLbT5GdhFMG5+S6G0nloSKBkI8NhXWwFKnL438TvxKcGDwneKz+gltYGz4D
PvU2zeLd0rH8Vi3rqFw3xckZrBs2OncxTl8zJskV/f6+EniWKk7A7fC/q1DYjan2
klNhR4I+Vod0zWihpmayqNNNFsMqOB8W+tcYUcoQtJaHqtqH3gspIEeAX6cxZZlo
avy2p9pqTIxu+PjHRElQuAPa/TWUz6QW1caP9xagXyxVGYIZUf8YSYjjjlqkBEzs
1t4B5FwxEBdbAOIoolSpEyOLedE/VY9sRdLq/UT2x09D8rKYbKGq6vbPidXJe8V4
BYLm9yAGApbkxXz1ShHvxW/hN0U0VVCtFqiCvyaISXZcVDSHK07Gkh6FOdBg/pCx
jy1MavHapWYL0tWBV+sHzAfQ7IoA9sgNFqG9Y/4uVW0elKzw2hCLGsMF2ouXUwck
Ps6SxvloDVNe+8DsrW/xfKeTeylbdxy+AhYQpibG33HEKWpSb7Q47zBytYvXpHi3
8frIsa0rIIq4yu7Bw45jgPwauNKYSCu99XEO+54fa7l0XSUejYKUjoaU8Rw3+h6m
+PmREJPgEV1OR9M0LrYdHZgzkYwAWyaRYDAW+WCHa5reljUp1v1n4HavHH0YRarZ
F/ocU9P3pa/HjMj6nV7FSoR9+LgYgo5e4nTURTsPrKuTPyxbShzSuEFGWTeego8q
Am4YT9M9T2DFQbA2Ll306LO6tc1eb0sjgw1K9q7R9TEWsNkYgKgdN/YgzLPYw0T8
XoVe9C7HF9CnyZgVey6fN52ia2L5qnUrvp89wTDL4LnJNLKgI2wh585XdXPC/y2g
41gOvAiwK235D3s4V8XdY4RgKVURz46krYxNIAT608L6xKJchaR2djdYLdBhmAQd
z8U5Vs16MyG/1Dh6H+2LOpNHu3RA/02jJFyxF40PW4XUtleZS1S+Fiu3pYe4fPIq
AK+TiYXu6vi3JohpenqxHpG8t9EFcvAsvwboNBxQLb6wYBUFGCgmX2wE+MYDH9g8
lS8g/db8bB+mKfgMdWSLrPvPaKrI5Efo+gnOuO6IXAth73TYaCs84Riod1R0eXmF
nr6grzGVTqN1kWbNp0Lrib4z9gHaluW4HSl04LG9xeu8Uj+SRXhYSnFDYS2Tm/Bq
D/GaBAJWMUChWOYJRniMGQpenKBPnewqeQzvTfvGPK4cXfG5nGR0Arf1LUm/X4XM
JD3l2PWrajuaF7sGsFVq9jPA0+eUoapAyQTDDPiS+hQAb0+6B6eSr+pDccBEZFSm
q6JkXgGz+w8oG6ho/eRd+gp1xQwLPcQHCeFAPWX7bHDXhk16fxAdz2ICfO69xrN1
u6fnoVjk3ti7bPk1OrU7Ci+kf3cTPNLOYnue9oxFTe1jhDBxMl1bRQECu4SsTmFU
6R5txDPLTbRzWTlBZyn0ZnC7k4i8XQQnSRrbXM4J/kBF59+ndc+GFit6GkgpLCUO
cd3IyMajVuZoqbXYyxKYYwOZWgMjPxQK5BGcULnpzS70gLOTBJVneLMpX/t4vyG3
n658WTOc9Wgkd9L7sCJ2WCsBDtTM1Wz9i2e1/mLqfHYdeFZs/3hmQGBpO9hK9+HT
bXeF4GQaaHjbSctMCG/I/eKPj6nqvmhl0YehXwzhJ9TBZje/Or3j/XQn6WSFGVk5
MSdSaUJl41jbAnjtavaMy0GtBbkf5274Gst2xpN0SARwrmXFSmqfRs1KOd1UcKWa
JvItPtWOYCR/tU67iDdLFnxPzR0tta9Jo1Z9Idh/M3hy4/45+e3V3t9Sapz1G/xN
1cTF2NY+kF3/nFpwLBNlBceXhuhJPxNw/TVFmu789ntdQY92aPBGT1p/6p0RgAiL
keQOjlnMf1VhgnI8UZYCNTqdJWn2lKrY6cig3tR9f+Gxy58/8Ei+SqPQmSvsYSBw
IFO5XFi+IAoSbGgEFd3kLVYPlRDjOKtGKZPL4AHya754nL7L7UL/YqxU1WM9ULV6
bFpOnI9NICSHY4+3PSConeannxvzaldNq9yhRfuZSF0CyU2eTTlY+Y9BGZfSewHz
adgSCaCRla6fqh2QDkaM1az7LYClVEztRBhOlOYGxTTCqrokucLnjkfw7595l/i7
4P7sBCxDgegdsfdFH/aqgj8QivutKdAI0khfr4lWAurY8505DyBF9A0esosNWFb0
GQe7IsU7VeVGs8MFEfD1eGE0yB3gKUqI4PWEy/5ufOn4DTTRpaZbIVLpCHUdBhdq
a9Hw+6jsC9BXosOr5xOxXWn59ELqXEFMOjy8zD+g10mDQR+8yK+Ku3NOiN/nc/er
aShhTdXpJ6XeA2VEKXutM/QKhqi7n/gTK+vEB9IpNrPF8rUcjl5Uypx+Zvg1/EFq
FxGXlm+9vMbhqnfbKGVVhUcpLlQg25niqrVNDMNR8CT+FharIx9wCjL8mIprHf13
e1lnbJcB6thHpZqPk1SudpSG46htv3IbdjC0nwfr/6VjtjiPWjYOoBlECECDquPG
SC37ea7LIuxv0DYcwynh5mApjbMPHXgxBNphhmA1gT/kDtgh9c9vtNMsjuEB+44q
9b5E1h1YDhqaHHaEyMr8g4jFiAleHGqFaFIRFKcrY4TbwLIKShGx/XGk4aTx05i8
BPCE9bdQuhv06gQhoa7o6KgpSIOEIjzEt/Knul/QBWGuP7huFerrLTOUsjnVtoSa
DM2Vgv91oSpYZnpA30FKBPfHQd/Y9ayH0mB67zbxmXqPSh3+HPUPnuHXUbNosAXi
bxThi0jNLw/HvukbgEOiA0YRrhi1idakamrw1d/uWgrGxuCTBon+eFXh9VgjoBf/
PDi1ca/n0ZgGI1u+37A8hySpX4Gu3Zg086y+bDQjSk8YwvAJhDQd2UEGLXJ8//kt
/fsfxXZLET0/r3a3sYnizna5I7FFeLxMNez8RN9Dl3KYVMAiGzQxgMMAON8mFh3e
gGPVyO5Cng9fwCUQSiMIs06Oa9amzbSCTMU7oUKP3NZvn6Xi1zXId6qDMbupbApN
KqpjyhkJv+09UaDDkAt9taLb5fAVUXrFXHaAvNZaO0qhX/FBTljxtJDm+oM7oZGU
ODs7pTF7baPdH0IUQqpjb7j9Tkw6xejIswSJdri2dj/ZTfrumn6X+CTFXkoBF7hu
wCdOueYo0ziDssnRLfc+cySFTSJjIrylqxk8QxW2vcWam75axeA515rQ8AiL8HWC
lUDWxzSf+TKY3pqWER/EuKHhcST710F9zt3Q2F0kfOK4H2QkCZDtzdHHhDyzqq9e
CY4KsRhUrKoA/hfBEh2i3ybhCT1nbJHz98LK1QBTOPhz29i6p2/Sp52Jp9JafdNU
dedXq+REQtHvyhegc3vRX1jubzE0My79HvPh+hbvbn9zh0KfHgZJmBH239D80ERJ
eSRVbil1vGqZOpos7ac4A21bYOoLlNAavTTUoJ5hPJszi8nQV3YQLZ5WCEtRqbny
mVqv3cDh3m01z34x/NXlrN8/InigDn07H9kSVkkYaN182sc78dILShba1xrKqFnp
KdkvhY084VpargRXDvZ0Np9jm82g7CWQAsyh/cusr7dCpE8i/PMpR+RnDsoudbCR
jDvScS1sP8rqYMAt6Bqx2eguzYlJD7ZOBDcTEKVjzvAla4hWxaZzSh5jVEbnX7sG
7oV6kwClX0vAGzKdyg2//14kIAiNFEoxRSJKXFSoOu9zoGjAzkeMI0a1MQwja7kw
ZT0atdq9kkug92xBlD9egZy5+5CKb9+CBlYKK3wud4fw6/llbfueY28snY8M+Lvd
C3AWfZSRqm2FhX4sbF6wceShXPw4UXnihzZml9mVxbDvnzGQkQqvOjX3HZcAHx3+
dGhDl6+/STv2pxVJGhnZlPoCgbuBWA5W8MLi+iiv+XKBuAAEDdnfAPDPigOg5MiV
aixAcfQ4GhSyWXLr4Iq0AXUQgHqpsb6Q2oYfP4hqWSrhA/3xQFWHagd2BC0rbn9M
8sBOa8T0I9sxgJfPhpdNG1grmae9UKWTpoBgKNL5UakMnELrezlujZ7BUs0un4kI
tO9OmOFUdEpn97yCMPDYZyS9T10zfnxQyovVmapLDXix/9inDYWNvCm85zWIsBdN
39pNUFeuai6YQxnO3+tUxWmxm45QPlC/GnTWy3CMaoV6ZebcVtnQBBl+WZ0bp1LE
4p+aMbDvgB3guz3cesOCh8wvvpYqZLNk8NXxeWEMxyA5xcbL8KW7Xc95qCRqFR2n
YdmNyNAMC4Lq1Gv9VU+BiLVKd4x7wIWHzPeW9EW6nYzR7FmhoeKi7emfyD0VOrL9
/S6LdFRXTrxSLP61aQLYyP1Kx2PEmY/zs4bGO5NsE4Y+Y5xt1W01JOxse8z29nk8
NQL4ul4bSXJBYvyqxIjSb6Eu8h1LZJcKjWJbFGnhoksLYqZi4Z4kuMnRIKCcOBEt
SxD+V6HaUZkau3cIzCvNwP5JsXz9rgki//3TGZwG1KkG5nLSe2SlqgkXlLjQc1H5
niyyft6WEiuivNYDKIr9gapdVYOmmwrGqJ27lRpgZxgUbJH6RfmBIGYa+efGUAcv
Ob+OY8IBhsbpJWRITLuc9Lptn/ubr6XEzXSqRVOX5ctWGpO4zbTFeH/zeKmPZEjB
uEZOV5kwh43pQD6mNwlshN8bo9+XwAVZkhMwLw3JjOUKIw4YVT5saqUhruahHzAg
W/iCkpZ8xIClmgWFfpALA8iVaUMgiVF1fhy5SDtDr9E3s0WU6TKDL+fMyPtEG5kb
gB+eBijv+KRTZNuxUiwGLOUfNcVE/EFeTRuvzuHFop6yg5/UotbYtxKbuWVcRXXL
EDX7z7v8ia7odBJME8QeBRmBK0oV/RsxM0qbmgCoQ2koAopfCTp2FzwgnUZ1Qh9n
q/qGLA5nd5JxccUq2B+/Y+5fBwA9bnsOqN6mamri3+WD38JXchF5X66W+QQ9vuAi
7p1mRi9DPwNOfFT86IOxFYhH9Z9v7uh8Lf3vrU0xOtslK8J95B4MN54FIVn2fiJS
RS9IJuCG4gBCQuvQICrDNTFIg/CbU4UXjVJUu2nmdVJfJP031makyVhSIr75T4xd
X9A/fKiYUgKXNkUgljaa7iQ4syObpzGk3m/dvEQL4Uwdgb5TgIKFjRoeYmxwARcR
Gay1/5uuEWIt3Awjgt/BVVuH/7VfyZP/ek6LumlQhQRfRU0Q7b7gXDtelkzwHtPj
2tBV9T/TGY4kXUEMoeSHY6jNtf5AwLERQcJeBfXyvKKzMryp07aMNKAXAHW5nRFn
ZtA0J3j3uIkf8m3IDVQG28N9ASqSia03i3dEIdS02Mnj07aD5z5U97pCHPW2LLS/
RUz+JO+Dtj+Q6GdT79EJ05yw7sWESrNDA1moXJhMqZ7gplm6lDIoD9Vgl1Zweyry
9aGMZN6Nrd45r6qcKVzsemt24QQjZhEFjJpzXM0FwyBprThdLOBJms4IkDp36bXk
aAQlHmLFAdd8NDzUda8PsPJBb6CMpRIf9byyjlMnZ4me8sdu15y2sYsVaNef6wf7
17oVF/Itqo79CB6NSSYkiQZUiS9Z9p62j3I85bZSKGQTUurBF6qEjhRa0Bazhgv2
2xjDQQdnG0BOzJEQvmeWmTKT/O0iyqGzRC8zAeJ9j2guaId+Nh+MXHQhEAuN/wkt
CgU7l8YHP/DvZn7mWt5yTJdVTN3kVhztZb5pbqxjHbx0AQi1/3pvyRmyO+p5JFl3
e6CEoSDOhrsYR7z4DcU3o2pvkikIUazjvN+Nx3efCDQ5ZA9T7/tcnKCzCE1PR49U
tHtwbWsDEIHAW0zn9bNtAGhXDtCukHRy5VHgKwdWdObjftk5iVWEBJTDke6JxcUj
vVXiLkaQFaXoiZiYmhutVhaTqcdgRhCOTXc9P1dnNGGecp02AFGaIpFI8vXYUHI+
gsF0v4IrfvuagD7QFIKEw8EeiT0YNZObm+GKD4j3dDb4vR6l4bgEVH9E9oGsYT/A
pKM4cw6gheqMElN1/mYRmDIv3gqFjcFFXScb5kBinaw8mnutkiSReRQR+ZRqxQtD
hDsQI6PS78zazbO7yAZxckhdlErizKKbn2IPeKvg0uORsJyPZz3B5Fs/LopFWmEn
VQIVlWW8YEqYGvOn2ZkVf+wfqLjk9FaErGDIs+sLw+7OHp9fgfV0MJ4r2Uci9kXv
qJf9HnV6jOlZVh1M0P790uhXzZQi5krsM+e3rQbu+S/BjY53+tIGK1U6tN4WE+bU
MOiheTLco1NeuKZuADX7hph0JksmmYrShvQIkAAUBGL3IcB0Zl5IJeqTTR6S/YVR
eV67o/FZqXDQymqaX5vbFhLgYw1lsmzxINMnq25Va8OG3coCRe2m+Oe2FHq7ILxO
JiBOuxxmAUieClGPlTC8HIOfYwYCowX1SJd6csL4e7tug3xxnQ3sG6Ii0uccEL5N
h8+Lh2KbtYE8MavIjKJGhvH/u/KiVpp3S6CHxQUabjiUn3Du4SyMUDnkZj80lsT5
++yYAoJ+XRLj0CROkbAS68lKiXpqT9+zrnWfjkenfiECWDjHegqgleiTIy03X20M
lLF8foxG4MVkSceJovcsMKjje6u6v/XrKzO4778zWLiAvj47rb9h9UQKcDu+KUpU
Es4aJFUOIvxeODFxzyVLvrRoPXLfWRqMen3A6utgiIBhlB87uZ2K3q0S3m/2Oarm
Wdrxnv45fspEh3c7l3Jt1ooy4baPGhKrqpJoYYyBX2vzknWXo0/pO9Ww8miFIj2w
kSUkZw5DEZR15+8AT3rKYXexmn9cflvim8Y7LFXnnWjPrivX6yh3rXedcBKq7X5l
zIGR/x+LJInp1RYshAbjy5Cs6VEa9GEt8PtVs12xWsomj9d799MoGuUJMHMdJxQp
4z1HBaeVLTvhv7OgblUIfxpNUP0gnvbdRXomn9QDV1/rhMDwFrojTrgcL/7Je+Zs
j0jffinXCj0nBxhHs0PTv/Y1oSLVDn+c4Zpe1oJ30LAhD4FpMHWP7Z6kz+ljD5aZ
8m+3u6nJsuY4vAvAbVZnOsjmQ7xv/RrxJPnJJouevkEUtSqE5sOF+UnBFAd847lY
MSGJZ0pRu1QgaQhdmc8gJl3CRuy4wFhOtUF1UMKyCKCN93gmcstYp7AzlJMJII4W
WV6kir5Whc8UHIFQpmhE4LBt89+b/CHPD8vDR3jGRrMxvZhwRCLm+rSYRkSTBhNE
E37T+JZly8qsC4G8mxxK021/XidQoIeSbNjomRB+sQllpbCeFeggQF3HMVXDtrWs
7SHF98mW3uIWZax8uB7Pw817rF/ZZSb9dv/mJHVnMx07kkWKNVdw0VgGdrZFKCV4
ztrgnD6uAW9OFEgaGzvSxPtqzOnbGu/yx0c6HMXDE56xC5ZFwW0J+qr4rVFCa5Ah
F+xpa2vjZWdVbgVIU5w2vQiKks0yvhqb9Q49lIgoiEYXFRKfrxDHMvkE3R3ourAS
nKWktkgIm4YP4IyWXCu6yoAC4Xp4tyfr/pOCLxSWi0yRCyW5N27SEIpHRkcVv695
rYyR6sAEbgW+RgxgRv+WUtXnQ5nzirITz+yvAftQ1/Hyv5PGNuYthQraNvsrHGWM
1Bu2MGRZGT93otI00DjSkt1NZ+H1rwN6rG9LRi/rS2KwjEw0BBXO7Vk51lS6SAIV
EnyyXLQ9Oj4IS5QOgv3oRMOxuSg2UByNtnG+AdspheYyzedWzVaAVAnMMj9ZQ6dE
ogGyf6jpWS2u/m3ZPsEDvJhy1kErt7Nuzbb4YGjkCgBjIwxfXFoh9sl9jF6owrB3
X3GP59+M6vt1637p7Z4nsH5CAUBslPWX3F3UI2lqc2CdJ4QKwBSfWO83ULZS4JQc
UNR3TVY0NZeoBpyNahMWTpy+OPTzSmSeFTq1Mbqxt2xV6m4K5AhvXsTDdHGaAver
0NWczrR2Xf8tw1ZmDiDnfknprV8CqiICcP7IKh1acLQgaCr3MjG3Ez59R5DEAkvl
O9tZxNZH+ynpl/ulIgGtEKXDFeKulG1NaRjQ0EdY6MyBOEONP5GtMTbsX/Hsvov9
bhiM5UOANgsAG27kHLxSE01AHzsVGCDHDAgq7A5GylhDB74hTH9bPqHMivPd2MQG
EGoJuDQixvAGkRveejuXB6emgC2cGcia2LslN1p9zMCZ8rM/ZqZ8JI4UDh6IzhrC
+Ep4GXHQhagFGZLlu7gZGHydTlRzWLmnupNM2b/Dz7JKxXn+aTr6Icbj2BP3FHJ4
cZXlHypz4uNkGwj/eHheyWJjwpzCo6BzV8i6EjzzBJ+mBNxHm5Zxl3CAU9Y8Sedr
aUxF9+5Cg2AHNze/kpWVXFb50YJQuFPQUd9vv5SRl1lFFOkOfPy6AfdJiGo81+XJ
J4d05iarjkjNmBDWowYBlHgc0B/ojs6SX2ScHxMIj7ey0RLQg+tYy93pan6Dd9ob
iCMpuJWye8IAlMiXTTpfoY6nrVtUA628gkInAEo5Vy6yuc2fbXEDAhUpDibCav9z
7bLJrN1OhaQyMltgFfdwHeqWWMQolUedv/KPwBjpxdKBuCXZUoBpCOJUeSyN3Qxa
BQGtC+poJpxpp/nmKPQk3nzKHq8wZc+7PWP0agYmFNCW4Plx8DAtak8uZ3yZV98P
wCmTVhBXArTi/vPDUS4lrOTUktO8JBqXpUb0EdpXaLN2zl+AwUwKofhMV6qwuukz
MCNVrzY7HfEk+8GPZNDIDW8oKmXeuuF31gEZnfXzBoSVx+ACK/iYu5YI0wFWLxqW
fPsAfMTCGz5hiMG9Dtm+4N/UwaR1bPumuBoZcQxkqT0CeT6WNnVzvCZ91RdRbv4V
qknj6w/QEEDtw/nfhHXN6a2eJp8uILriawCQHPo1wR0YvJPQbud8rsQrKxQZh1bU
7u8ioaRn0mdh20P5SUjFM3A0sR29sKsrxAhKI6kzt36d/PMEieySP4VehdMFuS9a
ZxerLATPchEaRlVGYGs1y3Sp2LlyOKLyzvTj5pPIdOAMY8yXHjt6PF6oqmXoanip
dfunEReECQG4z1t3//zhQ8B8QEzPvrQxLaEweBA4Z/uac3/awuXrRPGImtuZPRff
0Qia/DQ5gGV+yWenlM6lgoTIduJUE5Yj6luMrlgqSx3SwuxEikX56I0k624MDn8m
JpJHjroSbg60RfXyO1bzasGuH1n85U/qGBoj14+8RuWZyZ8U7C+ehlIAvH2k9YP9
DVXp1xkV1wIuEQq/+EgARpdsZKZ3Lc+8HuM7xUFX5NNYTD6p4pCOqhp+YGrCUCDJ
9rq6ra/LjLJBZpojTAazyn97l8RpA+yX7w0nPusZNHMi4WI7cmP8BLtYYvyhwSkq
wgDq3Wcy4Psga8gIDMMDcAN/QhJjBN1K9Asf9afQoG//MgmV9dpl+DnKjLW/t98Q
R0GOngxDjT0QSsH5NVFT++5AzxJs+2lEIduchYWc1V2dCEd82VWjChdrJ+djaq/I
LGdRy/Fkv0QQn0vK1x8GrVA1LPdf916hY8FbIFlIfc8M6WdeU70kZETjpDtfmIw8
0Gky1Ch2xPV4nhmdHsoJB4FcB1tWQBCCCXN9wVIzcYqvYFmd9xok7am43xBhTTpn
rlikNEZdEVnXUrnBM42rvRXt2/K8YYlhGV3awVEVXGAUmUN3lhtv2+xnawZS0tO4
+KxGqn3O/3GJ4KxpMiyoqLQ4kNKUONqJwBNMUthc0aTH+NmJLEG43TEA7W9P8a4A
lqomeYk8d9BmTYp0t3gb42zPY86NNwAfQ+1iKlV/u/enG1nrSoqNNniVNSi1Q/71
8vipyzRC1Qxx7O+rOTFv/uLVlfasp3UEODvNJmXT3w7p4+H/nDMb37k1gUflVREe
5ji/KFxW7m9q48hU2lewqZaARtLD9B+E7idVUabmO1eFRbHRRDyAIYDBbOHY7ls2
c4a7O/ACPzcYUYnFhmpDZeTK00BCJ8ofdJVzFrZAatbN+US3K/7YOZVZvI/8SC/w
hTswHFIfUrnhyPZM2mzMtR+UIKIJ0s+/fbKpctUDhiqerc00uILbfMD9vgtuoVG7
FOe6y1wcd7N7uWbxFqzWVKe2dYJCRf68Hasdwq97Dw6kAMkJbVTVyg8w2rQz6cnO
rQMhUH/YtiXKeNxUyYxQq0qPaTskwEDa8092jvoQk8bF4tZ1LHRT1Voh1nrIXZEV
K96RiI0pXOGEP1UKotfyps/mB3T0ffKGrhXm5uzqhcqDras+d11toXn+LruOwbHO
gE5Fe/qTEBu0xwe3qELHZhecxso4VtXaSnzmg+z6K7IP6l17Hw5CItXGW7Re5VPh
lT44YTRMZXI6qLSZiy8PKt0jphnrrhcqYviCr3dLayoChxNcR1oLNADVzHyOM3D+
MCoQOpA9vmlPkKbKqED+cr4Amky8Hfnu8+8lFfk3ORBLURp/jFpw3nvuPCPthEYT
TNLdTzf1HtsRm3dImY8H5KtzgglINItHtWDI8rbDV+cg7t/GNVNM4u7qATcvJXPi
4xjSs83lS/mPd3tpmoiZkhq0lyKYbrOKd6krguAcSNY56EfM/yPqAW4DRHpj3EiA
iRV24ygqFEw3D3qA2wYRGIPmQ87zNL3X5K/RJhcQb+JPvVomDzqTYhgszOcJ6Xfl
4D9KmRXJ3y0d7TPiKVwRbtEA4/JeD9T2CZEEYqE4sL89eCpw05gXYAsRytmnrrf5
x9sdytLy50cWkCzT9GAjJCKeE6GmQlcvvjitNoRR7lba4/nLYGiwUsf0DTxfzkVP
3VTbdWEniL72RoqalkTZ3wG6Bda7K/bSzlbUC3gQSSz248pwCM/fpVHLJbY7FC7B
LEfEkDtubx5ERqM4hIdAHkgbaYftILV40YczR7Kg/HUDlgPfClBb7QLHhSlN5xiR
IjD2tmPfGMlPzSy7PJ1JA8g2KT8cgl1gn//IOfi4l49VdWJLNAimfHRa45sZMSMA
F9h4685/jPusklwB/9i3R5XSVsFLbllFvPQQ8OOg0iELbnxNqi75qL5YMbHLbja0
0vp56uXMqNzNVNgsMTDGSo8Lf9GaBY93R7aN4ZnFlLlmQy3aTqnsqHWHXc2l/rxa
VNgFAyXkPEqryjDtKXKJQR0GnG/QJ2yvlrJu2N8GK04TdGG3TS1bWKlJKKpFwcOo
IFI/pE6KtHdD1uyBkkXFSO541jjSwrl7dm0KgojYbmQ57ca5luTrvbrm2ZE3ENBp
kc94Z2CTdre8rfR9qYVoCAKo+74sNLM1VOJ7BAn0HLDH4WhQNgez9YD4B8IRnxjh
xS06nJUxHLuHO/J2cZw2jBfj6eBnM3xRPXq4XNQhIcRoEGX86AiWBCyvdrr/h4M+
mu1A4qjipmOHzz0k1FwOQHJBCJ7okV3vcH/iMaQrWSoIvJZVhdc3CtftIDcuTzQS
C5r/JzhBBymIW+tlvwvQssp9QZKdu79u3uaHR4iRJPZmchKjURil7rCMeWJFEk2X
HVo0xJP9zpdxdOaHB6y0Fs71RBT0tnNdWNXFVmOI6G5HZeEeB9Qbt/Gb8fgtCm8a
7g9FMlKM+Yy6Cuaq/80XcI6x4J7qP9m5c3lcUyfkQR7fqV+u+lSBMuU5iADHCUUr
m6kdRQIgQOIJBmMm8zJaKkw6UwtP4TX1wyLwtSGeDMdqPWp5N2npHy5mwk4Kaz6p
8STQEyY5Q/WxOc/RJVtMAtv3W4hq4ozbHnfNINHnqmpPVfshSaHguwQmeYbig3Es
DBiGEljV4FzPvVvBzpIC+9e8UpGvW7862uVumcdM9WQmlj/Z4T+xCCKnenQBwu2W
s6hlHf5B7zJY5SXxpJFEZKG8jUOsT7dScASHXoBerSZJ2Bbh+AkyxWDdsrbmpHB0
E7C/DrYak1d4q+90Cw2TAQZyj/IudwmOwMNbNB2iC/ITcQrOAyNW2qsgPl7x3T1H
Ea470I7LW29B55H9iRN7e2+SrgeYf8xQG6RTbir51jsquLs6RbISowmmzkENIvOA
mB+9jdHNtJJGs+7czrb/Sb3QXf39LbRK5mJP6eM0vkLfGKOcyI7lsevFbhDQ1DSN
VraOuhTE0MSdGjy2R1JojsqQW5b6HiPYU6WWqghDGHdefpuWAE+cLM1oAJs7XkAK
01yBvjh/hT+oyWCnh4mhLTHtKcBqlju9QUht12kQQWCjuxNcu90HTw7cL6u6hTXz
+4q9Oyu/WQFu2NzmNBmibBv0p9bYMzGtxkuUld/pvJ2TwEzYn6WPM43fPTVzmP11
xiEyFCTWt7+5I4TZWHIhK+orwZGxixJ4OPZVqiwmvbcfoES3sDtqmFo7B3pPG+B+
3wiHmiW71hYnWYcSH/4AG0AfgtdvYyP9vvX/U+6BhPrr3TezzOkexXqqQKFHNr4x
rFcZ7ECICVqm60knwP06gKNn4pG9Ce/sFjeCJ9HtWQYHUYUBAZMMvO7Cf41n+M0o
H7UUSIEoBR8JYKZdj8koEpUF5UAEBAkNwDuW1PZCxnLTczXw3c3cLrDL0f5sNl84
lBSFz6bBHfQGSNMvVfHUXOUuIzYn2R5qK/Mow+NoX/5PHdYGw/rfY6IiIUnITErS
wmDGXvxyVJaxJfBvu/PEp+BgKdeSffq/N0loVIIvmERvfPCpKF7SChVvl0NsF2aJ
qZABNewAi1BhM/0G4HWECQrUs1dJSFzCfCpRmgZSRxIVx/TQvJzjm4xr+ZHmdhPK
hmgF2btA1lFL+iRLHbx53AJw3FeNe8QvASqBlTiqAWd5at4sBZCbJ+zsnrYds0/d
W4BldrutuKCpkar20GsTn4e4nvuO/S1GIbg3mElY7NZR2pog+B2ZFes+kGwDbax7
ccCBcS6sZGfD/d9IsOvTCeSwanJDUHW3MdN7lkw2PVMRvgE338oL/yHoHzvCT+0J
CXB8iHRpnhOQ5GsJ1eExRtU5tcdw+cjX7OQkEIQCqbOwYzp9QEi7YGxvrqnnTJGR
9Zee/h+KMI5JRljlFh7zw+6pU92wU0UKP28rgFfbCJThIXxB8GImkWXACcPktwSR
lf1PqmiqOqywgoJPF6ACciAG9n4tPHfVACUGrqejxEDxHqzH2/R2wpDfVo3a5gPN
27MIRxtWJ+qPWMNIvb7AU5gWVlDnZmeKI8QuN+KlA2trcvJDZExkI3FYVcdznegr
jCtVcpEM3cVMZ0Q2scBlMhuHNIQE52tsciJPsgK4jWj3BS2EquXwQPKvmyf3wu9w
+flq8LDo5P2ZqKwVuXH+ZpJ2nMAWGEwIi+JEBwxcnXKrT7aCswfD01TlPzYtIjXK
nI8OKPLgTNCFUP7+H7TPbgaXYO2WDJ1VPeEs0ccTv1iILPOUSvo+DlT5aT2N0j7z
6d6KbLeuG45xHASReiqSxPmUwQ+8nsrVUqqSz9DPY+GDcGMXxwgttkaLGx1+kvZh
rGruGN3MQywlcqUprDY255ls9ykiJR1kSc2OJAN/gGQ1rEKLFKhHmR5TkkE8XlSs
dR0aKfcsiLbrGVaC+x+QPsa2Ats2eBqimNM5AUDKj896cRysObbqIldtMta9EQQa
T8a5tSFbTy9yIMnspJ1FUA9zkCwVm2n2KOnfLrM4QGLsubWebBpW5VRJMwYPFgAD
eo3BN2Q7B1n4nEiiT4hTgTfApy3wuDhPt5gFXeW7YWrLYzDge3A6lkpIIpqlbIDp
Gqpe/NH6U6jVYgf5jyWOAZi8kIZFU5/dJMzvjIaFox4z/ktFBubAX0BKRYF0+7kV
KWKzFM4yZ5FxoShkZr+eQabZuesYwXbr1ITptlOLibedt1aaWaHOU4fSDFqfz4CN
jb9yuq2belC9Ud68WXZez+owscZsRyp9rZtmyy02wTmlZY9hcpVMap/3lC1xgaua
DLi0FzJODjztyIfxs0yskMj+sYagCxjxTKEtrWIRuqxkxbfA4SRmOSh/g5HHVCIq
37JDP9tATs0sU3M4ZeHmPbMQGWtYOyJXYtwI4PquvvUsP+GlJCnVB2gpddH9r7w/
9ZigQhtj9Q1nuaEIHm18TeiXbmVEShmwQDPoyZ52XoMjzgxB6cXYfOylMFG0p0Ld
2PkqrGC/0QiJ59Wh6eHFw2WiEGtSd0hKxxR6S6zEarx5KHnSf58Cbdwhv/UNOhbK
XtrbUMw/dIcAM3fFrGJXR9CNDDuaU3moOEn0OyXPeqaqFO8Eht8CuuivjIzsWkzO
deaJvEROi2VlrkvE6JXDN/bTScse5l4dAjrIGcbJovzlViVGtiTcA1lVQOC58Bak
u3jyYszTJv1EotZgd8avQ3lG1Wnm5BuKdZQDGiXnnAbCiJ6dMe8pNdUxLIEBtKAM
4fZk9S72SoUm+dzhShAqVSBr1Ymrwl2Ad4buaw/5MkNCrHmJG/3b64a6rW69u7+d
IbLbJGiWtiZUViVOi9NQDmRCBaFgHWgUmEaBT4mK3xyypg1g9KqHoKqLzZWkzE4H
3odoPkHq3cd71QNPnrRBvArtDoxCMeRN1oqG84KB9+YU/3WT7ZAN3dUdy1Tg+2HK
OEqf7NCyiH77NYzq6CmDDscVabEesjb3tqIgg/e6RtnBwkj1sxub+ZqTuEX0yyo4
J2pXNMKWwjqK2cCA2mHrvYZvrjRXgnvgwSV7I+ClcVDKR4FctiX9PZ1JFGR2jIn4
INng5uupXjWrXkVwdICRIAk37VB2WHT6M9iOH55RSOY5q/9PfZatR7FC0PtY0jM1
2NWeAGkPDu8UhJQvdhJAVnbAVNpSRrIVCeTvE28fp9ggdyKTN93M/y/853iyzArQ
x3IqaBlqH7gBSXuipiM/ev9AjVOGAgdad54+oUyO/vRsf+rLpLZt5wjcK6jM4UZX
gpm/o63okZ5Qzc9cNWDUTg==

`pragma protect end_protected
