// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
1REFZPhHOZEZln6sFtZF4NdNe9lYFoNlRv64q31zbbRI/GTXW975hSvLpNv7zLO6cjrJ+4AAeSyh
vq+dcU4jpoBljQ2czlfruCLtqBp7B08o0tq/D237OnD5jtZqo0Vk8xrvREOsVIzaY08ohmC52IQn
wQ/RGq/SNONX54WwA2OBImoI7X9LyGO5yOJUlePgxqndTCqwusjvJJ10BD8L/iT+pZNHIM/mphSj
w7NwwKK7w805Eqlm7N42Dh08aE7y9hfK8t1yf2QgAGCjWBgJ4b2WeZx+Y8Fj6NzA01A/UmhOGRAn
dy52E+jMEnrhHscHLoshzsV6NrJGjM+U5DIGog==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6880)
D06KsYemCmt4mHJWNgKmbz+fDXCpDJTCI6nlpVS8FlZYD5WrN3cEGaDvJ19gRWX5b+khoPXozAN2
CkLil5CH3vEbgcle6WwUeaNYv+AQNm8ZaBTPMQktjlQxtUOr9OYhxYrOz3n9L+4R2gh//JQxt9+6
1K7X3iFZ7xxQdDVrsKL2sULjq9zIgVF8AaLvWxOvz3vH0QSn1mGQYzuTaFmFrZxmww89R1pkxWjO
8lu2ybwTrHdFOpI1rvAKlm/7BCqeEdqMPSNy0tEG35w5JBCMlQ3C88mmoFUski5mCxdUzWRtx1ab
/vLUPuzijaspsD/G92DJk0F6MRJMjYCv7uyIegbs3bOH4J/8AwlZhEsjwGRv9fm8rx7OYj3P3u17
8yPn8FM88syFrDkyAJ4Xtooz1lT5ozcgJcIBp2CzdmbB8AE/XZX/2C+Ux3/2j/Q0uXfJbf4ZD1z6
vhf7Nh7wF6Eh+DSXPmzTYdpMea0+FOv4LNSIRaA9UB22l6Owpk0RuzhekdszASBhCYJ074JOykDO
zyHsAcKMU3Wy2bh94FkmtiBZHpnYOXyernFG5bwUbyU5hs+aZQjRqMrjwK5vn0tqzLzTDCpfz03Y
KcfC6UlNtDo/E99WRN4LfQ3cH+0vWPtHuQ0hxjGk/E5BCUx4jMG6RCF6YNhzj4mMcxCBMU5HFa8H
svrCo1HPK6J+7lgcOflJUhBPwEQgB2oWFVlG/03ATKDFdHcxTTqAdFkbXDa90dm7WzbMPgGYr402
qzNP8nPSHrzQCwFRc0Ln8d2JakqnXxhoAgdhFwad5LHmWgoe+hOGX4OKTo1cXcJXiJ5ycBurPFg0
3flms91Uo1jHHx04VFiEoQ8Jvd6iigkzKxBhSO8rnu4STms94bhxPfrCHfkuVtBvVg1DqGKK4crP
DFzr8o7l/shUeuoqQsc2aI2SSfM7RhnuTtkvZBOJAKqgy2P7giY6o7hSg53E/hcsba2GjkeNOxt3
Nrdzb/fA96+u1lvA4xNMT8DvL7bBwND0KDFYgVLSNkjl8JItBDSA/Ls3llwOA+TNmYogo42b1Aak
1RsE5jcNikzvg/JlsAjRXbSdM//z3v3RZup8kxDyffM9+NCGmgqtjtnvkq4HFcD5rEdQtuer0qPs
Wl1p8tPUMVNg9NsqNHUqtdgYC16r06TGx8Xjl4PEs712K6QLNmZ3BLc9UTlu8IoF12sa5YEfSr4S
RTV2SJJV32KGsvy3Q1P+h2zkVTmwSSufPg5rE8UJjPnvBd+NPvMjmFN8GlJHsR4/u5vG6h+d+cqa
0bJOMVkykEoSG0do2o2Uqn+7Z22ZMyvQRjDQMjfeBq+r/xc8QSuojrK8awXR4nkdgaTIvwIGyluV
OdChn7tDIVlqSOwzv3MTHWrvei0tdwo/MYZCbJ+PmUpew8T9Bj+3FbJYdh8yIvXoDhKJd+YmG5TS
BlzlUqazUEB2nOkI0Sb6j4Jgcb36kNinZYa1pQR4IaUYUH8tObLmpibycMJ3XFQGpguZPKsWTAl5
TlNle2Rjv/DESau3noR5EbwDideWCsbFrLZ/hIFsDbwf46FKiuVoaiYGTRHkObwBUkgpu3YwDbI9
X9spCwSSLab4cLd4etNMf5yclzbHl+3n8MO+jysHcB/3en6Ve2cHuOo8Zj228uQhHOnYz25NEtBe
z1ivJPdXcRPVTsmo8FLXHXORNrP+JDFASb+DKhPQXBJsYC07bAeuzYvyszY4TlfuG4WHDG0oIz0G
JoRpifEZYjXhWpDG2SGyrfNwc/eseTgubDz69JGeLjfFxqFF+qB/i0WLxDYQKknxDzyghWuwJuoL
Ga6T7JMipKG1ovHBbZhml069Tf52fFJSWMpEYkeTksAlk47lormn8DdLI/y4SPZlXvnKDWWR9A9y
qktOog+k55uNpBHHI49MfgDXO2uugZj5XUPGfLB2015MrbVOVhRuWoUmkEFcT+LLSgscNWNg7Jx+
u15GEGVA+1axIoi9uWcZaDWnQ6ThjurJAZMaaPwFOSYrpFiMplT7xzQz66k6aOVph4WWv98iMfbh
ezH/5GRsbl8TpqyNc4h1pNH6yOjK1YE9lBtauUJ7bNoWyTASvRC9ARwPSeUqh5LV12WptZjtRqmG
DBV53u+Wup3VAhnGwGvA+IHo0ZSuYDzSrWi+QRgtysWBnkIvKXb63m8HZKqBTDfFaeQpZL1vroCi
U7jwnKmFXWwY9/js2jUBBrEyHbRx/91qgQuOfNLJEApKdCQGj1LGUJiOHfYY0wLfZrMuOWThbRt5
k5G7Au92Rw7750m0komJTHDXvUZiEj9nrqBvufkMZMJFIMmk+DWuFOgewUC/2+s3xp9CrjpTd92V
aHrasRtTpKMRKb5RKdQ8SX+7/3OH1DJ4kaFXqTDTgfF7q2DH7k9oyff8S39PtgPEVVYRWGjYgbmv
+KRyx5tr+Ijs6PoBVEIWakjxJWS3akxfmRd9Cu3Kcel/w7dc5F5KCN1GGN6vclfRGTNHG0YmgJ2d
IO9U4U/vWkMQ5gHETk7a9vSmXc7h47kdkHXjshHDzMxnGB+SuyeH3iSMw0Ok9PcVvs/nhByWGM5q
VNugcXPlybnRkaPHBYhcewWzmGJPILbuv3qJ36Is424gvm5Bew6C6vpT9NxKcSf/1/BflXKEHmY9
1Dh0bOuQsWSpGV5JPLx8As3yWkAOgnCYL05PQzK38IocGRIiu9AXCsb3O5TmSYMfwVAEgePT5SCl
sncUMQXgkoYv8LHU82/VW5hh00zPxM9mp1p7TQuTPxjSCRrVStWGAO5OGDSGJT/k5pHrky4jzgO3
FmjwboqRDE+ikz60XqhilOfR5WLQEEIsbzIxaXyHmaXm4SlVUBDupidZzYKcOpaF8mrG3UXW9AaJ
2LHV1Z+jwHnVUCYBrR/QKPHv72RC7J3mjn2wpzEdyoTezRu1o/nxyjDaZ88FNnA5uvXLXY4ouaxD
TaGS7QVJt8ZgKIabeET5+e6jYl5ZVhwTla/hLfuo3mrJTP2RZMg27mnv999+wrvpBvxaZtHE9XPI
R631I5opu4yj7yy091lDGlC+8hpusT+mU4+FlWFsYm+Rtiu1K8UUSD5rrhQoyAjeBj8tf3qJiohr
PuM5Rv6iIoPtUeiWmX8/0Kr4q58+SwG7kDL242RmzvxODqU/DYvXgKnyuDkZEoXNXkw24dIRvSe6
tXjhRdneTAH7966TiRQ6yxOUfg26boT0JdVacOA9T0wfqiAxb2AsJmAO98Zf3aPee/fUAcn/osZR
0kxIgmsgfuReglEfOz312zHbhA333hu84cwxCgKjD1sx+T2o2vh3VIyNPke/1rAO+5yyqlsFXxSA
Z82ro//Z6ijoIBFgrglFf0GAhgG9+Ug873ihfuLJFkaYg9ShOrADSVRxTKkuK6lGrQZ/KINPO1jq
m9kGjqyeXonekwtzp6JkBpPR5rMKBh2OwxYtwPcwu5T+nqaVZrCL4ZRd0/cc40eQNaJ3ieMWo3Qq
jtujAGkal2xsa1wNnN4ZcsRu1vnTRFSBkHfEKKgWBDaVU0GLKEL52vJjdF5UumIm2z2XxcM3EcSy
WjrHPXUABO4v/mrPl87gDGw3leLLHtAyQcGj5lY9vNr93s2yOJocbvMuGefVXfC+3jYtnMhcRvdn
YRSHv7tpPf4DnaMc4xypAgMT70NM9pSPIyWmaPtoYio4c3mhmsUs4ovVBGZ590HhJLndrRUWxLaT
6zibyzIUgRWNUxQ2LBmEo5Ss5uIs2lC0dN/tABmxMStDg1BMo3Xuk3SPvXHngLXjcZ4hH35SzjKu
SgJ9E0LcmGjz+fippe4rEOyIJohdvAPfVwwMeKs9w1T5TGCHiaMeImay18M3wlE6ovARzLAQVyN5
ruQFj2lJHRbBioPKR1kDl3EA/SgdsOxbl9Fd0ktDYBmlyd8I4dnsbMboMzLwBNHYGqnOtG3dsa9B
E6QYv2aGCsKQp0YytgOy67VWocCV25NXrbKA1vmAaKpwod8Mzf8TlMjw74T3Pki8GEz1vTwENgu0
KDdOVedWGa2dd2BnfMHEgvimBdBGxQqaEg4Op47U43CzqJQy4s3GKG8e3qs5VroKSv5yrccMFTMH
K1JysXRHXSFsiSB5jNO2uJSsJpFlxUmWOkXVnebsWw4vlqzFYIQ8MnresHKEwETVkkQeCUqJk3u8
O9zB3IO1xGG2Bk+ufIBDJgXvEIuv1SzadOBRvI14zDURuZ08dwG/9PFzTusltmHRr8Wg4xCq5t+W
vpuXyCMPohiPZ+L/ffst9LBbkvJQ3vW3o380PaSjYpnQPQG3XSgFm7qkYjKogx2ilG0MrgASYrw+
+oWpgkE02agZvjm2i1EQngQDEV7RUQmGEVE1wV4VXiAFxxRhgvUKYcRg5uGCEXzykvVOh5rhayS5
ElNCfcnGqPaFv6dhiIdg3f0BBCmEGciK00FNkNFASP7Wa7NZwD00l2cOt/WG8nJUGHJ/doQjy06B
inEEYvs4vyr3D4sWIlSS7BMgTs3QcMXbw8H3dW90xFU6SiOL9TymvFMhcD3XYYgIyIyJZZHdXG7R
8/AGzkwkonyWbClomFxZcttoGaq4Gpi21Y8iC9a10qKlrp15YCzPWqxS8I1eg/AKvRdJw2x/JFhb
7AqKZanHhn9aju2q3dslgNv/83N0EC+gzw3MzYQPCH/DgOW31nvejQoyqHWegLAW+yps43fy7I5s
Db4tiwG0WhuZBCOgrxClPaz9PGdN/w8HTrKtIq2A1L/LC1sdhX695ohA6WPcgnU9hS3sXBFqs3k8
TvJ3+ooPrVROqkAhx9zJ2Hr65jk6wqHj2/FU7/IH6R4xgd2sPyQIieifXXZl5VP6ROYAPLGqqg9b
UG/SqtIT5+9TRD2QR8UUwKesEf7r+9Gz2ToJ8GOq5z3SF7T7GSaH/Y9Jd8rnOD1T+GpQWX/KVPNs
cjr90xTV5U1PQQlH0bxX0LZymn+5eXGuZPI6mde6X8w/Yqziu/U0m9drqmcsFYi8/jJ7Rs6eR4m/
3bvVhjsxj4/m1MLGjB3mwfhi/5zkUEiuBEkzOGX0lCVakdd73yCXW/mRjmeccWvQHVEhpkjjyiMH
z3JfcS3JnWJtxz8k1yjzr4pjkhpu2e2YUIhB/JHmm+8TEia84zPTsck40hYYz88Lde8ynswOzTNj
7Raw05aKoylUWjQEW0J0Vofw5upD6zIMNH3dgUvsuiDFOO4MQGB8VyjzaLP8vp/N9QxLygUYGOoP
NdhDU9NK5MTH+8JPfOwPuB5xBm2xGVmZhZ6301j60OHT8m/vw8Zch8CWLsdEXOJq0Ip1SgEjWFMn
6+Hy3rVOxa7TfBD3tjxWkl1akwe7A6iF/aiMuPnFDSx490oQkWVieGB1O/AMPpob2pezDYha7W4P
qKv/fD2GvauD8Q3uZiCthVy7Np6IKqbhlja89Mt+d59tllFPdRQ0xSwnNhggMqdyh5jZXdarDC7m
oT6umxltG12KqTHkCbiuzOTfUOkdLeVFwuo9GKR+yPTf773OIOyqPs53tDuhs3yCI/k705+uL6bf
O55OWF1hB2CPrmRTiUqhK3N+04l/oDLnOpB6PT1f+oMJoyJFDIOs4HznIXJVMku9uTfVcfeT/svF
sf7UzLlym8FI4mKjfQy90lN8Pagb8SglnJs/6TC4pqHvbO/mESTdA8vYbMdKcwnt2rnTh2vHDxuR
PxXSWZes84Yks4qaveCNr4vY4g1RN5FlHp6zvwjuGQsYZTHHQxt6scCFqBBXB2S4ePApZm+vZE9A
QgXMw91vOAWDIU2rQvQnqCIdQltzio/6malO1sutaW5ceosaP/VgUlc2Dq1HBkcBOJZUQ6akJGsd
TL4IKr4Pcn7SwCh/j1YQL6MmndPQP8Pd3ymLuyxgw5KdyvD3TbG1kI3guTHPv/oyCA+TUuQOhHZC
nRheY8kqyQrKi5uN9Rtl3LDgvFIabvlICc77ejGT4UUu0xlQM587zcCVE9vFidTGTogB47GeoDZ/
lV103+qcAo1KVTPXDOTnQO26eIqHN3IIIlizzYluUVHhPtWPxuqwXtHhvBLSIpFxScQ8bnnzWyUo
SkRm9hP2J8xvDilZEn1P7NqaCJ8zpeJKwgZJ9aEA4nQYOZei3JK103SL51BmWS7SidycDVl4bDSt
k8Yo0awdbY3qpLpZSd9W0xZuYvvi6JBdr9qxH7LMR8SkebOsfrwSr3nnJ2atjE7/oB3eil9dIaCS
Qxlb8otLjnAB5Vt/lWcQCgzd1l934fYvWzuYhSBO/8PLUD8kZWUxhugqVmA9cad6lcpT+38wVOXp
JbgFV8REBapsoDU6gCJqFqWNBmq2kohHZyWTwVtejHVexNKjZ73/Ls8YPVyuMJwvSKK0NwseKIix
9p3tXD6bsVFNQUWrM0Ev8aGCct9r0p/J+45CdjzJtj2YvA/jZvak74LzA5WoZWRh/VpP1cTkI9cE
qoDJyaQfuQ9pbYa6oRqtw4vEPj4DeXqHzFVnR72041PV1exWWeWjqF3WrHHC1cuZli/I37LPsews
ix6K443koxrBU+Pt1Y10cqE/CQA6vyxqaN39u449N7AD7mmPquhzIHUqMg7r8dWfyKonLlcLfmZV
pLwFHli6hHoNEDUlkq30qFwOn0c6RxbyAQL6Fo86/+hiZcWI99nQvLJPKFBF43/USZarMcLwrnU+
a4VYS7pY2djqsALzjQuUasLd9bI+F003unGulgeLrOyPqKzVMMBLpuL8MkLiFm+WDE4NykwLm1Xg
I3yhM8EewpquLnDp2QMTuF/imbVF/a/1dHqANfPpDm6c62xwKTrKZT/Y3TUgwlbaDuDB0DikC3u4
9ASZjPbeqwGpfnahU+jlfNMzRYAgdvP8Vo27r07vXUbHLz+dlIApd52CvJ9v+4AYlHRTfY1+UrIE
g6Rhbd27v0/BN8RQdgeHdLe3dNWaebmQK+xdEkdbeprae9IK69G1AwJCcm7Zn9d9rxBku5reRcKR
gTQ6GU5LIDRxAP5Io8Pi6pxpFgLO6mrxt7+hdm4qiNM178EekUuAjyTuEikOsJCO609iPrU5gZ2Y
J/sF9esbLK4F0mFhcBimXV7ubVz3LZkiS/Tjl/qvz3U7OQYP2VvdELcI5Z/gr9hnV7BUpIXtfDzG
lhoxtVzXuLKrcZHYCzJm7G+EDzBduas/T6IODDrvgdtKSO49Y4oHMiL4twc82eAOfa39G9JLbwjI
mRRNWboQ6OFYkP8rRrGLmMBz89fTilXfxQZsw0vN7yTgdwh2758DBaanc0e+1f6mfKRTXwJT0G62
aYIuIhZSrLkkH8onlgeKh+1fYg/INJyBAC8dn9tkOw539aqdFOZVMRg1CB8JuDkNZXmVjtabnTQa
86YJJrv9pHSwId+dC8C8VaBwkWlp2vdMinXasxJChgfQoiPRWEX0BeOF/fbXOhAHYSHEtpPJSvW0
LmpXc7Dosq0m5hbxR8UZ4CZkz1u1cIUKELxQkD3pfE5gzAVom45azyFS1cXxrqLTVLThIhTztz/a
6xv6otqPMxXTZA0OiyvQeDII4Oy8Em2FcNLK5DVFiFtMXqFaB1jXHJklpCwHAf6VYnBLjVaD0s9y
FaptLkwQlHr7Rq7s7cop1olCHMYVQkfuQ2vzLgVqiv2c2vMJEcHVyyKIBigRobwKiSe+IaVHNTiD
LdXRUbEJw39tMtgSrfJ0Mkrb+FLKGwgh7Fg7a+Q0X/nB/qGyy2O8huU4KDV8xVT++KpQTnNl7Sf2
tRFPqPWE2Vn1a0g/D//IXt857+N1AJPh8xo8lnIqM7G8V2zlwPcuz3SwrxkemBAr8jgYoRCaP/bc
D5hH2sjM5GUGfmS0q39O1YRe2xnVlg2byxnbvFg4EzSxvxEzbjwke7bvFxh+3IHCzwdR9cOceiPg
RwltVEJvbGAmdee3Vb+OG+T4J3oztw1xj92mO8wSM2f6x0TV3u+kqSCaIiI+oOBeV0oOGkxNXCYp
KuPcoIkBbcbJJJQjRikuOo9BRZo1JNc44HFLoR0WJdGZ5umycdWO6TnvjyLoEA0T9KoAggBUuVpa
6V1PssfTkWLgiTdqOEzTLFoYSzgchlcTy8NF66lnv/apJMqEByFTQ9F8/DBAaeOCOHXETqKvwQGz
GiWxU/JyTtycuLHnUF9tafMhE5RrjDnfeA/STc5iHupShAaqhTq4H0pAGNDlfxHeTqH+IVnmo0WU
B9NkCMkLxczgSljI+1i6Qjsvi1QJ37vbDKvWMOjCpI08wlrLtwGZv83CejSwwY4YM8iuZDSammyQ
D1trcHNzdluuferJJ8VQP0oxE4f2+Aa6Y/XDk62boFhbJMPmLrI9KF7rZE/4eRsYyCqeTxZ2L41S
yLO1a17Tz5QuUt0bDi2otY26Qj2HaTy+kMrbciouZVtPhXv94GO6KpEX+c0B1iYjQDUxOP4/mzCU
NKx49xiURzGmUqrbHRhD95vMJnt0m6tPohJuwXnTusxXbl/FEGjz0I4EqhPh86TtnGOK09fOTpKw
l7LP0uk3/4kEK3U3DS6kCKK4tdeK6NPTkWwTGx7zCDwRM3204JUYAjK9IQ+IIjSEAO/egpDWkW8/
oPL8fzhASM3D3h44yl60KI0qZ2U9VfzV25dK+MFGzifUcydxl9UFz7kvlib45obFZX9xvMTYCHxY
lbZG8W1WAAEEg7dWj97EuHHM6vI/1b+RIRlESt7UjFNMpaCN4dibEuwJTXaDLrICncAxGTzcYAMf
cFnXQxXC6yraFORnmxbtkKtUEGceXUvSshxH0c1y8MFtpwzPrfvyVB3jy00Lz6Fe4MzEm9UYeN1R
POWVnufOciApUoxEV9sX5QgBXNNa8znRZ0dV/ZBm6AE4sKnNdxlO7k9F+Nc8SlzJhfosL0D/6Jj9
BC0uiS6K4XggdzM2vnZ4ICvv+9hTvobtNAbe10Oljc+UNh/ZB0L3e5vFYjI5DJ7/3F9QGiG+0eCw
CYNWBl9MmFMz9oSimfTLsiTIXedBrYK1wX4kagmganUWRdp5yBgnakzRWobPAVoAmkseRyZ14qsR
xcNS/17M9s2fSSgtlJcbnC8EnbgvJk8mvBipgLfeeWfea5J/Q58qcrkY4nbF5lqAdz2Uy60H91BN
0RuTrhol124r4kvjfqU3YNb0NMl4bJ9+kWx4ypuQZNOmxtilD+yr0A==
`pragma protect end_protected
