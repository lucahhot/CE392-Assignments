// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
IiPT96KtUzP93NCuRNoUenekB6KSqsLsPbMdydy0uxpAJG8pdTKQ8gAs40/i8lq0kdmit6uVUEOc
2wQ9HI9BkB0fr704boG1pgJ6tK6SCjS9aaaQhIKAssDklPcSCMA3/SjZjXLIbKc3zI+kADUKD+W8
T1GsE/bKNeufLCzWIxgkhARd05oXYnU3zPlyvu4+ObzaaLE+KUdMqm67lH7ykL73vA7jTVOuXYWe
vNBscg5+NjUQ9dakL2FwnWcTql9rr4/j9Idr+MpCJ5ub6AM16ADZnJKyHDvDjeQFUJjBpuN5kcm4
um/VtUUjFBbP0TBpCpWeuVG2Sbaz0itCxOmWkA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 108144)
jpc/FemdzQlu4col8/yYqr9FWQgWSDdDqBNNkET7s4HKryeJshdrl1npSySwwCr/RqefCDOm87Nn
R87lYgJYB5EzNGmSMxYl17aNDtNFBVwI9h1QSCvGumtfX1EZ0IaNwnz5WRhV3g0blP45iqBwbxKr
ybJu1x8Mwdhk1JIBzTiitcLLy3h8AGlohb4tExz8SWwX1TNdjn+ONKpwOsYxuPrmDnzVu6clYzn+
f++3NysNiZvway2V+SZ2/dnE++shJkgo1sYNb91wNRnp6HWiyORJFErpMh/uZg1Ioq2QLv1Lq1wL
hxsttsAh47meBUs7jEAkLsr3g8WKxTJLqatJ28+5Jl7WiYOUsAw0dzEY4sD87jj4VNKMkhm3Z2MF
MmeWrvWJdNfCOltlaGKv7QCsuMSnfmoQJpbRWfU+fOUnjuKAz9bQURr/9I+jhS5aHvst8aIZuUw7
M7pS43EgyPkGj58RpPp0HzrcShOMtELqBAyr4F5vIQhAsWxAagFCOUYUhNAEu9XzGV4NYPpz6wGi
5gfWKkW7TJAa7u//LutcdxnIKItAPPNtT/cMsQzs0rkJCQSz6Wuae+zng1Zc7d7jzi+8r04XKiIe
o1Om8BvrOzhcPYQgzdh7sPjPPAKZ5KUmHO2/yGumTGkudFrahhcQtTFl2bnlvYxn7f9OIXaPnGrh
7FA40ItCaFvOLBsIm/zU2ednotxkNXRXp4CgEY8fQtmLydDcsidtJvTvFFg2FnbzTyjsLdfTmFwO
Ppo4TGOAla8fFTSZK0ZaNwlJ6NktnVHsEm83aYVwmsbW5kVQxYAwOG0r6BquyU3s0o6wO2ih+ecv
Yj7TyOQi1JIeXXT8Jpd3LQViL9Pkkwi1ZwFAbs3IOVaFSt07o7qFg06YGV93gFP5+D96JGTcM1ra
4HPCoPfbTzoPWS2ZRaOA1tGJ/a2OhduymNegb4b+JZkroHTzXExKjwl7+o0s3jtpglritt2rC01Y
Qdw+64vAUenWIIINxhygmpE95SEOl/k+Gu/D92hP6T484024xhi24lhFCHxh7wtGr8K7DhA9kPnC
lMs7vlfcF0fKJh7PqHZkmUgMW2qsOTzeIyBgdziijvPBoh+4E5UpRX9w+2S7spBNC83Gdd0l7j4r
HMpIom/cLbSEm7Ol5DkZgNctc0D/cTxxsLUXQOMlvbw6uELUn7K2d74uY7M1abzJ/JtFkQ6iFF48
i/20Bd5hu8v1IGne21ukMzDmWRROIPFiwVPW2ltG9zoKbgunm6+CHY7Fwc75yXpbAGqGuoPWmlY7
I0Z5cvyJWWj7S48xJ51JOb7M4PFff5Z9qX8Ss9PrYdOwmwOWUa2I5AJz6lB1PGliK6bkT7yoGUwY
51vosBhXw6Wns1kvfj5nMTDNwqQtifIToPucJp8alWeVDnLSI144QfL3nsZxU4DlnjX23m4UE3xT
IhQetEQ6T7X0DvVQIutu9RWmaQseYsgFCSq2wZ4k5+7Uila5NQEH3fnEq6nrS/ohaQMVxoDJk4Ka
HhEqgkviOCOiwNa+eC7KDJNKJ1jWis5mnrfjrmxzrehwUtNyk/q8uqdf2Cp0mQSGlGXSrkid1WK6
hO5vdNg08yms79yEiWq4REwdvWb9qdXiTX0gcBtd+/WVRA7KKep/2jFSiOnTKgOCBTmnEdYOJtoR
V9FiaOnZk1Gv+1uWOCG2l9kVabJ9p3KnEbjIToJrHUjnOHNHlmiGUqzlC4zLS/Q12ZIx5U2CGpSe
F7+l7EeIaYOaVt7eMelVy8kxP7YdVru6rqmJ9oAH3R+Trs+Sz/dgUe3auHA3OIhS1GPP7dB2lyTE
hPKHjWkop31e0zSObkd5vfgq6BTXbtJOYfbLZnr4PuKPtccJZzzpncU2np8ajtkZ8+rUoFlo+OPf
mfvaoy9SA9kXt2dOaXYpk32lFkBUEQ/Kd5myfbNRbK7lnHsEVQhgUkj0BQ3mpAz03J6RmcRMw6gC
REgFWY3ri49OOFknAtgzzJWk2lUwrnQUXbmmzLZkyQB6Ds4ydnz5Ly4DByMcschXBRXXh9Wr/+GA
/IYF4pKh0veqPxNesraqeVt783RkwvBWOvl5Q5ivkgKKad8UVNs5Mq99Dkzz76NNKcDB9COKzb3G
xptyO9qaR1gyljSdDV2Bm797aEuqnrQh8B8JziJgXrIsCk6eRLJhYeOrEypkSS7MkDAkjoL58Kj4
g6S5PtMOUuYx2OSC8frppLQjwccZbe57g/8u+RsdDluRnjUCj7FP08QvfRywBdAQBTv7HjxgwCt/
Otym3vsm1sSZ8a1rRoF4/xbArKwkQElTp1GsMGIFa4Iedva6WqDVbHQM/v2wX2dYsQQc4HwzLfQL
vOK+1td9urUAkVSkhhS3ckHhz26EHjqM3V45k5t2bB9hMj5C6c96rfCxpZuYya0C+v1UQmGyTcHU
sQAA67TRJE+0wQ9yyoDOs4k34L2RBqaIgqGwToCxBeeojLo08KB83v9hJ8uOaq3j0y8bOChANICa
jfnvq7E7JCOEwx4ChfWhxmP4JYo6/5sJ/dj/UK+98SubKA/Zop5JOKWqlbSbzJUDyasI25QUy1DB
qAXIhPKE6YZKmAGk6sQx/9003rZ3quvpgRYIdexJg0lo/D7wrS7/45OzEtHl+b9Nj/z7Gydyk+aI
Sask3oLmHoo84n/MJux8wI4Hx3eN7JG2QDhs7XBOOEWDYvpfvZS34GqVlrEIYnLTpWGZ1D0tm6zS
RIRneJtjMiHjsvi0+GXCyfjXV/qfNfCjx90DlW/w9bxjtimky3lS+BvPhMNfMUSI/DM3g7LhIwjW
0EtUvkCy8QafH9fSN+1TsHX+reuZ5Mp0rn3BJyx8zjLsYIrhk88K5OEky3XVcMQFwaNzTQvrHWgb
fAP82lY7Um3cuIvmb7zRAaLRzZgzqD817VwoVjUSZ0+9fOkDaFWcrDP3bXxulHwAwcKmtXckK9E+
bhdwdU8wTpWohJIU5seYBCRkNh5Lriu/Xh8y4DkGUvz6kNVS07tyNpqVeixQeaDDHXoqx5r8RPGU
PJ6TZ8Szu7pvWWws05psG39KfKidvdsZ16NkUJDu1yrlWCD1JF6QiujI6bQh4ywMwJsenqDL7HPj
/jVgP1OqpfvvnSa1M0VcUDYiHur7qAO2hQDjTHY8NGRWsVE6U7BAqeAt03LndvFotqLSHU8o9E3p
xoWTqOilIuS6UPMejynR9f4nAx3DKb23+Y98wng241TvdFnY+r+Tw16rlou3qzdNjy8FOYZVyC38
kQAoKcnusZFuExqzln3XfJdY5+zd93bi8pnVJ1N+9YiPuDScUfyahFGaZycbobVUZG/yX87GwDAh
kMSxcUFGWpCCsSKZrhaMhVli13x+10FQpL1Kz3widWFfHVwuEEK39rGhDksQjr7Ud6tfFu5yggcE
Ze075R/OQ6qwWLBHEFWBqlr5IdVMG8Ti0LYj65vGqGBqHK98Afze6UfrswLQKmYmw01VyKel07Mo
rqvn8fYiXTHIpnd/nTCf3VrmAws6U5BHcmAphZDqxmQyH1jP5rYbFA9omp1w+hQaw72a3bWWX7iK
TqyKy9hrGkbdF1y1KpnYkHC7PXF2GZ8h8WzgQ9iRRmte63jGNy880EjjVbAgrgk6CXJ7tDmsqTOO
ZCPuDMaK3FERDFOUFTT4WbeXtmVccuqkLeyQXD04ahgkP5Fq7ly1t+kbULwCKc3yd8990MTbdDZm
vyswC3uQ1XOaGbaXpHnB/JEH4Y0PEq2wgbugPNKchmw9+Ot1PoP3r3UC6vv+8iAm19P5OQ4bsntv
JMwb+KPxH4iaCKYpyti6dwQyi1pgPFQUx86rCqEc58AcMoE7iQ43D4ACfBLKZ42v2D9GEHTQqvgx
VCtDK3EBuUVvQQcdtZD+q3/ExJLGjZOC5KNtl3XdQy/x5mxbqlY4vVYojVkoDhHqnaaBWWCzNFG1
fOyHrrkY0VQKQ6hJy9ia0ImzAMB06AfpNWY9k0mNPa3gJ1FKm7mFq1sbh/5DsR9JkuGXmYlolOhF
kWaPomkrMWEWD/4uN7dcD24tk/pYEv01t5ag8UOw0tGDvRhhjUFuVQFnkoqLgMGqOS93H6mPQxBV
DvDLOuwEV1ImsNi0CsEY0JsctMaiMSLhamAFRDsZz/9GOPWmDmkF2CfcQj7b1FwcOf/YIvckZDwu
AzuqjaLE5sP+m+Wg3qv6Yy95BjsTRs3xwniIQuUn5cjjiXW31QBJEpWlrdUjoPdqD5DwZrk0yrbc
5uSssLaBMF/jvoy+pysXsP1NPLHneRK3ksgUWYl7P/PKWldgKmUGQNgsIOwSI6ihbx0of3iiYKP3
p2Kf9YFl4ccOMjjYJf4bTVBxNG3hLEYUa/NtEibL/Qt64bOw1i5lmfJMxaxePIBkFSMh8DrQz4UX
ObzffM1MNe36VnrtAfR1MqTZw51QmhH90lSKQ1Gxzk0a+DGD0q92QoVOjIpU9OPfUb5zKxa+kdJz
JvHKBhIoYhOj/maYgNuMHMgwE4twCQRPhBQKsZYkc228BntEy5ei1TzruBtaFU4A5DxalKHskOgJ
+c9Zl1Z7FM8NuuwMUuvJG5ujdP/Z6QoOjn7rg3nl9gOnb/w8bhytYn6pKZobJSOoJTEwrWos2aQW
1Nb6q6HyMnOTY1ZUMdi0vQHstBvCNp+CP+2ZyR6CQGzEMLJXUh2Rc4qJo1FIIh4H5y9Hnm8x5pnj
ok6qR6fD9VwwvqkBrBqBl3iR29wzz3ebmlKr0vnSaKq2Q2wy5BjkRgWBCoyJQ3TQ84ikK76lJ3rX
ivAMYqj0LtasqSj+OHds2R/2FGYUdS/Tfya/2rNjz6RfGuPW1KdZAKf3Rc6HEEULeIqmY8dqwWWB
jTpGzO99SAJzQ5glM9buOSEXD0jnsnCcaD2JoDB0zZWoCzB3cakD9l7PinfJ66Q9lDko26sc7paE
r39bmgFy49n4/T6PVbR1aiaxv3Ub6riT3WkMhVynYUwHVBLGiOK7+UE64y90OzslP7Rgizi9vSb7
8wxyeEMADSCKbKn8n/94vwri9Wtgm0cDGiCyAqraRaDVKv9+FgdLMtdzV4jLPmusV1dxEgPV9Z4d
MyF4Rmj4qyXjX1UtkoglVuoDocl9oh/y6kLVnbcsE9E2UuMfJg8JMT4JsCLVlcApGW/sTGRxH2az
ixvPolr6hzKhc4OhdIpfj4FriTgpw9lwPSAtOsXfp5tiNO6OUlylrEAtiRSavqxtBdmNfoSsniFi
esUYChWuJnSRrfzV1ZTFNOFzvemvjMR67tSP9fXGzyWSfejl5Yu8+pUKeW1sQ4esmeQKXaJH6zot
ldfNc7lrim3To4X7+FZRMk6UWsUbGR7JtYYHfeyaU+XKTNisw4w0lZSXYaYB7jINl1Ny0vT3Y/yz
JQucGiQGYIHDoDrOCZhGdOM2jW3wQkmtFBjnC9X2mbPRy315JuIapRkivsHkrqtjVMwvOz9pDevY
sRn23CPp7StDOy8IsEF7X3VUdfSsO2oDMLS6TF0hT5IJvMY9UrVLnP/kFElXchI0SUHbMLK51YTZ
dGQyf6dmJlf8D4uTjrW9odB0VTW6mSVMRTEU90LPUmVoKmDxxzLrsTty/AyPs+l/H0AOMzPC0ens
SCoQo6MG3CfsIAxkDRRYcGCLZqlvGpkQFFwFMDRNIArUfSQvySRQa+/OcbzblN8xJzisWxufPBZ7
L9W/+AglK3R5jjsSVzzM0CXyPUQynHtZslwwIN+Ex8OG8VwMzORITmwNbeENNZNcwskA45r2ZHxo
4Qc1DY9i0GYzhLvJlcKcdAD3+MRrylsKWh4c8XbLzAfG1o0u8jfY7v1dkge2DGZ5rHLOB59Nlenc
k2t2KcO3oKINfxlUFa3UvvwIYXpCNuoGevU6V5dCS3h8LrXFvxAF1gi8lv9+0DReUo8Lo+bCPtEp
PC+8MD9Yryz42rk+xenf+vuHdo+imJdEN9y02PFxwK+Jy74cSlsUIoEs/Dm1erlLOK9I/Ci2+fYS
o4UKpWBA5u0NO1CdQ19746txsqR2BH3jXVIlHMUJCPD9988IBNwBXmyeX8WkO9A+Su9O0DTfY74X
ipK22O84IYUGvovIOmndzW1CQTynOG4YwAqAOTgUZOzjw9/M9cPmmn+WQxr+5QVCzF8nKFLkj6qS
IJkUl5on/bcyqoqoQHfQClNdIAVesWySV22xH6iJIJvzjaih1s4vpmPKSncqUoD4wbd65Kyp6F4+
BxbG0ReG2ZWQ+US0A6WfijrqOndO33e4Q6Rlyp7zADk/Se8ZNSsUl6IzV4nPywfCSp/Gm6CZvDVB
7YazsLee4BmNjOIMjGmidzmOclVOZun+vSmQ4RUxDOjEQKVzdkMI2vvtOLukISzRM6Kji2KGttIu
2QJ6qKErDtuLrSl6fR9IktR0gIb7l6vRcIZAfD/9+do9+WSnedAIOiFLHihSHf/EF+Sp1IV/2UYV
89yqVEbo0FJoftvHI+jT75lGzbRPiJf4rSGQQ5uS5QgaGx3SjBvhxYl2TPzZHcQzl3/MW2bAq4IA
pjrEVj1q4JWdiUqEStR3i27uQHH18P6UhAaqqeYTp0QGu3aM8vMQGUayRCdvgCnYm17ca/0+I1X5
1/jukerz/gNPfdYibOCtwYObTG35d3GsUSbqiE3RNsD2crkEqeUN/9mTaGTSktxyUXZH7ZIAm0iB
BF6/QiczdvNZCRFiGJzTqh1BYxWXTMclWckLeMFt8Dhl4vFLWgUoN67nBCLOB9oi/KQBlZAksBcd
upuEN/thgoDmHnDfCCgXSVWu0dMZjDzz+c1jwohk+oLPRVoMWNaZ/IsjAhmeCJNOV33JdwXlc+8/
nyfLpSPfCB4Zk5cc+NR5kK6kMebWHxrVzNzgV/ZBS8681lF10uHhZbSOQEPTT82rk0GfBJjYuVcJ
H9yW8bazSPAwUjNhoeIjqUB34QXRs+Xyh9juH7xMgH6D1yOZyQ8zQzxornropPKJvMzG8ujvUZVo
JZnQXWnGCblfhdevhqdDFyJcFqFVAE6yMOi6nPM20rAX/toWOMCwtihFNn9ULCTsoaT/FHXEyRC8
AAuOMsBjPcLaoun/GpNt/ooLguQj6E+aN7Kx2+REljksqgwLlzwB5bK/zF3eqgJ0MrIS902Jx9/Z
E+u4XZmSEdqgri0ucXLCXstSBRI1tmp9ziL8jRghff/5wmqWpNdC6ZCj3+HqrN48Xe/kz8xFMpiF
SqohNN2T3mPlnVV2mBBFFZdQLKk94lV5mOEhdKRsk9v2sG8cS8rMy2TcFCFwQ2ePJiRahRHKIHFT
yqiWKGPqLZun4ExrOydOGEwglvdsUB9/tQ1ueU/+pCHpIs3/yEACscH5Fcrbbte0rAfCp1prxC+I
JWRMj+yNoqTjgFoF1fao4vCLOZfutGJ46u7ChMrBt/DEQ8Eq2mM1gjTyusve+QegMVzBpN6mj7Fk
+DrPzXFwBWqwkwBetP09Z2KXqtCprDB/wuaBgFow8FiFdmqptAkiC8Hg41qw+PSX3jzJuy+UW8fO
QOwg5SrfKDD4E/3sVDcO2iP208ZsL+SV9958rCw7cFkTFzyFuknai0TTYcYROZWsnytvzn9tKdAn
2tvsqZeGeCbKUV8Akh9OduUyzcz5ljcrVpcqA/IIxFT2j25J5J7aeWgYKYSCP5PepiGjt7TC78dt
yLmWPjg8j2QzASUkjvt3oNkYHcTKc0LP2JgVTfJDJtvB+xqadmRyXNhHTvLd7R12YXk1uCz5U540
2DNhZF10HXvxIhz0KJfqDoJgi6jcggRWv+BVaDVUzkOIRD6hpGhIdQCFbXohpc2gNIBugBHmmIQc
dnVA2mFehC7DgWMmP+FdMGNgD8gL0rWgjFsZTfPauX+4pN3DPm/Djvlj0S7opxiqrL5gFaS1KdzU
AYxVQb2ecJ9u0meOdJXQYRVGYUKOJx/ESNhljjG5SRdFfDcXzqkcFV8GI3bD7iPmlx4s07AT/Yo7
/OCzLu0A+TvpGt84InIyFhpeVr7+AoYcIRw6znXOka9+6e97OqnLDI+scABUBRqfdflLn6W6VlI3
SsKwFRggQrX/MphAIZLaorZlIhJ/uCES+pinvUiiHOVONsOotsC/v27yC9hp6N2As25J9AxXgKpt
3X4O5qHOyh+VUVjiW7GIKjrioYXmMmtMRqkiayzsM58Gr7vIqWni2aBwUC7b02GX0fJ3P1aYwhHr
dx6FMIaeI7D+zl0Ufawq33kgb3aO4/eB/2vZPjMY9pqvW/RFZSMHh+x8BaEsoBuEbzPbEcqSCWlq
bsqU2WvcChti/w6yhzTvU6O1ueZTcJCijp1FJvEcXQn1wQhq7fOclTvK2BCVIgFMFciE2G1NycwY
frGeqHZwAA9a4aW9js7a93HrSD5on4/Q8BiO7q1ZR5E4D4fg4bvI5g3jLxmdPH/jvteEViNaziEH
aLVw4sTeor4GzEC5j9intwzN9dXwhGryOWKGowcQ0PIyxkg3WuyroeN8hZG0OSikl4MiCgmhqaOT
yG8+bVyR3D2zc8juwOK/hc1H5weGaCAoWWnlqcguUwyZQFzZLZga8ef39QNloJ6G/AXG5Ds3yuZW
BqFVhAgMuAjbmKDQEXxS4mwVh3Gauy6PpsTxsTsd/X1vF3WvjJSCops/un/2aM635gNJKFxCgkw5
R7REwCe7xVpCMoiUlZqFjMG7FeWy4qHXXtAslrVgDVtEFeo3ZdVIVKkH8uO0IKuGL5fPJHs5Sxcd
y4QC7gPkPzLhfkZInqK8cQrVyVqnXDTIai6otsLiSSut3XZYfKOdejH/tup5AHBI0zjXt4xLVolY
2nLo/jqldvn2KXCjPfPufmfbFl0FJcvmn8f+6fLQ9wou1Fb4hNadnIzk37HezK6heSRWql8vhTXh
Qozt/G8TkQCAmD67+WMrLKgtPN7kY58kkxmyTZCVJ8Q0N74bYOcD2/G1Iv4ypoHK+8Pxc9WV4rHf
mXG3XK3k3sf7IcvBj8ln/op2FXpxZPaFjG1qyGxSk91mEdwm+yCQH6tPiPacFxZdmbZ7KjBc/4Xm
LH2k7bgyxr1h1AtELVkohIU/Wpr9bKuB/+iILPbSoaJ1DAazwX7wRzrJtwOUTkHVoX0rYraG8mZT
V5Chd8LDIl0efNCXIDUW8bNzId2bevkcG4h8bFM59/1YXp0EBPYq5oPuJGI6nyRiht0X0NU4B+PV
9C+QMKHAczq6bE/Qk2oR3gPrN1XKnI/YB0Sup6jU+eEa/5Qj7/GJnNq4LQBXyM+yaSWBNMwgh4Bf
EFMpDg/h8HNUUgns1zGsy6194E9Fo21JUHN84/EjceA5qaTUwkGQfXIlwDWCa3PrMfVIhe4ltNyE
shS5E8zwSePabFCaNh+qcbCKXSsQ/sC2nmlgp/eAGkTJlaOnWPONKg/OiZSl4yRX7TiC1L5zbOVD
oSnE4TajIiaXSp8mfkGQnxBDi14v2Az7ACzZJ0LwFgwvCw+GJfFzn8nWY6M0DiLXsUP02z5ycos5
VrB/e9GjlWG/qEO9YoHCBJkAE+J0HvoHPyU7wL3zY1fXKHwMhEfw8ijwKLTLufmB2rKkJmyW2435
lf5EY+WNTm92XSIeIGcpWk8mp7WJyMBCbxO/46SxoLVPDHRGmy7Ff0Z+d/dmY9H/YoeDOkzJ635k
0AGEzXLOq9cnslbJ2kBCRNDtlJ3qRk/pMJZdVLI3d+QxPIeUYYQpEcJlHd2wh2T6SWyeexr1a5vu
dh2OOjtYImwDsy2yc2tTAyK3BuxsTFWTaWuMd8c7xa7RRbodne3TspJyO8etx1TPRsceygChKv1s
nJHsbyEaH8x9MNYk3lRMms+fZZ2IDNBZkMa3z5sqS7vhBkBgJgwv50mBKBdkmsmjBWfPBKP8KaS4
CE+6xDQxDi3BPj+7hDHFq1XHYyGHxQDVmt581+S0KhPCQy5Gr8M31DAAyZBcnCHp84AZmYVbJOkz
bldOPESZye2STWmWFV0qH8ZjqDyZvD+D6VoHGv5merXKA+gqQufTcVVuGDbkqR7s2k02+DpIRMvR
8Dhgu34zMB+dG81jl3q48uez+eazdiD9WRfnRzkfhjbTuEjxwn9WvgO2n8ztTgk/JzmZ0xdFz+AD
+Wtt9sR/d77GKSGcggwu11imb/k5+Er6dCC+HDU3d0dwHv7atR2m9mFK8Dg+Gdf9ykJgHiPlmHA/
6gOmT57vg2u5hk1pdGVqfDyWZTEJ2jdGSTGuwGFMiAPf/pcskcfnHiSLyIJbr3htLzSjBqbewrqD
TTljqQwVWFGSwoR6BjSBAlFtX4fjqGW/ec1G5sCRDn3ZHA90ZY9Kju9cF/KpXIrn8UqyhcM3BagA
m7FDtNMQMKx0q/jgpQEoRd1f9IKd4uANJxSEHdlvvpcgcIEzYXOsxaXztvhV+g/kLjVLLPD/xAkT
ADnVeaZIrwnQlJk3EXz5TXWp2HZHtX6AXRGphUDfPfnGGyzGW5comxAQRk+E0yMqEgSMrdeQtnuH
oGS1TG4kFrsTVag3xpMZwNzhoF7+H6toxyjrx4n/BqrbCfxVXaRPbXfkM5l9Wci0AIAPAcB5BlJz
MR38ErmIojfFitbhtmUcTMt5c5ouPUP0Hzw6ucXGcFuCU4ljEQtuTNIPKZkdagj322ypOLKUVevZ
u6a7meHACIta4hA40EljzT6JTz7H4IeNlh5wfiomJHIftAZ4XvYyNSVKWQe7bRWJwFHQc0cCxuOq
aaZmVe8p6P3wE6qJiaxgvIk1bs6xPWzZMG4loQUC6zNpm5WVT0P0DBpIvcdD5s0mRX5FHa34qSN7
DxxbwXd1Kgvx0nWYWeMVHDnM1vrZs6GdMOYBRDRpyifO3lydhNN7X0zb/ZlzBcdKMiEOTfR8Wn+q
Hq8Zpy9ouF+3pQRU4CbbJv0e+u50wiyePRKRRTg4vsIMaC7+IwL3Y4sqyxnr/7+sGLfk1cefv7HM
JOVBZMusRJE7IWaQgdtsIRYyokrJoqWxMGvNjqrMfXp4pBuVNtlC537BKXBZgK7jx23j/bNeKFE7
Jh4ZZwoAiztj7yy1m+68Jq1QcM4NI7ROSr7sggelM47rA7/cbTgRh+e4HP1Zy6bhEbk72kAik+MZ
U5oONIn8hGT3Wwp2TudvJXEQbvDo+jX2s6WIthtgUVI9fDphNHRmcplhQ8mMuuPeIHdLiwjITdzD
dbOIqtptSLR9X7T5mz3xJs6SmeKNcXO3Lq0la6lW99FYHclGbCKT3EtutB9kxoa2t0aKOrC5PJ1W
4qWO8Ai6uv3FKHSuNaHb61fJzSCVZL9F9PEoaQy8wpMYRIvxZ7E6NKyyjKbfVx8oMGYzCeeLVlS5
tqclvxug96pv5AvBX4yg/C+Pbht061EGdxlKrI89HO5JjAg/jePujXNt3opBSJj7cuD8AU6Fw7V8
uBfFZ4yuv6rSh1MF+AXrulZI2y7bM1VeMJAYadwKyBML0+QC8EVzBITKL4GT3AnJpMJoSVWuR93k
H7li48Cd/Zu13b15sElaxUzWO9yKEqwXv3X7ISbTkqqdbzLVWgxuADXgb4vlxc8Q33PbPVAJhrKz
lGI+2nE12iqWnk7wlJG22i8Nqt1u4BUwmWXp1ZGxySUkw5OSQPPkxKQJmAdpLcf8KqLZ0q4OcRlW
h2X+nI/FQjBFz7ZbfASUykkNskVXkJtXYaynEtjgNEW/VBgUpFMqHfgxrAaPRoagja+aHoETmp7e
YKgVB4JAzsWXgY06y2nwyFLPzC+9U9XeuLgj4rSD3F5dKB1JQZ/5hSfGhEb0PN+ULqyD6wk/RpRP
YtKfZO0GQ+gzA+6btqBY085k7D3UTbxJCGfWMnudOc7DiupTelPoboQsnONItRBHUmhV+pDvpJYQ
3OtvdMSJzmXPFaDdDhYN/svSt6dx8fa3yD4RgFLepF/1/VSwgI0DyDrlcm61t533nAthEEA8ps36
Cp/GcwK0/bYRMUrLbSId1M/88AO8+bHJVhyHaDzyXPAU7/CWpkgIBBwQGurj2D4eYmXXoVS/ISy8
oHX5FxPOMIR/3BhRA1m22UlSLyEHMBaJSiZlsA0kgo2j2qKQpUfiJ5n+N0IZOESwUSWB+fTPCGbk
MPEXfKRVKkU6flaM/u6EGdyWDkkFtH7mcNl36l5REzmA6pBV9PNaXb2H/9eQVmWNejpDdbkLbrjK
dto8yA9aIAcqWAAnIRZgjRe70D2VM7uXQoVkCj/Jyxlnj6DOJrrOOegg8KnkK92Avn6SHJzYd9TM
3V+A4dQoS/xehfldJS3nhLG59+6w9Z9mYZSZByAO3+7B8h62ch4TqYLwYLY6QnkPRTplVVpxWedR
5yrAPl0VSy/1NWstxuhlhAJdeYxwXjhWAp1LW0uHOSoRD8smSBHp90E2pR92rpniKukDpLraYk4K
R9aKKOIlRr0Z1oxOPLZAlw2KhDzIvqcZaxeolPN6iMN5fyCqCzvt1dtehkRd+sq0MfNz1GJN8XfL
7G6+fynJJPZ5yS1Kq6uXVoIdWVYtSRB26AJ3vyGvq/QoHUw5PG52q0e4lCYKoGPTu8jiZsnWBZoV
C/pjURVwgQNX0kU027mAYCwNo1vAwooVLqVYjf1hEQk8+k3uB62lWLUckcGndwMdD8tqiOAHLHCb
gG5nH23jsi/nj7LD4PNBYBST1XhaKm67B6uCLv3tRW5gUOC5o4xj+XKk96qUrbuamMWRfQ591mjP
SLLg6JhIIIhKa/nJVPMF/5So4VY8YGV2BWB05DuBqwP/FRcPV+/Ah/bmRiSOSV9hEwqAitJZv8u4
3zhP/tnIgiRtxHvLfy/7sHdHTeSZH1wJmn+L3SaUNHzJyDIBxLKd9Kx4qoc1RqzDUgg+KMNzMgq6
UnzgpAebq0fdSnURf4c+YyRphcNj/CJviNs9rleKcSI0Sp72mweWkKxzPDbygPoHDvlVDPyvqE7E
rLVdL5SJh8DdoscIdi00jXsROmhRsgs+pd9obGWAydFGrM1PBC7bUEKuUDivcJ1PE6O6IubJZSFH
L9DtDmIi74KD2JXtP7OdEFfir1Y2AL6UtAKAOuk+eEkbFtIYpDxBPgAyC/xiNvWNyY0cb6xaTNe2
UQuL0gPphd4pWu0q/Hubfe11prpDDT2u4zlyi5EnjS8Mg0B+IrKcQBbugXm58Odha7cvJ9yKeiU+
6gPVZNapSRU11s9OiH6eFNsTiW7yqRi1+nJvh0Jc6CTOa9oVdQ0mIi344IdUwDftylAO4sPUEGjS
KRZbXlz/0/tZ/qdWCzYKxA7xvbgMUphvUJAivZyTmj3ua6s00ySo4F3lCVH0XAxzqHDkHCadg83N
0qp8rYDKtXnMgTDqlrcFqPeSCQjbAl3khsdJ4JAZG8wdPVug2q5NLwPn7qy5mewjhTZmQd++PZc5
ljPeX1MHczmBOo7KTdEGjrmDF7NtZeVPumUcP3jSQwZ606+bGda1BkprDQqfuXyFrlljSGR/r2t4
mfRF+eSSF3M0lW78OpR0hMtEjG3NT761dO0fAHTPZxAx4zQ1h2QUfjo5hsLAIQpAiiB8yfjv+Mvu
T4KpAs/g4DySOM/vQRbYU0VNsO3RmUVE8eJqGK2y6M7mrTFOFr2PggmUtByysHVjhJbvdnZBdSDk
8Ua4JoX5h4/4DVtAuRxbf4k8Li5sZNNF4ekxjK6cvpgWr/xRM4M6LOa1AS+FgOu6AS3ngpuw83vT
OXyr1vRGuJ0+keF5Q0K7ac4GLkMS4ZvLG9WYjvhuziLoypSpLIm4L0VqqPcjYKFVJ8CgnjGJMZK2
yaf9jQAOqYgLyoz0DqpPcMX5A4CfEdNAV9lRb84kV30FLd+bQLdQ73dY0j9dOFIS6SQ8eIKM/jOI
w3QcYKQ1oY6rQw2Yvw4vLDw+FXmZtKuqnheBtCfBt9vg3y3ozMj3m/aD34QiLxMVmJPiZ87/N5x2
YXIlVfJxvTddOai+ZAVycQoEQMNbRGOL+4tEE1S3gROw5OQruTnTZ7lEzQ/zjD/ssjuT+L01CCiy
J6EfkI0ZNJNwVEAMINudprcTvXQTnIO8WOeewAH+J/SLJJMunmgkg5YKjBh0W67t32MSXZpavJn7
amwMQK2DUotzWkKOe0KHZ+2ylONGv2/RN7QpKZ1zo0tncZTI8MJWn+sEgue8CJKIFkHV8isDggPj
SnQCGab/UcixMMKTloENm5G3dM5QPpG7rtmucXl0Jb26/oCqU9BOTYFzaqqSfaXj+N2ckEzfvxt0
WRqfZiHxNseyPUMb6jHMjA24Gs27VBN7QWfmWVMba3lkrJcRsIlYsq3rm4SNfPwcVkh9L7HASAz7
Bk4AYW8vtyVXCQ56qLPpVS54EfQJP8OIedAO8LdvtFy1OiLzHhgwwuv4sboTZui2HSKbvA+MhMZr
Fw3SgKb3zPtKlCmzMxJSMX74BavH8UCLmw590RcpEP+8rWsBOEObN7WnyLyqW2oYs9Ky4oEq+Ae7
6DImtS5/KpR3vFS55mbhxZuJWGCx5HQjjYZvVUuJwq4jMPyY8CCs7CPhh4frxhvq7E8Oi7nIHywA
LPyQBtFQ3Lqrkp2MYOynTCeKWAcmLLAJNBf8ZbIitV/FzqpI3/Tco3kAWvq5oOgYE9aGaIkXPMEC
ir8LedhcIsgog+rH3OI4yXy+L0dQIYqFZmMVmzHS3zLskgJ8LcOjNZ3YEnQL8e7q95ZFXklwRtHp
ERdnpT2j3NX5/7rvziYhVlcQkie0YqXbaECdCuanRZTIRrb8SQ1wGFXChAeGVtXCHRgDxwqIPR1g
YCa+GEIJ+T26zfmm/K1TKViZyuTkUwYObwT2mCD46FuqqeZjoRh6kLzvXFRZINXlpN0faNl9P8Ad
hkeVcAMZZi9EcBBXlTG7u9WkvaNsHV8UK+SmEkKrrGq7vAPPhbaUrObJpQtXxVaGE0KT+HOiOfOh
UlHCbsi9sjtns9lBWz6AbOAGJbxoF+JCkmcUnLEZMZfnHeYD/u35ekLDiJiYf8nd/UugMmgkjEyW
VZR+oXSfJkewmjYRFK5MKcHAWCRJcAT2hfnuSXBKM7txLVxzpqhEzv9UH5U/fHo5O3Hrtf5geHco
7G64fIFDe+oKU4VxMJElJ15dRodcIZ36GW+ruBdgBHACl5pgAsfAMf2r3G98GjtLmSYFDLSJ/Wrr
sU/Rc44kgTZKGNIhL9KRlq9QhH53W5Ts9EznLnHEqWChMwWUn8oSZHA0jhiGOnZYkfb347QJiOmr
ka6Bmp+PqYu6muhcdlTeTqKj1w0CvpJqLXHNCzsjuz2kDuJsKaaFXdap3ShwA4WfEOBY/Gerw3Vy
6Gx8PJCbqUS+BZ4vMje26lKVlaLzfBGdE3pd5dulHFSbHnbIw33oMfGSzbFQvQcwdtQFh1AS95HA
NtjCDSzpq6Ooep+rJivw8wYqdzQ1MVvwcR6vT8g9QNRNgJ4oaZhs9IWcXBvC+MPKI8xvdCDNj6uD
qqkLjV00SoWImqDfWilq4ilC0EeCACiBmXkkIW04Kw+95fqXm/j9qTFoKD52Z4piNIY5uCRnwJKi
0klPJbOIF2WJ06TPRbQ6P3lYEI5wWe2L3znK7GgSL6R+sTLfw5/qo/MTi7uNJfQ9ivZnSB77hBXP
DYxacs9EvJpfvQiggF75WCVKuF0BsIvo2qdOOp8PN6POt+Xuo/mujjJ2ftA1q1aKpcRgGfLm+qNB
Eu1u+njZoVQlL8+qEvvL8aoR3S8HV/9dAQHDGsqiNHcQpo70YASJPybt4cBsZoWMNDdkVgBg4J0V
2xcYtkfhQKwdaBPgIz3q19usIMw5kOBOlHWgmRVzjHSbiH7fbuZM68FGD9WHdn+JqbLYNMtRdozM
PzPEYyDcd4vHuVKkO5s3Hv5hsi92bwDkYpWU05UvhsijSg2lqMh7iX6CnrYCxC3qRKdXt+5h2Uvc
mG752NXbCTzYHnu/8CI+AgrS0udy/mT3eXKC7ZI4sd+5ghqoWUfxew9nNIv25nbsi+dWa3AZgreZ
U4b+r8jm4r6+5Mln6Ql/w8yIpCC6vwHKj8Q6Orob5o1OLRndsYH8EANwg6xNQ9xS6/jbtXRNMtuL
SY2CD3GgAjxK5iMks/jZEI2ttN/oXiNalVbQlrPSDld/5RtHXrgaeZrTGxvBvzAgfYC5xDkETxHu
3LTy7WXH/Wr0JLYh2Ed/iK9F1ZEGN0qw6YaX6CbNaPysPG1FaBvg7QufPB+ykF5aVT2vXJtTNtx3
0OmFQRo7POnSilps9OMvp5Y7MUDn9nhMpYCmywr8poYjbfNWdDS7UpalnFq8OR/9Yq7tDicMX9oa
ExcdFLrlCuMR3Av0ILg/MMi8BZVXy6gkj2NCw9aA0a3q/Ls+rJMP4xaBlaA6uCZ/J1xlY+jB52A8
UU9HZbJsAzZL6eaIO/8auBRpsrB0r0Bxi9ytxyy2Ax4KsfCmxxCpGZDkwjfX0t0hkeNh5jgnhmCw
SuyC5k5m9qF4bJnPLJvayeWl43UIBRg4gY6DJe55esddqz9RvvMMrD88AlZ3r3zDyBx1xqkN2+lt
sMzruG3lBAJsPqFo5lcqsJPgbNoJPG+3pFwwsWXuubaMmyh3562K6COzOY6ln1fTu1URrku4vEKk
80FFANlEzw+5fMmN+2EM1D/Uo+7S8aQKX5eaR8wUWwv2H0YZySv2xm/pMnvmYNQt+LMprKVtuqox
QTo0ejmHP2po21RTcMQlHt9cL50OUPVjOTeJh5PdnPocmVAXTP1PDnta0G9/8fPRjloT8iQrywY0
5Bhbi4Y3/sM//crYlqfNEYHuvv9h+9sIjnio7e89aDusd6upbFSE+hL+Y9q9K948O3doPZ0jtWpV
Ow8ofV+HUQFJU6EowyhWT8ZmGA0ULse9FdUzt7b8sUmFNab1IDLX12ff7dplm5DWMZYFmH9A6SxP
xh4tGbNNsoMJIjUqntMBdsRVTxgN9Kgvbdb7TywpBVsCtUPttIEKUqiqj9+8Uit2ZVEmcX5JAnZJ
R0FHIl1HPN0INXf8epVs8RGufYznI5RfWxbZr+6nu/VgM+T915cbo14F7+n69FGt0grpd/gfQOBx
CPrYA7Mea7TxG619VBIiwDUlkwv2oqTII12Ygb/v/F6TnKAZGNmw/8/7shUWrkMb/ykb8kLXHZg3
hhlHolYPNAMbzweSYMIG73iTY3nOulXEOZBkSuJT8SnVLqDh605JluDyb0FZS583Pz0dxQyynHLJ
hMnqLoAym012P8QESYxun++Aqt7A09tcTGGy1h6TA2hEkywoceu13vTvTQ8LQOUBZCibh9XL/6Ma
OqS0BF5/9O68qThGbmiRm3l0gtDlCYGJQNQuKLdrN1Be+H7A5leukpfqIKneZFB+syvxlhfZyiwm
yhFHdfOHja9ULWIn1HWRdwuqDdmu5HGp/sc5setMi6TnzJW1X+kEi8vpHyib1jii6I7ayUq+r+jn
qCdkqfc/Qh2HJSR+cPaQh7wJvKvGNG/C8ugd+9rHpWYsHrgDn60BTACYtptEudlVovUvSkJrJmUE
ks5CAkg4fx3ZDlEi8O7NxzbwUT7QDxXTcZZ2ELqu+QrW2nttWnIvx6ejOaQfgpzdCkbYLamuuoXj
wDZTw15aT0nLmlJIEpoEhbxJ+evgAHt0nfGy8ltkZCXk91A5K20eG6ZqiHWp1xjvy7n3+WzDWK0/
R7aNg4NObK7BnxbvxTluoxYP5CgunnpMIKTYr7cDafufl6f7OXlUeuv3swH3pfq/7k36W0sW4veN
9Y3IBHXQSQ3hFE+DW3CwuC1gElZCszRuau0+zZe9mNdsdji6WcCAqXaHLNx8Ml+9NuhPSsZA9f1c
bmGsYhkdKaxbg4ENPOQBbPZkVPAQocnlQI5U+DW3ump/cEr2qKNBF1Lhdl2JDP1dpbluZdOHhUNo
Hcz3n7IRi8H4tDCd7TB5uA/75LfS9vARs3zC6KujcqlXPOzg+atYOaVo+6zsuwWbin8K077wb8OR
+6n0gaqiMHVqhYFp26mfZiaMXo9LLuVoeboNaK4NX0tNYPXPfIhQat6T0aJyYNdSLAsre7IumpeX
RA23Q2oXdIXZ1rQjVLCIhyjiYIdVRcOuSdoYK/e/9ea1FMFxxovhJIfSzVymuZaXmfb8Wa3p2XnH
23qeeLozZRxHkXqI20KW6aXV/SxNfsSOi5Im6tPMq4OZIB5ZcleS9KcLtk3/0UAFUecai1ZhPl16
ifGpIuEl9CaF/PIwWR4qShIII8lz5eRYDxotxN1Eql28AXvlv73jogcgnPr8dcrwvL3iOtjAZAh/
6c5MWyUSvVlV4g6b8iiVsZM+bNRjqSu+X7+kzExl7IepNpK2fi9WevEM45hyo9r54JwEGIS5Bmvj
vDE53RjcAoH2IO02N1OmoeH/E0cqTGcPoC928aW3KwHdl2AincksxlakPeT4JSX+QNo3f6GjNj2M
CVa1yiDrIJyJT/j6Mem+TOvaaCkLA2/BIre2R/vZxqQdiuwjiQ8qdLhZPzpXuwjXAp4jsf7sXxQi
zgg6F8sEo7GzmFflZsFvysOVY67yB0qKYamrS+UAEhheToOCyQJuB2eqESjJbOAgKthKq2lG/Pxc
6IChmA1FpiYjRewTaomBWBX8lxfWojPED7ID85oQ1UwhRM+Uf/doxTnxgIFdd61jF9gm91ACdb2w
J7spfuQ0IEeydoqhW2kiFO1eHvdyEoWQrs43pgaDf6iCSM8h1v05MLX0Q96pWKB0hPZGYuSPXi1s
w3S5MPIJ+A6hcin69vI/VCBJgYI+iH84JicYqo8gBOmiURh27F6TPGyvawq1Svy5nE2xtCBxQPd+
ptwPasQyZx+ORycwC2cXrN+6zQ2cD3g/TdVXjbSezmJDqVwxfDE4nEbNu208bNVQMr+cLIWG1DTe
Nx54PWWDKm6yNuZl4eIBLY3/hAOUmNfFAHyKPgTgIcgcGEVtKBmWpBiudZTNnXw5BGqb1rSFEabQ
h6zxuJbgGAxdoos50DDbfYIo7S+qrA1+pZ6IQuOKZ/M/VtULsnZF9DChs6Pdl4m1CWh91MXKzKIr
vMAzRu9DPIH43MBDVjVLwLIx+MBC8gsJ0RoCTBEuFlc5sCku9LvF1zOgy7hMQkY8fJ8lRU0cA735
ooCBeEt/hLKfxtnxOZW3mpxQmBOG+odv3FSGF7SJo51boQopn3attsAlFq9LzTPvxv1c5Kw5tNR7
8on/Qh3Q/c5AHAcA4TD5px4OIAPJ/laQ5q5+fSFaxyx35RKAQiLXdHQ8F+ohzTCjZINeXE9g8V4L
97G+oYpsg/UYKakmxiEJvjsSnpqLE04zLk6RjB54qDanHIt/meWe19aP2uLhOdkRdmEaG5MEMHk1
A4CmbLLHfl0dmP+zCoeP3CXwzBt5UjsNA0S/hBXu2RRiFaRFkzW0Xn8lSLXtRHHDxjq+oPqqFFfe
gYUzTOx9x/RYf3T13YMEhC20bdaqRnafNL1rwBxGM+p3XfPW39AHkZw/fJvgLBh4lFXhh1hiuP7z
G0GjCdpBU1GmaqpCFSXuvmfkIzasbRs2ExvWPFrjXxI8U2IdoikQ6J333NHSTtbtKQ94U4HmWc3m
ZIgU6HaIzSYX1iL6XpyVSlrM6sAWVaReJLC51SgDgJMW0uZpT9BLyl47eSqfD/1u+2rXMKzE79XG
RnucHyUrmhvRHofl8H6J3EzQl/hDZZRL/gwz2qHD9RgJCAoi0MFvDO4DQsREiXO25nLvlq450xDy
8FX6O6p/KQPTlOT0CvJYK4nIAFugCAmbqCzF5KaglVioqjqDqP3pOTgM8av6igmrsjrVn3vKjD2q
ZjfVEBBgUGrLoi60oNxUlzdJnxdfNfWPjQnFlEPP8hBFu/0ItUh52HfoIHIcHJPwRHz+arkW8sCN
ZBiY9i9HxTMx+EoOb6dNRzJfYg5tNz1AxbWFUUcBgBALrJQL2kuVH57m1lmUCH88p0t+qqlZB9U5
XGL8jKPloNepYCUbgS8Y3+wR4TgBG2mewNtLemAEyrj1yMg09wrx4EawEgOS71vI2wpyhxi1AFPl
IrG9C57wrZXok4YzOjEP0cAAKwwNSJ6LwhfAfZRdQVC8qcV0C+F0suzXEVvwqo+Na+3UFPQ3jkV5
10rvZc+x1DOjNK1KA7takxhxQV7yPmg0T/jsEAQGv+2WuqDPJupcmq7EccyQs4JRhL04NRAs3OGv
/fpgLJKXqgzG5EZPGAsWT8xFMeg4BrzHdYMLrqMtjk5bII7CqG0Q+9C4bM/+Nu5fF0hlSMlzqlKq
cgj6cbpv1H5p3naVK7UQaPG7fTDyG/dnzZ5W9EKmruTPcRwT9L25Axd9RLBDheqJiu5YlewYf2xg
7Y9quGUBE/+uLlCZ9WBooMQcq45uHqgjXDldHxOsM9pjY8f1BOKcj3XSnjf0ZL21CaezUxC6eKK8
lBgf0qPSQImOnxU+sZPRrUvSPOqcy3wy4OZmu82oDKqILt+WueWpfs8M/XWvJTY1Bxq6U9rCjYi7
MEwnt4FMHg8XunZB5Y2LkbsRw91FEwnyybQ1CanlaiD26jcJlFXvc8+IPBAyO5o1bVEaViIdVZ3K
V9qJW5Kj8shACQGWfivP2n2rvWtYhX1v3DgEEPq8VyIOoCVUnTyKUDdQE4MZUj85HN5W91lVK4Ii
Qxf26pSZ1buvkYIiXnpufn8+2QLQ6pfZ678gYUtRNt/zo31hLXrwfXa/qi+FwFSpUoi0vxV3QDHo
ds8Bo3TT9FJ4d4HZ+rDITaCVNSLlapumUkGEyeEtpBTNgGHyhkNIfmmmkKi0aAxcmx+DqrILoI85
76UrOEMPFdRPzHVZfo5S3QoMgOgQjrO1SzitOSAssWobwyeowh7XNr/vbRlfXJzx8ue+pqtXDjuT
c39/mx8BZ4y3xcL6cvuPvJ0YZ5t2Cdd9oDhUwrcUvScRTdjuQlkn+JRJFp1WR+VQOtKBAx40MPdb
CMFpIgCZSV393zK427MpiVjylA6hdrBSmniTIh5E186uXkM9rd0fbZOX8nCtQC1ES0efVBfrSnQO
0ivYTI3Ow16caH6B5vRjh4N+a3W9Bo/W1JgVuJcmcRiEt+vO+LP0YBda6tSlyJTZ4+JuXm4vEMzg
SRk2d/IdBOgo1Sl0zkvXffoxOlvC00TEBCXpXS5RzSNrlnzYk5Oo36TL2zDlRKHQklox8ClrQ76j
XSbqzOXqmoqxLT/8WZsHn8hwtCNUN58CTmvIvnLqKRvp8eBhN0SwhuwBUWBRUWtmzQ107CfnI+nF
YFv8dSUs23mgs4avhHRSQ7R2lbcYmWm7TROLXD9B9LyqlKvViVNgDPzPM0xhj14dPcK+r1G8rgx/
aeJVetvmcTdM/6cef5WYOXWewfl4iujDzqq1URj2ONQol1zeC+sqkrLM0FoxwXcJS3Q1uzJiH/dK
P0w4ToAJmH09bMv36nyr6HXCyaL/ylFIibrhvibleydDabPehuOglmjqhl+Uz3D/5tmeIwQow0fZ
KPBRbOAahwTJtxfAm5oE+bloNwewMHRc0dwb6cNy/q8ieFKAZ4KbmUFOpTb0Wkul81BSExr8CzlI
N+hw6s5ESuPJvkxZO+1bi3npXWx+RWpkw9mrxWs2CtKDJKTDB/OmZZuaOnL34JMuq4gY5EgS+b2/
p8jrybisXPbdaK1i0KBx/rgL+XDzEPbozSihcgJC5KCDV4tGz0OgLOw4r5gmKXaf9POrTkaiE20E
GpZYn7ujY/a6xO4AuF07kscjMlPOENDwI0rHFzs8RyPc0vB+S/DLU/4CUYQbJBA6EgXXYdkcQR2O
tl81GT/pVFIl2Yo3PEqkaNebgjTasdQkKmj7YtYpI/9w0ET2Ls2IlnSIA8h47l2xAXE46hAUfMtL
VDoqbNrMfoSINS75mWwZCSD0wjXde1Myt2qn2tEKV5IBw9cpkbvMUiPRfz+LBvk8g6jQvWOulxci
0IP7vQuqREquMzqkP3qoglAJxp+dKjWMRA1YZNbBSYwodGfOoH+nWc0xQD5/unx3wkoOz7hI+/jF
kpAUgCW/JAHxhD8iSXVvFqR+ojLg4qIBUzWpDe+cxsRuVJSSC1mZHra4X6e+q+L51dzPrc8IEh3m
FtcfJYy15nxxP6+62ARCJurDLK5i8LHeWbqNZR1GKq7a1DNJmhmHmUxW8aNwon8kolMuQKeYMb7y
SnUxWs4OkMAbMJpy4tccuDVSHll7OZ2niob7CRocZb/Awt6a5vWNsurufH0uYKVDaIdmcMts1tFV
QaYtzbr5MiTxcRXxhI5c3pUPnDUmAVEz5cC/NQy1Gfujtz0PA8pKUSZ42IV4ClMielPTIVinHQcZ
auazi1yt03SBYLu2TSYONS8o+vLcDuTmtJDQ9d6wyRLIkP57poCfweSI89p4l5uzUOFee7y02A5m
JkfB1N4ae7Y2GBPSmkdwzWC4Zc3zQq/uO+WTPIOUJqnoOySceOxTa+Z3wPpU1ZUOH535LRraHfba
16lxNMPt9+Wm3I/5vtMeEAWZD7iBbqy+T4T47OebSq4qFKik20E9r9DYqv0alVUXXj3ydgwSQFXn
oRl7f14QEeWCmTW34GsyqiJnTdRH3osAj+PZQy7qm5s7QuUHrHDS+9wK756/ibbpqb+oB+BtPjf0
8emGgbaKRwvCyo661SNK6BetKn8rz6umQkOFGBY+5OvgpDkeQDzD3DgNrpLPJ3yP8fo+ZWegTI/I
1bgjpJdmcx9XYLzZlW4mOgDnjHNqAiz/n0n+VYc+FPxJV/9JwtnDy1KiUAtVx5bs1Q1uhXmDPgsD
ZxWol0OziV+rK7szwNuqlgRUjlNL8ja2ji+QDAy2GKSsRKJvqSpYSmOSiZqpY0h8LrBn7DQ9T+W8
SFxr/lN8NnilUtGfvNloThpxbeqb54U9zHJGGxeSDzi8lEdWx/k/Rks4lcHEx5CJX82pvhUIdreb
GXEeuu/ywTWBsyHtlMffdaSi63Xm7zdqVnO1ymC8PDtEKeaJosSvalpkiK8f8pFVrqaNFXzxSo0A
/tB8PAfc1IKk75rAGnAEBGjTO3TUGPTNEtEOqcfqNY/Dc3kQyS8O7Iw5wKOcZN+ooEbBb6tlNcnR
himKfwy7Is/pVVaK9+tfxDed90LgFXmjpoSdNhzv9/2zH58oDdJScBzHIPLbd59+RqDq7f7SYWVi
Tmee0RzNXtS1jufXNYW6PIairgBXV7JuaxoH1A4OwmNTTpVaP0V9w+hf92zZf+Z/fOxG6OFsFmM9
cCNA0+pplEvjGhS2B9dGAonETA9mfMWoal+VKigQwENqPUoEDqIQUMnLvhMXttsgONU82/6CgpsY
UbmTy/cG111vTY8UUo+7ZUrb+zWq6vtHJ5aQrXujZrku0xCaWk2R2/XmJmniwzi0m23LDmQa3Svf
9w4Rm2WziTewagFXCyhynkYeZJ8z03UIih2g9kosL1qDiPCqLnf/Od8JK+yF0S/EkoN2inhcZuGI
E52F7rv+l/HXTj4zK4se9ZKJWnCViNCS7hy/9W6AfhZHKyUecFWUQVLFcHfcnwIETFPpphcNsgFy
CfSu3XJ155cKTdvclX+Nto0bFpMAoUnSiOUe0N6lJrbwkQVQxwEMAHh3vXnDwX5NhKDtTdT3WerS
KnW5hNCSSubzq1Xz7nOCiIwyJOL2/lGMxjGEBbOW5AJeQbIS8yWGsGQ8DAuSbbMUPPkZ3wJfuxym
YoKFDgRhXLCJdPHmGMz0Y1YHlZSV+rATRfyjbQnJXSXhIxbN0xnS6cY64ar/LCqEQ/X5crNvE6xm
08+jec8sLNjjSemgFPmS4p0hdvNSkDTPGUmLiDtTWSPb1T1FY2eTNe0JNhiMnYkqVCf/+abrkb0c
yystx0KZ7Dqpf31ilBQG+LGk5WRdwuOvJz9vwZQqkZvos3Kzt9hdTuXdc05RWrpGJlzvHziBI6cB
igUh9WywtZ+9N2Kh+F4nuX3NsNUnjfGKKMtQjZE29EgPHRblFkn7dFXYd6P5su5c56JO7McgCFbC
Nh/xLsBJoPp9O+Ytof7D1Ai4+BTGthlOwWwJbDbToWPnLXUX6mQJ+p8ClJ8f37scW/G6k7nYdU+k
UkRXWpyLb6/nEjm9ztGNsc2TjzytDDSN8uDFNmlZ2BdGkF7H4BYRAsP4A+pRa5eOW1pAFTULxLhZ
gFRtrHoa7wO5ySOy+Dl9ybxTqyyUnTwWPTfZV91w5DLHzPUEEou2CthZrFDg4t5VwQEz2PhHOha7
ebmCd4hKmJjNoAJfuVSuF/W8SQy/Al/HrboTy4PK5LXzRITBUPeuf6lq5ifj/XHKYCzf1E1+BgE4
9u3gBbQ4fTHp3KRwtMbskAHtZLRSO/l+DBFLMO6B8hqSr7gP/P4goPAhuHwDmw99Uz6PX/xPACpL
TbUihlOv6yOTtg2pvBzNwoK+sCzwWypGIz8wkGDer3l77T4C1Z+Hq6uL+JHPYMvfk5ApzeV7P8ph
bh/jOxlfT3z97QnOAnQ16Dx2DhP3S9DkVuVPVtyuiY5fIio1ZrNjiZeUkDSqZjH4+L0W9894uXWu
5SHXxrU35z+V2rMwmTcuTDEAp//EeHp2PL4lErMwWc3KamtUAsAUETLF4akqdqsgw/58z3xgY1RB
1epu3bijguF7Q518e78tu3mXSw4StKatHmlbdTmon546r5OgbfPXpNA9Lvx2WcbsJhmwFc0VIw1r
NfW9mhEUKE7XEbm3RInylDpRjCcDsrwTibbSxZ8j+d5DfcuDUR7bEccJYG/bjHn6gm6So7xAhLNW
R6NDg8jCNibRnM4VzKQA0KlnENq110FrNSiMmHQqKBUB+OGY+ibk+hjmeXYVVieJnuUqI3PLDo+v
tWpLd9g7SsOLAKx4FFWII6m76lD5utqFzopwg/kOek0BXuLzeHJ55uC1HHzxSgLb4irtF5ISDk/B
DQd5pA7dreOZaPUVI5gr/NFDOISgjcnj1tiN5NFz3fQrfQMEcZfmqoe/puOq7vaz7rSgWtzoPDh7
LBUksdo0xb6Vssf+t6mS8HNaVKxjUJWy4Zj1F1Glre49IGCKQ0+jyxXf33HV6W/8yofmko8SCnir
tAIMVojlKZAdUA1aDYniuO/ojMbr9lW8ZDXOF9BqoFQ0G6iBrWIa6LxqJz1SVCIYkcQx58XrgrLb
03jXa91G+EbrhV0qNZY/eElTP92Iwvl7Fj2n73zAR1YSM1UsdlT/JONHwlU4stpXxbaEZSyGFkgY
5Ggtk7jhpWRJTPJLs3eFRLJ+mWduKyx0G1YxUaJnJ9FI82XvVLqvkBI7+TdaqrGoO07IB63JLxC4
DyLphbRh1msgw5y5i0o2d9hB3aCQ1OxrcZjxP8Sl97XlkBcHoutVH9B3T5K2XNbODZRqnrUUlqyR
tXHIMHCPyyqkPvxqYPeeEttvlvZJ1Pp4d1sboIepvn4/sbP4ZRodfKjy6/Pe5tsVgM9s3yOiuOGH
AMIejHCcFPvEQFtbCyiaycNcABdShay5blkPTIAXZ5XMr+ZA0j8+ScfggDi/mL7PImjQ2syqmqwL
8m4Zf/fJnQlca7Yg5Sjj/veBGVslUfb0qZtQttD4fJddN0knxCqfxPW5dkAGtv1cIDqayVvVQROX
tVPgOvlAss3cDqVmg2g7B237PNAh3hMQ/UrxL2hXJY5lI2F9zMpwXHaI54wL48iRsEtiDfS6+mAY
OjoFsKXWESGrvyk2Cucasagvp2hLIPm3BTScIVP+zNltt/7g4sEnIFAK9diN/3r6/NiedYbAiWwi
7XQBexT3UG6TP7z07gz8T3+EMjDdh2OEoEzvpxoyIt2y7jUfDrLMzQH/WoObyk9u4pQHTh3KN9qX
DCHvTVh/Y7umbSoqhJsKSJmyUnYcVoyPRGm2rwN4lLenZfmEdQ8DrVNrWmIUN76J+tqBUI9CEX32
ufOcMFdfIWjAVSLq8I9YhGKAs49wFaWRMe3qPe+FNfVH8Xr4ExzrmSwija7MamB01FwqiKbydl/o
IbgNXld1eB8M7fWfYD5c3X+YNgXqQtGyIp2Qpp4c9Jdlr9UPLn3zVNBF0dt5Qxqc1gWYnkKpIQYO
0BCmY4mPQRAUnDGfGDYMUlBbKYWFd7Ov6Z2e4TfFu0aGRzBGSZVP5yqlb59UyB6aCT+yepNFc0l8
gP0m2xwSOSAz9xltkrElKeH1MXGCk7veFSIrCd7b6VFWS7Bd6PdiUNmgv+lwpZCEf9XYdyoihzws
l31Db3rKJovD8pRpNublp6hHvz8CajiaWQNYctEYxyNWPFry/P9qm+KWBQX0Iajbzf0ifvq4CaaV
fUONn+OzBzXR5Yp5DfkQm4h0AMXUOuWWr2BGhctupu9JgXxlo1L8TbPz0KpvaGBFvykwS+m6WCBs
pAX5qO/hu0JjXZrh4ctT6+ZcrzEZVu5/TqUHirghK4PVrOT1dd/Ejte7gKwV6nV7Z1twRHHEeK8I
L/Fq+8SCpWg6R+WeLzP3NRBKcL/1Z9XNRBrl5dODx0yWDNhXGI4PA++bJlXlNDUF0VPzBVAQxvvi
NPZSgfqGR9lTPtIiCVNNfsOjawgYo3DYitR4bgWDj9BMoFd9xsPhBQYjW5gnBfMnohgeH1OfeNb6
4X1ipY+IzaC4aWhI1O2E2Idj70b7BsWmQs7LWDKLmRLVvIR4Dcm29KagXMhBUhRTmizVV11r5oCj
XIhBAjIMPbEPOBWj9QNAki4tKoDujH+GAbXc+1v3qzSeklF4Om9pylM5pUaEJ6uoK3AR0Y7yq2fw
1wSj5yE4WRX0Yjhx/Om7tM7kQLcxDPstO22n/a/OtrzR1xQSxsiP+fFgGtwoVE9h6qXR0WJLwAsS
w1uMYw/ex2gnMqXU55eblGqbFjdGacvfmQLH5nX18NozKwOUgxdHivumpfqiBlQSY4DPlEXBXOlo
hAlipwsu4MrKup0O0l8v77bT60zq9tpiNlzDY0H33Vi2HvFSYDJfa0Omgrw/BTJsPNjGyPNeKFAm
MPDD4u14zwXTshDlWQdgTeJqSEiFoY6JIjN+Onl5ijXRUFqzWdLu+vVIkM9rNkS+gopFiStkXb8Y
F02VMjmkYK2xkBdeY83l1uvMKr6o4kj6VW56FpRceKsvMBRemjuQ7xWA5nZkhN3MR9umTYwZ/+am
eap7XV2SIakKsu6FuAb+upsKUCdb8sPVA51AeOdo9mk50P+ZZU+AFEH/ZuIWq29KZB0a4xvRQDcd
bDARDaIqq2AecFXI/SPPgIs4S9pm9Z1+uWApR6gA92xaQYd0yfimAovuRrEy7bEvpAnWPrZmfiOC
1xQeCkcVPL4DwmdQarvfhSpzxLzEL7qGDOiFa61yi6s0ZHbj3FjnYNDgmOzgWebAacZuM+vKOQwm
PyK3hFe0ZMfx1Y9oAfi6Y3XqFlF4lF/TmjBlAtXziuouy7r+043jqKXyp35ezIJNMRoqNzjrk/mz
ELkRGFrtUKfF/JyMHi+VORXQXaLTKTHdlkAi+OgOnnhMcxMNDrzBHXn/5tW/eAZXmO5O03Y9GLcr
k8nw4eMlzZLscPihDFeYJ3pSdgC5M4nednTB/Ud1mhs3gp+rEjPTFcnFkvVJ12hxM2qjbRunP6GD
fOqJin9ID855jjidyRYUuayf3vOkWRWzWPjcWDxpOK0dEHjEgBe7FyR9Ekcm3ZgDiSree77ADDv4
7qWZcoATC4axOFHON2/sY4u2sq3Xe8F4X5afe0bQSod86W07BxHjeKO+8j8/Cu8SrKArc7aIUq+p
rCkyhokEPztmFgg2rn2JhX8anEeOaEMOBS8xQi/MNpWb1bk4U3G+H77+NeQxEp5kbEdthkICqStG
Y59Z9vZdrHzeIUs/PGvL352Y1Drck7NQ4KsNvb9f2Hv79HisxfbAKCTEfUmxXa0W9DPW6/JwgI4O
ps2IBcpFbR08iXDkt30Pa/WT3nnShgUtyrNng39pHT1Ls4FJzRDzmaFK5w4wB5yyegu+ZGuC+JG3
HIxHHka/GCZmmJ2/7X63VY0Q3b41N5CXqE0/VbLS8kAZWsan90S8wsynHNApb2NYHM4W7YrtYpIc
0c4RMZAYQ0LsE08I1K9cg7fnDXNiNPyRV5//fGOmFDHYZHMWmnSb8GFkiJy+9FPvEk4M2u5rIrj3
7IpYqx+6McbyxU90/c2MU8mav56wwxzWuXQHTtBs6GV3QlqMCZmd8nvQ0nSAPIy4hhuxhMNZf6uE
SMmJapqdUotJZCmNoU1La6Ad+2SbvMCpiZ4Bzg11Uom7ts+ngQCDN3TTUrm1KbxOuDp1SKECKOQe
ZsHLr+pnBuqQexL83nH13KWd73m9Xcf1bPtM+CIR/ugzTv+dOhd8JVoBxFzstm42DP/j4EjDD9qN
YsNiCVkGfIuWqNhu92zuAFu2Y242AUXMp5z7XDJ0xxWn5X1vRFVHsaW8oef3AaHb2I3FcsvKM2GC
03PdoW21Y07Iu+A9AWojQ3aK6inlM/esIoGh8qsm0CKm8M8T/SLd9BnSwwCoVcpn0ar+12ESzR1B
ti9awFxNctyB7Trz4j6sbvn7Mq5sO6DjqdheyTPNCogNyolLWzTM927bptn9T31yK9kA1rPijmiN
Ae0bOZ/DBnbAleo58QP2nit8Vj/nhdRuRzz5Q7plNuB3oGOKu2CaUvtOaJgR9XiuBRY8boW7CrYU
fJqWN6JK0gAbtayMpojuRcaSeHSGyG12lMvDx+/EgYzQUxtSxyisuZHHVPhArpmwn8gwRRtjo+Ix
HmjRAbyE21ECKmhX2EyCyHqBdtaevr0moignUJQa+7fjLtMrKEEwZAnvxawRuRqfpbNO3aZxKqOh
jgZvcdZRDQt11YzC0oK7XvZKViyudzxqEewmjzHG62muhXdm7X51iyVVLZ4rzMgJWzUaRUCFtw1C
o61+wQgX6DapBLol6cHj0qENAA5xeMR7c9UHtGnbgWlbxLjuH67Cazkn5jFyJm/UgqQBvuXNB+ws
7SXikivhTj5LE/q5fTQOaMeh/9k0aoz4pSq+HIkj5cnQCSD8OkgH6JPlamligzc7XDduJHurLAKH
V92ZNzzF5x6wAtYjpaDtlUt3MubLJu4MYzoyTTnb7cyP/K0QpbCA+eHF4r21bzzVdR4J3viNa6GD
ERCnPozjtNsCm61HaCBGNYciQJS+RgkVv0Lu/CKtkdGnUR7Jb0oymUIM0z6kLhq895alKQsZB+2q
/mfWPL90wLvj53rcmuvPY2TpHKIBk736Q4kLAdsKRpizEnaDUp3yZZjpzkb0n/RudEUtS4xyotc6
rKkroJP7wOkiVMITZxKmW6BWt7kh7/pRs/FPf6PgXE+V+zIN28TK0vZMiQCIYleAx3G1wa45V60m
2verlonMeYdCMs0G+p50aWGj2Z82ybgOMPpf7+8u7b2yOfQc6V51N5SkyzL7DLq2cgTPjX2Hn3od
dZe1xyiS7w64uLfOEKyRJ+z45q7cXxdC2hMMHs9rLhI7/Ju4Uc2m5PMzKYlhSx8PMf0b1dSdhh9J
6hHbusivRrdrfQuqgky2bbN2wE+S9rVkdW9u5Z4mpBHdFYUlylMn5ZbOP/6D94xrv6oiK77Dq261
kspj+lTL38mfE2Uz856Bew/TMNB+njUkPgbOTemgg9BPHZSjjTw+fmpCcIpkb1IciCasZTZ6ve87
84jCOmd0QU8eTTp841Tfjh/3Lm0g89O0rD8ENLn2ph7/mPIePCvvwCccAfk3EYHSMo6bL8WAG0sb
SaBY6XiIrboMRF3XHuhwI5Jj3f9TkD4w/Y14Snlpm98YSfLCjNvkid3Xlna/mGbMIw2li7zhVe0D
n3chhNfHFwgNU+3P3oViQb45myrZDyIWdPsfXUhPJbJoZ1q4Zp7L01RreZrvQIh3ZHXdwemM3aCK
P3X7Ti4tEutEyVs9FsAeM6gPRZYZM255uQkTrjv5AnoV+ArVrVgGeaDlmUYys2Oub7Wqpa8YMWuh
oPXRb02E0FOVyWsNOYxMAMxzuRZFQhsG5gLQ0SzSKJlyDi5YtgORQt/v5vhwmJR8syyivujGw/Gi
re365h2J2JbB/6Vtgzojjp7Lo9SMyIarNkD/xVVCwkfhyDWl4vj1l5WoOfNFQwSBXSVmSlUrP1z1
by0dVSAE66WapklhKsPM9K2jlisFDJR1olbk5CxN/Y9t5I/NAQsVXNJ/cxHy82j49SMoJInX+AYD
b4VFBY6tzjyrFDllPqdC+pK6zoJ5UTdiRwFDMIhnzS2gHOoFIZH1tVUA7TB0Ep5Uxc0z7PFOZmg4
6JWBGi1Vjw7Z/QnJUSoq1A+LaeblPEt54huYmjy5seg9OA7gMnHUk9h3KmaF1umaD6aR5AUeidfQ
vMNqq8fbrnGDtEeVihBAd9E5KrnVtxa25GSvJbY46WslBOzk/Kvctkc3XdDciXUOVqtqfv6KR9Jk
BRyVGQJ+NGB3Au2Ao+n6r8kBx0SMG1AvlLwEWaeAiL41/P7XgL6UM07tJe9s1lyBRv2nyyLNUUEX
78lbWVtFIrB87JjMEwvpSsQ2tNtopcJtHadhKHK8HmeYAjREGI0nxVK5hyKJm/bET/rkqaKAgOs5
N0rbZH/ikLcm0BPDitSOFsjZZpLFsCw5T5AuIOhZCNylglEbsOGIcM8/qBgmTMol793MVv8X2hZp
eycCdYC56k3uGyAMlPcn50sFMzf8yFXYkdat8s/mFumjLJj5KwcGXZd/JkDn8X0RaQeM+qbzZnvQ
OFF5YjeK5i+EdWAADJwv8qgnRXSpV28hhpuM9FANAx656MAEBQ1kpkfg+d7mbw3R+8I+8CQMOSMH
ddNlxqcotesA/huhyPp5lmm2qTEZgyddWnDnr3ubk7Cga7yCiVFzTaX+h2qP81dhkWBhARsYfmAK
BS2TVCeIvPpCCILBxylJ+/eQAJQpcdPGG6v7pLQU9E5VgSipYoQxWIwcV5EPTvZHfzhhV4tbF9/U
dfCPp4h5WAG1mWQJxijkZTxjUW841CM2Anw6SHb4hm/q6YY650IczOD7YrHdOvjRxUj/TbtVoR1b
VSKC48Z1UaSExZENbZLtCfiW1MK5Yg9+XewnU+l7SgrOwdGM/67/psJNKTuVOpsdeLycWkE4nfFn
d8mJFcjl3ZsxHLnIQs4/5gdSaw+Z/YJjhdc8AH/cSmeHnwdLvmLr3cNLHElxASZfTOA80cWmZRVG
2Y3mNGa1UMpyLJ4jRoI5GzO2CrX+OIgC0kWK+lyTgsSFEXOOitRij8JxLKw0Gn+5kNI/K0V9D/Br
9pJfnrv0xPMTXoLiIURTxCQMj6FrNIAvuTfrnUWf6n9LYX0k+g9kGUKcrvb/XekRGmiwt1qr8xs2
cMuol2Wk+3rqx0oDf707mbh290xPYoieOYPkAzlnRhn3dPq12a+F++KK8QkF2WVEpiP2vW7EcNE1
0HIahCCol632KM1tQri61fgOJUud+8z/boB9Q7AnCKyy7S4R2A/oBGYvNTb9QHxcYOQDGApcTRSE
ihq6uoPxAMI26AJ9O/QlnMOzIquLBaT/h1xlS6ziKINJCagGaz7eaY8RdK9PhyvsKM9Hsps8gCNo
78FZIb+6o9E+HaHdKaVXW8AasqYntEz2Pn6jfX6UGBLx26HykRcx40ePd/jJCuNrGl23G9I9QMTb
25Sk2mZ11vCUIQWAEkva7DU2b+NP+u9VWpxz5fGASgoHAwRMWvt+uGU7qn/S0zEI23DFkOD7A1ss
jOga89PMCvo3feV+Htba1flE0VpbWEZ/snvEQo3INsW/6t4CIQVCZapxHDiypjfUN9wmycLD8bmM
cZR3kTImyMhMgyq1YJNkFNhitcQeTDzA5WRbmFMljWpW7ZCTg8aMRZ57oWWOXeJ8eTxPYvoHzpFT
udIJ2Qb/RTBxTz6PYnxURMQGeg3AN1wnHbvB7+CHkKRG3BtjXVvhVpe/Uf2MHzHQftnJsl/3hIbL
BLfEYoHe9K2lN3dJL3dpWrIT5PCWBtK8gjOXrv5JBndqWTb6btIDkhKP+iEiwECyOk/oG13gmSOB
HFkqj6IS8p1uKIuqJ3BrKTEcW+8pExFXCLlzRcQUhUqFirttxQcVFgum+39SJndUPiOtpGQaRilc
zDzTV6PEUQcpZG+rKkTJFVe43MTSlAhEEzuuCnXe1XaLYo9fSc71GAJjtsjcco1PJFMBqgu1ev1S
5nWKh7ZduxYAbrpnv4sN/KboBci1asW0UIO6nEjBS5/Clru8Ps5gdqPo4ZWx9rYL1OC4QkjpURXD
Kg+/XvAzKDIzxstBdLzSgAC7r612nNAfUg3mCCmVLgLyCxJsbGomjnIIzQlQ4/UcZZz0FApTgnh9
8mc6R9w+HxyzYf9PKDHXsMyYV4DHfc9RzSYVQ0ubYMwZ2Jd29DJxrpFwenD1SEU+OrSjng3/LQIs
rm4+RrUjDu0q0tjXyWLERfWAeKXmZSPNJrzvadRgX20SrdU8JdpWtZyEXpB0V901uJ28zCT/4cJx
pSBX0FH8OfpYHTjLZOhFwhAsQKr3mI7Es04RxWy/a3uYo7/HMxBlMJW9ed6q2fsuKmH3O274KcFl
FcuCrXT46V22L37SnUv0kxkSorRNbmFA8dnXFWpbQwaMfhw1mN+4nAggG+tFs75SeKzm1WTc9wjh
UZksgPftibjkCUyGgnwARq2OjFq+ZHT1rPBVbBG+RPs4NmUkkPVYlZLNdfwL63gY8pVNgGBqnTjE
kq8raMpVFxb+K/4HOJ1vC1Hm+lNbPF2yFk95Jgk9C1Mg0LFwUcpjek8/hnfl2vIcGq84VvBt36t5
HGe8qPWc6WcvV3ktrMex0WU8VISJIbrd3uS09HwulGQVLsqRde76OM5EDFXt7f7UWn8AGyh09QWW
K09r6ecib7UPcTHu1NSbQ97bwSERS6x7N4tGqjAEPOgoHZFiE0maN4BArO52ibKENtu2wx6u8aP5
NOBoGfNiUC5UWI5HbwV87/KVgCuddY6nJ82lHu6rSQUDL9eIKZS3TBxErPooPQuQU+Br1r55mK37
JG7LRLLCvu+e3Q00+JLXcKSapNamj993++9Nh7sFaiT4p5vt/z6Y14B6/o/gu67R1u2/5fVcNEje
CH7RSVCkUw2flGJz1BDOWzCZtBg9x09lBxj45GM9yDZp+3pg0b4jup7zBaqnc4195a7dDvN+rA78
mKB5bQI7Vkw1RViZ44zZQkgSIt2Xd/7blJPh7nJuA/mFPj74sBTvTogBgIN8IHHMFe5nAbW2aJR/
+D2P9yoHOwbJAo2hCxZ2X977aEBL0BoqkmKaLiGVGnZxqkbRpNVYjRGJf3Vv5OVa6s3DCPeCjVou
VNho4LFidUMYHgilMPM+hAV+dhN6nFvrABbl+JbcbWXpJt6aefx49Qa6Qn0iy4pJH6Xo3LtI4y3O
7ah8Ee97Uont6fWHuoUmjYXaywFdKLUAkkz4/EAvDtHWpqbWnBGT7npO1OPBVLLTAZl/izpeuKIZ
IvMFNL5MNIg8reb0M0lF7C+u0OJPyWmmnOEo30rUv4wY4Zt6UxjHjN3hJTTTG9HONG/8pS3YDal4
Hq1lOfMOxe/03kItrqcJ3jAyG1mIrbto3fq6ILSD720JTnOyivX1lyBvc55ayYHKXE3SguTOQEZb
PJT/qFUhyc5YWNxtTx4lrL9v2z/1NNOm0F/7ChtJzBGTLHCw2V1MxHRQNONvZDPrsJob/e1bj/mJ
+QyZ4hF7H7ZBrl6WKRwC4NOBavOuhym7Lan6H/esoUK30qCKtpB+N+OhRWhqS+wjGamT1fguKVMz
lPbngdqoFJBKsBp19pJkboQ7rQU/AsqjHv6ng6L95EF5cDtLm3VF7T39dl6C4Xt3yAn1c4eY3SK4
xjEuHeF+tjgXlD2TFMMs7tfIRSNtFbshQKGJvnylZaglG2UHR9VbEB/nPhh2j6mTSBqUjUx0tD4c
v3mHAQ7CnsacDgw1LQLzSSCyJgMyDSYsIn9LOpsm+WitPNZ5BM65SKHtFUlr8Q1E3Fa9lOWtyhm4
ULRvGjU0qe73vO4AWYtqTNE1s2AG/cOM2sG81+HQvi/aP40cSZKndM7KiWv9cik5qBdQ0LtD5ynp
wzZ39UDFSoFgsQ/seOOk0BSwcZ2BO4YUC4SyMmAHbr1oh0S6ZmOHzAtddIBVSWMB1KgZcT06BPV3
GixW1ddZkHy+x2aLsj0sWbNzZvArzU6C4SyMkOJG2Rh85PSaSPG+2IAmq/mYYOeGKNEsBQY4vSxn
12v7ZicItxC6CUglTRcFr/4UpmY4WEXepxI2KNfwD+Q9w2mrq5Xw/zyOtL9MtvSlS1MogZRsOZ23
Iou96+lAA6UHnqNRp1iubWmEsT9Xyxy2jbN05s2rMRgBrHoFUwRqVjKKlSxIF7EcRoqa5nVnGQiI
v1wCOH9eGX0tObEpS9p3tgyQ8Oe+xe0QTLflmZQSBnQ5ubbDzTT88R/9XGfHsSNK/+RMhPGIKVri
c0nw4bjo5xd8MYIeCrKM+JKgsX2NjZ3MYZrFNwkp5LYak5KSolnsVtHTb3WbtPKNyzE0viUWJL6b
J7jmPX4NKDIIx3B7Vg9u+5MyzgZtiDJwH90HDCqJmMkR78eTLjYGefVjHfyUYAj03WIK2DhJVrwM
KHmsyatL1XFF76o1uN/s+btTViBGmPcANtZhcT56WyANlSPiEs3a9O+uKEwIwdovYu6ZwfJAwfUF
plcDRrDekPDrrEuJ3TCCoh1PMRzlX2zlNRn0btfMAo9Ir1BtRQF9/R3SPu4JyBp3xKRfeJIC2/R5
q7UnqgUJ8Qg2Aqbl8sE1xvYc8yrkWr44zH1g2tETAGm3ooO7his6zkQeiy/WIrIwuOgvS2YQOcy6
QuKHh/5q9MQtIImldW/ZFXrfx8XZEzUzPN6eDbKvSLsjT9XX5TV9XcgoJw5R6d0gmanAoTibVsvS
Wq5NaNVdI0Ujn83rlT33eUYiMPNkp3lrfwjFfZH2pu1iXfWTyPOcwJu/Bgy67oog9UTSGnvwMpdt
PrMxVzlyL1zK6nl01WK39ms3H1c9z4lwpIK0NLD+zRVueWuJqP3PFtK7I3UMBKisIoVvu+BDLP7w
4a2FDzxaQqZrj6N4M1f8tEPcHc0NBGO5VT8rxyel8zO3frYp5i+QZJtiuytFRJZtG3xjXeJyJZSz
e+5G1RtM5x9SwXIHugsH4tyKrvKI6EnRRH7Rlx9xjtQ4pIQ43jGTQYYz5ahn0lwhL3HCmXEysnn6
abD1WmgScpKL6MerzWXQgbHU4qkbLa6GWglWTi7W08hKfB/2oa87I2t4JrSfQACUc5MwIfrFInQS
GrRUv03l7tsNxZvv/SiRGwPaVwFjXjYP14E8FoH6XrAWwxqqQiOFuCrnZGWlVMpqZmKt0LiGsVeo
AKqW9aQLss4guwtuoWcoB+WhN/3nsHCvPpNvVrnkcVnRGTZAxElUkgy4AdjyZbs6Cqlc4iwsgTx8
vhcNwdnRyaQJZLz5coxZdCClV2HpXT7+0nqKUA0i+vl0EZd9oYntQQ3BG3tH1/Lz3wxWf5naZ1if
1hZxDdxP5cO2rE9El4E/nZwwJ5wb6AvVRinvd/KOow9d6Ls+BhVCApV36ku07Yip5iWg41qsBhzd
X0BuqWD3FmUtK74NU3kyuP9oPxPS2fNhKkNCnDDKDjt5iyP3If83FZD9ZVAPbcyIw8mXetYLk83w
GYM9aGT+SWkxljpivYJH3NQ/CR+O5ikFPQSlTuxa1/PP2gKPXipBAsNNGSaSju7LA6rMTvYx3dWg
W+9Fxuv46lttTZbYyakRaGnMrIj0WNGN5fPLGLknrBuGXEbQ/o/7DWYUuHY9BavL2Cb+tx4dl0cM
Y4Th3Sm99IYKlMgZHPtDryVpT09pjXbh+kuWZTEctvxwMtfVHfbOmb96IWhm96ebQe9rMnTuwYem
ZGTLVwaOI5mi4IsRmAL8TuuEmBPndg0TlhEmncFvTXfvn2HkwDExo3HbOgcUqzOuojoNFzbgZ22t
hW6C2KIg8lMf85pU4xAfnwP05c8OJKLfnNrdE2vBetvqnGukzJgBK74DAl3Aawty5N9pGP3ZYW0S
Mma43e3PU4NRTbRYgw2ggEklgbfT66PkIkxZrTEWBKOz1SvE/Iop9rQUt8AXDzkJiNmLoq+KJIrl
vqWUAQSh/JVlnzOqY58hyzbKEBg2U26oPXO+5TJTnHKmqDxUS98QhQhhBb5wZ5S3qiFJlUYROwoz
t7vDyBtf5bpr+rFWLcpmOOo4JPEu7TrNRTd/xzA5YxtShSwUhoCBUmNFBO5Hzecg2LWw6HpgAwVh
VYnwuck1aZn3lD+5IS8YxoMdceovpypu4E1osloTBcYRduEgP4tjr7YWdxmV3oe34rSvfYg5KOES
f3AeNGr5v5X9vWtXn16gSUoPGmWoCFLnprnkpirlL/kiVNJqT9bqOYCssa02OorXZeenpgF/irni
cLXSuoR+wAo+zLhaNmr4rggFqXPA0q+JsDukRD+NxpUEWK6ACd+qA8oKUqtRSxw5JhOYaPrXOLxG
FIZowVSLd07Maf0PGkJs267a+tr9toybkTmAHXI0DCqTlaLf/x6DfoFZ9IvRQFodYGuFXRsrB/8m
4cyJznZWjQ/9PFTAypvSPZ71ulTwuaxPjwKWqJqdDdKYwkvPcvJfMNY7TUX0qi0SyvMGJEac6uW1
R2R8WNov85Nwk9fxnDM4VssZekTh94g0asjq0P/3kYK28Xn1HiHzDBOyMay8kB8ksZs4fPMOSn6S
HR7R7lkJxUNLgrw2700nlZGMFYsxZ6/yqoVfNKQ9Dy2sWWgFA4yrbHft/oMA+z3rRVEHJ8jjCnd+
lbE82CGzV6CQF2iLA1DQDgj0Ld8mWNXjIjthg5YgVIpbX2zflChR1Kf9jxXwLdtxZY9wAHsyRxsE
3WniyrBiMmoJL2PcXpiVH87mItjA5sNT3b9cM04MqtGtYKn6UT5cwJ1r4vNJsucXQI5xt/nqFy/E
k4xoqRvZSK73M9aXyJY1aIp4tJGXby3EiSazbeXsM4s+iizBeqsHn/QS4530Q0Dkga6MkJVKffrE
2qg+7hN3Vz8azKiqJQ9CTPVh00f/eMZoQIHfzsgOxnxuF7gspXMAZJCqwhv9Kx8tdS+/fBTMV7l2
mWbRJt3hhlb3KENSccSK6l3uO1/c+gN7Muam960p3nCVecH+tcPk63aQFHlBI+zoQpTp1/aOhLvS
krihhTdw3ohykubUndj67AJi0CweJxoClRvDuD7kT0CVQBtnOy3nCztVAvDajxYmQlvD2diy5Pun
cYdfLcmpGDFxXA8g5i3003r9barJ7Cmq6jw/VuWLlvXiTn3WCt+lP+y5ccrqwiW8NWb86XZ7ga5b
O1n2/2d2z3AgIA0xGyC9YDcoi6dBSwUxmb7MVO8ExylVxfnEdBSANwoIBv+O+njMFqfj23gVLaB+
rLXMYtZ48Rpm9LenVsYq/8nvMjBXZF7NEuiFbpjl8J6Vnif42Q6SLEiOBQbaZq3ui9nPEqILrBeV
tJOyNSZmTmNFO0TDSPsFU5bn7SaLGMa5gyG3/OLsxTI8lvEhGrDjKf7Rq84rxQMayxs9PUKYC0Yu
7cL7gL9VpzOu9nmldnKDWWi2CnjbfSRj7+4FJD7gzv6C6FSQjcDe+nP+Pe2H3C61AUBSKHf/h5l6
kwh7tvtJIvzGNbIQnhLdd+vyOSzucf1uPPj8fucxFS9lnsgJcCxoBTv/kKO2GOliE8bwo31tmWOS
CMcRsP9cx/kGWGJnQlhW3zClbBcdNsgLJbh01ENJfgqrPobN7l7bA4suoB6PBz7wpj8vXKQlNiwK
2guq2igxr13nModmeRcd75z35BJ1biLWAYYtmSIwxc561boQSJ+m838eW/xMeNRTyF2Vv228Hdqb
7x8MC/k7zrsvI0Z+sKyflGGtrXWR/lWhfO9TQlfWeqVhcfOPF08lTTPS7GefC1EbsaMLSvnqbNS9
I+lc7RbMavk2RI2riCFENjApdNzGddCdfSbUpMWlzAsaMLGiXpYsPVdRmpWCulGyUFnUmGFCq55C
G6sARCKVvU+DVE+j/UKHA14xLeVOtjra+F56r+rWKFAql/aw7zgRCIgxSsiYYKo4ia1kElXy6ihq
JtkNxxPmR+QQ9Joqeo4Iw/Jpplb8LVY2dA3L3hNq9EfBnDuYpatyrG+7PyrUmZnpWbpHVMP7OFoO
8IxV87TWrHr1asl/ZXOfD6RAOCiGb7UmDrYMA+8G5QZhihUL78s+lmMU/y1aGOg9k89g4XMJKi3H
o/hP6Ihp9XVuSFaAWVZioxbcF1rX1ptXXIHzVgR6Xo8+SeLnDrINCvRbJFRLTovKeRYk6StLuGY+
sfMbW99k5kg6yGviZBxifDsiafkPeXfPP+4xTlySNOzaC5r3DSLfn+uq/eZmWTGcFDRAbdKRggCg
UoWwwGP42+CeaHhBcel4aTLXsWPhta3eA6pWwrCPEcVmsAwcWSbrh6fHVxwBXKgAzOfPgcx3JQ15
F7PIW6U6twA0ZMw2H/0GcPt3tnHFRFuQ+DRuB6IR5kB0Rw3tSfOL6cHLANUpSl5Rj7NY89W7Q6HH
bov4bP33/eg4DTE/fsk+fDXaCQ3210e0w3MQAitQYwBg+2O3XsIVrVlEzz8Q4dhPUTGXEZ+GNOv0
ctF6XAKMwwgEnCErVE4a2egkgIs3AzEuvtgtgA0kgirkNaQiIDPZRAzEHYT/obMxWWWnDSmp/fdn
FwV3WekgdxjgWRpZzZmYBfAv1jRbxNRLaR3VHfozxXaqwY+rnoPT6LLz/VfgAixDW81PG4rZ04io
K1UksZAOvI0z/c61P2tbRbGREP8gSFbDqpd7zEXEbvDp20ch8nULtOeCL4lA/EygBgIpXVp9khWk
2uslVf/el8Tkz79V4+tE2XpsSc40PnLQK+nOfVCBvjLv/vdMP3IFIc/lMmHW0kE9hTLUCFcNCXJD
c6zHcIv9ku++6YJB7WkMDrIAg7sJFaHOa9TbhjiIytUeyUNxGfIoLDS1ZqmsPhcitfSTGhcYfWom
kOltnu8Bx6al6pz4/fnMlPvJDa7r89SwwOhxJoQVV5csSxk8DPDp6pw8M8MOafgDiBAAqUrUqhZg
2NFIcd7BZxRTHAJ0bSi8fvVat24jS//c1XMXOPCsxy0dNbMuidR2xm5VZjeSYw4AwaDb/8rIq+Sz
ZyqU+/q84//UXKSlTBjw8A+U314TypmITtLye6kr8TCf0TP8Bif8mI/r8u41IcdqVoQ9iYtsoH6J
yPJ/cMS7i0zVQ7Cm6xusGhHwtzK7Pu65h6QjS6CYrwfVrlIFbOGt3bT0Ko/cUVBoneTYo6WQzSZ4
8tzMG2xrQEaiVy+KbpducJoChxgxewjMYhvYrvpX7NNcJuz3Xr7xROZNEz3b6KxcGzrZejxD7wpc
chRd0giJmshq+mrYkdL4r4byWWvhQf+i43HnsnQHrydrXPBWCNeH+fzpoNOqrTy5N7xfSu8+vZla
V3z9KzF47VkacEaMKw3fqZfJAvOZMcMCbmXO+Lgr4Td3QdaFIEQ22C89Z6f3M+bVOm3boJ8gyOM3
wJlYdpOqnT/+3DB0sTN9CWVuQxFplenyxU0eZyub/dFzO+9T/eHcabS3+r4kj80pgWRKwisulpXl
4CPx+Hxm6xI8D7ZLjgFKiO3iGQV0eDoJNBMeJgaBbN3ap907oMICdcVqnHKPqCCb/t91bfR11GR8
QdegAZzho8DaO5SA/XCr0ICr89G7Mog9XaZ7DMZ705b/+qQXb8zoATgdq5lyXPn/B2zfvSBJIx36
PzRFo8XZJiseevzgrRiGSuDRJ3d6zHs3PpQWxW/RiEcE5QU0YtCcue1cJcMhik2JLesqEaRcox2F
/1HhKQleGqeuzApTnKUYHc569XlCFljIozDlOtNE/8E2t8CuBAUMvaSDSDvx6Djz1BCBJ5EOb8VG
8Zp6IftNrltA2CCvrYjeF08YgYYQMlcJvg3GzkZPyl7AKV1uKFPAcnG5FCoVvZ9gwFfNd12iue2W
K2TneXPcUHNsi2Y7V1ngMOrJuB/TNpCagZqt342VckhRjXePY+fJuLxYujOhYKNCEmSmxIqClnfD
hPDQdMqUs/JrCv+pllQStHqEVTvTbsVtIYoec+6CBPqRLUfSVOuf8rECrJCSk4WNXHxPqgDk078Y
5rBQUVWPyt2Zvj1BGfoBXAO2EwE3plEvLFq98RiUjbXes0EQfDDlkz17ltujJIvBou/uWO/oyLAu
MnXZemQIybjE9H4mTt8byRsgG+/tTX1l7OFvVSOfwDI7mIVyYlEXLZDEi6/mcE+as0gRa0iHTGY/
ljwO72N91biVPCU2ZmhYN+3aPl+oeUwNkODLPTPRMS3e2LIBPx/VmuehpOzgRa1RrKx4YPbOjOW1
nADPEPe6NjuLF3AM2h62YSl2hgj5EzOPASj56xGJrmsiJIOxxjRoL1i+HK45CbcjGHPFcJCQb331
WRhqEBkcKHb/yolqwnj6tObBkNW2Wi6keXOp2nnxKW/LlhpXIQN1uNnxFxHB2B7YcA2Ctip7ldeo
2RIO0mvs15vbr41vGl6jSGmOmh1+S27AXhEq3147yzg3g+vgcmYY0MKZmzVhAx/PE0BnLtGrhWs2
Fbkkm9NEa1/U04OnfHtbJjyng7bJgXv4L+c5TU71PANdAN2A62CE4xgxzKZNS2Y80GUfM3YaMc/P
huIbdu0KVpSEXFBJyzDE2TQMQlBotscsqxp5MIaBenIPwKpyrVVpW0mIVNejBUuNd0MGzoeuoevC
hpTi3gypCA92eaGy1dzrclk2prDClzxBuQECAmzQYGRVGLUoHqL/72aLpiOK6Ct10HGr6GSAI3Mc
7nx0/idrt/nVaaGDEcsat5LTX4BQNj4wGCVXJti5XEdOws29jb9Rtw9jI17CzTRLkSq3aCZW/xNM
AnqBgplONOjCUNzFqkha109bhPtLPawWNlucaywjyqe6SmXeRoWH2z9e26jHOMHFwGPfpckkmucr
6/Bu0JG35huQEAFcaU8jdFzgoSYcV6uLUn+lE4A4qWy09QWltEIfr1UqMR2PGW+2PrOhixMz3Bef
ypvivPGq7bPsb9MYRhfH/Z1CvlxWkcEfKHm58rT53Q74i3lB0JrumV1/LbKeJJSWudlwHLkFM2km
K1Ze/IFBB11m+rixceVMxqMfBH9ZAnTqnD82LIfokLCiqbjP8Klfx9Gk01Ma/UwpSoY2j4ZtvDSS
2O8T3bzOkV6UyTw5WwNuP4sbsWveG1NG92AH09aFmkA4QTKwY2+dM+uw9CZ9mbDcblCJ0sLmy0fe
gPSfEHCHjEMg+vAUBS5wA8k381b/RUZA6JhPWeiiaRJceUqn6m64Ej8Se8E0iZdVpsGhCP603X9E
ZksnEoLCrGWW6fH/DMpdhN5Ejut4tUTr3NbrMmQ7+GcFRHWqjo9C5J1eFZjSX8VlJUyHa6gSdxdS
wPpzEisVK+kr6qVWfLwvf2QvQMPpr+3yfwfpAMRsMNh2IznNomH5NcwFVslqDYnFq9d4vcRrWdTb
1YTnJoNJwvNuv5CanrGcYP6d+duRHBbMHVFUOBFzmQ9COz/1YqFxxGsene7APRnEoyD2JrEjVOZX
iaWRw9p2DdNf/B7HSlLDMtystp4EE+Y+iaahxMzse0B8lAPMWSRPzvclyobbTdoM813IGmHkqkBr
JygfmYCgC1r3BvUhwMo2UQYGzXQyeZ+mDoadY0LxA+/y7QBzl8Ywcn39AQNOPFJj9HAPHpJG1qrP
FLDQQk/ddM48DEW1wlwfNGZUoL719jiKUfsv4wl6oQ+3FP7Mq8tlOpdrpG04kI9Ul4PCTVikDawk
HWvndsilBrR+Th9y2ZoFuBT4PvdvEBuFFodC+xilo1ABQiCZIwxoKjbYE6eAGG0UzJp1GcbLhh4/
LrCVPIjwbWbA4E0ZC829c2vot4VIy5bL0EppTWWqSAo589v7SOrbTDJBgrFHLd59Ia+PTEOGG8lz
q/ZxduSx53tVu3FhVoiJJwZkqc7wl0nDWLVUBdIvOjvR1FkzHnjsHMJFDDRK2Z2IY1uog55yaKO/
qbYZQUt4MQg1SHJZLMlRTURM926c3Bv75vggJB6GVpn/uPPVoj77B10Yb2XoBUpGkrnB2nzQmZ/y
BenmZbnoZrIeBzIGuzvRedMxhL2NJd78ei4cY8QiiPgxQs+YB6LZzLLFdi1Bpf5pasuO3of2usHQ
LnfJu52Hq9C0OEFsBriwaZFP9YYC4bmAWD/ayhnYAdyE1yA9emaAcNYb3HEclk/T3I62A8T4+Qtt
eY5hvnxgXfV34H1DlCCSJYzteXsux08gx9rKrXkpfluiiD+x698smInmImbyKqG3SN9q8tqOyBVP
JLFl1pn4NyBdLtwqfQYlhTXKvh/tkmAEykqlCcM2pf8AuPtcpq+mnJgUa5WQbQomA64J0lkDtpwg
tgC+Etba2A6VFq8DQuQdpem5XnkMcNFB1MPOERepX/8WiydpgQi1XSLlcg+GOUFifoUVlx2BBvp8
7cebJMDbuKOYMHkHDes73GkW97iDDNjtHbxVMtxucJ+Ud4/mgLOoHSO3AVPpI6S8LMW9Bzk7ADJO
XMNqhJxzy3kkbG6bSXWBoZC8khaJGpy04jVzRjN6960HExkiG5sD8L/KaJT+onbVh8D+gpmVAZfh
S6TXKJq0wA3FMxff7PUrHLn4+5vCGU+JXEJ9OtA5EFlp/Qt11JOnE9Irw5IBKvj+8PBIJ2wP1VDj
TR0qiu99aU+UcjIhHJlLngkqKWeriC0bfqEO248vJwraeHtK/5G8wFx+XyqbTzpb20yL+VXQkTqk
XDxtI0y8zi0YgffZMaw/gCfLlC2pvW2W4z3aeE15j5Szgffky/v6n/2PTEvSDdEyPVk7nGjLl5FY
ndS7lqPQPthWL9tQ9C4BGFTxznIua1FtgPqv52RXw9TQ1onH/B+AkDAHTjX68akBUQyz7WvJHn1j
Sa7/MuREY8kta3wWr/pyQxFMIFsJawo5KCaUfRffy+NLtHMEFBVupLoDRgeTt7aK6YROSfnRp70D
WXHKSAcPr6TTGs56M5BCO0TyWj4PCtA5dDhuaxB0yT1ZhJdANeRzktJ2+Z3t7WdfaJ0XHSpxww4W
TUus5CbfGpmeeSzyXanUsBTvL7XXYuN3wzYgFmgaveZlyIUbIFVYYZDug9V7NGvlCg1FYXmJx12h
3wD2DZ55qE+rCgN0miawIobbQ9SYisPTtCHnTa5WbM94DsJz2MidbsAPsdDPOYCYiQMtEuPcykgO
ByteSk54r6pp5RA+CL+uphMkvqhveqChMzCWv95eZslA6NCMJUIhOtf5kYC/QsL/tffkaqtZRHsc
uoODv/7OrO8uPezm4stLi0wGuas42ukY5tNZhj4c9SEKGzyww6iE2nfxLATM737J9R6jipETPjsT
24JzI4mBqaVF8ZC3FX7IuBPnDR2b1aEErkRnQmFRLkMi+ciuwTtLK2EwJsrC6PkndbE4jRkLcsWe
L/uPKQpY2THNA37hu8bqnqfGU3sx1vHpwVxDYIgoTwd3RxrdEl7Te99/Wxvyq3X2FxnocGnAJJYV
nLolaFhIDc4k8JxOpUI1q5xEU7QWOiqy/Jyk2PwIks/jSfX6Q/KV5s/FpPcPzxBaxFgBRDgph/4W
kXHfnUNqJ9Tyct8kZPCLxsy1kodore+p7iLe8xWNtSFZ8+IgYBgn68DNgyDK049oxu93cVAv8Ryv
ui8OXB+2WSo26JlhXhwjvc85FdxoCoVM1GhFfnRY/WRs1tmWynb+Om5tPeor2ify2CWXXGB4e+l9
m34/dM9qoBlC+kozCAYmdGM09cQ4jiV8XeAfjZF/1/2habTf6tOr3Mc6aTWHsR3BwF7VbnzZhU+L
K0cCAefGGw++Hr/OFDRRp6KX/D4EUCbcKARez8qJp4xpxjxCLOL3R40ThEyyym/W7LfyinAhrbMx
NKFfp7GY5GpwKOkLqzOb0mmwW+s2outwhOX6wHgFTGnJT9UZIpfAvuzc+K3E4G9N2CQSLTGxDlbt
OCQm7sW9RF5Ehkl3UglCTcmI9+6xYFBwxr5ntZvoDx77YuFv2jwCyJ+5TJ8JalmS31qwJz0ePMOT
0BEL//VvOz4TOtv4lary4DWOfX14AN3ON7WSdbXXVWajGCZ8WhXnwp6EtljT3vW6JfkYhAPpxPKl
vmReTii/XHuznsvle63GF4V+i5fxl8YnjVsG4xgPzNk+bvsTksbJVQsxAExomsFkzecf0Od0jkNE
BQOtLMGYrsP43AKSADiXxj1mD8XGVWho0341Fz2Oh3MO0b1uC/d+wbioUPbRHlVwKBcat95s/dCO
bvGUF3Albq+Uy6VTumpT9+DGFkguJRt1fG1G6WzyYVteHlpegipKwmAgisE3NG77f+SD70qftDz/
C6+TYjYFFDhu8BEELwqmkCMq9P5b7ogIZeaiOBUQtoL/61Ffas1CC5I92kk8KYRg0rSqzNRM76mG
fPJ6RFrOjBjRox5nL+WFjdt1+D68LPD8Jumj58XwtrBnkHQFAeh2na+QLQ9iMYv20RSIkCxIpYdT
04M4GnvRwR5/dbopmLiIjHRIm3O+mhn0vc6fds/jxT3jV0/L30n18XbzD/faF1ALAPmmHh689MOB
j84hgZsvJO7n2/8st4DTj7Bq3N0tpeyYRDkiCZjwIOIe7QsXX/PbWzypTuZPbUjJxeMQk5K0WaTZ
3lX6aoKe61PqmAXu5xaWZmn+GFtUlq4kJJMX9wyxfbogUdDKzeI/ND3zPPvJS0/oSrqAnzYqFVlf
r+f0pDMFCb9SL7n+jxMnTYDVOo7gtp34z6HrI/FUBp5CDBAhhGVikaTEyLknH9iKfrRqMkBDVDn5
lk2BrzyQ9bHmMjpi0RK89qCMxGXxouxZA8DczVII/JP/f9QchzP7U2nHaXqlMZpL9xsLvblRlMXG
69Wv9y9BFZ/lK3aJXi7YuBJOa75i50mNyU4qE1eyKxHOqlRdtraBu/v7M7RtnR7XMMnt4nQp9keo
obV0c0Ow/DB/WOjR1npszpFrM4UqY0Cse3gwIRsdY0vVuT7x8XVT31J9w2T4vx3DKPnnK/GP3Xv/
NcjChSdytOrrHZFiMwbYtVTKdBEjMK3MG3Dw9dj1SRwsc1LHpJfFNI2+qAGT5NPj/m7+YmMfIynX
j8l3Y5u2hJeH7DB8H4CVngP/lVG+By7Cf02pxkVMhvnOyOBP1PdKzpN69S1M9AXKPO8ffZeYVpLu
0KCszusbGenIsGWXkItVQ1R3WKKcc9M2HN0rHqEgUNViE7zpKCQAGCLaelHX7zkRCysIjTMNAnHH
pRzZKmABjW7AnB1WbgEi9dUShMTSvHFJ7Ic4aTuh9YEjGi0i2lbslOHY+VREu5PD95X4afjZLLuy
7jKJ0b4FzaXWVYiDW8RDqyDoGudXRtrJk5tW2c8pMzlIypU6EzcqKRiFMlQBETDg3GjB5WgvA+0v
RWMt+LnBeffbpa48ZKnHPHYnpSTE2FRjqa7n1PPuqj2SJ9THPCqm40UOD7z5U6LiXwsOjimpqcWS
4SUY5Qgfc8pTiRtGXDfrG2ObP/9tpZ0N6sMBjYdJBJ7xTVs1oRa5w7hpskmbRZ8+0C8CjVcIXlXL
Cr/ZoJDS22RpTPspLeYLls5Yd+0/irHY+SGZjYPPH65lpN5B42JUWxWubPjAyug2OhvHzLi3jxZg
QZptSpWwWT8bw2WlzB6Cs4dD+CwAy38BtqS3q2DvbGXhx+J6XjemlwaNlOs2ZOtWCI0sFiDBTRI0
jzZv3d7cbO3s+nhSnlkopPQH79VM+H76l8Y2l772VHQ2aJRnAiqhKm93l3BKAShGn9FZgJer8O1d
nqBHXvP9jP7LOoNfAF+x0mZWY1APYtEk3b8CjX3TvGK+SIA+jrYZsFgXNqgLmjEfIpxu9HXE4uIG
5YFSmEFR6gFfm+Z9znFFIsebztIHJv3VY98QAftDZ7GI2yF5AllJqEbHC1XWGNWkTn4rxkPTFd2S
v7r7DtHgb0imStw2Cf2Q6lEDsUr+A1CL3mOPFxKmx3l3DCe7MyfF/4+mZMc2y+rF3aR4U2w/OaHl
UhjdDjjldj75yW62EcJayGvpl/XTQAcq634y7qITLtPYSg3umMu+Jn/An/85zK34MRbX1nSQAwOs
JJC1ldmuhZD0IwlokuodN+8/LM6PM+wa451snBUuv5DJsHMIWyH8MKnUbdV6G90k52OdV17Pf0YX
cx6QC6YnoBgYdAfklF2+QGx+ZZf0u1Bo/rODmPeR/fks+gyKnCXDnd9p7j6sjWpmQW1Ovjw/2zz/
rfAOnxxd9rH5TV6eZB2jS331Punmcxrf2JJT82ndkUJpDmqbjfNnO4H0oY3Z+sGUSEVYEyP0kvCZ
PCFcxNckD1EOGjXJPGjGuqwLFYk5XqheYDEAshDTtt0LENH5O1ZmCeJRDFMK0nahTHD/zs4JnWLG
qZ5dJx4pQTNd31Osp1eFQELt1SLfaQOW9OPSX02LYvGn4CMFvHpdblUl8tyEjKY6wkaKxzgcF2vW
/vafpPjVeQ+wGs0akkobBGaQVONLJe9o7lI+IIwSHXg0cZQZ7v2i29loQRcuVc/GskPMe7Z5EWBT
QNoYzcHbwSx90XW9+5TuhLG0pH0Z1NQEG9wNnfiL1NUTHBVLvcShRZwnVCRZ6Zd9JIaXV1ugQoUJ
SwdO43TOzsjpE7PbTjww5gFZGVUxNJH9bxqemfsxJz0CbuA0UXFmwZqP+5Jl7wcWuyQ8RGc+qAF+
gUXE4dsNT9B0SMXznTk+xk1fX2O7qELkM5Hb7UDjwbjSloW2CzNGZDiZIbHwXoTiQA8okJyRkeJs
r7tsTFEw+MRpOpBdS1YFDlENEJav2F10n4qhnt+Vy5P0P5zMmPEncxV4zJCx8hEIzMfEpHoxbEau
01OLsRQFU7CCrFxEhzrUMQEvaNfRcqJrBI2egw8iFRAmsW/S3et46EEID7ejQSP8NjSs4KWZdJMn
apYGRukjl4gqxv03UFylGQJ0/2q0YGHwAA3V6uVud96g0WXGMrFHASPRsPQH2d8ziusYNqPuFH3w
vtAYm5ID54yYaoTrfEEbLik/qTLZKtKxsMxuK64FeBzyhedYzoUG9jjSNI97va9PpWKjwX7NzxOl
NDVdat9t0vsRTuFYh5C+UoWsq0mdc00KsE4omfLmZOHMIj76L/6xoGtbki0UeAgMqJLkBbHIw1Bj
Tkf0/8xUUFkYigzeDp55pfJRG8VN9vU6kHTT/WqFczSHHa5sQjEPGqbFtnN2p+eKBv1PQYrL/sYF
/cVQhWyBosU0GHohhXu13tyIJ/M3Klj1XcNdiHOtbYmIb3KqEVnVfb9EiRYMhN/CYbq9ux+/SCWv
+DeM+/8jZQtTPObEAvOHo/w0bf89mivhwJrTLGYyc1IE9qgbsMW+N0B1SkUg6dJYmP/MYSqhpHtf
7cchI/mCbkSjkwme1jxpAPeumxYzYmXx+L5Qu26w6vg/D6E7xgKnl9TooffTni4o6e/lzMsKlevt
uS9WEugERBuBOMkUp8f8Sktt/yQpw+YN3QDMbT0C6m074g38JyE6HGY02lQfpqyKt0Q9HCb4/0lT
oRLXJ+ocyjserEaCUmG9QRzGSCr/TvFDLyWXlwd7O2eHVfH/8E9/RE1vEbB1/v263/dGANYR1IQ7
/rf3624MmLRnxI1kaq/X0o7eBpSimk+g3O6xd4rkplQ//IgK7DjSjXdT+4TJYryXS5D/jTFBT4+X
UTsJ3tmW+g2Abm4n2hvik7QjiHcoLAMoMy1NhiphQ9khSZq4GshONAN03g6+dRP9Jet6U4nIMv2q
SSAz8ec1fc5VXg32Zdr+lXRWMCNhhTn76+CHO7ZI9fsz0nB4w7fgjqX6nfvjoPLAvLGSHP3O2MnM
GtFRil6d9ti+rg5hXavbDgeZxbco48eY9JG1EjVv7Y4q1V7U9W7nxsZtvvv2lnT83x6dhl+1FK4/
Rx0mhsW3wO/A5vrkaspE3r169bMJEn0bEU8KA5CPWuch6ASC4WVW/8rYqQLSS+lfJHkOMfF/7CAK
hRiBm9oeyV+n4gxSU6q4GpqbpBmN6MXIDeKPjx9vRAAuWRjQRYrI/4DADDdfCHai84P03HUViIiw
wbmJSfs2f4U7VZl4DwT4x8vSE6+Js/F+ZlvcifnZJToGWDO4oGCKVjf9jEH/VBGsjkcptqYmkOsn
eS5wxJjKh6KhX101r9nu7NCloVmW7fh2EhxeLESOmdZttgflou7JU1a+MBDr/f8sAZxk5KMVFptx
0x6FhnTNrY2bmDZXsc2UScDXgxpQ3z5vS1hBWgG/+kMbOVedwJQtsQY9TBYRvrcuDBVDs2ha5Yhx
C4AjqAwAdfwwpGvoUx5S2DD2wUMNQ+f+g/uadVEss+ww6oPtJSL3Ae2AZcy9EzLRgK9kTtjJkudy
lH3KDIxGmBdwxIzVtutXZG3pDxQFNpCeLF97AcmnOJ3gpUYoNdsw5k7J6Gsu/4iRj9QEdBRlNN2k
uznORw4mDHbbGKPlAwvbfjJKCcrzANiSLI7wWARHO/bKSKJSSd0XwxUd1XPJcycw6QntE/Y2LYmO
V7B+xID0sg5Pe6LGZnWQ8pafrHE6zN+z9I305GnkQoTHHxrc2wiCs4bzAU6pDG0gff0xTWWg2ZSK
QKnz2uQm5kFl+7TJVI/uwpS6mDn6RkbDgvYsCA2l6u3S9noY4B0QPPc3UR+7HNz3wJf6bvhljn/r
lCyf+v4Wrp00lPv7x1gpPM9iHUZvgS+ej0gKsPRQRPZp/7VJCxgBDO6fG+iuMiXYwDGhh7GVuLrl
TgGpEkcI8QkSr/dunADtfvvZUsmkyPsJlNdyflMB2moaeXWqz/hki628AURg0/cZUzH2b/pAW4jb
/bHRbPNX+o0a3KPK7ixh1GizPEXDmIS7gBTruS9MjZQbS4BpNM1E0SYmoiRzA8HYIAvu/PuICDTC
eebti3vvYFmdSlFtRpbQud0p1E0vUkjkVCinvzpiLW4RaxbaVMso1+SdrjNR0vHCwzy4NmuBja4i
hsiJVY8DUIKT2VEQLlNk6zv3iaBsNav/fsj05CR0ZI7mL6XilZ16QAlAzTEjNmx9sNoryQmdLhjU
7Q3o1m9CBE61soHpnHwzFvyT8k+PJ4/3nlTkaQvGo9Tj7DLGLO8yOeIkJ89BZXph45NeHmvM3u8h
dLJJgMF1UXe+McYzEAnxrq0p25oSgYWhfTrICLXupZsZZKadAB5LFNBmIx0mEf8f/+srVaq2ysCi
+aLuteB6vF47BlgRFnx4HxBRFAGRRSTV2hIoK2yQLAaJwcp9v4YKkV/1wJ+PVnLkK0RbXdhgY3yn
41xZLBjuYEHxZxCcNsTY796x+WcZNO3o7VK6nwHmadi9izHaFLAmzYruF1Yl7lnyei1eWtJwI4Sn
DgQydvQ8WcLq9rx8p2ZzkP1Ehtf6FIlfbKsV4mxslMSMfLx+znRnylZH8WuE20N+RZhRgunBc2ZK
yf0Wg6mJMbHn9r6nxn/hStMX6Ih/H1tXudqgMdOnxhJKS80AxF/wUd7szKs8OMphoMWRKYVOfsn9
XtkDi1vf9mlxiwW/V0f5BYJCql1aBHDGvoe2r/mIqSOVmHEoO4T2MiHFJsGmnDkCr6Z7ctqLxsho
oc7DQVhiM4YTB4ANOqyylWN73OhFt6MuAHTxlOkVQVSF8QiQ1Fh3tM4UNrqhr0GbIwhk2nPJOMsi
OSaQmpL7fJpoun1IZ7W/gCNTseQuYeXVI5T3FeFxuEbOtpCr71+t9N4csFW1dDZfGyohInfmxX1O
FB3kAbQiclQYk2Xk3ChEQP0hS1owNiS+yZxblnIrsWlMi1QwK9xc92yfnK2ag/jZgk3tklM4G+FO
qb6eA3VDNjb/oh+mqfODUuSePrQtsHH3kAgH3o3MH2udWl8VCvOt7iuZFvzCdwRCIia10SnrhTC9
xjhXFhzocIHaOCiUjV2c5JHrOKRvKQV/CstvWE0aNmobaoq8ynejwiA05ug5THzEWuy+poORq92y
9VeggIaTKHqDoxbtXsMiy5XcNkksTcP6dwn7JhcnTNkUdukTp47yySdIGbxcZztoAAozdRy6css0
SQQPebKTVBZPJ/ufpyNVA8Phb4g+sPxl8+2UOV/qBQ4QPxt4JATevK9Qb3SFb9UsuIBx+QdiE9Yd
3BoShdUfGvTjEOrtc2szY3IkN4xmlD9H840NT61ZZvycYffFhyTdYoeA2LyGRtHQTS6F5cLtXwRi
Xfj63ssOjCPVo8oT1BWmjYaV580vCyq6g4Jr7hnPwHdHIY3+nl9faH4O/gBdb9LQzVWVLDdpGpzr
xY+e1Kjb6X4FrI6lAss+2LMIcqv5CSEJSzU7LTmUc9c/Z0WH4ACcoUOc2v8DX3xycKCSflkV5S3d
XT7SGx8u8ioR/WAnvjP796PkH/Ost97rmah9GL2tcPxFtb2iQU4PBcy59MjrN2X4BKF8FNbmPV+N
VeDZ1azyQMSHw9EGu+VVWwtL7Bipx9H3IpaoHBDtRAeSDDn/uE17tWnuX4Bt3RZSbUZqGLrqRj99
TU6ua8Rmx+ZwUc+u+WA701fYiPzDBoTKqDdZdbCAK9HNiZq5kgeoninb8DR+Mf/Z1HjpIIsLSqH0
t82lnsVMV1mKWxwq0nU2sqsQkkwbAIlTxIf3ImRDe1bbhl2Cq97ARMOx1FwNlHE2O0nULUFYc1hs
ZZwZd8TuOoQsGCGjLk/dFTUAjMHcsX8EmFFEZBGTGXPglBPk/hfn205MLLBPblFWYlmkvlSaj8au
Y91Tyk3v6domo8FWnqEBtRje1zJgfakKkyMm+2QvSfcOx9AiLCEqYdDazqYZQSnrdmKqfq2ElJED
Q6ZPT8uiKe+nCui8fgSsYWX24Xc3fWvueYQVNBSEBwHENoBoQNmClVgFJ1DXaFpuDqUw4NMe/Bnw
HqW/nGSJeRqmE+XLM97hU7V6SVtNYX4/1tD1mE5GpnI8cCL6sqpVvT13Ow1DoW/BmnGQ7096WfHI
Ic6fUJRtSRjc8lhQ5aAjxsjalRTeGACjFRToE5iAD3ZUtGc5gAHUROlOEuVf0Jk9A9SZwAUFGSgN
cudS7vA3VBi1A2kXa8W5+QNoZx1eTlQZV+KuIFZeeIAPnBkuU1V5mlsEUlPnhkD/iu4235nvVU0M
JCpJyUVTSTkMmeza7ZSZwsQ1poyf7QZ8wqo1JOkqk5JBgUYVAbhpgnLyTUeQ1SjiHdH1HuNQ72on
cpa42WXj/x2aS7JJK/GmMfPiqrl2JvIQ48Z1qweL7kasZXzJ2VMfv2NLsa6SrMm9hBftizU/64xR
cuSRPy2zo5tQ0z5ycZM1Dqp+eEzgehEYRRqtfQuPU2yXGoYIcIjZS3p9DURCXwnERlue8ZsLF/PZ
MzL9xM6e8IQsLTlZSatFKrEMvNeYI+hhKrbOA8XlJwW22A26yHud291XPdCKXNqVBbaMyrqw1CX9
c/Klm65mrTKvSLg9BMoXJsfvi+D501ldSGP7VZC2hRYo+zlkxUaqQlCu5yTsoouUrCJ9Gge7O5tF
IOQSCGG0q1s6M+sWzmSkij3RB3Ypad7WFTLj/0Hl8PnMhlOwg/CCMrfhyHmPBUTnCmdXCA4Lr5C9
r6O6g8WWF0BXYx1W+Rh7cCvseMfxllzyNsBVs8MOT16odhX+AjdfrhNujltjakP63Mb7DsP8oN9H
TNiKQQeV4JohEIU+AB8uQnNKAyGe6Bu2v5K+mCFkG1UnYEK/vXj9PI+6VqEqoLw3S/zs/vvF1mws
TMS11sC1c7c4ILKHyH2+/B9M2lFnYK9aGcL0k6Gplc3GgZl0+P/cj0mWwC0MtHSq213dz/bHBS3o
puZ9XsLot3BL8NjT5nMVx3WKd+07WeRfFL6uyxYB1dME1kltCCjr1GKFbhYXtNzm0qCvFhBu76ga
d7PG7QcfiF4fJXG2GCKt2KXImJma0zLcGz8sRASxVYj+yfCNci/sqQM16BqEPXY6KixGGnadM8wc
bX648UoeCFITUwODI88jfTuVfdtj8vBuBhFIQzPC4dBSwu6dA72mT0oiUS42JcRYGWKWIwg43Go2
RplkE7ljoGqoVVxq7W/MiM01q/MK+NtBtWCeMiackMavaSH20gRY5Thj23v6hXwgcef9Z4G1Sf/F
pL8oAwxMpkVCZ1hY1GcfUTTnGemx+1DzfMNuD/IZ7kT8HmfNvxr/cHnCU71CTkOT3AZAM+QH9zeY
ZEkGVImwOeb5LwBWGpNzkp+knxIW/H9L0igNk+G0Z9YtyOOnUKY1uvJXieWAqM9Tg/cweFhy457B
OIc5+nG8uhpigziQqTzvLPBFOKTAp7q0+ZRiZrlDMwVn0Dmrm9qU2IzetdLT9bZj9fvhvYHepobA
gnk6qG/SPFelimx68NPlBzqe+klTXIymoNOcYY8/6dzkawv462n3+H+iQhVEiDzQ90K9TEj33tgq
ZO9sizEjpm5WPHqR3rfuU2/I9XEeDuLiGiQm07A1TTOva0DKvGyXYRizLMgQoRGt6zPnSI7a4spr
txCMqpK2GTrUkDklYy0KEcx+McfUhiLGu5bUbV1iQtQm+QgujFTX2Hco3/saD6UHZcrrIzH1GDX3
ZTcOWqmDovAz2j/XCfGKWJ02Lr9mtydxmVRSJIPnLuurWL5X/ladAIhHDuMbQBRRxdsDTa76ErIK
89rNJ3ZiRZQsDz/ZVmrHAaKC+0wgBekRSDJVV5guy54Zyoq5PvCfj7Ctl2iO91bNdysI7gdYqigZ
s7KNFj6tKg6ywPctL9wDhXY6Mc37y3Lz7Onbk9DWAiXVGaG1W5zhr+2v/1lzl5GirdZSgtTKHT0M
NmDnBjN/BsdDVSFlI50QileiXOgFdCDAX0am8lvGWhqKrhnc693tGIPfZx9wUAdrUoQrgDbalEeN
5PubYXY8fnwBUpGukC647QYLKHKgOIcGRf7cg+gLlWMrVT32Xb/R2DzvpKf8m1Gev/Of+j1MJNAf
WIYAJOeimDmpug7gJLxt3HJALZvcvizJwcgnexgxhyecYnpAmNvMvB89jJdAbVePtMo8lDkG6fhP
UoMwVCgqUoY+/bUe4eCDOxDjLs3QkJFLlVGzrmIqa6saghQUC0hVgrOUuLdw/OQpEwaLFUb9MHKE
1sr97N3bgTdXdIO66mtV3nvh5J310oQ+PLLgG0QoLC9+qZj5Acwd8hHRZLHFMUWVhcWt4pNdc8t+
lmuMZiodA5mKev+fFHLSLubbY++PI+m4+j8ndKjlHPzpXjOXVPNAO4HQRDoWtfYwtYxGj6n7SOhB
Da+cmQpcclsvB1ekPDSRVNr140VnoYCSvpCIFBUH+JmFEA90RBxguDRH7pWe+FZpFFiEQXFfUsFG
4at3NLNCP95rjMFIkGfRTHQuPn5NDd2yw/TYpq6iqFAcifFivzxeY+7w1qbtdjcNNak+4E+TMB3P
s1qG1E6vY3AGjG1xZuNWXobQyHF8AlCpbTL4Eqn7knY9BBf+XWgxPW97eCPXfE5rO1r+49arNjV0
LNvOc4U+3UiFkBZiGNUe6Ufa7LR2c1jo+wMDxTEPWxx8AvE2sz/AhhazQEZwvv/JnpGbqYdil1ha
AfWDIbVEh4uJI6HGW5UAgqJCY4Xz+04GnTGWXlYfcDbghDVQdNLvJhoVTx7lmMoUBpSI/NEEOeON
c5R1HOCzD4v3jIglBazSOltxOg/L6PGfeydDvq+yY8YJmDjbaUpibscT/pOpAp2q9io4Tojt7Uv1
xQLdbuRVhQWrv1rLPLsR0YQSB6ESi6s1yHA5sNKF8m4UlBNcM1dMBIIep2timrwrqMNmt+J5j5qJ
WyjQqNcyw5sKgsA3kUh01zO0RgIPehKN84M/827kx+J52raUS0mNjao6WPHRnk5bvt4/M/BZ8DLo
1vznq+HsQz09g8Po+tMwDrrKHWPAfQ5nmdf+9CtDB4bqjFXzj/UhxiGHUrCdRQKQxOGIN0c9d6vU
4Pnc6iNraH5O4qg0HNw+BgDZkUVdvbFcwIYC9mTAKOJ7i716egmu/IKwdqFoOKZSjoK32GvvgEWF
vyojrDAiNrrjMjozkTYUHBMWsf6cJw5mkIWELRBDATtVi0Wwi+8XyYol9xLyByFo25nMdcZNAllX
xQn0suNqtyVAMSRdOE/lDblyohOeygKqlfJ4Eea/Vjw4r1LfcsuWG+EmEp6LyzjcpW2f1sPfJ1+r
H7nhoDGd4/MNmSWRMn74zqdn16IrjJyybszon8Cpl2MQ7ys0eqGEbuMHEp5zf4mCo/8+ieWiUl47
xGzs/rWoWsDzmvP1huBN9Tov5NgyXO5zXyyqc+TvQwjm5YNqYrwpJmpUAV0Z75y0wl6svInau9uf
ZMjxH+NpHXrjLefJPlpQvGa0XSvhWTkapg/Xn3SH5CzNa99UHRVH4YhPg/Q+GhkJ+mFL7qYZoS9J
c2oTmwpxopZPyPNPOwA844/5S12jFkjALctMrHLe7L0OOkhGMKsF4+4upS0m/U/Cpdprey/D8/VK
EeYx86TPgQWBI2tbCDcnqVbnX+xqFnct3VDvppLyG//ZqHMrKlSoMSq9glpi1jitOs98K8esfabR
RWJVWcXsFiY12HSmD14Zm2ZpAp80tbY5YQZTSFK3ig+MSNJL3ixaguDyByxAdyf3Z4uzsLIyk21h
JQ3QJz617buYJSWBrE1hlwXVeU06jgBYkbJAVGv8nZZamNmmdKNw0YlyNtONfYQe/3BxZRX6ZbLR
evV+jXFrIVTMeqaRDP4g4226RkPgKkO7Gk4tUvKjKU9N4k6doArKj/ae6fxesVhah0eMjsdKJS07
uh1JAv+RPo9vx5kB5+LHYHZo3UmUhjn/hn8tM5HzBFskTwLpOKVgo/thddzLOG5zfGYInhq8lCYA
Ru722mLUY2L1GIRRVfVD13Fkszqc6bQt6gCpygbN7so/tTJsIxXb3FJ7E/K3Cs2bmKfOsNmHtZQ6
8P5WGQwCygFCVRUCCiNrA+CLE2E6jMwU25h6Ca3AADoOsDbt+uOXfP1jaE3XGvK2Totvv8Fg/ld0
ugKOhgIC28nkJJ/ciGK9TcBkgrg2WNOl2VWZRtPc694kf1EcS1yo7fln/mOx+EyyR82LHX4K+rlH
Mvd+wvcszWQB6UtF+4rzG88Y2nA3VGkuHe06F3h137rX7H0MEGnx7g2122M7q47at6GjBWGnRDvw
9Xlzpl+/sduO8KGkK8mTIqrqQswvWWOVfXTkgBOHXGynQMG2gSOEICZXQeNerqbFjuMLXYbJiPoq
87UwpIJmixZGWQdtx3lByxN1W35sy2hzbjiu98mOoVWL09w4YBxJxNkgvbmtsxVKCPPHJx6t37Na
YAYk7U8RB3vQum8NTE0FqqmjgTR1mYgwIt1jBWx/2ISe0/n5JjfAY2Wn+4JJeaAbbE0u0+PavqCS
1jgX9S5UPX0OnmlK84QvjHVOpB59O3vMGQOkoANg18MHJVifnl35vqzUGHB3T5tGmbEAh+v6N2Sb
mq1B3lYZPyceb8IU8ghbPAGJXy/dO8dMeUIge9F5RSIhB37/MK8XQH4SBANLKHj81LCnIALi5hQB
amHEoELuP2RqmOtVo9PqCtwSLputdvbJbOxiEw92wGSgyUtMhDnLOzlgjf8gX8E0HkhbdU8AryvM
MBDxiv3Abaslp1OIj94DfVImbBRoypvFlPzCtLHx7WBi54N5SnRbmKmLWy0TN5Je/qAy7OW+VkSC
3LTn0MOZ3QFL80OW0DYH/OXvkPZGVnpcLC+cowfZ+2PUMAwwmj31bw9FplSeEmK0CSuXFjCwbOXW
8pWexXT0lHVn7yGFxTfZ1r+e1BCaBcdDAdUG7v9d5EOAsuy5LIyxnBMwm+jvk1AFKwTw2HOiYmUH
kS8aiN6apD1KbyFDH97ShwnqwU7EcaBnLIn6W5aTE82HxBR+vKET6XVZcqhrD+OmVafFiQzkHC23
NwiFz4kH/dnKmeCzYe+0RvmbeXY7o3ZIjuWPOp17u/kWo40BAGWjuKCXCJ/D1bGtWOVGqL4weStC
JEMnWiUVIUGuLR6gtMdRhWIN2nbpfUbKijtgkR+XQPeBD866/FE/PBV7atBHh2MFxnUml2UMOG8s
xf1ckP7fHcCvQ4JD9QuJznXZfWz2J+B1JdALr/4IhWyo6adYDlyPKz80NS29Se3QBH2S3odEM3fP
33SYligieFujinN3Z8NubjhWi0g4XoNccGial6XPPUB4w/VcdHxmYXLHvDrI7KTdtohiE3tt7mrR
1BUJ85DkgMF477YfbHAT2DbkG5GvVRVapg1PQXb0Nh16sbB7tFGQMnM/hthEBOfTiVpU9yHcczB8
RU+yE1V/11BhWGmAWSLk/+uNmTWLaGiibVJLTGObiDyZ596aXvdWxzzQ+4wg7BWR1t81LLoas9cU
SrwHjzT1nTmw9boaVI79KwvjWeKzUobP8Rlm5Sb9OJYHfNREyxC9OuS/i3cG6VVLq/ZW/pXSPXX9
osizZfX9P2TNtawp2aVln1LKhk18e1iahWAdSxVZNYMQn9a5hfzWMDmuKTDE3yYAq+FWCb67H+Uk
iAsNwWl7TBoqy4KXfE3JfTED1aQiYf2GNEphg9Ij7oiPvMl3tjKEgyFh3fmziQGldVv5tFAnCbJx
3Lyl4zqCZEAjZIFrHNTiD5Rquanc1SbXVtbU6ZaXfKsSm9Dmgi58E7NAFFSqnqvnSvK7lHLfrMyg
J0kglbC89Fh08b6drAqR9E7LDjDSuQ7GTSaBWWRQsxuYyXTPUt23e4fdinOe2tlCSoafn1RKovzV
8nSuAJsLJThUEg41/GLSZOFWXVBd5vVGfWgQY9AyTxmuCu4+fUPJZ1eLcpP6H9mgAJPkxNj5fyMM
hGvIN1oXPGwIYLEQaSkZCFcZObmWx6t/DlNx069x3osLOZjKSVsXlDgiORyd6Lmgx7/i+ZeMyofk
DiPD0YybznW/Ksq5KNM53WjDmRNGZ7YmuYD8vrBmSOKICKPwfvWlW2fkseqbHPgwSC59HvhLAOSd
Tk3W+Efz3Xrr8FxGQlpLUmh4AxKreCavifupGFrbc3sntwanyDV65Hy+JJ6Bb0sVOdQXx92MmDKh
TzeM+JErdfEBmOedP4xGGe0eAM7hMuce3OApxcR8YeEExWNjkDsauGAvub4pNxQOZwti3Mu2LyEf
ztzvu5Ty0w8zmkoYsOpxBM4va5fxczqB7aLDfmL8FPj2248QTY4gVvSWbWLy9VvIWokIdd/pauBK
qAf9rVYIYwN+W0/8D5RYGosaHpd0mzdVnIuBAeWRkaVET4802L+AoE42c8e9oPoubbOV0s583I+z
ZKZB//2idybhq/BqD6jLWuuqBDkdJyn/3msNnMzNRaapeB6sPEdF4mLIT8wRQc55j5kFQ1dNxgpW
OCDlGq47HluiEK9VUkFXoyZjEgcX/1mBcHxNLFlG2kKMmK+RjmAqtgnE1P1ThYqezFNPRVI3K+YP
aUsSBCWCZ9klMhbk1ceKd9ClVq5k6T8hxZluEeoXhyPPkxLLTSgVmQEcXzjdn9m6ik6LqPvFfK7T
nFC+dNhGEGWfSGfacQg3mXmqa1yzaf5zKFBHztiNiw/H63+Bsf++BUPgFbfqb3ur8akWXia/M6A+
shgSktC0ZPHZoTBDQdxn2HJwpkD0ZgzvBjWdqQdyAqwD/UVmT8XJEA+N+F3LM2KZtbtvav5luOIP
Ni2PJaSHNON83PGR3e8Bwh5/p8Av3GEg5KB7/LqMdwODyyNN03HIG1cJGQqb74aR/my3WqX+WD2E
qQyku4bgscAiIVQZ/Og3i8QzhtiULlXz327axm5nIevNkNhThaQQ413HxXTesAtgFH7sTJ1NgFb3
1heOSzR43ZHTyg78+JX00yMKKoGtvHeNOgPtP/d1ws7Y5ptlbf5MVlZaujX7oqkD7jTw0o+ppQI/
WhL0xfKYsXB6ne0B1wgR1B0ncrUUmDqfq8T81zlv0a0D5B6CxBEGembxvg4ag1yR8G+PCVYV+87j
9uTwdj/3PHEEqJLIFu8f6uTodkd6M/ayTSGzUNhue1Bbb1lcFerSNnx1S+X1wb23YhjFmTRLw7+N
ydacYvPySg7WdY8ybKPZwW7udfufQiZBhanLJQBzrAwBt77Lj/ahOuBD++/m2DSJMqEDhB5ycS8u
PVlsEfs6zB9c/LxsKUwOwzkktk3xEBVSx3mCBgxvf9jm4hxhRGI95JxlvCQMd42+V4YwR/F1B/Ev
1lwJEpy1y3msRdbbHlhJ9ujb2LR6oRe0qzrIa0FWJrkVle0NrK7yNk0kVoyv+8pbRjp5A5xLyB34
d8HRWTUgRccAPPeR+oXjAv23YKm+g13hvFS2M4iN6u9tE9pF39zJeFUwmwW+0p6e+qKpwUKa9aJz
fap/Uac59/Y4WFIAwt/rKqr9h6sSu4FtXYlkGzrqBiHOopAIu6azFp4hwii5Pt2wJhhc3FwS+/PO
w/gr8BVartyVJvAkwlcpIYGPbdEq9ppRMt9nxwo5CYGGwQxCIEnuGu2wkDNl5OgNPnl7rt2YlzoZ
Pe+K3p/PZpMW5R+L1O3k5mFgb7bZABGzi9qcGc+Vhp/n5mJFEjy8WL5cGhEt0xUZypssWRtBcTKQ
9e0Q5KWrm9b5VjS8BrsMehRT+9xMF8UiV88vr+XOjA0eVFW/PjBrnCIOjTqcbLgpkAdsGO7tSgBI
A8Vw9yFp3wv6ZaF+dkP43xpl3JbNXvOD9NLl8mRck/TG/yS2ogU+BhL61+yFLVBcBTUl0v7i7KX+
ghq0uznSfOsXo96Zz7nfh8SFdBDpX7atv5GA2yEZ2A6K3EMSE8TQqIsbfVEYF8qRnHdyb6QzpGUG
eQHAIu7SBZtdRqBeCjvGblc6/5Hfs4AyA/dI5EcduWsvXGeIH/Bv2+nm01h+Y2m3raFFC/1t2/tM
fhWVn0PQchPNztookqyBUulOO/RQEI3ztWWvyZ2z6/Bz1tU3XDdz4rBCcPMn2Hz0DQC3HJWwwJD0
6/ErFhho7KhbEZoV+THknMxTI9lJPm1zemnox75muEcq2kuha3b1+ZwusE24/VruxuaKGO2cIL11
/h7avRRFfUamwAQLKo8ssnz8SPwWJadKIhINuA1somJUYA7k+iwFzS0U5Rmkp0pr3oLblx0j+fVX
gd3v5Jmkh/73HtKPPBby0dq2CHlkJWj4Ez5ohSUeS/Idhou9/cmgYjy0xSNjAeI4X0tc8icecnWi
QBK429Hjl7S99d5HeONb21i/0uf2ETDnH+LuidsCYzr985zruqSn/gWEyiOrGm2rNbpgaMFaM7FB
CD6HRO0aTSwZvmJfcutGUBVn4O7uwT2U9tOxtAqziyh72nHLGLdqo+ZjbXRkUNRkibpYrt2Elx8A
OD/4NHq/vXV/b3UVIKmj2SxqSt7MlmFFjYHPV0NGtxZU3vPYEV8X7zJ6S0QiYI9zoD0WE+bNWntj
nBTtGJAJ0+vFCBTapRu58f8pfVXsEDnpLbDkpDbCHLn2LwkhmYLsC2JIZ+4jy0dntQ/gCMjD430I
kG5F3IkokHRoaVBws/QF8QuZNe9V6IpZoPQtpQ5q+S57bkyVxxMluXaQt9UtDkklxZT0gBBxlaLc
0ThU5euaFdvHa4LC+m4ZwSeHYQkIpMWXw08CBLQEOSjPZfYiWgCQnGFAT5m6uf1y3Zemzta6AS+5
j6BfacQYtEC7EhVv2EM8D+PDa7L5ni6E3Qwe/J4cnyyYFob65zk+QhX8zVEKr0mF3MdyD5KLqFL8
MNpBkf98mPeBgTMo8Z3iAekzyh4ERYZzCyIlv/DIS4AJVk+vXHyGn1Lbj4CuHEUhq3FDz8HyXLOE
g+4BJjffwPr62yyqsqdp0WbzHI4eLAaPtN1inQEh0FDJkh1sfct5QG1OZiPZocz5HD0bHrLTzzjL
FuBHUmKRV5NanOH2KraLfsV7o2FvXRInzx456JE0snB8R9Nsu5YA0yWAmcyn3D56d8Il628Qko5A
Y+CXZmyevcQBLpYbctyt+nP1LipBzcYXWRHJSKu7nj37m/CPSQ6CLoqxhQlgiFnu24fhw8fhs3Bk
EcxggL77RXhTT66BDQHyglWD3YQKRIJIbd0An9erMrlnpX7dQKXrauXApHu3+YWihN66tUrvIPCq
HHVt6uCjle9PUDug4dFOQL8Vmnl7KKJ0+bNUcJ3P/sAO/F7XYc551iuw8Vk/bWOVdoqlBcbC56Gz
0mtBWu/90wSo1RZnZJQlNWxyXWO4vQpRX5c1uBsRHpzeyjzlBk4PQXsRLbusPD9k0na/1fV4OD2V
NRSXuYtk6mXgm9znAUQ5hP8Vj9IDsSaD7rYqh4+LnRklHKc3Fj3nSqcq/gbWADL6j7xxASOpSDH5
YXUIQrOnrXZo08U0/OGo8pIW7nYYrt8Ut+ggDRQyGRB8Wjb0Isn8hsQFMKjE6XQxgB6XyYjSnd9a
mXXKkntFCxIx7/6hsUre9c6U7j2iCav/U28wbJJ4yELWQIt5CoKSQV/eMARTjuLazpmdiGwPEDs9
Z/hI0gyu07v+QDTxhJ4IO3aX0Ihdm0swW6KGtMegIdp9x3bihPgJi26mmPervGlndxw1zCSvRocl
nIT/Y1mvhzOATIZRzXvhnmY55rf/Sqju/EirntFruQ1nfKpau+oEqtfQYZbFi1T8Vp4T1cKqIJQb
v17Gj+8VV3cqUVc0gdB/DCxanPOQzHHdo2yR88ylUtiR2U0kmytJ01FaoaDBSVVGfPU/K+3VZ6d0
8aDkD4GTwd+1G3uXRqx+OoGY2qJ9IpsGYF5y00mvTXfooq/pUIQkhH8IwDJcbgbsG5sGXnLflc16
SaWBWeJcw4L7VgX1GXqj4Nh72gBSMQKjwwvfkt1iHEOsA0NWauPBe8m226qOqTaffarMwEWTEArz
A2+sUseAKL+GtYEBAb/HN3VS6A/WudsYBaDFDRNQDLe0GKD7KO7NIx6VhO5s6w/d5b2emHIs5Hx5
XwlfnZ1roe+qLly2huhSZnDWYvYPOkBy41Ti7eoBhG7GLCYhI/qb3VfolNHxbyabslz1qjiWScie
CXQiy7SLSNPNQ/Ke8TeZoUMOoPDwHmKTPseHt9kBlw+BVnkfR0R7o6HvpZ6PN9+UKqrY3cYU2wEX
TgQMOQ6nCP1MPTpuZSD+SlHNMHKnL2Sd97Bb1iH6Zvskb/l5givnJzdnZ4k/Bsh+o9CKn/i8WXha
2FyjxrrTo6n+iBSLz1Qc0/RRhJwoaDld9Mo/R6xDFuI4HPcqwR7FJioj6LAEXQ/jMW5PjL1/S4Ah
UoHM/8NrHa1jK358teAAwLSrnSCdsixGE+jPJHE6x3xgxqkXjs1zBmZL3VsJfJg0xs+3zq3rR2Sf
rje9LQIbBoxH7BUpn6+4VhW1s4Opl4owz4FtN/27ARh/3n4ZfOffE1aH+DTI32AA+XfHKpz/POH9
AtpCMh5LDY6tsva4esgPyHpYxTrBf75lhWfya0eTeOXHlzrp/d3DIFFBIbogVEbuPYDuXvse5L6N
wGP37wy1x3dfIatePaUlVKVlTgnZMPElCT10tatC1aB1EBVH+nVbhhDUm0fM1SYIuA+ps0NrTuLQ
5CLAgPMGvC+momIH+oxANljHhdHbzFNmPLGBqHPHfJ3B34a88Z00LT6wvl3e2/I7O1o/G+QEXkbu
ngPF1ldNH1U2g7fOrfDT1721kqs1oS86/CovQS9y4v7cvT+klu1sBOYw8ijITjUt6BNawKQLvhZ3
GFjwiYSqu1jHy5KvThueVsVpyRIV6nCr6ExbMRaLih5qBCw4WC58PgEsLPhc0HpKRgZyQjm+iopM
QvI/Zl25kuZaMmjje7ZoRsF4xaIrtpUkPiUGMsXVdondf3X9OXgDMFW15bWYeaqlisCdLqWBvWed
yGQVGxDjo/OP4i32gXtPywhDB9c5EQ/64yhr/gZJGYB72Nko3H+GK6QNmAb/7lETwguL2itB5MJ9
G/Ygd33qY86usglHn/NTKqfeVlD15DfxG3mwTrgOT3CdDd4uy7Ops0GewxcsdP5b0eieYJNPlgt0
bRKK6MNXvVDuJYI7GNVzQoEi5swZrhlVK1vC4LavgJCrIeTUPvImbfAANKZKM4AAF8gY9q0XOeHr
G1qjJUoOFNL/4PkBP7wsx/cD3CygLnW6DQmbTsguOem+C6810mRGp4D6srbYsOvcZZUc0M4Ea2kr
pEVREMQMQ2P5DVcPaf8ShEY3pSSznWwqMJpWCxiL3Pk8t5oAoHlZYOFjBpN07+ZU63W9Usb3t8JW
SjCYNcTI/WazUiN02/F5FkStJvIiXeJ+CMytYY08AQQfR724KVtIN0K/RHgd7lljFLfVNV0IOXtb
BhtNYGaxu/ixTu84Aes3Er1wKbWsLviWSeXGflAVDqTGjV/VB7y1/7UQNGXgER30MdDtokwNHdho
hPdzJvK9BhyWXlnh+pQWQb0++C2hM887/3rfXIkK4MOOaon9DrydDwOcPlDwD1cl1+00qyHprjSa
GsBBu4gfw1MrR48mEX7kePv7ut2B0GS0dO/no0OacLvRJwWsN8klnk0aKkW7bFtbGzzdUhGIuSuE
HDkE5RmFCUWYY2clNofMCo9v7eRA4woHSBbLVLIjKm6FhI+9wg1/TbU135UbaVirguP8lsnj5uuR
dZ2JGN8X28yoVUGwIsfxS32rMpz2uu5a9N89Dym/a6UecF00ekcRPTxEqtYKzWZ1ZtW1ijED7C/D
6LI9LjtsYgOfQfk/3hCUbSg0lOonW0h5YlobAn+zBw0sEspLjL71k+cU+T7G8bIBaSoK9Ejg9b0M
3zqThrTOgb1s6zbHNhEENjvqJ74zU0Fm/Mso3epWJRGFYyLTSxjk+JVlpzE/xheSPNeM1y62qZt6
5pjlVm2peY1/5hQkD+dDiLlyRNb3zPxNgF7Eu2rqA0PGX4EMFECfg02Ep4w4rT4mfdL2/fgamD8W
qAJzSy8/nB67dSHqAxfTYEpWiK+hN7RQqLZiN5uWNZ75fJtMlf4jQ31spOQPN1YC9QHqivOTvpuY
ENtcupA9Q22wwOBmy1bO8NPtFj6LTEa9i8J6T7Uy9cTNp0JCD/9mB2XBR8ne6f1bQJNUNPpmbzIC
aeowVeeJifqMfyPkDGKvsDI6ELUQwCiWKcyQ8/mIbor/8SxlLuajdfzv9ppvT6bUhoyTHCR4On1s
D0v1zedo8NPoGUjZTU+WJGEjUR42Un39IGP5U9Dn4i1eF0hKgMqo+5o2CRgtAI0Y/3iiffs2DkT3
i7xDMM1K+9tkbY2rtt3M6q3/7ghcVfT+9kAIiru+bN8eBV0YzdpBtvL/AUuT2CpCA7qrag8R/97y
Q/gOkDljn0LB0SJ8z9EtWY+8vEawcYpftMQHgRRs8mnu4N0XJXAQJJt5Mm7oo2VxfxGKHG5qJSEP
y+zziMM2IGmf7LOFGG7iOPnulZvqVoMXaebaM5JP5KkAjbiRKG8ucR3eXJ4RFAd0k6F1fm4Ntjtv
9hZDtArijbEPvFzXw8wMyhLDVpJJ3YvERYT6HV8vLjw9flENe01LVHEwUool8Y7XcdtXF+3mc19t
DdM3jKHIqKM6axxmEA+xMTm8bl4CD4WCEE47jI0+RRovVkSDFvC9wgrZxSTcOB61QSDLKIFBDZ3z
dv1Wxwjj183XD+U2Yc1G8/gSiKVpM3OIzuCDAVNFVqFG7zpseq/SG0+Wgey6mDfrVtDk0uRynvEt
WsSXlWw4Go6g3MJTwewG94gl5isAC2Gco/y9LzyTKep3iGdS6D7x+loDsWIb39ccIgiJO+M7MqMD
pzxLq7ePta5dyU/vo41g8+eig8cM4peCCKCf0C3o9l+lrULOqUzmRY2b7MNDe6Oh1HuujxMN45R2
GbHzHtzhkQZ9EGVH449EPTDx8HCGy4LUmeZ226ojShI8wEG+GaM0/7K0DWSbj2p5bW/j1UUHRqnd
LzKFw12gX2Wk09X7WotZtG1bdyFGjRTQAAecjlBW2v+66UuQ+YFh6JdpcWBlWdWygwQLgE6zaeN1
xp/+ArfsEioE0sEziQIHfoe6a7lX11Fb34KA1VHdN0rV325TYMDO+pS8aw/g1gz7rvXYnHie/eQf
9FhWMmJiIxcrTknU/PMbc3jjcspmep59ezKl0nkvOdgcf5NjoO6O6CRtJqr8blA27fHArU/oupci
592+ebBiQj2kLhsBJ0A7O64I+vWbzONHo2hHaaJ9cm60OrNAcmHeqV7IjhD8n30Qv6jrqtFyld8K
/p0aaBpC3t3ROyj5PLiy+3XF0K3GHpknhgsNsGHeGF1kj+RmTVlR6GGjEGVvj/z0mLFVzNxRjUxK
FNyA3AAW+kiWNqrxkHA6Qi11I6SFBmi8qZQwjtk/z7K/5A3PmuGHz8T3zPbdZh88juxLebSDoj+C
3D7os9tV4SRYA5sKTh3Gc2H5BurgSlwtCS5Bif+SWzC677+VPR8PQEGwbXohBgLR3R/01o7GxxzJ
5M48KCjdzBPDXFeH7PItydeOkdtNWsGZ5gDf87d1q9WtogY8eYeKcHbDvfPzFICnVmnandlNuRxu
rE5KD+oMBKO4pa2T1UJTZZkQXJRnFygPisCJwxYn4OXqsfb7VySCyF/X/z+IJxKWkB4VoaotK889
WxmD5UbcTuOz0QMzxYuEYPcPHJcymf/HE335WoXVcsPzxldHg9hElySCV3T9BVws624oSyPEwLWy
WF24uJXRVmQdKVNBNT3ix8IyxVjQPkvfsFXYP1iAGjbyCc4DAYt/yZRd6R9WcbdJVbXj1wtRmonB
oQibvwPPh00AvaW/SYGnjjl7DWPr+FC7Ia2xY02tRBKPA5U3lfEZ+94mguGPatSqVGEUv23+ntme
UlqNCwWBGDbWNJyykve3ZLg94hWs+1iiw9JQFCAc6YolVXGaKjumy1V099sy15bc5ra018CMsUfb
sI2Nm+eDsH9RZNZmig0oKLFp22zb/3+L7Uh0K7FWfvy1QYzKtT3yDq5XHtBPmf+7GRjPKusTm1uk
5Ro28hhMenemZd8InNnSgfqdmD4Q7sz5j2eRjhAaBh2Pk5si7x3mTezUa/2lD6pO8WUk/exzuKFn
uTzoXn34WeYyNX0G6cewxB02U+/d58xU/Dxt0c76/Cy9k4bhhuQunjcTzk1MY8C594cXof8lwfAO
Agbvk2T2whD0D2W6Q0Dc9ZRaLRAzGrmyw5LI+gEjHATL7nMZ4wEDtvtsetBt9IXJPXhUuNMIQCjn
ntyurFy+V6RIBTY5ozLTcsH/aR4dqn7lmUJWJyJiv98TcCsyLjYQgC6R3jcY5lIFL++PwA9t5zd2
CRdG5FYYzDonWOVQSmhB1LxQqz+uqdbfxSphN1KG3gHSF584K+juXYcOa9ko4VUbNMIeGQbw1Omz
gcBha/B+zMCtAztX0X6Y+KtqO7FXcu1t047HvaKHPqExwGkGnl3vcQBKYuCFmzqTR/p3dDTTXgvm
Fw+pPvFcEUAQrU3iqeuy3VGcTTxPUjAgkCksGO4O5/1/ikdJjGuH18Q+p1Lkn4+w9aW6pquCJv5w
dRAt4rfmkWQs5kUgZN6m8Ik/M7CEJlJTHmn/qJWOWMe3+oqDeWDmfgsGLlNLUE1TWAArZiA3c9hr
Lt1aS2Ldx+jt/KWoF2ZoJg/I4qOLQjRYPVvCbdwZFk3jX4sCx1Io8zWV4OMPjpxIQ44MDqZop+rn
wpHQiAO6EPRhmr//5iqERGfAXd7E5oISLbCu4t5NqcEfGwbz17k2CUCFdH9oRY1rdzs8wsbHMmj1
RylBefhBl+WlUV04kB8W+qRWAs9mNGm86vXi6e/MDQQWPdt4ezopRIIVR8/5RBxXbRzechqz9Yx0
6unV0YEvk42QA3WaeGaKCRaP8qHO9Qi7zO3vb5N3jEa1FWZcfsMhARtfpBaxFQxlQoJHpj89j6fA
nqFt6U/eYxa7tzPKheggbLa6v/itCe/hxBT93jTovkGjVfGAx3o5hxUzdlR+Y41aYXLp/hDPyGZG
54sp20wbPQniNxA/1uHs57uy4ZemVAWCbMG3l0Opp+dEdf3gdLFaU/gh4y8/7XL+SgiG4eXk66L1
dNn83iwo97i0QBN0qR9Q8ydtOWt44uhsIQCkUmsjtVKaLS1Xk2OteJ3YVixgGTBrrMzth9+pqNTW
wTpqXPoL8Wt/aKaIOoNQR51Mv8SHROUEuKlVzbqK3xt0o7woJJqT4NpKEuydaIXlIuWexnYuJTS/
MKQUPZQcKmgDczqvkd09nksJhvDNpobkM/7PtzX+5AGYoewBTTfTRB97pEI5NDNcBwcutajh7aM5
SMBkTj5zx2+hgBN1pKpkWbCe3zxa/G8tz32vzVOn1iMI7xFffIJjXrX+bQ28QbhG4Kg10+eJTbw6
FqXq+XlV9H9jR2hCZz17/kiUo2E+6Y5FGPPpyycks8o35ywNS+2V6uXoQQF/3xmzjS5xfrfI6yTj
3G+sNfFfY/59AbBBbr8AOXscqQ29GjFkQ9D90XFbuO5mh/rizWQsvdmrA1N4GzsAIjSJ2pCeLTEa
xOvpH/ANHWnillnxkbFaaBBYtX01xkG/0EuUn+INziwV3a5sju6IfAOxRYzbO9tg+s9tboR4+sr5
ma5HFhy2ZeNUfCCiDzFCffd64tlbmsvBhijn02oqLTVyTAwd0+Lcyuo6X2YsxpLAZ34N5tfkGlfQ
uJpcVuLAeZ14CzWi5S361JceKSe1w3hfihrn6pe4mVe6SAHPJBUaYqrrz/i2z8EWrhj8dCNa26+N
vm6vMkMb+QenekXhWdVkzYq02+NTSEXAcRABZ6/2BksMG26nLJXI9HXdAB+VSugM6Nj9wPbbm8wd
SAIw8w5IJBecnaxg+wG20bE0zjOB5KaHxX8pzcqS0X9YoIXZZOrwyzXQ9bkmiB58UN7heWVp8/61
K3Xy1EzaRQB8le6LFnDOKe69RFvXdrNXTMiqAEx3epX3hTVXuLjUiKTtcOtE0W5ART+nwuzmEL7E
5eXEs0TeYHLM7teQGrvwQbF0DZZNFb6Bi2jnlHux7bBUTcCNdxjgmM6vngp1gXGEEfSrygHTR3h/
fKaY2IIAeC5oSaokZRzzGdQ/ghqet5PraRJF7WBPlDN9zXm+NfGd8IzGXnGTVGd2FBNr8SEuTgQr
Wt7Ph/hYTj/XvuSut0Wxqn1St5xYfGIocSO8ZpojZR86LjNkIC6CQ64XelPQqOn36uVcMvNyRTAk
Hsu9SwsCGmUKLKdeeC4ORPtRpmtwEfC/aQVKelLuAzpr3T7HPBcueOv8rzqVsfTkgd8zswxpVZTR
WBDeOStj/tN4izY0+0PqIpwtR+rX0KMCEaUPYPzrkngE/PJuGsoOUZSahFKc2gBa+Hxea2v0TGrv
gUrdZ8W51D8l5e1Aja5T7U93ibGnTWMSYASOPF1sp+akFevyeVX0QMzqsYgmMo5l4anxbHwn31Wf
UG0lRJIWeTXb8Vh+TgQSA/0rTejRV0a8+yvmO0M2ajpiibJI2MvWAyMBuWoXubiX7mGkGHXlR2wj
yyBxBZOlQbgoXalkURROOrEGOLqUcRvz4OVNi/pgVDIiq2KngpJPy//pooea+GMK8nIRbl5KRTlE
n+4uAtGWVMIz0TZllmrdtZYiWxSFr+hrNx911v1zS/bRBlKkmjA3V2zu2ofEXnkEl/JjJBJ5rj/k
IzfC4rpVNElyziVQy1/eGEiiLiQxHuCSlnsrRx7f2ik/zDH6qL9vXBejsW8D5EYg+v9vsQD/LOqM
22dMP+Z4ou/rOzS5Jf6ZZN8o8MfhciykgAfDk8+3Jq9y5EHNz2LXIEoDNpSHH5q8bOyeD8AZAe61
IA/0f4ReUlFWI5fmZYjmWA4EG6f1ZOj8KfIYqGm7Uc2tI2fsIqzQPpZectPp4lfNrj9XSaIoXwo0
Tlgc6BAsGaO1ytoEuESVFx3ooVIuet6HQ3WXREOehm/DSNXd22UkxGW4isbiYZHUIFDiQJO9pAu3
3voV+JJ7wbG98T6u/u1VVV0QvPvRKYSWHrHhYiN7vtPxjyfw2Gst5QKOlvCE4H/7tUiWxQMJ0XJc
yK1neB66NG5CR9ACBOVZ8Zxtyq/r8L77J/W2Gz1LWB5rJA9IHoQxJYAsfZm1mTGpJEjGwmLlsGTh
yURdGAplB3K9eKcXyhvZnPjimtZpC2HxYRIzUjPAD9ppKbuC7gIN5NdGpnAukZb9zYrSfCniLoEI
kavvD2H7Kbyq3LoFth8vIz7M8wI89Bxa36a3KvYIQkGWEBE43+fc+G4FRYZWHRC/FQwKqlH6nBpr
db1OYaEWk5gcrKMl19aO6UTsLRIa/Py2fYHMHDl7+bzS8XybRdED+jpEccVk5K+5hjqHKXxaOH0z
dg4HYwmvHv7DZIIZpoXjue1RYs1bEP7SuFmX/FSZiO6NrkT7HjLC/fvfHOaagQ/WHHjlQCO2DeW4
D26L9GUhuvMIX1zBIfIPFsSeebBdsppdj5ZIUPHrQtUCsuQBMEjd3RMuE4M93RnNE6AvqWyWdNRJ
+v0odDA06/88LKt9REcRhivIxos90YzpM3F9Fjd5VX/rZzKsP7AFmC/lxKi9kmCodbzJU8aoapr7
j94PiGTDtgVEIdgAc9dEGlSZUa2j8lxwmFD5UxVVL9y0rrTF1/FHT5ZnXYmVy8mGjCckAZQqd0CF
NRtZYC4XRzIjkEgsVoj+hrCBJFdPkLKBKsN+1I4NXEJxNijGSfpLwpc5ep8xVQSKySSRsjSd6LN1
Rt6de1ArgJGLXDmo55loJOjlOZ4SUsxfh8bZQypP4EWWR3q8WCoJe/ieaaUhQ3An8Yae8LAeBwG9
GFmh5cAQMK93g8JMu55cPPmPJt1HzPkjnEb7N1/U+DJ3CO03h0C5Qv6tISoefd3jooW/B4nFaK78
QS0ZQejSdElU5sDHW2Qu0mXYYoFHom87E6lcg6P5TqOj9ZaL9TvtqR/immSa6Y8+R/lwAn1hDIMF
P8kz2eP1HToL9nItLTRj6Od+6iyiIZv17RvD2BhppgYpYsuKMmvu4Eru/4BOQnp0888lDgyY0wnA
MqqApmsnOwKVfZYkcAC4211t6jSHJdmXF9SetT0NvE5/OObxus0tjBqqFH4z3l1D1G+FPusdEuSl
Jf/3+v7lOcjBwzcYRDPE8zo4FBAk1DovZfR0JiBTu8EYmKSNc6o6T7lKXhpAr/cr5zBHcgk8SoBf
yFga/7h+MCGcsjfIePgju8qPPhhFnaElbSu5UV80YYiGGeHRjapq/z/RaURxUmSmkvuHFu+Pflcl
YOwmPAERacUzgXW2O6NFJ/IynP77TKMA7+PWCgZk3tqUM8u2PSZ2iUWn/ql4JwIlkUusO619gW7K
OWzb4YP43V7fd1y6Zs0cDUr9DhtLpomVnfCqt6fsGEwAgQmsPQuHYxRCQY2P2zXvQBM9SrN/N8iA
i0mBWRbCuk7/bbc4wUt2bnO1EmygwUtzBSkQ/kwtxyii13Cs1fQEUkdu0q6iCi8B2os9+UFgLVye
QfAjtsslkbhvTVF4e2564KqO885e1K/wJr5rK49bM/d6Wu3/qHKu97XiRGhXRfva0ARX2I3MJp00
uyy/8dkamzNkG/rosWRETNxR5IHxgVnl7VY7xupaC1DkTPL22M1QrEweNJTZXXs3J8XCgHYOxso5
Z8tUXzTJ5r4GPKqvtdrypbIuFK2v1nMQ6DNnLXl0FSEcqkcyiFj1q+sY26OVFcpkII8oJS5QmGCv
fBeaBGIbkmkqNU2DfzVMl9hruzop+WvgJdCZU/kp8HXU2z3ZB9HefBp1HcN+ahF77bLnsoS8xzos
ZROj0YoGC9e3YBfd495DqBycKKeu46xyO4CzTXmQRoZ2ogXtkOWmdwb2evUJkqMyvCrjQa8t97e3
AnoXX/wFX0cxAiPeNrQMWnbFX55Xnos26gTXpNk8F4yml4M4apUdjb8uRIornXe9znXbgb6Ynnor
A5Stm+a3M0KnH72rH21qOvJ0uC/wJiTt1m87Wb4zHYvbbdvoZsa8UnDM+7Mxt7klux17U+fn/97a
7qv0Vr88mq4CT/J+SPUHiU8UGQFYt0v6t8sePDYddd8DFbXt+uWuUlhiopxrbrgQ+j8su2ogQV2+
mIDgKsGFl9uzBPohetbIhJ5LG0h7vWiw+QVF/Rz6n/N31uFLFYAu82IaXybPVS39NziKz/u4HdNp
ElIQvsamDaRpqRSrkpk5c65kLkDkjfS43eyYG0SGQC7u4vi37Zv+DEdoX59NAwbbaZfnyT2twq+3
yzgB4fbJGSnbOl6bhh+oIjPGAapUh/wOkNE1/hwVbP60fxym8c9nw07hnkCwdx/Q6HCwQ82g4V9K
B8YhGXPE9O7wkPbkLgpDCtzNXq0wWmNRyyRYp2yd2ysmJOxV1gW8Zpt4k9gkYhX9B+MhVEwUEmK/
C/VAAsm8S8rIn9Fiv19aqVrGwiLgF6qqzkxvVVANHS0Drkaf6CvzYKlIp4wyM4pDxIEXzp1Q2wAa
NVz7+caqfT4VHjUwliVKQByXC+c2sOAaQYK+Dvi966TKiaGY7DHEqrbBEm0wqjqLouzKshmIkdvY
AISGZHSGzcKqNRUI65TtCYjOQxYwK5uOqB4VfZcZBgCbla8kY2qss/Bd9ezJ8s9kG6jnCSitlZxX
HoC+kTL05LpU/QahUpEdHfz7xoqDtmunZ4QMt+csgebXAFdNM4b8MlqAGzaTyQrs1gqFcY+mQ8zA
zI1R8xuvMIkYG7lyZWMZ/vYMZ6+SS8hYvMr1buSgE2Gjod04pyAOc/Xgk3Wy8jxRj2mlQPHKs11p
vICAoLd+xPEdSBgwjykCF+6Gh3ygAbrLesh1bUKfAlqGlIIYYpbw4Kw4imR41cHeVjD6dPyJamdk
2GM9DuYCNP3IVzYlLv7s2SNl7Y9fFJK8k5xLAVYCOg/+AaTEjoEFKQ/0zUYORNY/Y1reoYr14XET
ZLlWgFOo0dDuMzNO9/eIReR61Aj2wWsPCcEl6D4aNv8rDtqvR34DbPO1fdsrBrF1JRjSrf4dIrUv
EuDev8th7xdNldF66O6Y/YI5xbGKIfwU0U0m0cMwR7LHyhWX396uJFtdAK3Xf3he7v5foAOCOJzT
Xw8V53le19VjVuC40ObOqqhmV60GM2+ReuZr1Ppr2fgs60d7xI+CuSjV5mSg/WH3x2O9ZpNYJpF6
X047IoJfL3Rd1khib6v3JCzE+hUk7YU0toDFsDVzO5miPu1gujVA2qC0TnarzA9tyySnU+B7xElG
aY5UKKaBHuI3f/P2C/pd37tGrB37tlTvvUWJClvH6tcQpHio941xgCzzKsDRHs6letqDX3rx/yTQ
FDp8CS//uWFeKNvqbqJLA0Ik8gM8wahG36n1zTZ7pmdA7iIWF/P6hcPerCeQhRnjbWVNoP6M9SXe
d+0amvrHavMsdx2H2cgk3enuV6DPh+aeDHh8mDkhMWTP4Mufm5iCZX6c2L2vhTzkwAW76LZ3CYHm
Po1FwsE377qE9VGg5z0iPBy+26EKF8F9Zpm120cwlllrhFiWBo3nmOPom1SPnSSDe9OysXHO37OB
w/rFMLunC5G0NdSX21kWua8AKTMD3BLhCsyzwScEBKjhOacjCTi0LdsJidtl92tUUqJUxjonZ/09
YEi2eVwsB90E34hVSKhZNUfE68XhYzGRh3PpF7KT8pSO7nyCilTtWSN82S/7v5lj8mPSTHEuH8PU
d9cySAxzf+dmJFzl8UETakBvTOUZ5CaUTmhtk7+YG2jzAd75NKBGfxrjtIC6F69IG4Job/4tUK1k
wZpAo1dIDU/EbVbm6uqzEzDzv+7y4gPdD8pYP1rjIUBi97ZeFYL2E9eBvvCrJGuXj9XuxoYrqoE5
i9/sMtsMV0d198STR3dhpAjbyICsgl5CwmBSwITl4MDI/FL+DjiYnk1aV73fBkvazm20TjxGma/K
/D13EJD6XeYB/PjaNoHkyLBMXp6eqY8DK5BX7k9U5PpzO/g2vZpTiw6L+ttuEuVTxAXXGcHvaQ0x
/YsHM888a04QqpikSeX7dWvpNawys3z0kFOx4zmL/VHimL1QtVSI0LX9h1hNyht+AKQD0j1GR3VR
3TnS32kd4Emm8YPz/KANV1xFUM8gJ8xlIwMRHWhMrRjm8CU6Qry7W2OotGXIvyb1eHQMLc3p/37w
WdYslROHOpM4yHmIK61Tvy5gQ87gfqrnXOYKO1Oi6idhYvpP5+wzXgzPdVrb56daHZYOK60R5dHc
pnt9gts7W/0APRbqiVcLSZswYzVls06rjKktxRG/Vr+96rhSEHFAEtAFfF/BydFXplkRy/8pk/4d
LS574APThrRFUGqv6OgkbfOxuSpG0xdh6UbULU/szF5nG2o2KZI37iQ645ynyNbhxyKqFeJ4teXT
z89Y9p2eFd2CxxqAcnfZtI3ufUSXy4leTF7p63/2HyKkNDW/WwiUiyRS/sZROyRjc0bmQE9nNiwB
NRKW5F+2ecuCsrkV6bvwWv3eunKOs3CKCaUx2yJmOErzW4gyDbrCqXhRfeVOdPmhxIKyK2oKorLj
QhS6GapJXcvjWfgrcSmHi+Wzp8j/BAqF/JUJyeYI2iu1OBlmi7I4K8Ry5VJTt6QJXvj0ih+uUCgs
NuIwWpSh3lYfUqtG7t7HM8kh4n9mhtZDCLQAFZCYbrj4vJ7opGkvf9CMBysdrVDqqqCXUh7Z391L
hirPyQcaAcDnAoU3i8XWkUK01PFNOfDlk62RUaAs5thdw0vwn0k6FiKG2fxtpT93OfsDytDLqpeM
mVzopeonXAjCT8HimUfYb4xE8hK0d/Jx4yMFg3gm9XjbZLAzHSMqQPW2ikNw6urlSVT9vd/Tmlfz
+8vJF80zYJ8fF+Fklhik3FSbUlvZpv1cog8nLFwk7CqNXqnuerJ7cpNHJfcVtl5D3sHc+wTfT9jq
YdlJS4BHXH11gDdLU6VAmHVJqys3WhTzn+wYCIQgtvfz/haTTeCVy6d2kVbbDPKnL/8DLdnQ2OIZ
7msHLN8PFmqcbLHcGUzu2HoEj0IMow6zbSZ763Ub5CSosuB3cOcmDrQkrcAHpTUKXAuQ8uTIWCC3
GsBfEMngp/muIzpeL1POySYIKG+2TQ2tQNpZA5+oOhw3C9fOB7+0QZvm9DMoKsAFWxjm78Wy4lNO
CVSIciaiV/pognbNW9yQgyIVMi9jxD0UeZsZ2dJUinIFr9FWI/JtuBSw3KYL3B/Om2KZk2ooXsMd
f5qUyOyV66Qv1jt1+OL6Mr3OptRSoCP2zf+TGp7QDZhdQyQb8Ur1UrdqpicSIQZgUmmxZzbjnss7
3EMnjIDUkiOcg944yf5UyCHz3dywfHaLcXjooGUF2zo92oGS2ELgVs8QhLM2WVIG7T0aBBlsP5m0
ZJ7KcIjJA9zd/VEF3KtAJmI8r570CUXsGBsC7vTcegbmOr8IRCrsrx30TRB9dOp8kPTehGxIMF0u
1OxWbXwLsJo0XmViT1fpB4EiPF7y6PFjeyAnLfyeqeyOQLVzEMfAF+JdYXD545hAe7lSHmGlXUFq
HKqD+b726ing3UGHGZdqwEb1s4ywJTMnerYq42hjsKZKxeJpyIzVlsccod8WiP/frOAMFlyPynXq
WQC3TMt3FH7QoZj442EFnzszJ/1YI1ZIPy/13XHPLMJL3IWAYqZYJfhTsxIkR7x3mnv1+kYWHBVi
fdfToaatASx55E8CIdaMYLaCeM/+79LJtzd3KJDyOMh7PR1COy3xzRZhY2woYgwTxjzjmZDbRdU+
xKM2SbZgtJdqOmxJuNEInrdGSA+xcGeMw7UHwrR4/0hjoEur5KX098cZ9OPl9aCt+7vNM0kX5pFY
JPklrdV64jL9SN3jD8Mwz2V6koDAztkx7dZ+kndRpIDlS1+luK3uhCUPH/1VqseOdqn3zF33D7nZ
fRixliyamvJWRFBXRPwG7uwbfiuJAw985mfiABI/MSBOAfANYbgUKP8n25qIRteZOqekxNIFsHKv
berb3FhVYVcr7u7d6UuGcead5/byLv5B4OWJ5OeGCPCfPuBg0aPoLDNLuvZz51D9gdafeDWZ1vhP
1esVF2C9hTGxip29+7ff4a7fnklIJIxmbukgCgvuKzyWk/I0pgM/sacFgArDHfw2ttAOah3MCzDC
TgFZ6In9McODzqfZEBAJJFZLT7svrz9K/tEBRNzhL5XGF+mBOfzjCmVC+BAOkzSqkdt8JG2HPdUI
3879aSPOP6+HIo5FwEfppb7VxV8dOh1ODyetV3bNTSt+o3vg7dnh41lmKasUIQ2qMOJBjDm84hLv
7lik/DKsA9RvdNpruOp+3SeOjBa9REqzhszH3PT15LTlxGXmlT5jiiS03DMqFYfqArcWExLGbw9b
nUNhuIOlf9Ugd+6fmttXzsY5Y9zTPg6Glq9gGACC6UZvAFdqTpR6LDgKRArIwbuoI06+XjPniSUQ
oqYEpzuktRDGjJrIET46x81KI/+pFas85hfHmDHxV+i/R9t9aBnCiwhEtudrjTHsQZA8OWKOWoZa
gRc58fSEycYCd4eQvwcmPv9tunilXaBhMCK+WaaG78pFu9PuiO0tY3ylQOmsoi9RZXumaXb0+mgb
fUPgKT5o0Z00nIk40PLwP25MxWROpiEs6RSyZtVqjjFgg393NeBLvBBr1RjpdflbtiOiVXe9/N+g
hXxyrYhAtdOr3zVf5GDq861d4FnvsKtFrdUrsxYZWu3cy3miDqld6Fuy9sTOw5P7QCKU8DjruY03
n4SKFEgMj1iYWNO3nfEf1luLWdk+PgzSBF0wbyzPfnB2ijJBZCbstac7WKMBsfmZK9rLIO+BWMGp
dFEOfyEMC9I7Ad2zvGF4nEO/ENk1XL7OJDhLqZbYmOICnae0Et5TeP4AEj6h/BOlFuhtHQ5Dg9ER
EqGzq47Mc0qQ3K7bjAT63UDV73fbE/xRcgUU/YqgNhv601jq/pfn3dt0W8sIk82zpjeHfjN5CTbf
22Iciau3cTLeEzdG6hFAe+0vDdqvChtRIFKGcbVFmvft1X6x0sj29ExWnt6YK080k/rYRwTwayMO
r4QO1F5iWGttvvTO8pE4aHnAGJF/O1Jx7vxvIgnSC3rZnHLt+4jp2LCxTyQVHBrYDsZbqTuqp54G
KdP1YEnO6wpP7igf+94uWJAl4vOzbaxLOZj44v4kGOvVJDUZ6Uq1K+gCHWhOY+CxhZ2zbwOoCQTV
GraQh+IdyXifakQL+EDRbJE+gOEV0DliR2hCQ62M4KNTKA2EVAJnssDuYZuZF5Fc7Pa04TyN0BF4
KxYz6oYVWSJQAHL/gZIyHpgATtor4sCAEnGofS0NF/HHqdGPvPJLKd0Eko9csnXw45PnI+UMDgjN
Y6AsF3e8smPUCyvmp4aCjFx/KVrv1fztTCu5E94nwxcYPf5kb1vOMFk3nht3vHMQm61zW4ELPP7Q
4b5esL952sN8s15CPO19njucBC7DwRRqXL7cb6Brv7NQMWSIQYAolGv0qLRMxLtdpmsuOO2KRHPa
2bjE2vvPjgCzP/vVx+sATQRD9K+1ZNbe+3pyUCq6zxyAFjnXKei6FlTLKx9PMVgNTFjUI2PomOPJ
GLn3wQIu7sYXRnxofG7HXLdmYPGAqt70872QsWjsdQXsJWDREMdN4f91Uouw0FcQAWlm4WNvzvg4
/iL4LvSwe7J7wMKCxVoH5K8KVRCnUZpMDoMHaL3oUZBkA43oEpCPSeilS5bBI50O7B7e+nKvCwzA
mog8vY3TAxMDkHQQ/u5GRpX9UN+e4fyPg5W90d6fQ7RHB9WuqdEp4YSJZJW9gY7bDOaIpcLHQV71
oW+SDjXjdyUqHRX9R/WzWx0cwiwMi0expHB7tl5EzoJcHSm8nzMnQkOwUC++DMdhg+iShSkKlgRL
aIMG97snHaQV4rQEw5DSn+QSC/ZU/lhA+B/7Fglna5vMHTlF9Ml76BLXhF3KypAUh5qxX+g7E8Rs
0QSWUg+V+XVQ912nOsXJZhdP1LxzhsZEIXJdbwRLzYXsnA+12d0S2g8jhUrIzKOPGGNwe1DBhN+a
iXR1BZRSsxFZrkjATe6Kb5Ii9u0axk9ak9WgHkAPx8QxOilauguMJ06Hva2m7Wgi45BzJ2gn/IJP
zdvhPzJn/A3QWwD0vEETtatn4edC5fvKScVQPZ7Qfq64GiQ7pOeMT/x/AwH6Bn3PkUudvMsg37V2
ZCoRy7dDHzubSi9CjxvOpI/XuwKJCdoQdFlZologYMnKoNSoMRWr7UZMLQqp1LgxUScrxW/zVUcX
YL7sQNVcCj9Od/SDOHYHX3HJ+e4lhDz0AifI+2JRRLS8pWxS7I9eBILBEzescItqZfNtG8Nfs89f
WZOOZKP3mZ28Xui6l1qng3Tjvd3UnwxHBgP/Xd9hc1SyFwrOyn8tn51LGi4YLWloAEX2E6Zpu2OS
qi4frSLOCUHI8OOzyJ+4AODOfuxaElk8woU5xmg4cmRdxE17M37J/QmfugpzUoY1sRsf6bXjqRKx
xVc822lAik2wmCSrxJiamevIpiwdT1zp0FMQDrUph+Qt4EDPYB9tZHtkwTB2RivsyTGpchoCF6Hp
4PtGPX8xDVO5H2TANBJzx4qUmPr3ccvIjKiq36ZDZ+o9C0Toy3KTC3QGmN8OLhrwRBDrerkKUHTu
td9Ov03y0Mn/pk2KKpXYEP6te5OIGRVa0IFes/kzv6kyi85qrpOeyvuD1uKEhDVu2QYxfI67CxEC
e5UM4qYXq6lFelbDjgOitKaixB7FlTPrGSyNyHHWq+9l/rsb+/hAmz+sgrIqVHBThkTAGC9zcL9h
6jIl62dXxJGTglCwQD8+Vx/+BbVWdZdZ8znG9rOLErEyPmi9qs+w6z8HgYbvOud0xxSC3B8LUU6M
pioneAIVqMIXzyPvE/xgUHzkW9WJ4EhMaaZjXC54U7GoHVXyniRW+xNyJ4fwDEmsy0aNvYa8ms/Q
2AFt6VZY7ArqK2HG3PCgDiNXqTTOK8uc5AI0R8C9BkHTWbQ7ACzx8AhRTvdGG3jD8Be2ARbOrgua
GKJPGCf7M4z6toEHBXvjSvNiWxCtp5zPqncBO/eefcomTbZUxU8294ZqH6mH4cSlQBYx3Y89cMST
+o0if6ONE27ADqJo3CTQz4jLwUQcqdrekTmb4BA+o2Vjr9eTS37Bk9ISab33VxMHdcJBZetIqpfd
l9XCu8Eeg5E3fhZoYXiXdiIld41jkkmBRj8jW/ztW6Zi3YMdHkR8BUoR0QEp5XeBwBNUfxv24yeR
9mclr29zT8L6QhbWh/Ue+QRZIsGafe9Cuw9abZhEulKpJyh1V43HOClewDOK/t4tmxY9Nj1Nnk6x
SPh3dUqwSifTZ5wKJXtGeM8H4YdDJPMXtsnkq8enWowYexfJFLuIPQIimQAnZ6bYI06eIYw2/NZ5
hGtLm05jUmt/rXiNN9WoiqDPH4ye7US9MSba1q4hYjdQOhtv74O5e3FydFBdnv7uIDon5C3z/sU+
cIA0U9POZrFWG56MM7GZUG2dYazNvsoRWs8iIme/TXuhZIEzRXzPpTEELbitpn/nNMxi+ApkOXFb
7oETTvxmrNWVDdApAAmx++w1EOJr8Hprvoo3MF9XFMp/iIgvjuWSnAw6tAhoBTalSUQxnhrGFVYw
IaZq1ETq7T2h3370QbtNSnuu2SUI7c14M40sRzXCy1h+qajgNjpbcNQnnGgWPb3GWNL8vut3Ms+5
C6kOc3yk2wRce5n38IzLR/OgWwDYROSb7PeZa4DUqTvZCpmEJw+UlQGMBax9Efd8DOPBoSIWE/IH
0cmI6ADUcxrouj5iWZWfH8KdCMVBsjCGwPFsTqvF1OnKnOHz2rwXtTef14J3og0ed2A8CQ+XycJv
UxfXB+CCaFkLvwIjdUhPgxi95DgRPQaWz4IV2hccC8JDVYK/5egYjX1PNQ8jKurggb9pAmNj6EVu
PU53c3zyrJ38a4B9w10WrLrfqJMh0g95gMdENT6s+MBO6UN3+VCSNc30XkM4ySjttbVxX3fhFNZn
Qd8BshFZVbn8uqdqjXxfXN9JGxY8qSRPC8vWtFo3KLcz3Mnyu4aIWHt+AxE8fGDP1jbGO0WMWspu
yPWSD+OaElH1RaYlheeVAiQhEk7xEjvSWzHED4DzStanL06wjW1iesx5dq6Vjmdtj/yZVAx5wCUc
yV9aMkBUkrTd0HvDwFUp9M87iVN58y+M22GBTSTASwyDP3SW0+SzAxKr3F4XlQKniPcVRBhvTX4T
hnjrhNFoDebIgabNiBIJ77pUloEXvzjdBK7oOJvY8Rt+MjozDTN32Xc2OfxustkSXf1RBT/Schsy
ROePvgkUFzgMqjP2bvOhr/9FEQAQNKytZ4lZyk0cdhJZ8mU4iKKzugZtHv6snOb7kcCYJ5KsNOxl
oe2jWBN29zh+6wCyiK/O3asWMvFh3td7DHNYVjXD3xJYvBfQxEkYppeaXgyBqJ+hU9qP87ehhVVr
EJi231cH+Hhy2IingaJJjceh9EFw1EhTDH37bf4FPYpVNjn+SvzESTBcsY85xwahJyAymwBMZYjF
oS3Wnf72mLSBj1eQ9therKRGRhunCgEjQOgc1l8qyNNhGd7vMdfIKp8WwbdU0nJUmMPyBcrcJXKD
z74LQ66fHaU+J4PFwKFfhCmc3Q+x5XrCir956yIdtW91ijgVLYdAbr0DVJY+2iGt+ZtrP4eNJQoN
P7LhMNhHB6Hp6I6quV+MkWSzRyGLZZAY60E5YZNaNrOoN81hq3p9MIeFZlvIFaWsOHCFoiXBjFFp
H1UC5Cvs5a1o1Fc7rz8zdUp3SGzECRJA3m9lJbux2oAkxw7VROKo5KAutFtsU+kNmY0kFdZpopHG
ydtyYOv/fChlHv6QkIZpcBhgY4AENvuqcKLjaGvCzXgJ/dOMyMU0NuthhlJX5WY7lL+Y/kf17myB
xUcZZtrtOGN2hrEmWkHzwS/ChTQoWCLPFSYu4zB6cme5g2xBe40eDCCTyfRp9zjUnkXAjpsyKIso
s03n1eA1Q2Ao2OQ9Dk4OjJgzDVOVyO/TTPRc6Rh/ZC2dFcw3KIp+4PHdgZPuTVohL8RkR8ySr3HU
AARm40kZ2agArolssYWPbo/IkyAQVW+eOcTx9oaMGhkOtaHwNmGBZ1XJlBkWPgq95zfjbMqn8Q7C
9w+WA1WKRu/aGja4hGd/Niha3AA4T7MAcM4sN987NEf+PEJHVVCmqnzpVDeFKX3IlX1ButBaMrVG
dfalsJJB/Dg3nHJ3mSZngfG3S1O5qhW+YY1SFoxV6fmDUi+klMSG86OsXDS0SdUQVyE9GTWa6AiI
fqRGmRlrR/MwMO0HhXusgI0IU+KEK+kU/C5CPDS0jFl5EgjaAhqBDLWlr/zWCErLuiCOnaIcxzfz
LSmUsgX6uY3YjLhSCCr9fIS2Z2cEA2jUUrROPlGQOpI5dTOJ7AIqZzQoaiXw76ag5OVURaDCvwmo
TETcHhOnG26wDi+xRDfGVhdTMzAKHqBZVwFTBxHoBKqVU868yHQ1MD0OWokJ/Xz/5tRL+e/PaZEl
vdD7MxLUNddauz3pcpHSc+xFy3Xzrv80dzp9gvvVwdFLVVrsvzOlq5XseQaUYYrBUmzUTYcJ1Mta
vZUChmMw/0B1g7F5E8lg3BR32l/krbEwHx3Yui6TKoO2LHUxk7/rfGieYgTVvrIcEVe07+ZQjcSi
CHDujddcHx7X7NGl/C/2VYFVGmsIXvRk4sUkCeMUEgfUCjFFV6oXdYwaWtFPSkU5hsDxDYmYAEhE
y12AJb7xvgE9T48HvFqgU9OwX5O165KzHNpVoPnbNHwWqsSlUSurvp/BhUhz/2IXu6LP+VjKRN37
qSFroCzaknu3okGKH0xrmBUlmV+xTCNa6KI//h8wL1G9XcRc2uEmDaNXDbNsgAut4Vr17keeYnqJ
tf31LmdkwtrQ9+QPXyYZIVbCynN1i6bsNzccJa4JN7Cn2KZSL7I9kqCOD/2wZY+aP4w0Er4rtBkn
T6G3UX/FwQmaIVy5gc+aWoOwL5KK5PpKrP1P9EhN9y2A25O9vekh+pfvkyFEq2vfo4crjL+Dssyy
Ct5Xs2uUIb02GwKouygiRa+hIXU7+sQPrqjPPfPTAb093qmmXBr9Tux7HCCDUtBxA+RhN91T8IJ4
XeTSwKvTMS2wNmmPWsHOyQB3dt1cvn3rqI2kb6SxL6tepfdTUboEXlp8Xs3u8UokIXclUN4jxqar
lFuG86bCWNvCLxiNRquOQ1vNUrJqhnlREIdVbzVVHlASB/ZJ1paW1NLus/eGf+VEJwOYYij6fNN9
qVRF9ysh2Ko/mo0F7YPD48gQcRkLVsyecmCn46egS1iE6lJ5Djf5e1g6EP/b3+wW9IWgMLELanip
8up3SZLusgdq2qn7QSTc4enzmLFWDOgz4x/v629xPqnGWMJv7Tp7J817qztQb6N4d6La5ZjNCxAk
hoEWC7nJlKAPuVMbjCPQHuYQZXi0lcGJTvioVuBQ3uu1YVhiyM+epU+S1dN5yjnhPyxwtVYV1w5k
JOp4d8JnRgwbJdye9tPZpOrZ0jyvgsIb3pCAeC89P+q493oiegGBpdUbji0OYR0Ju5HCzRqa6t8S
fw9JlUlCdgo9qj/ZKT6Lqk/9PNoYZ8LudBZ9/BcqCIWZ4/xLLRe5jfTKEXUEATdEwd5zX9cz32C4
bpwg5dfsCKi0FizCmmWFEnlTZwxP1SjDaUHqmAE1j3B8Ui8Cp6AZipxBUU9vaLtZMgiBZ/LAjuVW
1OIBLUDC5O/Z/G2AO3OCdYzIWu8dbzBfHLXifkdbZ3uPGbdBnQwYsdP0mSiYCd8kvhdW20UexAOO
b1lZl+/zemgPBrwqOeASOS8w4ZttEixLTAnwGqJJIaKh0ls/6vld5mQhcBzp/2OPqNO0UoH0AvUq
o70mQmQ2kda3rh8+n2U2oQsinbIOlUC80qaG5imUCtcQFnH1+PjTaNF2W+lRdLCASOVDHukURJyB
N39n6PELv/l7HJa7P6yYbp11tupKZAdT6NVLmK9tK69ubj3CBKBOKF7Sw83JSlIYoyeY2qHpBkxn
yfIRGOjTy0ipV4maFYv/9YATBLhWsw2FsmZXFVktbvMsG8oc5Frvp/wdXQRmSUqb5/U9vBOQ75hu
6pTNE5pD5KqPIpKK9uI3Lfz57vwcXJB3ev3EIV6DKGpXlhXre2LSUQuMFUmo7+A0RE0c+1aNo3xx
0ZGt8Ff6LBA9pZYjHJfLqsZr/nlCGeSYk4Q9Jp4ckQykGuLnBXi0klDzopw3qDH8ZAOXN52Ua2V9
mnF/dh61nApZ10ZG5XZfDeqHAoPh0m5VK1ZFYRPZ7EiXXKaNI/1zaJZORSDL1gBupgTvtJpiWi/p
yUV9tFSqYIxw5f73QrR2yU0g6DGCQeT3KUSo456SF//qQrGSkB37W/X7hmoFSpzxG1I4IxTvaYN3
EvEKoAebo0U3aTdrloEnzzbl57UJrCO/tuVs//B0HBkRnrJrDa2xRk5peoKrcswCp7LpgE7QKqCa
If/83KVr9LSfskfpv48CEpioZLx4erwFY9tV050mJembnRN23rSMxBTa8acG6gAu0PmQeDHl5HnO
HLPormw30n/VNEn57XBPz+MCTq3f338j1NVWuPN9TKxZihSpnmUvCstsvMB1SVSc1q1iApw+cskr
N/KguVFfhfP7aL3+jI/3+1tcq1E8K4V7oYJQvZUtDLmDSz/meN73rc5LF+UHSC2hxFyrkSb7fyfh
aQ+LlGE4UK7q0CK0XfrPA6zEnO6lmi63AfNivh1eAnRm3ZOxX1TdUK0vfF71NHGkrBHY7IRNP1h9
dX0lODmUBJfbmKiUIUDTsSNzjWUcfL41PCn3TftULGB1D811VBELh8QMv/bDtzqTbqR7CT+husRM
OfPskWGemWsjsP/YaFFZJg64qpbE5pS+1FMgW37OYxVoVXHghdyIGQoFvfPJKbNzbNsJVsGjpGH/
h7lV+bFhzmY0Z6dDKrKH0LXsrqYSH3dWMtBtTg9aln6V94ounks2Y59SvqQmJ25m3+FGkBIHcl4F
FgWjMnqg+tsUQD6XA6yGR6FE1kjF9wYFbH/6zpWOjKLXhGHz+os1V0jdZDCXCG8QKLxKC0zxYEjV
UHDi1s4kElQpiGndR99YEnrGyknrLjN24xoMrzTFPmIuHgthUAb8jZzjFrQXjId2AnYOTfu2r59j
MSxbyY/U28mDfwQ5pKc3Dj44VDwikHEmjTg8NDfSSvCcCkTm/AI7VQsl2wKvDF4aLfzgJ6GeX2pa
U9/MV60reBc6uf/YDnZUsf/MG2kKNeupQLk3yxuEVvmsQXqK/9tub16oSLO0UEg22n5wJnDoEDXB
07MJRKKUo3QNO3nOnyStx1YJdj9/qbKFeEbToSn0lQH+mFlmsAmHki2tVVBBhJu2L8rAxUjhkltk
BGF0G4yj1jKM+MuZsAUdf5V2SYz1zTeq3NYwY5ei+G3PXgx8OyOd1cQH6wYD5KBZpAmdRRNW4ZSo
N1lBbqw3rG/D4ofJcSByrM2nqDY6HlTm7SdVUiXLxpHFCEk6ExxpE6bNzouA5Q5HAfwaxo/LFtIY
GqFndju/vmcK8JU5YwvJsM08yNUd+NcGaZJybohdl1v1S/uIISgO8ao2xUhyBvz30izsSNBngcNT
8mP5du+RLegNu0GjazN/UEKNh8fLqBPNZ9ZRKy8va2v0BKns/Z7B2p4iv3vEI5ml48O6X4wNds5l
jVHYkWqqVmWMKdRtn8/EQwcuYwvJHmxZ4nhiZDZ6IrTOr9HcWR8/1trxeKwK+997PuOw6OXBzRI0
KlH5KCCvOb0p2JCalGW6O5Wo0daVyGQ2TRpCcoeVooVJyOoGAf8uIL7Qjfk7mKd5bkOEhXjzoFGz
5S6w+p9fA7Trar5ehTZRqf1rVit0a8irWFSETr3gjHOQOAYoBIxykSJBj90ZAPXIH2WIx50E0RNJ
FidIkS6nbq5g7Ge3i0rDGV6J+CtFbyHYfAjVtKG7tOAKHRurom6/0SYqYDTqiRBRkDs8ksc9AKaq
DiaPrQ0zkvmzoVav5P9WGvtruONqILo/Y13Oc1JlAcj3MBFwrcKG+oCtLB3TKUOb9Gh/3nRKaZx6
QTe9t99UjjnzpQSWmnovndAPmZ01UhXXRYyG4MetJjdkhTmLX7MOTTArv1qHOObBkm77xvArSTun
3nA85+KejYSi2aLkdXbnf7EnjX2GiziSp2nOJgzZHZ2FD+AiqYl0Mx71u0ihXJ+TdS+75N4HVWF4
1E4mRT8MWcnIUxs2JiQoZ+PL4r2uJVT5kPjMhPzRo5dMuhiWUyau27mHKe1ub0Pg7y+t8vvhPiFn
CZjQMxutvc7vqq7oKW+IRyXFbPPVixydiGpQDqqs1uQujVUC2I1HzTlShuWErQElvynJjwfED5OW
YFWOIyW0XAOka6iFRwfRYCs63clCQ8uToqiiWKqiU+NOKQ/zhJ9WNGP1+0/lYWFenx1jBTyqLswR
ab0MMsIW9EQ1Q3WXu90VHax10MQl7PUu/nXT77sRuW1oFoOVE94HZ6bYdl7p12OfvSEqVK2O27J0
SL+3qXl182f3K6YMzy6z50pGkxkm/o9w3k6o1uvKzEuTT9jzB5mV71F2hiNxAmGfZ8Y7hCkV7lWM
2Us9u1ReHRF/NELV3zkfl7UZH8iclqXjf9vwz6JmpgzyxxoxInZ1r9IPh6M73UZ3KUT97tH9JkNO
l4J7SPepT2HinUZmLcLmIHhPz37SLwugUiNzQi9/5VY3NDv/z6iB4K2nXiBeRrU9E+wzENGb8vqy
eY4RoCtFqjEaHwz3zM1HobK1E02NC+5pNEg7kGJYy5EX+XWJCVaAdKI8/I+rxF3RgWpU8dKFAe5/
vGiph9vONFL6NtCsS9s9AXOL/rKe+yfTsoPkFANKmWeCBfpV97aH/bsPQ4sCiHrJYE6l0qJ9tZ//
QP7QcpnmA0AXT0SKnC3A/3ppfcRlg+dt2jAHZY01Pf5uMI9w0EqytDDac7XdFNCiTQtWxxZVcRFx
SVFz6xYDIr/6mmQ80hQF4Z4kt0Vz270jCGYxq9UQpUqdua5zJiAkqAACAykViZbovpW1ia/MY8np
sJhCe1u7rmSRvISkCR80//K58KQ5vfMBM1oIFecVJ7IwWW9NDyUc058Yfngb4R94vzwKzMVkplNc
/A5oghAb4TtpDrAHKHmnkl7BgS5P/AM4L9ectuyyFmg4Z6mAnaUWas3DpwWS6oGGnyrLW2492iMK
gjb0V/rJ3NJUDZqGgB8J4qSAi5HDE7n4zS4vDXGMIV4xP7XEBfpfDDpvaMFOSQQSx7bJm9SdsKdJ
8rvOT3NQMJ1qH2kJ4zBp2yWjCLdSrDYrvEkb2sVDzduCww1Cv7S0Yvid8nQOP/TE319nRa654YUe
w5Q71GnUt7vuuWN79GspH76WnUbXphe/wQrjBKXud7lIOTudJ84HcM/X6IDu8dYoSfSTAhO9fgl1
nKyEhHTPlx6VgjoSs3G+tyO/NOkle/vf+sAq+t0a+4IV6dwbOd2Telsb4CKoa3TeBhbAab5uNVtf
+ndHMJTCy5/c6vXi9bVCaQFVqhbRQ3lODbVcFov6fEA0nWEs4n+W5IeaxKueKE58P9h+qKhcTKe0
nmPVZPuSLstlg8YGsuqveGYqcgq8Da6oJx84cytTwhwf3tDDIqm9eTonC3Q6h9tm73x95Qt8cTTB
lbL54PXE7fGLoPE9Da60SMWJcKzK6l5jcaJX7XiWQEsqTpP/RqT4yP9ExcXFfh3kfcFxmFtaPfLm
dsyjwWvocvCJ4DzGWX312bWEEqL3LDm1oKKkUbSBxcWHhvtb0u203q8FgK5ARnAjTQVgf4GwdnSb
hAiVa+coAr3bBiXYwm8m8qg1emIjolMUpSA1BKIzDIqWQBQRAtcJQOAeJSxoXJjMxtZwS5qrQY+I
oeLOsIMlLGGO/FntLdBrIHZv3BArvqAQr5kMxUYW08iTGLJfVFSGXJImfAhdlqK0dHfvGBiWTJAx
GSOA0XiDPQk8XMhr2x4HyL4x4DxpPRDL4r/uIUrFpuidOce0UdV8L0N+azfEGHvU8PgFfeZpr8iE
ooBjD8pZoDDI0M1IkqfLBeTJCFJ6txgX2gvhli9bjkOCxN4z1zhprTQUSqC6uXh4ELhgteYbjdmY
uL4hCvUnzmHIdgaHgK2W2p3Bjc1uIu296wHI5JQUFm70eAdC4Hv6ZfmLIKZyQkbhRHGSk1Zn8BQ6
7rq0bN6qwSXDeO7KBDDoKTJ9JalQ64LtijXz4wOZMemHXIUj1TtlVySRidKyRSQ+QJ7K3w2rXrRZ
5Il/YqAUFaLQcp0UbRa/TOTju0IQjt9Nk123fpHhEv5BKwYBKvFHt58MQ+hl6PEVAn4ruS2Xuw+9
2xqYhI7inZpn1NgWSFTECg5hbcrutQOKtkykAsi5dJfetY//P3jVoMRQQnQKYCGyCcFc1L5vvifB
dTaNEsGjiCrsqebd9OxWZNgBxUO5kbDh/UnUAP1dWIRqSQPkBamI5iPh0xz/JbPGSLLLBCwdq+Bh
26H19iUxmPA0Vuhu8U0KMNUYp3Tgc17tgaF5U6gIJjleYxKVVr2Pq9Zg5G6F58KwAZlktyK4KOKR
90nYYlfrgLyWdUu4GzleARVxidvoBp73ggIM2qMzEJdKB7YuAR9hKs/zmbTSZ5FLe3bWtMr6RL1c
gnsu4vmF/SNQ8XpUAtv5m2XyY996+xXGiPty07syj1JJXTC4OGlB3EsvWlNMLPoQ5NWMV0Xkrchk
SxzuB0yauzaj1DY6U7GSUHFwPtNltz0m7kmt2RyrItRYzihqc4XlHP43fLQFuEjiWH8EzyiYD4/Q
R6WY6CxM3HxCbh2n9qDyO/P1E3PYf/YhJAweFrAJIka7TFnHE6OTphjp91GWNGPmqW4RhWfHJitF
6l2tfiTDgizGI+VSThWDvgdLNt5Dx1Z9p2GaWEeJQeZM6BFLMJ5fwXiZCxRkr3G/9aAtWm7gLdZD
naJN5XIA/y2u5W1fFjXmOTEoOK50cCgpdsp6zYe7zmFhlu0Q/rCNJYCD+8AWG7MGSfQakppabz8l
ZIUGUVCyW1/rnhakG6jyqD4Vl2doev31d47IcJ/Mpl3PWAMsnL0OjnHJbYVeD7p/weBuPndCDudE
sjmoVWrKUEAUjXpQfHowLcZ4PxAjYHV7KOadfNkuF0esYSOAbkqRdMEmG9B4AC1UMCTZ9LgsV5xP
McmRyLR7rTSRBubP979aMdKGDa6TizSMptSwtQclURg9x9BGB5sCyGMMhu+TmwCAO9hjPKm6KPHw
B4hjl6Zcd8QUqOLkXSOEQUS1dOhPjFQOlXfcxjo2joifmVb7U9FIz26YKkRtBgRnSh5Qs/7AzXAk
tYOE+Z/jDy3Ixqr1BJBRbtqEqcOQjUpwsCYiUmR2IF7vcQ4ziegdZGcE9id63sVdqvrTCFumku/X
bBclB4bUyPviH7Z+HkSM+w+hNWWC0V+ZVjWVvxEacaA8Gimqdeub1GcPrGP74/h6Hx0B0e0whxLq
PAqM9mfVD1erfYwh1T7qIuCtpkdU0JTwyMIIGMiEkuzXQo6xMI46FdKD3THdBoz7NrW2NkO0PTc/
tzlKeyHgesne0sF5Ty1/AFIGKx1VIpXpMUeknZM1ShtQOVafKSN1JfWKoVSlCULe1Pl8bt4+02TE
sOTNp9eBJ2Wp7Hx6I+eB4GlHvoz1pvcNWOlt41jjno2NuNo3sYTJXr/fGj/pg1ut56167RhNkgsv
d/l9kjTXrdxBIJKFMf1iQOQDSUQvCWxZO+qo/Q1AOZMnbwhJ1YbrbYJLXvZF8GOV7UAoU14fxqIu
Edlrd49RvxA64dYEPH5zkyY/WVsk/z95veU6X4Abq70YrlYpRjlVQUSglMrThat4dh1/RN1NC9K2
BxV9fKzT//tlAdYKajQOZirV3QXT7CACAiX8zOpxH8Sbx8KHxyhsOB9l2lH+32JQkZm3MCix3Sc6
Xu1s32JH/cyQIT1udvYrorzVJrvrlQeJOBKtk/Pf+JKLNeOGi7G5ZJBoUJpchfk96SQE9IWooUMJ
c4dmt6OxqLYT9bTF/DmLwXZmIqaQkJuF3e+gC8YgTmRf9WZZohuRseW1L/pYIW9C05WzF2uWvh4P
78HjQWhqLTjeUjVJR6noJSGri3wQitXbiz73BlBZcUX4vnq/94+tZEjsmiY51wm+C/TU80wW30yB
Tmta61CPFdnj4pX3CB07AAQfa1ATdSTpaCweNNTLVQzZX2ZcumYAM+FuLiNrG5UB5+qsaLbk9Hed
8oG89dl4mhjK9E2a3dZXLEri5nYI/9j8D4Ze1D7RpjrBdO4eqAFP3KXg7RFRMs86efpOxaRYZ5zz
uMp6Zflrt0ZA/6x0BAdnGuOXaeS/Naix83bO7Hl8cb6CQSKBkT+hMOfcyuXdXxgM1dUC8H9SlQQj
ETRNFg2VcCOi8z+OEH31PNPxRxqhtSG2MKGqi/bvdBbF+iC7O3hELuie2vlyVLHhdS7fWGN6qp2O
BOX9rWi4CIuH66MT8YNHHZGwJ8psuEqmf8uQYYAQlkq0E1iM++eHDTljj4yrGjVenFLeY6aODBMe
A8p2hw7Cmee1WXqxdbzYdWq/jdyBtLFjtazTaH5IDEE4/zd5ZbSenMfdU4Fm3iXpbuKLexXg4RxD
9cDWBL0lGZwUNDCM6ZUbcbpAPcgu15cZvAKk+DiqBMV+VNetms2scARLE78eNe3A6YzkwONfeNf3
geDS367M8QzcKY2PGWzqYTALpq371Yvj8XivdV9TJbH0ZBZT95fHFxG8FBP6w4v1Dv3bS7h9lnsP
J18vYKyPwN6AD7iGT8NyjUNBVdaUdvhUwgi/N6MmK4gtiBkEaemDMeeKgZIt93XnzyOuHxzmSUXX
wmFlVfl/1JI6G0JmP9LkKXC9Bt/t4lCK1QYkGPEffj3Fpi4TGl7bv/dm78OuTDEWMu7hXXA3Fy9z
o5YBG3nLBPYZFd/5cb9RmzM6Pw2ryiagVb79q9sK/lX64h6SlfAEyNGpBxOgQZEuAjsnWmWIwqXJ
ImV/C+bmoj8GSxgmum2G5lFGcDSnOPrAw+2KgPfgdxDyuoJkSGY896NepTfsvniGCpkHYRexAi/3
4mIof4wDGh9qg/niamXPFwX3itnJLV+ta7dEL8K3S/wPm/bYgUM0Pe9eTePNAfWDD/ZbiWPzCqTh
Eyh63JdUeN4Hb678SVKuiounGgL2d4fuCKkoo9ocA5ygs1A9rv7U5P6brqi9VnxgXmPHGtHQFwEA
EwQ62UwYpOfTywyrAfhpIPweXwS2G6JDPx0NkEw0ZXxGmyakdimgZ3qXK7A2/eJkuPt+4Vd6lKX1
SYO+/cIC8Aa/8obQWx/0rdVu2bLWgD4JlT1HO+n0PHNvvD2+SoiobiNcPbPT2bpRbMKkCxK7YMno
hMuG9MxUhjtLvz7kbcWRjtbINRAFjAYq08Dpbf6pyXakGyoQCQ/ufDjHuuknmFUsPiLK1PpelopU
YP5IjrflZZFBzIYod53H5F0fHIjqleRXn4SuUGvS6fMSbmf/cKxjxtfFi85eTmfJvTKnEb//wVHs
ynyr9ptDb8un9dDDVWKvY3RYmq7S+edI74gdtYZ+1x4avDmHwfOsWKEkk7Dp251Je5M7BYNPeFZ6
AnhGfv5424hw+ty/3GshnElbaHd1inNO41IOHudnE9wtpFCj5h26GZ1KB5X7kJVwn4Bd4jeRLSca
TQ+qIWQ/sG8wnZHfyTiWHPrygpT1BI5QLERfDK3M5QvfZUv+YWPZL8hvmmvwstJZNiUYa1VuHaUm
oD04lUVqUEQQ+YzywrPjoZ4BF9Lb5XY4xYdTcEROPxRKa57r97FyxjRRn/N3+Xp4RsfY6I6Eg7hj
E7qlTyAlYkSnFEVOvH0PJYlKyRfxMSD1Qwi8M/Cz8eNoY09Yz0dBeZaTjQshP5wn3hNDP7Y9O5Kp
nj0YA4ykf8W6N83yA52QWJge8wKFkshzjtmfeqBlYA0zHkRbp8JokA8MwJIz5YA+lgQH5Hh8FgTw
WIrWGEb/ef6WEKGQaaUWehNcnUqrFqV0nkE6oe9KVoALFUIBUbwTxgKHLG5YV4ezwAmIJUM/QR6h
lTxBlAkAuHVZA3IhViANCCTx2vNADgVHz3aSmhHrDI4huqe6qkonbaW9Wp7NTmg9kBplhp0hqLZ/
BpK37sea8qbo0sCNRfrR0zvsRJZGVLinrL/WpDWvlLwYr0BdHMktWGA/DEUSPKe4SvxeSZix5hKG
unwvm5oKwQyWPg5C+qoFbM2NS1koilPh2LHHAHEbz1X3NGZqEFmDDnKzuDFd0y0oAejrPnuEXcn+
xcpmI/aDYyxAjjMB95qaQYtgm2CNnEw9qgD1rCvwvyAPko2H84ii7oInqjCO/eLiw14pvg7708Ks
1lxgdHRvYqvaOSVTHsfvvg2u6jJIIhSbapRU3LrOtTKi6su7Ir4mP1Pp/peUz9rnWf3nZHP+mNuL
yaieHOXrlfG5KjzMk7SJQmOjHD+xJyj+TydHWSlixi5w6C1VxRuF40kjdCMxZoLMGH9vG3/dvQ3L
xLEKmQgy1JWUKkSBQih77kJeTw46Vpn5deW9cYcJHJuWsh5wB1eXAEsb3RGlzp6M5sVCto0aqvIn
BAXfBnzIWmXDzcUaGJU8K4YhPTU5fijMVjbkc8mXdx+MMXeQrtEeTx27f8RVmOn/QcxI48mJE/rw
Y92jItx3K478ZhzulbgFbmsign/8+LNCUIrZ+dVHfx6emTOQ87eiiBTajfnVOEDuVuZ3WiF0TfU0
Dd1lCVjR3R3L6gNUOZDjQ4XEHrf5imc0aE21SRCs78Wxi2GnTjVnuHN+JcopLstuRVHwZtSrHILT
ergCTRJNdaWPHCU8uN8/GZrLFBgoqHp9QoZtN0cBcY2BR20cRM3IB61XfkhNKHHMmWmowTdG5dSC
vWCqIdUN4jjgg+w9hcEubsJfYWPmWWrOsk0sExY4eqSvOIkMAnQNMgQC4WtlHK2w+ilSFEnOJXqn
uVH4Ip4MDZpI0j/nQ4gmB8jkR/MqBexJ9lJxJnvX1ICAyuxtZ2jFK4ZbMfZIXHA/QVSd+qBPUFt5
mqYIlf76b3y4waI2RBeFSwrPZiCYHxA+RVxu2roWzxrBt2NT1hhxYP6Auq1/yoNNtyx0AD7bdu0T
HCkjUPlMmWmZoYliapnEjrJoeovkq6lgSjHoRzxEQrzBQkU5QanypA7qjjxOT0ldAKBnBRg0dc3q
Z44l9bV4IzyWTkegrLATYL6fvIdQmRizkWErpQLIuTwv8fOUDg708XEs1ly0NATazQDbZrLEqsLZ
UmBwp0Aj3teOwrX3J3MqUU7EBGZaKXBBsaLk2fohyU24VzUy9lrY8qr5D3RNdIPLgZw1jvg1/s0q
HRSAPt59YlzCeBNa4uE+EFiGLeADWDfyYwuMi/cBwlBjs1Zldbk81+ef3pK1S3zgdhl7tqSPawpw
k+QYkggcpAuFcPZu8rqJTdUigSiNbn7cCFEGLUPc57wymx3hP+jbJBmrnKcNUL2x7znLzBYUVlmd
nYY9hK/aIyu+tIYYQxNUXhNhSQouPPOgrqQQInDH6haZyIn2tGLY3hNUUoVj1eT6xodYCWUMgj0u
MV4+jTXJCaSxfwz/N3iNXO5K5Dsozc+PjuSwsi2zH7UWyX4ESbdlNLhHtIi7T0HR7/V4udLAJB4J
Sg7+uZv3ExjCQKASIzlprFS9ekFdDnXnrlMKXVYF3g0X0TJqGYhMsbQqDd/bOIt/8cc1p3SkewrS
2nGx2ja43OASyLT7dh2rx+mNdLFoRxETY59i9FcsYfZlH1iJ1QWST5aoIz0yWxW8luZAbLwBArCQ
f2MBYWlzADGFe4YE05ehRxAWQZ07hxbJT2kpV0zhIzf5waqDQdTolWDx7NmW4VXSYAVfDZoSqWl1
nwcXRTwRBn7jek3cYxHrGDyS4AGayU3q2ay3dBWKEAry3OYLYwdq7h3RkJxW9r6+VE0p/ocHQkCv
cs46BZOK2CgBS6gnYc8IP3jcJ3yfr0hM641uJ257DkadvShFAfntFTeNFYGJR8Vaz86HQqoATdh5
8RtglZ/+QDGagUKTVOQnKEInZ3cPCI4WkFyMupSbsRHcHmoG8T7e7TbD4tqNXZLrG/5iVeUKYUDZ
YND9r9ZXYGS+9MYCExaIg0bt5DqpGEFquH4Q49Igecx1bnZZ7oQYSBu8QeVbUWL9j6ddB+kfYrn3
nhb1QhUt6dc2kjHsJ8oJMSCz2ogdZZDkU/p+AhCc1O4sUTYkxussf33JLqjBfk2JFMGVq/IIic6Z
+KbdCI8bsIaBjn71VgqZYi7bNQHb/rgtiWuxcg7UKyTkep9whejAUeZ+kHviySMwebkUwRF9S+w0
AGDf+HHf/s+k6QTc9EA/MkDT/kv4XswNIyDhLriklQAnCQ0KMpT37/jHBSPVUlDqfdWEovlhYUav
iBH4s0Uxn+uVPKmgtKbA9cbdMoBjPQzCAWOfSTwpdDqIABq5dxcNzS7Wq1gnDLFR8x1Ot9uH/0Ij
KQoGYcothctxaRYd7e2eCBMaGPWjPfQm/tLYnmp+KmclhyoC2WnL5IZZbITPKCs/bAf9TvdW2oJd
3mCwdS+yRQz3f2SGvDlQRcyNKZNCPg3TWVTtnqBoKgfggydOOLN2QMzS4iKYQRKfnb+OHGOQGvVN
1eks+1LcUTXYE5leg9cqDDm+89nFIZFy4IOn2f42cnN61Hqcu8w+C2FQOIjcnk4ly5cdzUbb9Pfy
NAESin1HRI1SNf+dQelXXPNsxLZWFc3msxGh8xZoIE+gbEIzzmu2eRUmNU2aUUZTW7OTP5KXz0rZ
QUOioDdY8sYH3EN8/XJv1/1ZJd3+jXsjX40ZlqMXe94fiI3J0inXpb9Fuw5I7bzB/A/5WzyvLuIK
U5D8JFCl6D3BqRZPqnWIY7N4V+aeerPVsvsqu4hz91gQJ41S5lOnLYuRSuyLz6JcnqKGeRO/3tfI
S+AJH/8uTfVqEbs7dBmSm23wt3k+9A/KjqMK0lQu7ebOFUUG64xZSayrvTkyx2C8rdsTOYIK9OhJ
0zY8LZIMUEODXEKiAWyPZ0n0K0NfKl0JjOGH/p/Mppi/3sqxsEpuIJeHcNoiosubu3eMkeIE6/oT
R8hEF0BYDK4bvzNgO3KSB/Q0PlHXlzja3QoqyH8AcM0rp24yPd7Cq/BrqRVbFBdngx7VBs47O/p/
8kC6WrddR306zvMbl0TqdXbhathAE7k+TzEgfw9wJpTk1Hh4Mv2Bcbp3Jnmwlw+dYewnaglX/+C6
O6+jl+I8PqBHVE3a034mwCgTcGBgA0kJXchDJo2UPKAB61tvgsckadhcIf3a5HYv9A8mWAxwqn1E
pHWV8N1orseV75D6YaUsFWDlEK31RVwg/l5/iTHktBNRo71Jn9uxJbmeQ8Y1fDaB1hWnaGZnZdoH
6w6elhcV55DQHvAvkQE3fVL/YIgfDVhjsMnEjjskyWU2QJBIoyLkiQFsdhrdiz6LegUxBt6D9lzG
VVsfBp2Gu+Aojju4KYTMfcQ++cNCciPU+s9aAL4MmKbER/nStvbK6eg9WLjoZcDGJgFk6bAU6naO
73ICfKzdgedEGwlAQtd/dSh1uZbMyxCplLbdY2dERXksmUjtvrkRn4Ok89sMzx3QopDob7BACHUG
7itNqrR24yVNe8OfYspUSZVLmmwqFsD+flXhapnfvL++LhT/IfLul6kMwEQYwWfA4yLGapQzo1Zz
j9Q5oTV3ATRMKntIIR9zhcwJSx8w3JqnrLVdzan3QNJ8o/5C1gyVzSh2cz9dYI85yRtD5x3UvDRZ
+INEwPJ2fgymRoz/ra3O9OSubU9H2hAcM18ru64+qhCm52fguUt0N4rfM4MNqewDe4Zvy+FD0js5
bs2bTTq6aX3oUW5Qv3VZ6tAc6DOoGVtcIERF4pDXXEX4HR41Im8BzC/42u5dkdk8/Grd1O5WDHpe
mgRxN2S9pgqqxwlANjNMO26wYpFXC/Kvs8upg2WP19ATP96pIwSlt2pDoY/ZplJJGKthzuhI9T0U
XCv1MC8OCWNXQ8hLWuycmYYrQh1J+rn354lyn3Te2CHRutOxRVeL7E0I/o4DBUETldb6EK12sKZS
OkPHVVtztIuq8r2FE1uH4hzK+D3HXeL0FYQG2AneKskQ65hP/6TftA3eOTHJhccssUjzFhqTyIHZ
zWzDvieTRCTKAuzBcMuvEoU9IQwlH4/3+6qNRTgj+dDzg/fOQQf5LL8+D6amKrXobOvtoUUj6Kd8
nhif9Fz3Gd+uGvO2nVuiMEQIyJjJ77K+uupskQ/vyFr3trvufZaZN2cLYUs+J5LrwkDPmGhEsG6w
kUEQiUsSeFRrpciT20CQVHTuGC4TKoJiv5Qnyy6ZuctFtUsd2BYRJh9CWZPBd2w1SB0Lf+nIGESA
XxiIP5bAt6aFpZy/VD8OgHJaY7I75qOB7oENuTYq2pBPwqbsKa61swpr8yhmYe6hK3iqwf62P8YH
nWmiCafHLfvVNcqIrYnUnv0dkCCvm/sSS3HUnDEVGMMN2rbpCsZ4UY3QL6Z8xo4DX9C7+ilXtyxm
flQT28pWn/rzUywShqP0vq08wb9sSym/uucrKruhNSw6nzZbHLI+Xv/nGM2pL3p3tMGJ+JlBPRtt
vVXThjecjoalbLRLf7jkxjT5+i2SSWsO0EmFhG7vyJOpu8BwgbxMrtTYKPze7pesAXgsIOgrZIgZ
xA5advnIq0a5dYZgIfCZKVteE0CpM3w4VdAcqjkh1x21uCxqqepkEfFbvskqpKW+3HD7BD/YCkJY
lOvr1M6f+FmBi4l+DDmfh+Ktc2Jxy5bAyP1B+Mp8FK8WrrKI05WtvGL4okztxOxWiM/CesOmM1l9
f010ymp352TJfLQCIOjj1fxKzRRY00VrEFOwyL2pL/28RppkqTy9+3tdnr4ec3G/uWohajY6Bhxe
xhxExVWTTTn37QXn5LEUaDhmELK7cZsvMCCreuF6tD1yElB5oaM5YvLLbnfIznrA3OpyN3zHZVWG
8iVh1X4oA+q4q/Edvd7E2kyDsgwxv+/u0YvHcDAeTmvzLoHGk+/K9kA0l614Q71fNcgWjsklvovf
SeVKdJRpL6WXgfzGxIBxT3hpwu8jfwIIni52UCKDSTZH4p3b5iNhRJryIWlWxqaS735dVCoetlyr
RPljdtAxLh8Q2KKuaNeBYyAOgPN9xSZ5lz5a/QkcOBtDuEaQ7Qpb1q0JjKXcvqYqv6HpnIQxDApA
H1wBMGXOH4QBKhH8eXyJz2bexBrIEyMlsuj3Ny3CRKSvbNekIC7r7sVzsCIV1Xx3D4Fgxq8dcwCQ
FHs3Jp4l54F+elCIJrgxKjdvmTIc0lxFHRCCkenx3kccQnXvpbaw8DI46hlruKqB5W143Fb99tyS
s5pwRw3boQpPNA+d3ZY68Rp/hNE3JihekqeTpctU9o1yvKKJHN0UiUslIm4zrx1XwLyejN/6kFeQ
EfP0Id+BJ3IhnMxKVIMseDQdA1pOE3NXWNbsVX5yzsnCzbK5GvXDr3wHZMl8RB5qYrL7TSiJYmYt
DrG3JXvPEj2MS4A7coc4SUdx0xofLyqIVoW1mdxLiPYZZoCgPLVGb6J+SmFtuSdmZ6+Kl8O3QsFG
z7mQwFOveBSnRFeOVAaBTFc11whx7J3NxJZ0oLumTc6egzWq2NNudK+O+kGEyHwNyeAaW/GgDBHI
DKgOVok2+mWV51kq4IrdWN+VQpU700VqKogODT5a7y1mKy8663rfRW+e1I1tSvRMsgwsU4SlQ5U5
djcNZNQsGFCdq8BtrL+xMp2BtBGqI34vy2v/EWGmgM035FgAc7+x3OlGXjMCe8CzLNCp5SoT6nsl
byRBFfiyuGuP9aUQkl9gMkD0pPeaRThrNqWO2FDKf/jRJ3M9wUcPGW0rYWY5Tffja0nbM80C+7FS
6QzO87VaO51wcOspsszE5ne4QRWlfVqiJGrN/K038OorzBLH2Ecv6tEFZSA2+0HAZIoyzwH4zFz/
lItsg6o4pPfClc+52NClJ5eRdwYHfWMmjUMldinBP2Mdi8Vq642gyEGbxnH4Ue3jCBJne22jRHkd
p9Na2f1cZph8rk8KKxyExRvgJ5HhMhHCCGHab5kigbchtRBzuOU7itLBNkt9CxRk+C+bRQmEEWpV
TlPxgWghsUnEIvmZKhNvtn98fEbrVLd3w+8mkREVVUuE9vB3Y9bFwrqApdSdh1y7lDqZibxV4h9H
7E6PXcmYraIffJ7x0rtA31NgkD+bZRiPx7DXzIBSoGa1Xm+kgv30I0IybA2OkwOsEK//0M2Ya76q
dcaci82Kehi8EurvtJE1ja9EMYH8pXY3DZcDQ+sTqpVXkq/WK3Q+QzWl/wsV7JwBv9iRkvyk736y
SPVVpuGEjLyv7mcOtnqe6eBhLcgfDTAyTyRX/h5bb/PPh696RJTB/CfgIP9NrOs9WY6Ly2IeBMXW
qAXP64TnawDnxOzn7G5XcxSh+fAkilovpqSmDuBgGbHfHux/WqYFFbWZg2/TGeUpm2b/3t7CGfAu
UrEEfaveWjB6C0jepBU2F4JXJ7bzljkcXTag8i/Hk9lwUNEtIfBn9gBlH10EONR6O+ABM/+3eqiG
qoADaT3N5B90P/MEYMPK/BnTfPeUllo6JJ4vDMirWmg1uR0uANSW/qsgAkJQd1EekOvGfWZBRzP+
oFB8MKR4NGc3wuKu9t1Zk+26ghjk8M5SUuZr0XTW7VdJStWVDB7Cm7ihJQIbFK2iS6gJKpr3gx1K
gX97vrQDi61wEzrpLoskIucxYHYxdd6gU3inXIdegwsTs5UuLLOMhk+SLxn/wVjfCgkeS+Xs0KVa
DX67BRscztt7yBKPzkxn/RfJ40vS0hyGWLxruRUkKBw9rfbJo+E0apn6OLYdiceV3lTC4jTr/TNX
yBzV+ajQmfWbG+O5iC/T/hCOqNeCogoe1U7/SFCSB2VoS59KgStXqMVmikUajhmRCVoldPV7C4Ek
gi8M9+uUJ7tAHTdkNTKuWkQtnYMnuoMxv1DuP78c9ANV6unN0qO63haFSkL5QnR4t+1geVg3bk6K
h42GXi1G5K+oYOKTruTo0VznQ0mHA6ezGUBSau1VeV/KILTkluyZGYhx+MuHDUY+bWy86DHTUHEv
CDz+Yd4QOMAZwWztB4slreFzokUO20qV/CatlOuSx08HfNOltIdZfaBKkv4osE8BE56QWX5gnDXX
iK9X/wFmTDxUp7Mg6wC/ck2jPD6VPmUeWktqTdic+xjkVLRyYifBiBrxSalYA1a+rwsK1bhM4e74
l9uxqA745uF9xM/q0yLfdI6l3ejqCKeXfwvqUiVWW6YAWWR8ISkvgDnwtfMNkYu3hYggJEuZdS2i
j4/fm4N1ePREO1uDuTLQ3zSR3WZsw3Ypjce+9msYRbrhTwI3NoRq9NC3GPGZLssdm3qNlBqF3RUA
smFqznmoLHUZkjSw/zV/oyTZIUAzzSMPNXiT2VpWirIz3Lha+qSr/dZDo5ShgghQ+bbgfhcUqYrS
C22i2CwZ8rBPIgyjzjajRoGLDAdwkdPprM0vzlgy/soF+zYq2faqxJ7/0cpceUuE/eWY6Eh2GKTJ
HmDDguY7+isL1CyxW+WDZjMuLU1YY8LtMnKz/WRu+izFhbCcsxKxXtoLD8SAzXHkJ2J9TN8T69Af
KJnaTRcZ993WMEpIijqZ4wR5Ad6LYSilfiuo1X+5W1CenIy2ohhQ0QGQj0Jo0uHmGEnwZHmTqb2t
p95UsaK6W+uoCVRrjeg5p25Umq6fo0VHFNdwNtlQd1gZl7YYqmaOO77HLhhcGaM8JL4EE6P1TChy
XwpsonqRc+GnImFsV7+6IEXvAdeU8pvpWyArxz3YVWbZs5lF8XLSv3eA/S2R9+zbjRpKkVhGHaDn
IQPS6WbOcIrscoUwewpukf5Nd6xfklOqcZgBi2QTTHX91pnC3wZAH9xDkc7FABFcSA3i5ZquiaCj
u+VQv/X1WUHd2ZQwxSyShdHPyy7W7Kgonm5ZGV4JKzWRRMgtcUe1uyouq7dNAczyGNSrAGQUnXzh
ZyFgqiEReJWadZmnbnrHU1TcGyoDSW6ZsOs4zHjnrBLEQ900NVCnU7tzfVx0hEETBXUH1z12WAZt
uDOUNaHpIFB++Nas5DRorH7/kWbPf4DUAKae8m5RWh8IbJfNTCOl9kInDwcY6hcJeP5rHlEG2lch
U+3QQvnQYVpvf0WG21bXX11VpbxtOayns2qfyUCfsw5DnsXbHCR7OcPm3CEJOzR5ijr86AsJ9mIe
h5sg9HOoHZvBYouafldBiKWJRwS2UPtrOUp08UdVgkyGih1eOmXrPtd0eHWK7ByI1F8thCURU90c
b8Yv+BYR6L+CeZ5rpIPjpnzM/lnUBZTe9pDZylzFjSK0yv+UcYkS7/NtaTm09CZbCdEjBQeKxfeY
f6XpktPAgiKKBKXJojX+OmLmvoAxx7657d3SaRZnWO6X3cePy7+4/Kdn4jvdkrWWRg8t3JMbNSci
kvXUkup65oYj7TazArET7guQqOuZ1ekPKkMRs9W21UWcHixdeEn3/1vuU6T/h97mI7ltJ1v2Ql1d
V6XkdlBBUqW9x6R8zNZevTNxFfuDRxNVkDXQPRguebzteo5Zxl0JY+MDFPUwst2raVlyoM3Kz5mA
zMnBzjYQWoVhVeTiKIEyteXH2RitmXHmDn7GrJP8AXKrDpu8hL3IkZyl2RDi12EGv1IJQ+tDAUnK
QK+A+DBGWX5WYWY8VXIDB8i1ads0z3vJzcAcRTyZfbM5xuUcMM39QEedCkFVsOprKxq+EXn7ZLBj
JY0GGG+awk38eC5KT28bu8o5yTG8OJkdemybBccZKEMHh7cyHkn7QpTXEL1T1MfDNg9hjgtz4we4
Qbm6yI7Qc9tNZyCJ08HYmuQ+9jAKFSHdRQHnZYzcKTkenOlP9mIy+zUsCY2nc4TjYqJTT2WvwAZ6
1mhI/XTz6wJhe8IwkjMebr7yQ2ILwlqHi/NCdW7yPmeuTM8QJO30Jakm+Y1vcM/2mQsEwIRY78Ke
VzYbGpg9AcMSxYLtiotLAsg2/n8/ZOUnqJKJswaQGIY6ZE5wqv/ZACXhow6DFLr1MTm6ShS27VLB
AorjiiPPcYTtAp8xT4iNs650M2cFNMePP8jtfZdOT7nZytjWZVYcJ9DePguIv22VnW44ZbWPXP/2
hSbb8xl3yDm2BOPOSi3ohDxCx/1k+jVX6syQD+ZwqnIEGkFqThoxanNfA9ZL1dJYOpK66u2tCMOB
lAjjk7YlYKwwchob5+SNgpMzTmlPY3cFAKWxNvV2+Kne/lbYqHQm3yLgIQ8m3TqN6mqra7HcglEl
JorOCmha3jRJrURDIebZGb0jDwXBZSVCI08u1rYlHS6Ugs0YAINi7+32XrqK/LRJcIlTfuB9P3oe
5g/PLqDOyNLhVwJ9I1S+S7VoWEa6Jeeb2cOF5fQ4mNi3WXEITi5B4wEG6cfayGDJFArI9GqWohPQ
wEr56eSorGlaBdZ5SOuwPO9SBifwM5zABEsa9ysHMCpDBa2Ri65rRnJIfaWQpsUuLOpDRGXet88Z
4v4OTQ/vAyZwJ89r9jy3KJp/Qeg9LtxGtESR71CoxEkLt2uXU2Y/RC8ihn/dPzBRR9j2OU+fYZEx
b1nJ4n5LSScjMUryroU//1KH1PXXXzbaRsS0uqt5mxxsVFGHdkW9TfqaPE52Jo+tm1I7zVGyDJvO
JKCk5NWUY+E1nYRPg7jj1wqFkxS2EDgnzR61k+ZVGSM5rw82MR9fHgRF6VOWLjOqawW1UmovYn3s
z2vNqtjMRyLW0Kz9GbVwt33ICn8i3LqBN3NBJOTbGYVxLL2qAGXlKXwjD2JFM4CYfm926zQgdl1G
3g2u03RnfadYHhoT8FgFIWrOUL+9vMXIpFc8rgFNKX7I+QNTdmNEYHpypr8MBqxVjkyUSd8cI33O
HxcgViqrLVxH7P+erLRFFMRobP9cG1cwz5IUnBv7UuK9zQGsKjyoRmpsGeLyMpf3iFwiMDoj+1g+
yEmvmiZQ7Y/CDVgApUCJcthiaZRakqyQY+2l36M5tVDsZOSwfaiKyF7ZZbQ/RnscKHnLzuFY1++A
56KOLjJpHsL5i8hVjyfiPCibLZNUeU/tqqLaKigQQpuztqqrdk7aGGZJWvt0D3UyWMTUcvH9vrx0
/Z1FbganP7vLM/4VEQmi5aaGfZXZKGFQQY4nnMIijTAKcVU1hgg102tc+BvsJB9kpLvdPV8d4U7p
J1LrGGACs2DDeIJF4y5COpYgn7iJCllmXL5zfZbbGM30SuucoOw5zKVOEoySSO5N7I1Tsw9QoE09
IJO9kUxQRh76ubueTnQiocT72pp+eHtefox0yKpE4hG/YJnpPf5oarTJyjEyDQHbdRvAJ7ofhw+W
eOmi2nrjyGXPN+4H1CjAvwi0wetKk/1z1np/u3IutWFrKsQt0uaJ6UbifSRaBF1guGVoDmkhkUby
C0PLpX+Q0UT75yQZ1I3F2kZ1o9qg94fV2rbeO23kNxVYhADzIMml1rALLeFyYiia1jXyq3JHpEZU
JHFqoz3fYSI23xCmEsUxAVagEDEXtOliX/m8hP+vT2jI3e3GFF7PA4DfI94ZC5arL9fKP4+33Tt+
EEeP4GlRSu3/aVVDthkSKQGxbcy7qiMbz8ngbAT8+xha1LZUBkVsuA+oOOpjQua/0dUD0Nzm1k6b
6pStnh6Fh7lxGFWqdoCGvzx6NM7BowsuHjtcRb7U6Ys+TvDmeYMF5+FZr9jlkp3PcT4cmpqQtznt
52rlopop7cEB6xSk1sIEYAiwaxsmyha51VRfhqW9Hq6lofufpZMbSqX0O77dCQAnjo2RVOdDv6b8
A5Eo6SlXjLwBTfq4/cXT6UIJS6BWEfbWIiIpcyonUZ0Wzak4/UA1pSDjw/eyaPpdmHMH/7V8tvL5
GFmixiVINN/NgVyNS/Cn83Q7mO2jRAWe+Ksv+nAeqFRxM93+wk5L4CJFxiL6b1QtkzBSk/ZgyODf
yxIQKbGMJQLUK0nyBOohDpjUAE/tH2BXZt4EYf9CwaGNYBkERNlF1jbWtI8fwHHlldPetK7OoGWb
BTdJFZcQ8wDKiVJnlJ0CeGBd/55LajYeZZJaAlLjc+WQThzMSe3nyib/bFUDGgkas+fEPprI70wg
PGve5aodV69vUgbqKfz95cCl37WaFhqShsANDtTN76tTrHNe4o2uuHAr6VqaMxNt90xaPbzin0NS
5MhXdhKVKxNzZ/JAk5Hv/IoJiw3XBYGACuA4gaVQapxucicpVHb4FLSQL3xNM/66UDYnWQEX8Soy
WTXdayZi77yrtpYtVEZknSN7qc2BqqFI8XGrLp1h/SNweaKxVmKYsfNt3uUo9wRiJkYrhIyC2f5H
R/i/Odbz1/Tn1po3nPY43U81QDdBH1prBZzzAsnewO/1E8AQsJ2EfS95aVt4FlA/+pwQEeWPVgyX
DOC2fWi0ngwrj7e3B1zVrWFjHtCOObUjIkO16UmEcq68zUVbRgxJ457HJOAWI4lHWSnFUjOziCPB
HlDe59Q0K8AtYLO5Sy8RVF9oc7GESVhrC/lvlpL1AwQHmU096eqEKqLC/h+jFyshbgZBtdctghr2
TdBYR/8yiS4V8/BFvTYBcau4NwyFAFfVmS713QbJKbxzVBQzBRKS7S10jfn+RJUKF4iOnwe940H5
OsWlEABxd/nhbJVU17Xna4nqtFGI/OazRyv1amcplitROY3AuS/cvGeGhDe7Th7h4S/6N2IW+ez9
UW2GavRaolFftORrolKxnINDTNCzlMOLn4/VwM1KVZqbyi/TSNou0oZOLIZw4EEtLVCrt4VAJ4aj
GUNGlbKNkdCdAnXQW5OQkJ9VefAH2jappo2s2JkL1X1L9qKLFMeNywiA4wMi1bczYQGEROWzV6GR
ycRmTMHz0Sqt6WGp/q0y6PmZGc/pyX/Sl8yC8DeyHb8bU2ImCcpmRZLDvKEP/PrFS8v3E16O5e8j
WD5D46M5KpMHcxP/pmOb2qWCBXPVKepvDwtFK5akDE3Jl+Ff4whrQKH0RUg+JWW2gt5vOzJBoZ70
Uv539KPK1gTSuve80J78dPRWshewkRN9MZ8qSrgPRWD7gpkSk2vKgHNJGsgX5NaXO0pPr2wEReTp
EfEQD1u1sd3CSkQagL6mZzdxXXZf94sZJ00sHPuX25uvwWAJjCP3nlr9LGea99PmvnO4gEFaHNa8
Xb+oWNL+uId1l+jDscryTpBlfHC/raazH4xDY+VtLjVYqgtEdnP8DrUnN0D9Ez3IOIVicXJuthXx
kaSBBs9RullC36GVeAS1IW2xAqtQ8sKNvEF9CHUyqwubkZfExCh0kslouwOus2s0G59jgd9i3qzi
GGwGIG02oN8YjPML1RpL7vyupkGFmPlWK1KkMWUrKKnHmI2pX8801OxKfAfeKyvuG8mUQzSiYeuQ
2mVLQ0XvY2oslHGsE75OFg0lf5TyZPCgIke71xworfowYZx2Ufric0kkf8B9SJEULt5DC+nnBdgM
gtCnWzwwWNtRRsh0oBXL9q7wXqyQwE8t/NQms6auOaqNJeyUDrUu0PcQfnhp1YlLXr7U/Dkf9EVZ
X/yD9gLfkJ8OJHQiipWmNvLLAc+nE+AGlccADJ7iSRwLsYfemPaQBW/E5Wu2PHtN52JbCJNk0CbO
Ue/YdfNDjWcIAlRBgEWKezruoCfyon05hP5kxdTa48EvjfaEJCaSF0e45qoCdaMgVXrGLhNauMkL
UVeslneeNFfe9V9m8BeBX5WOxdZkWllTdhe+vGCPCPL9dfDfr6VFoHhwKTSHLNU/CBu1DHDP5FUw
Lnuk/b0LbddKHgP36HO3yS8+VHhqeIyBsQ58f7Mmiuh4kY979Qu5ph4pGD1ljp0sHIpY0Uu5JICv
o7pIvJ0AUvwhigr9Gvtv8ucPmWNryr18mU5/YIPjYxb3YHMMjQh+XAbVkqMc0G/sJvy+BdlPWWaG
W7HgY0xKBEDA/PgguESyA2yDBlXJj5zRG+/BvcPyFG47+R1fCfsKY6zADGJdWB6jKAh7W4zuMx31
Qx4ZpA3HJQF4hfB1ro2mlgsZ3UCjGZh1C3m5KqrLOm3XaLe4g4r7QxbNW/QlZlJ6lAqFeNqxrRUB
oxekaOZWTh8/GAQewXiyry9yo/fMsdQ2aEjgDduSxU8GVRcavXB4c1ZJv6ePIZAAFI8WF3fvWXsV
jB95ZoqS3gC4c1qVdjuq7IGTDK18/Fx0BZbkK91lFMEQZcHfF05IgZ2v8hfWN+ZMMOyEHJIeGXLu
iFAxxtYvCW5q/0cmGN3nXSkbj71qCgpe9xYe1On35bEdBDSrp2J//x4Sgd3YfC0CcFaF4IA42XXI
NqV0jMwPHIPARhnFJf8Xqm2IqiSdkHiXK+qXhOv1WeqG2VyvzKFIvWrFfWbHGeQzPj0FhT2Yotnl
xGMqTmZZg5HLlGBimb2JcTfzesDRj0xVwOWKvRLCArtf219nnP73xmGhPkPie4tdJBgtIvjI5Byk
ktAvJPkZKi1X3M8WQHIITSkZwdlae7TwB2B7uGhF3SNml4Px+oHwsKK6XZeisvmWOmLgRnRUmN/Y
IkOpY/5aLlfofuEF3ECfb5etPnQXR9orpjVv+ygT9U30pU9CuXG2yefI37GgWDSkbCtvnrrvc/dx
DNlhdi46Ml8oaB5PAnSwCmZnkIAA2XapIChnlIj39qRTo+Q0V+Dg32q28VdADYSWaIEQTPyi1Lef
pztwRXiil2fvk70l2bab7aO6mpSWITPZKxgCoDqGHwkQyckmMs1bjjDzr2NwZ2y41BWvOXtX1AYx
tE+hCPIqtqyQGrzjqHunjEujxN9Fd3g5aITdmwWgVrVRckzKivVRaONmkBh0b3+UVHdqwUGp0T6S
6ZE+OQbT4gR5J9wmNKwyDHIPpWf4ixj0atppGDqJYBKLle+1akKKCmaUDOPFHYPFWAFmroSXRMYx
IMlua4P5v5aFW5WeD1u7Kg1v6iBy5AuvIrGth/C9mKoCG3Q6udT7xTfwcZ5A6kUIyrejXQ/IzX4u
lMo+UpWPp+PmDUZtyej+nXLT+mTEbDVgwO+ek/6R/COXlYG9Kuq4+dO3WX9euaOHwbzwt4CmZlcZ
kXPS3imdd7VFN2VduSyDT8x0FiZUHPB5k+yr3Jwzlpbfup6bUclUYPqU9fgRKRA4H4jhaGRDUwMo
IvM3eHUMLkOIX5hRm54N5Y2UYJuD7Va/yhcmDe+6Vxd9ngfbXH00BXxk5Th5Xw4Olapn+DWyhwsD
gB1gYk9LVTgyR/e5JRJ2yjOLjmp8k3s3j/1f6UuXYp10IpsSynXtpV2NGYLh5pkdpPkLDMpKnl2S
/9e8mgRm2HVqQ/xz3syFhDvHpN8zcAeSxuSLSYj8UwMOUxgulHxJ2K7isR6lu3RWmnqYduI/+9rD
5e30lvNZCxSiIeEQEzdghfHHKrTv5lDDQSQvmPKEdscNggPYSdKCsWQMePTF6HPXORnnvylsPT+m
P/ofknvdU89iUmQNK/4/6hu5NQy18obcnSyXfmohA6AFa0q6OOZQhZZ87hr6eQErScznsm4yPagK
j/nZOK1GYHMdbU8YN5+XLe1OT3K8FTel7tLN0elTihfruHfliEZmeMcA6z1vsz0TT2BWzTTiHgy8
BxEv88K1AjUxlH6c8tmhJvtP9EmCIi79FlEvOUylfz1ZRkKvw7bFjuzslbs6Yp9MhaeFP7a0zXsX
wmp7Kk9M0d2+yU6ToL0QRhrb5Fn46Feci9GYb+W4VWSKaoWJEoN2QhuvcTLUIv3qC01Cd7dubOjc
YQBlureeY934kQPo41w2aTjLZQeg4bv8AVbOBOqn3VYsMVzqofLY+UBs5KU4EGyYAXYwZcJAnMbk
04bPEj4VrrGeCe+rxRLxbBCsBBY8ku2OFg4FtudmTK9JCXd6u4KMmDoer1NC40L6fCCE1oVAO36p
Cuf1eoh8FiAiPHzU6oGRGXvTbA08LHgGeuHX8fh74YZiPmDbqOtGNuTRr5YnZUVelgo7VdjZP/Ja
Ej+fqXGgS9Hp3cn/xsRJ4V2wdINBktGCZKsqXFZXdIqt8+1RpxdixCbLRhcAVpU7Co/aqjIdMdG9
puvsrumB8vxnUWwISJlUDsOeuLKDfWlUzh2ru3OVvc9RyRTK62uvIzSxcIHd770mYk/axP77yhRk
KEyDhHojUeLYudlS7rl1cPhcDNSX7MbrRUasI+Zw8PjPAZ6c1hT3mmm6qYVOf3P1fK7ZlB1t217H
trziydcwyFpxnzINiUf2kbBhKET1vnIkkpagCMjX6BEJAFRxTfCW3LNhHmtRM5fNIGEf5i00ULkc
dz9hLTWZM2za6bNz57vWMRqYkFtMCHcEtTMA8cdXyqGg3paoKD/V5F296p5RV5u+pBpRqf52rru7
U5RKZazAKYbn91xXk9z6l/ZDb6QGzCGWp1yAJYzxn3VV0i0XvbksPx2mYu4tmkp6QdfGTtG/1kxH
TwfON+KqL/6ZbOkSvUHZhNIhUVlFcdK4ux1wZCg2JdQ2QAk2XtTFCJKToWZEZrIxtWttip5tys40
1f02jyGM44z3vljE21l2n0NFun8njop4DAZAyEBZ30eUEf/752RnHyWH2EnS3uNxMGlZ2wk+Ysgg
A9GACVT/er/J5zChXxVCKxqgtMN4c7RExQlzWeJbeVOxEZgTdXn8dY1vp2TCI++k5aKE8UxHD4Ns
ZXo/vaYgBQ2n6xY7M2kmKl26hGS0EZnOdJrd8CkdQz7bw2XIEgS6PoqpxOJeF/0PFEybAkQdjmvm
5GXozqCC/WgkntXdkeSPeSARYch9bNfd0Jx1ZBT3NPXNR3rjgicQ0pYDJJjCwDGUom5UtGge6rod
MCf8bGUNOkbtydp/jAiKQrCx0WSEd+VKS/y1Ai9IcYtH4EuZmF8gzzQX5agQJR4AC2tp9r776jnw
3/HruZKk7r8IMGeDn4FuV4yaS981hs1q8gjhX3JQyvAnIz7ObwaWUBGj+QqZo0TWoo7Hh2hK70g8
6n+66wf8ADj6JuqbIvt+wQeqO84ygDTSotHCYy4h0tiek/KsSpFuJyPT/dZonCHkzvQ8Ipb6Fsvb
XKUmloC6W5Meu5rayJY2Bjbwqnx0IPCJYKyyw7fd8qVYFpk4h4nKmrKxJp/y7Zc/R9S1jrSpbHQF
XhiMlFO7tIPM0DEPuJzftyii3K4zvPl8q3H7g+tnsZMNCQyminpRSH3ktcg4t2Iv9klxB5fX1cY7
+2W/pg48CsoVvH3t1K4pngIU2LnjnaM75MbNfr6zJCRU1DX/0EhApjtdZJDQMftFLxt4Totg8jlj
kBa0mAhgUKfoQABME1sGBxwNxm61bYZCjdcMjLaZg/5oy2tOqgk4K+8NEa1ZgPgdLEVzryJYUVak
e125d9LcUH7yQXHWxarFcMdpmcDaabEmGa5pqvU+tHMwj76gh/osXz3YY4ic+UCkQ8bCXHVrAKZq
mMaDllRhqlavt4Lpzau5WDhyDD5iA56uzyS9ALik1vpE/EDnd+iYbCSDN9T5+lgYUrHRe5CexL+t
MpFtn6M866eKVtCe19ry+CFbdxJyUuNXM3I+lKbfnIdu/pTBEEL2oidGaP+oOK+BGmIuOs7EO1VD
5CPBbiukB+LNLHlymGjzux1Dq+PADERwwbiCDKtIMhtF6aM6Fc5iFkEtmWdPZ/W2+VGBNQZzm1m6
NOaRkSlYlWpSPScE+II/JqW30rx1/HcGcABdrd9KagRpwM4OU6a05NVFLK1EJ4eL7FnnpCuBHBoF
Cl1ZpL1foyCawYixLQf1i968iOdWrOSVg6Y40ObqSwj1Myhkg0poytbjU19ov5/iXWYNDXj4408J
VOiUv2mtYWRJmuUtN4I9+jrvlVvR+FVw/y3+kGe0JCCriuL07zpWE9lWqC6cG8ONlm34iv0kBV/m
x7WWomhE9mhRXcgA1LT0KU45v+/4nvlyEP8b+lIeG4jX5aosp/4AmQ51NSj54JHhEm1alWtwnQ4R
LEpbGXf7Ct5zrWRLjAAEG64o6kwMywMbrTB85pftUtM6dcueRC/OpucgdZcLdbIrQhfZsdAtsvc2
Ucif5hu/0uC5l2OC9VIt0uT+ZKQ4HipJDVTLubPeKhCBh1Eifbhuh0a8N2H1VsN/6ua2YH3d3hEa
umHY95KVVQUUif7sJRdXdAdZkJCxvQhMXUBjeQMZiZ7E0Pi/09e2KbIoVLMxQazHZ0pdI+V8EjAH
9TNnqAmzWt9HJ/yrycXaoHC1pTu7SnUzUDzVL/lVRMJ4EFl0w9Ieg3jdY/6FdyKgxjrqTra4KzJz
gahDzQtMi0c1mz1CiWbFkdWi1oKXs8ZQ5rmvTF8vBJ+snndg38mLqkK4LOp9v1GbhBSy/DucI7s6
SMCKvtXsmM2Qi4p3Tt6WbzXrF61pgy8C5lyRiBm/a6jZfHE3RCSyH+hdnGVjWii7nNEKdjmrNXiE
hp7oRA2xQXkvnlK6+7MVcnsVsLlskZyZtEPvXRPyeiQ5inp+ysZIiSFhMo4gU6lWBX2lu3oRYtdL
1/BSKcQPqEn05eb7sUUeUG0TmwbOuVIbtfTlzfjS8KC/gVXFooWmHCLKkzYeRQ6VKx5EXYED2gbr
7FyAZW80Y8g5v6/i4qrVQLvBhVuxdVHnv78TPk2uzxcutulHpM6xVNQnmtextoayIlsJK48TuOEp
tt7yIp3ACFQAett29wlu/K8Y4nrPKT0zLrENbCoU+rDI29/8/46ZT4TY9wijFrNhuOcFyNam3O31
HGSzgcNdLyUeitLhiuPKcL+o+v1/c6gq/4zvltrQqRzN6L49FrZuJPz7HVTbrufG9sxXdDXjru+K
s/D03VDJhL41NwY09w9c5Rk+mG2+G5jgHA+pwrZICt5QKwefjESldktJBv3+DKumJzWKCKWzYPCs
u0EsjiHJUfx48DzY+GAF4PNZnGyBSHvVK1I0lt///MOp+deZI0kkbfOKK18jgbtmbdfWSFTMLKte
FQwbXZiXVz+/EqJFkX4HXNt4RQtoRoJl6sXT8gSnH6dW/BT1yFZcYLBmfEsFuZXZ+OogWRGHVBen
j0ZFb9HDh0uc/gZhE5LUa+vMDRVjlzMTEs5oWLqxhdvsFufJU/eQFZMe9XFvW0QTswLoqWuBczb0
2C+LF5MMplEKAsjREHvn9LWyToy5xHtwKMg4x8PGReHC6G2zmScfCjQ93ORugqThsNsBgMCS5UdE
wnA+xcuMRgqkteK3xD4kwmk9qWXUJS/2HBNkGoBO8qBflfx6Fh6jSrHCMMw+0wFTiFT+4flIvi9D
nDr2pCoVJ5GekfUPh/nBlhDWuzu7biU2kd/G5AYP+CKlafc8drtA7DvggmmkgmvsUkULotVh4vkZ
GZO/F23lF7xcCIWPLzh5ydzoqQ2p9obqmRRwiSB4nB8KmKGMJQOxZBjfIOLuE8XGFbOn71E1IweO
okU0sUgO+VzRqI5z/BY2r+22EXGtTX7TXYzJGwPCWc+sex6C9ZEy5elBNy3qmx6t9gHvZoA3csvR
pjtt4HF3A4xKHJQr0G47V/zXEeWQ3IjgEB2OeX+pTXdWa9fmKhN+iIb4iCud3kfeJKiPjtTtsKIY
qdyuyzA2qfY2k7LtOh2HVV9nGViw/rbaV9MZyP9Tcfy1jhRXhyP6/qU6LZbC8PsaXkgo+xj3LOqd
rIYjmmLy/wJ+yqGRWtjGeXWjTU2eHf6Sc8K0tyJPIzqTM7o3wqPibc0Ym2UnH6xLthTVfm5NPMqW
umoQvqIAyMh/mJD3D+RTAEWF8FeE8XheWaHFOAsyleYH1ndpj4fTiB7Tl9+sWOs0wKL6+uPI08VR
J9NEDGndSJuZTBYriT1PSepoIJjCgaMPwSRjiWhhzbt2T3sEVWkrm3oZEs9GOeid3+srb6wt5IPo
PCMSQYrRHwB3UUPNveJHUwNCU28saY4r7Lkrpm0Ny2oFIBc8APvyjxmDSmKdiuRY/nJ2MGXPySbf
F9nI1+CqNvUC+gvIpgHPtUbingWvbs9fcsJ5n/jGPetbpexJ56mPl5erDQyM4MJSdjlKcvWheo8X
aXWOFUC0ZJxSDj+rtS1oj0d4Qkw1WP1GiTAyvEcF8UxchxSfbSTVnN9PPVX9KUVsYRCoBTbp6RWc
7GmXea0eKQIkoHDUGv3uFchZhshJtAKXJjwSlXuYD7vNwkXFznqCj3CcbaYTf5aDw502SJWRxU3J
U1UrTh6hXcqCRjjbYr+ZCSGpbmyNQ1Mt6FkH87L60/EB2kYk2KCOK9l1qw2eEy9XQ/rjNK/iAWA0
e1l9EftBlemwH2SUbog3ufS13qwAqYLGUyDfTMnjIps5JfJrzxVvyIekDg+BSYfMvXlidRFq+H7Y
7Oq/4PMqPqOxc6chZZwGpYpqgnwPR+cP3LfOzxE8H0TtB486dYnbeITRVee6RU5vIUchyhoCEuFu
K3RWvNpGavWfoeWAK7fOP/jr0axujSOg3Zzlz17sT5xtgpi5mWcGjJV37WplWIJc4YPT6EIpuvs4
UL1M2Ca3qnCoyXZGtBFahn11r7zRnKvnz7KnbP/Y3L2kJ2x9PYyoU9eeesZWQhN5CttCDnSRl2c3
8lLfsdJ7HHDJtfSbNkfFQeZ5yrOf2sdLSLAxzg63wj3XSmJYBzFXvy2ootcHOutlrYTk0WH1PIuk
WQHiIy3O3g/Lwj9OZ+xa0DuV19W+irdGapfAPu7KGEpiVgW3O6lfo2U+MHqpJXzDGKXLnHIFplHg
cbvSsNhqd1ZLVg62YO4LrZiNKHlD3jtYMDmB7uTu5MuOZe+P5e1uQErE4RFLVp/81Y5z68mw+TRs
VDCYPZdDbdeY6kSfiqg0znKhkHR7S3SZNaZF3BMzpDEEFH11uoltG6o66I4hpvF56oCJY3yDnyw5
mAbmE+UdVK4eZ/Fks8Ovrt/d3NUPXnNHt2qOq58TF81q9mgcguS1W2glnS48Gx8L/QFOK1tjxgQJ
/VugEw6+fZH6lZhn8EE8JsV4WGf1mzv2Ii1/IUM8d8oshonAXmrmDL8STMYDumj6xnHnjNilptFL
4LJz7xkc715GtodZkH5m/kfyEWUIHPWLR0izQW2Y1u11TaRgOgIIfz8eg0zfFDzVpQfIdgaxr6M+
2damqxXInWGZjifpzxTM2rnaJ/MiuLmpRGpXWbc07U4G0KO5LVJm3t9pIQW0YfMeXKl+5Tg2m8Mt
X4vlvQsMtxHEIHjLWT4nFCvD34ZDn3lYGx7Hxt38WJrlHaeyjaQGH1nMkEqGmtcpodnT3GOlSidm
iXlo27Kox8XW+8YagnNDSW8DvZT28+0cSbL+BeIUweEVenogRM7QDC1tlB/rV/ankFwpb76lfR6G
HrmU0UkArto8EXgrsjWrVQH9uLvQQIVsJvE1jPjnDX/6S501TBBTnPJzREWjvR5bK+jHtejzMGF9
pjXUrsSl0+ymyuRz11MR0lb63IlXUmkd0WTj3/GTr762QTPhH9nIwq5X2bZ+SYJOQNS1j7Q1kauk
IUsI2+Mt7KWovJST/3Pe507hCXvBWdD3gDGUMWIoXsW05eJNLz084ziv16pYwZkpoUb4co5a7G2/
KZDyUY4ETxCi2O3si1PVmg8xJnDfZ9DZjKYJf2UsyJazCmvV86/oh+QNCIoDEGhPxUCYbmVQWG/a
MSh976+c8dCwlr+TfyBTmAB149IKydcqY5lj4QcCEqeOVtDOQbD+vP10ldygrSlZIt2jOvWnkPDw
UlSCPT2A3hMjf/uvtqZhbtKhdKeNMiGW/WDz0oAEZaAxSFKDoj4dzrgtLMakR7yJltj/Rfam+BWS
Jm31VQnbn1e5i4J4j9KpipS819We5y+dGIfIEHIN3MCfsHug5YqeBRgMkEMgvGk9+Xy/1Wp0KInh
V1RE1m5kBHBNhwuaoabaFNo5uECyfcs0Yr2fHe6VlpABJMVlr+1YbZpwPFYkHXy46iorwNf2zOHW
PmcYxCdDpdcH3+L86/igK1c2eVqtvfx71nkEmZ0MHqGMnYmsd2iLJRdO1zUy3NSgzHC7o3//J3Vh
QdaeNcjF5mMq84k/U1usW6XrdMICdv8WZtB/jNZjUYCx4pTijD6Wlshb8Cdu+F8eqii3DKTMIhyq
LRUADq5/mwGv/BLsLH2DVn+T5UOA0GhpmUb1oX2dUusBJJG+MgZvm57MgFlnm0ZXWHFDE9cjQIpw
97SIvO1i4MR1XhRPpbzfKsFq9D7+uyyZ1FAypELxL0h7UmUDFXzSkdgOVWouCaFyvE4k855GeEvu
X0muBEWEPNBxQe8S/kvuqRqkoqvGuE3f6Oe0vjVpvQltl1LElAG4s1TPghiPnGxSkUcxVuNok3FW
ZtMxT1Tyy63ajx7mQ01zVDigLV1mqlsV3Oxa0KKUdGrPw9V8XSYIa7gLYxLaWpPKLrU2dAFFSrbW
mhdJCb3Sb8VCF/PmYSUBSU4phqHyPAQVVlsFMqc/EhizVOEF96nJJ+tNFCO7R91Efe9cWwLRQQLh
xRsTzpHrDMPTwUX0fC5ZcaWkQE4BixrNasDzhEgmvarPAUxAHRDkmY3/zajXz9U13MOnDMcbU1n6
fPO8SJnYEom5Gzt6wiYfb/7IJ3GwIWFisjsnIuBUhykj+5MzqE936LNwQoFD+XWlmfYXz3GIC/WC
F0Fl1oCj+hRSpU+SBKt7wzh/ntIIfriBwcSMHZNtzPUsVmLO/baJUqSkeuNwGUQhvSTZw7/2aKbV
eJYoMPzKMZ18syucKNCi4BK/I+dkJEpGC7Khh9wVcyz6sORWrlhHqfOSf4T9ehCx3Sbu6EToUbZl
xIV19dtpuAMATH9vHReifpqbTG1y5A/NZJMNmS+sS0c8mGrozIhRgBzwWNgGVKyNORDz7ugF96kV
BGmWloCXPAuDaslQsZaF4hwbLkmZqL9LwMZLlPzOSQjHMc+6f7fAQ8mvbU7t+xWmfdANXf5WG9cC
5dcbhJUNyRZfUrfhE6J6aFG9e9s8/UjVuMRGPDDn/gbtZJkrUPym8r38i9w2HrGg8cWiWZ2E2JRN
oZw4q6v3W114MONJlxZx1k3L4qHb40Pmkcr/doGbY2S7XVfzGtANvpEEZ+7+FmZxSMgTIuHXBhIm
6kmh7B3FsO44wili8/eC74yw3/fuU41TqWyqKRN1a8KmUad4U6/iJUJ6gZVxJzJyYen7pyqtLC+T
LxhGox0zM2cdu9cXWxc9i8SpAJwKoaaRfrztV2pdUaKxfCBW53IzTnl3ANABkZPScGi1l6TmcVdu
2WYVNvVRibsDOLbvUfKpaXOWk75CzjqX1LRx0MejwpsbjDPI+AB7tJHbTq5BQ24sbv4i0FXZaXO3
EPC0nAN9QdOcfOjzJ4llPooEVU8yAif0bNcYvCOujrgWdo8uqZyPCr7oXSqI6T6aZbR/0RfWFluN
SKUkttUYD2UbLHew8Al/hcrFH+MN+BLwVpv4gBtHfoQ380Io5V43vc/Fzex7AlYFEeTFOfj1RWRx
6kBSBFdHInC0oRxOsr65O/s/37FrRLZ/M50kULsMp223Mu29mSQYYMkZTZm7QBLEieMF3dMDsiG6
AiWo2Cflggk+JdZ8mdezyn15P4HRNhLJdyVpJ7AQJpzU1VeSaT/lrDyxgXO29ihEes9n1CE0rk/F
6VX8IXiJyT0Z4yqq+iS+CS1jKK0prZgBgI4JwrmRKLYnj8vFgJ3e68cFpI2KqOgX4Xz5PDPIl4qz
5aOVXQzoHNdSmR9KVHD34TurD8euuXz6GtrC4mgZ0hUhxu4u8uh/HTKIUD6rce9XM5m8YjYEqvsf
bYZ1j+MpsZuvvETPFL6IzlhCP7+CWWGQdNm6WKFP00M4h5rHB+IszLaz3Kv8dt8qOcc29LSms+mb
Bi3WXxMysz8pizcO1AEvNAFUlWYWngMaRShVdNr7gC090zB8/IZF4oHzja2x7x6/uzolaf6qE0IR
w3qDatDQyfHauLjWryg9ChA+hPu918GgTh29m3prNL0hpaTh8D+JLLYIrfRSKwCZ80QGUyg8rfcO
qTMu4+sByeJzu3/w5SZv6DKn3ffYDLt4iY/z8xrvUeBz3KoOmEb6GS+ZbGhY65ttqyeZ8gC6FQv2
HZLmLoOafwOtKFY8izFiqt+HAQFANLf2tJd7mR11zWrbtbEC5RVjfHWoXR/hz8FQnjlaeLldu6bG
k8YvhLCB+EzThwr5K4+E/8aO3dyMAt/mi2/X65daLvpAPcSeBx7Tsm3UjV6giMuMJy07UmUN/Nqs
xE2UvVuaHIdwjVBN29up3oS+NdBQWH6mncIOW3JE8dyAdxGgmJWamcLKvMadb9G+WjvXv07LyS74
4WTw+LOtmNOyTdV8TWpQ6Cc9wWASsrbCUN0/CISi1mEJIRJcFnk3aPBAB5CNQXNJ5t9YAPCAnhMd
zGFHYGaNDCkOfI2WyxurnG2Pl1b+amwQFbeY5Cf0wYIBhmfo2xA3E5ijy5qukXttDNXDDuzAFqYp
Po+keXJ/bJDh303BvDsDPg5aNBZCEW/btTeP5tlGUTjrz1T30qnUjapbt03V1wgsNa9RHXynyVL5
3UCa0agoXznzuoKuI3VbCkr/+TK2bw9AGv7gufBtQiU08UzDsNMbYCsOes1J7NURDYKUjp63UdxS
NZNWCOkLGk5iT/2HcRBC9NX/6eARhcesTQh0LMYT6WA/botgSlVvqnqarttdpKnoEC0BAkGwCzCx
btPcWcfIR8BLL+o4Dx8z7eju5F9t7vFtcD0NegRNrme2TH6JeyyKqzJhajZ2iqq9LK6kwJs/YTQT
IATUn0Iik5ZNHAOpVgOrH41QTZQ03UzZ4ty0cu78KYo+GD5VWm10nfMzwedTgsYzCdgbPpccRM1t
MFyV4Dn8oDn33yIHZl1rMqpgshuJQyiRsihW7wUu5ezeryyqlClaji37WAz/qxrrtbV1e+dFfRje
nQLgcZDZMCYvxo1UAQWV9eQGLCAh1vKtOe6JrbE0TpRXjoB0L6R8hyjnutRAqsRphTNO64Nl3wXA
QycKl4u34hrIBAQ3++aymCUbfiKWXWWFQoy1cKh8FW2BsTzqIsnajLYHBMA4sNyr9V4ud30Rmygc
ym+exBT38L/c7kvESKBotsl+Ds3iGsjE5Zrs7X9XJFsUlDcrw6bWDMgNWRbPjrzVY8OLX0ABsXVd
ZIeuylPNWTCSCKDjnlFuKCL5L5yojK6mR6YSnFEWEiYpC7Kz0wG3eJ2JIoK4JpBTVqoEaPDlPzSL
/06JfN/7L4TlYrzlzkHxZrY5QKkD9d7wQh0CGQTnGkb4A77U7tvIlBIIY8bm5a4my86ii27WsyJ4
VkcR2pUUMniX9inQMAkwrr9gRRPpvxa4d89eS+MyaB7LAoZPYKaOI1OG5WF5HOlMDhGlT+MDP2nN
w1tZTsuyLDrwGDCkgs/lsvUzWxZpD9XpbrlNBgnEEUVWoBHU0DWNFWte1jGTt26tpdoJJ6M01bL0
NGyDMvHHhTvBwq04GpxcX9K1LXzFFINB75RkEIboRnDwKLE7rCmiuNu+EypDjG8WsUeixoMZCMr3
2kr2y06eAWXX8511iXSFdMEiu7fSg08aAoZEKW5kVEUUxOMqB0P1fLPLFIlelS3DQs9BIgu0Hx3t
sDLNvfd2o0eeZ9F6ThKzj/pbjaQDkvEugdm734aUhSM0ktbXUREj+SoS9uPsX6dbRq+/rDLVv8qh
qa4o0gjBD4j6cL3L8ZLArfVD7W/bzxArvv2Ktz62Y8TRqrZboYWGabP/wr8LPnPN7I2paND3OiRe
ZTF5jrEMc4pGtB3OFw5A4iGDfr8qOwMytsPa2EsID7noNC2i3hNTHXVfwFuk6pQSO+YqgD/6suMS
MiYCM3Oj05M2pkpUFWApLQWzA9/YYcH0zX767cVOr5RPwBjxN9Ciy/Yi4/ISdIdxCpQw4mCvLx/w
YBEB0oWyhZ8HBIuzKSiISwhfpBbmcdBXnINtbyqr5lB4Utq11M42LlmeT9FrrACCIFMflI3CTDx2
BR7U42R1i/NSWcohZHQMlpbAD8dDsEpTjjP3QxfLnEI1QsbnA1DNEd3XZ3+TZCeQ6tIqi/V3fdYG
XPFAN0k/UFIZptvpKr2yTGuL5Tvu92/gnu9S2Iwsbk1WvxCpZYuCOVvZ72KkWFYhjpcUHGKJn5is
XSJPxzZyVm0Q/awaaCyZd0NxC7exDVD7iKgC9xf9/hBj7qIql6yNXJNq84wunJMsUQS99/HTxv7r
F+G8AW2tFxa8Oo/l1ELbse70c3x7BRoWAlDbapzaHij1vRlkhItfpKuezmCUZ1/NmAWhHRqQDZBL
vF1AEyz71jL1WMRZjGj+WyuKgKcxClTMIogCWU+pPsza9CCCCUixIxUGVtt02UExUDsTPpaVOfMu
4+9j6dyoP3cJzb/E6nXpGYRgX0sDTYcdUITJFOtLfVo92vLlxG4aZjX+hmSG8UQjY2t5xnetGfvi
14JOptvXJseFvGl9Ghlkqw2e6qhUtcXckR7TgobHpkiHc4AKCEeNf+OFgPZ6oJ/KcOMOPSrVqpru
PPa86FpgDFqHihpIwc7gpRD93Uk1SnJSNGi9IqmMO4ml9Dwnkz3gtn7xxJZntUrG1wLeOws8+1HT
WFKuraj2MoXC9HRdQ+xPc3oGrmr63gWCLJB47wOM11JM/Z1KTx+aZSOjHsPz9UTOK58HIW4bdWWJ
X0NU4sjhoVdphuwuC+xuqxLCKIPDyx1M+FjpjVUIR7SrF/8PZ4C+yldlj8yx1C/CdfAoLoF2Ahse
SaU5eTTEg/xwJCenJDJjuyIRu9waO/6r7Q0sdr7HMifoZnU+6Sye5PFhcUpq/AcbOJLMJiXouLkz
iNqNtLPGZFO5ukFZ35na3AsTdJVGgbZTaGxbBQOAMUqvPmbJDdgFqjYPzExmr9fUw0e1TiFOSmDo
0VTPB1oHLB1GEn3aGxLumcizGZVnJJNSO7FIyVxZYsZCpTIAwopBagSRW0+fu47nBTBjYzkderDN
XK9Owmjb7zA8Fxnz4pjMGi942WxHBwnMdszApCC2tVbep3rR+prxhdrJf4hgr0eEhovoLg2arm0L
n5seqD8WEY5V0cIiVkv5po2APoz8eggpcsbsoJW/E9afzynUEGEpGOD/VjtOVepdDnqekmDDPc6q
I3147FRPOwaJ5P2/6boPKniE4/UErXD32gg5eGsOgHJLc0+esoLFw0WGJcO1i2WOjTGwDY5goC01
rgRzxWwLpf3TbDdJGn+gB9qEKRr1rjMjYFrS5ysJ3VhaqN1uMGGs6IKFgkKYGr9+VMqvp8T7OpaD
b25KT0Qs6hTmwIR+GD/tHPd5H40wElWxSr/kUtUA0z1y8h3zDmJBA3uGaKFutL+rReVRk9LUAPY/
o2NCoHFOfdbXb58f1akUJMD1mbVVEe2bvuIJqqwzK8oW0LW3L9KW8WRpL2ilploSuuzHeU43Krp0
IW5Kl7m+mxLvAOmeUYxEN/C4IE5oALyN8Ik72rpTEmOZ+ZfQGQyAmqoXkJYObRsoSHehDBzts1iS
5FQD8hlF3fKfCI0QouxKvV+UjQsUjzsvsde/SHw2R5/oXeu0EJ1KKxHMV9haewOAJJWxSYWIifps
wrauGV8Y4W6YmttbU73SvD2GCG/R+rQ7n+HoigcaAgwpWukPDwCdeIPgK22aEwIUfqahQv2haVFs
LIH36Otq0qkR/dCKyoBa7i+u1YL6TSNMU2RoAbXUWEB77XWLuwJY2fgdhbI/AFoI2fx2Wo4pfsAm
JrmjRM3IcSCSI1Q7T3MxS9n7o2gVIgDtk+czPT5zElszMFO91+hbJDdW8wlKmLl51j2QZa2p+w8c
Mz54SAzNtjFhG7+V8B3kSMgUa1l6fufRu4GWnpNlAh4N7nGsx6gX0cG/9olVxiVy8JGsHV+jfAHW
DKz1uZXBvaOq+hQvtJRlQbC1Eu8nAePvPIjIgDJ5nVmZoZbiMQnY1tdrtR6q8McPp42eAAv5Va8o
Dx8v1HU4cikD9dTwPlE0t3RqaqF2xAhwhBvp5xgcWOi+Oks4h220x0hlWu8mRRxLMHIjtScJak/t
kPHptIeyj4V+t3dW6rfi2sPRXYylGjlSJlwu/Cvt+6L/OQCJkhS/wADp8lDwgySRiItz9pyNz4OJ
0VzpgpkQtpNaDVaeHm2CFplhJQWejyGgOF8ScG2UpxJymRv9ERDL+UZrC8RKDPyUOdVhWoJw/Hvu
GmnGy0+bs/1q8RnFasX/BsTgDa5sTH3EigkzbTUwWek3gjdX4+glOJEW7au4lVthkXh8UGR0wONJ
1UZSnllHIg15qiMj7OMKUtYk84CT3lsHrTXfzIFJX8gizmkrlou9Kvn13QvDyOFwWs+coM/yKkOH
5OAoQwQ1GPvc8wVfiW5chUKiHaNm4b7mZ8tA4nDMvW9riMstsl3yvxBlG3oxpQ3ZEtNYN9gAzF1Q
lg/nxItPeTk6o8yExWhsonAGCVm68VkkteDP8a73YtDhwsNJULvMWZdk4Q74gbCMghVZh27KGxiU
kIC0z7TV769V1T7lm+nx7iJSurVv5rTSfNCpjnmnf+JDEoerRhpxwuy5JupiJRhdrWEr8A4AJbmR
tNMFOnzBut65fnoiSwpOSR42LOPhu8bPhdNtsXeyCxH+aww2e2tuy8myP6w74ErOQxJu0xBMOKqW
dqsK7lx5bsDojM9j0oPeI4aOlnf/Q90yNEe91B7y7vkUpwiYfxTlxTU/Q7jKME2PV2vAN6gNgRjE
7ygcFKaRtHbsURapi+0HBjaEdVSa28GazFKEYr4v4PqU+r4lPxdh21QhjqiwyPQWhxItLRi93mFU
FdClJSDTYk6faHgZbanY0YaBOrWEO2XNEEuL9Q8L41IKc1bMVP2AddcljM5R0H507pH7YAtw2ilo
EWZhqYK6uQdbWOcv9xeqzbxQPXxIiipQ6gebdrhIu/zT7kCAF3KmPGVwfEwvuesNniN7hRrrFjFJ
hmPL+kqFH9XZJX8/B4bjbeGpjk5YWgd+7Mn5MNmHjVx8NrawF4dFAgITfJHQTwJX2ldbSnWkieuf
1MnE+2LK2xiLGBrZJ5t/hd/RhxcrYqR1j7VNco6MyxUezo8dog549VUPLE7RWuVdNd7BHZLQthgp
DZyGY+YTcgV+d74/kQqQbzZpcidBZRuyS8Sd263npaY8p9UG5i7nIY28fB+raZ4ZsCKvYbJcQwdB
hpNVhKBtp0FBuAyxUMRPpG8a0RtYsTILtwpJuTmITa6Zzf8+7ycP9WWDE40YPs0BREnAwYBSrPsr
FUc6kgiMbsgJf20ZBcF8BuE8f7cTCRlLeVMPg2/AWrLXYlsl5cs39VGQHSU/zvolZIPzpx9Rrs7e
tCfLZwvKbVcc0ej5MvQDVZtqJWkU5mxs15MMwgkGa11BSepvG20ANYTmhf6FmB3KSuMwOH+9RNK7
McsfCC819rAfkt4MdWRTuY5Q7Bbb5NWIlv7+YE5BSO/gc2Rv6Izks8DMmNg+MhliIV9BCx/wJ5ow
B+bZJ1uoXsIAM2p47XtH4wHGPVSyffRq7UgpuG5EmF2654lxngjnERGMXOa8rVrxI7UOka0hAhOu
KuH+nAzBmctR2neH84WTeYXFADkDlmDcU8doYoTu59JxRVyJKm/BbVPiwIMKr3tTUjrqZWpEA15J
/JnofegqR8SREeZM0HauTrn0dvW2+FfX/p7T6w9NUL6+VC+L9Cu0tCu3bJ2F5RFhN1lXLk7k4b83
wLWUS4FDtMO0sCEZr88Wo++euFJEPN79m2eCSFfC0kz1MIXV1I4FMyFxvhJHvAx/+3HI76czhRmP
yoPfCNu+b5T1IaYYLisAqKonIm17icqHIEHBe0hftn5Asw/r5kOx/jfWDhIV3Ob2LDtuWw8EjeDQ
yrx32nj/7t9bWCjXQlDVJIGt82qbgVEvoC8iDjiVxht+jO2s6GjlBppQYt/LTxkUnaO2NegPq0wE
azdC6BcJWmL0rYnf2Zs9mRhNAgJsOnhG7QPfrfZnG1X7O8NsAhIHwRDGSV3mqxY1kE5+jlnft1qp
ySTTiFGyTP7Ti+Hgy2k7NFQxGQRs3ZIXlzSXtJe8SGx60SC65BGQLCd72vU289TLcYehDQjkT88h
VfmHkIXyIiDCAhbKL9GsITkaM2ZnoIoskaWKA8cNm0mVYaXe9aGtK0VJjbNczqi0gK/WE54ks/v4
VtRRwEZIXKdlZZoj3HrL9uKwL7asPnEriQyKTj4T2IoOOl7Dz5p2efJ9BMAZ9ILxforuISrB3S2G
x9TuJhA/7+TpxXjyzxYxlie2rCVBekHApfcUXCsJzzmoJaGbg1RU+MUoqu/7tuzBEHTPM76AS06A
t+13xV1Jlc1Cer/HmVm7gR+35Da2zfH920lUwOJw3Qt54bQ1kxIkFT1GfAhfxi4hZ8j8wrsdQB+u
NqRNpTisoClZmHAPfa9K4UmJchgsp3/Mp/t91Zo3JHR/liCrA+QYNucfn2GUNmGg+ISZvhJwNKHT
5T7hqrBRO/EtjkZVybQM64xfnOS4mmbuOQyQ+ncJyupHVxXOJwhRwi1/pZauT7qm/DZ9xJZGym64
q1nUgWFJabTzFxeA7z9wWOWQFVpm+6MrlHBqk4juPeGAy+g1ZvupYNFLAiSukZrpuR6eebDjmG00
h9/UlLdDfMdbCEIDtkfTtEEy2RZ/PUz6PFERxoNrt3v9nMxF+gQNDMZRFHxQQ5XszFnv/0sXSWWm
/7XQDe/9WwJClNlxrCKxsaEl+CLX+bdlVC/DF6x7KkLOd2BDxcKgcGNhzJWkYVd5VGr1D14D/zPF
vVtYYafm0FgK7Z/nX/451t5a82JPjh5Oz7JRCLS7iz5BnFT9Gqj2fytasxN6Er0qb/d1ZmFUuJB8
6EAHeWne45yD1f06uvgzqi+TdD8eSfQ/w/sDdHUdeKc+O7N04dfxgBjKZKjGLwGM2B2jAIEt/jYn
+rKqASHq3WMBc0TsNv5HmBCPQ1WPKMtr3hTamDEE4W+60+hWbtLgAOqCD/ufI8Jpv3pIDTyBpJyt
smwk9A/TEntNGwK5gVriEWdcnnA30jY6SXvnAFCJCUx5vGpctxx8HA1M2YMET7cXY+EZFZT6yI05
zphYitRAHqAD+I3vhKSirjmcAuYNrMJi3tuSSce5uF1G35G3/BDM+sUtSS7Rs4jt5l2xTFPeEDDo
PfUF9Y8UifyLuHb3xmRMkHs2tv94LILhLhIi3Efj84nD+FBGvSOtoBn0Rqf1SMmD5ksCWW4wpuON
XH0im7SGhDH7mJ4UR2zQffImZXHGMzK0iSZ6LefFYHFQA8bGbqlaxzZLhsTgNdTw1KOZo3PdgcOw
yoqLUcJn7uHJwOSXrs+XG9WQWk/Jm44RCLF2Y44WHiiAlNiCRcCN4gYQYOzvIpBMynpXCSxOGGWz
Q/N/l5AUMGy6ZQn21t2fLFLk1Pd1IH1E1hWM/AOVqCfRagv70cQn7c+PnuqGFU6JNrtPjNuOvEIZ
KFBrgI0BLo/jxifmVOeN+prlCFRgD50+3yWhCkT/3+m9ZbKuxLeUdUD95HTIctgGYFK0f0GdoJE1
dmazpkd+nRFmNtcF24P3DwUDGUCJzqs4qMC0PSR8+tHM0CeWhDO5Fr3jb4Y1z4I9kv4aVzaIEawz
Ag04PVHynGH/2c0OaHamMQOXTmtIXqjuGp8VRF7/uvzK9C2phqHHyrQ0qoHMLG7LKEaYInHIY6M6
mvY0BIccjU9IK1DkMhBUVjlu9oojB5ov/Ihhdzx0zk3xBzsbd4Rwc077kKMvIai0gON7l88jMDm7
1x8TBems7sUJf1qci/c6JCj/alSvYVzEzKPAjdddVcGe+E2c2QuY2TkM2QosZwPRuLu3uqlW74c1
b7F8o6ta06PPRBrBCyCTKqVSoAUu45A3UqubbQzHtveq28vrtQFtd6xCaU7UnpijDQgpzcCA986i
3TDJ/DVrjXz5U6mNhpmiYuZT8NepZysbB4kJxT8PhgRxf+xRXZkQVwGF8D6vz6MBmyMTQdr1XV1s
++5g9Kkk08OrPoKGzZIHKqPPFtgRnrPeUBN7GQTdj36Bktkl0qOEAQE5ZpCSvvrz7yR+2m231Q7m
tALg6qHtyL7Duyqa7zAz+38yk5GJ173yQIkfiXTvzOh/oIUjFeZXxOv7ODqWkSfGH7MfQUgFweWI
ZdrKRlB98MFWzYBvxO7Mo+TqbkN1sXPbb9t4q3GfMwwly5vphNjHIeQ/owRIH/CGf2H3/dTV8nm1
a4Pt1tRd44ehJfs/JhZwcysJldAnmYL9h9AVmmEFzsvZYgAoXEoersmPc4GxgCt0Iu2CQFJKkEbl
JVgLbps6IUN6aF0zEuLzMDrzZwu6V1qLP/Lp2o9bSWMzPVkUwqid1V1ZkYxbSHHiUspPlHPh9jT1
jo57ODBbGVKetOb9NyC8t7WSvQFe1skFc0ET3n2clLGu3NQ0oiq12vAw9wNfbqc1R3wMdhO5xG/W
jRwnE12oOrKcbLAMu1yuGMoxiWQGkTlBcDWfTHKWzSws0Xd21mSx7W94kAo4BPuyndTDLh/dF+/D
FZlsaRXbrAVf01r32gNvaD4AkUjIiwwNhlZmo5i9cVvYjJTlCQWj8t3MhZVbr+y/Kkx17CZbjYd0
nlmppxxhbGOilUsmAezVKdzbfyceylIzWFDB8cDSqRwD7yKcDfV3ufTaK2co2Eu6RNIF716bE1kR
khqVAGNF6w4/nT5BQjOOK1zw6KTcPKOLhDK8ibIjcA+unrCww9AANSamX9GW1++GMIXEhvNSL3ps
LhTvRMfZamVVeH0umyJJ0+A+6jjbEpCze2pQiPCob0D9nT+SRovDE536T0cDTw/7vK0YjDkUkmvi
Gtx/Whoe3Fy2/C1vKriv2X+LrNpy71n8FcYH787R5Dw6rL6nFIcytExTckL5vlVOqyl/WM41Jh/4
7NDEkP2KVqc2HedoBFawRn00/f/O7mha80/DIc/AqoK81A+B9YJXQFuVAIc35vLxSrGm1kIpde9y
Zyks1A+RLCAVHDjlk/EMZOKvfkmuxAU8WBVEb9GGM0af0NYbOdsPQxGBZtw/oWH1IeoT5Khd1jyv
o7TyOtO8rPc9TXVwqg3WzIdVwvJ9Bm58grUnPkCEWS28K8UzughYboxr6LIygjIzlcBxDPKcbHeI
ynjHgIEhDsPB5sKcGWlBeMuadM6TkDs4OCLwIid1KMn49N8DgTrW1mLIdlhOQlB8tNAEn5r+KheF
UeLvlHgae90Ssu44u+mpMcqsPD10KavTEduekaJFpM47w3Xedv+GVIiwSY38Ys2EXBYXUxqc3R9R
uUrl5mCGaK/cDEs85zc1tGCRRE9ys6bqVWFV5bwkZYN3xkqa1VkhbSoIqPqAU/Evj7vRFGkyq5s3
+uvP4nwyMEIo0U2WdIeI5Zf4EzuNjw2va86vU8ANyf5cIWHzbwPbJgDSKKgeLGfTiCJBoM4wJeVZ
DOxxcPiqaW8CxKted+fuEwmba0xjIYBUO/jo+u1H6ivT46R3vCHnxaD1xoE6NasjrwSvHp9gSQha
tgg1d0nCAES85e1r9PytEbLAT4QSdC2mu3cq5ZKH7HLuziVFDj004f1YFZxgtoWIauI6dDO9uz6i
4YOSxuudJwQXrYonD4Ag6dvSw/YIbdWOIEoA6wS8ChELl2srswmnLKKTRoGnbgnQYwLuSmtureSr
e4IIEtExnKKy0AcQK0CVwy7RFTkew623oNvA3Zf6aJRucA1qxjVxJoWvc/aJkBargxY7ErvYRbHK
jDsvTT47xsYBSIwOHrE82MxhPfVna6JMsUvTPC+N1C2cvQKV1eSqfih+27ARO6cfEMRFPBLHyV+Q
qUoVcKwX1oZQM8oETAKDLfwKOPXsO4bKISLBzzs4GoshxPYQ4PacByOSTP5MTrqKzgA9yBUh5AsD
lTP5so/t5yYFB7C3Mr47pPe8DeVWCX6AkxsGjtRdXY+iWQ1dgONY2BtYMgbJD4JQOYqkm/gfEbH8
NojbVnBw1GAUxjReEjlums1oFqjkItjl2dziGEDqUH3veQNUVI28qdRf974HsJhNG36Bq5YpUO7w
GLt5o5a98u1YFBBT8WL5u/GvqtYTVZLEK5wRoRftiv1dpqTEnthiLMh0bjv80kIG4b4hNzhx2+tx
Oo1C8Wa2bxsQgzhHV/YlreuPQt8O/vJX7888nOssD1Pl3KwPsHGNeDwTOm/T6LrRQXXPpIy0Q5bv
xAbbttfjv0eihaxGL6QrsVjYSTOM8eAd/2G9EoZwfZRY/kCvK5xncVUtU/xitKo4yNPXC7dqog4J
5bNj0jhSrzIJnUQj/OBCgeK9K5vMhyULPc/mVaRGSOnj+5Rl1rvGuU5YcO4Z7M9KMpePAlQhVye7
gaGyl66ZQlsv6MGVGn4QksqzwOF1WKHR/O24PlpVnlazG205wGHHcEyqJKyb8wSfiiQfVq5c7fF2
uSgVJxlm1fepNvk5YOxtCgPASNW642ZdpPx35kH/lfHAyOSAujCXzGefR5NS3dLvo2silIjA+Gm7
+oigsDk2zP4fAdAfAd2nl40P+4GqKcOpFy1vaPxpAC6oCJ95+hnSEAlSWCbJytWa38dONS44crzr
qMWIG+oAiDrS6LSjEVjjVbt8SQhJ/iWJzHOOoAT66Li8pNFOhcQu8FGsFH4mBGDNH10XWVL1Jq5A
9e1WEsMB8JmmIVTSoLnK3Xh3Z74pRGAN8gdCSB6XqiqBB67dEHAE8Rc+zZLFiwcGPsFRKz9j7CtX
OsE16oM5azBNl+5ZpnNQmgZDDU7ksGyDvtvG6dvtXABt7hgSgOuZc8MGyW7yQnBbgnla1lTK8K61
OzyuyH0rcyhzqkZD+HuRXAqGE9egRFN3bMvKkzXyjxnxO9Kk/m0XQ0uTtxp5TmS7ZbLnQvt+5dfh
SLkY8ISAcl/H0zC+5kUprtXUwMr2moI4vhPuHEfhWQ40ja0bb3dbAEvAhivfnYI2Liab6n3ruPAf
FBWfC1DHlXWSYRrnYADS68z29g3qZTYg7dLZISnJo88C8eKV3ULffGXJwappgBlPXdMiAjQQRVZt
0hg7Ye1e5JPQggcVtx4yCdicj4/1NwSzhqwMO+vHzbG/cJ8TdJY+8834BQs8D8XM6hd87krI4Mbx
kH92CXkd3Pz6SzGBOPiCBXCKlDoIvRVC7DqbnSqosCHtwGEDcdlYhaoW/JWv3g78+DwQ6g+ZJ+Yv
y5x1pLKCAaYoaqkEGlZ+rZbvSk4K7tCllU0142vjvFEwR58T4vLsMQov69zaHvFJ01657Nj8tALz
OEKajx21uU5O6PaLkCaDs+N7LWMqsxmkEbidqGLdik4fy6Rav+pOsXyUvtbKRBJV4mPre43Zj4Ap
aI9DUfz9ZD7lf3tYbYeoFo8TDX35LgckhLl5L1hGB+XB49GYYVBI3CqKnQiZi8b1ESaQG9zE+p3U
TYvnNF1bl03RQlHX+vAsPg5vMS9Wokh1jcox3xl1amNhKAIQV/YnE9Wo37rcdvy4OrJt/0FHzp8k
pMq/HcPCiHYaCIyTm4mI/rv0jMSqATMOz+Z47Hm9UdPbI5nsqXYHq8La/UI0iPdx7gZ8glD4RaOF
CCc1do2q2tbp4RjjdXFX6VjKe6RfmOqvYcrIQ09dNHquAyDIk1mjpel8ufQsPbl+LGdd3agVKBZE
K7gaQwhdHrmUFLoQHPWx+G0emyO01wbysu3QoLRfqvmVOkdDDnAzxo5UsmxTgS/Yr0zL/Ck7b3GA
iAPbFbSDFeHPEtdbwSVW760PyKfPzYz93lZYV5EdTO5nChfJWQ4wucSQLjCNmf/CEhk9bpm0LRLP
Edp+cGkljZeFgpeTsZkjydfzqSqNrWIsYR96f8+yhf3wq6s4S7OaoBTusuOawqXSN5QSedUf+/gE
kE991oGIk33m+qKS1sUcWt95qqT0y4EzJ7Qd/CrVk1/tXe+9C+d+9TDALqrPWhJqu8KoIZV3SAk+
OzrB9A4t2Da+8cEDUlx9W21STC9MC1d5SRchXoq5wWYcucLalGIyBHtuIkEnvjjjd7QyILJkAs8i
fT2vmbGKdo35UVIjaOKl44B03I3ZJ5UMFM96nOvnMq5wPosWRKPTnEZs5KcE/6WxBBegNHI62xX9
eP8aoEtMdFzUWlgGUjVEDqWJxn9gDXoVdRVSpH8ZmNeXPJNzIEUwNt40f1M5SnHp2Cv/ScVNzZ88
sqo2WB3K9AYMmNhtDLa9/Yvh1M40JIEsVcHwisrueJu1Nqk5edGJ3WEQsGILxfm2HgTJdgZC/v4z
aLzoJVOB8sNnT53hqAxaI9ivWZUOhyHHQuW/5hDk3RM4ajOv44YwtQ0hRcbfIV9CmpIBv//lx4sQ
4Zif6ahrAgljy33kF7J+xQn+VRpFhHd17I2098XJHYtQ/F2x+JDDH6eQ5Gf5cUSyhiT2UD0t24xW
9eXgMhxssAzds2adU6kZmaTORubnghlSeNz7rwkkCLPKxxihJSNWCSogC0s6zUfCuZKTv3D+MFj9
eEBVOZdcs/MCNuQA8wUnQmDwQ/wntI0bA/w6jwRIyW5Wo/9wB9Y+hEW05NRndcIScH7kBWVwg12V
63/ZTMoJRGRs0cb8P6wsmOc/SzbDr0dpMmSDF56fByZft+kZ02jo9BiYwggcpPQ9GX7Ba5C1UibR
WL2JQAG/o9otlW9FlFsKHBkwMvLIn6rKiwYQMqIlsF6h7gRtif1b9Qp+Kgqkiv1pR9cMxPawAuy0
+rnz3UqHGyMN9SxOFYAs0rdHKUzbuF15LFZWLrNwrdwR3prcWhKEW+Xg3V0pNRldWn3nGjjdoNcV
18S4vKfrrxLHwGuKZVBp8yQinUq83XqocPY64/fJ3+ODAc6MR0ULhMZOwIfXP2FNNpBUYzZY2p1s
NwzpEwJQsseWQReQenkLl946wLXmRx0MFAi/OUWiR78BjWqH+dhZey/CtpGQt8B330h5SzqjdKnp
9K0jU7jE36LfIGym2/EjgYMe7L2ZAeJw4kg+3BSyYdvXkKKpHxxeXbLddMZxwhnMINDowMV3530J
XzKP+G0t4/hFRTeHDVZ924P5SE8IGKHwRQeRBFp8wJ+EII+zUIulhd+SE2yoN126KgOBr3jb6pof
J7Qdwwv2jcUyJpAaU8Uzr/M5hsiVGy6x8M4LflXZXQgRaTX56i2foLt2b887KKO6kW7WuLzYG6BM
OOKSnNn3b12xXyb4DvzaSjO6SndmrtfFpJONbkqWgHT+JmYE6Z63jFewzpw6SOaoymytyH8Dc3bp
wz0te7KZD6K9vxaC1ZipyyINU6ZQMGPImr5u+JbAV7SUjoO6SGIBw3XC6ik+KdXn93WZTMt8qspJ
anbE27nxCQmhbT655S/mxLd1RX7Tdp952UFPx6iebPg72DDLtuqSpLClscHhfoAgLIzTNCNNZmYY
wCpJ2ibJDFJTUlinuvVDR/xM3BKvITvnU8cUqTM2RMA24XvNU4cOEqPmzR9Qk56sEVl4TdTJSDgc
agmlk4bNO+gKriRsm4W62bkP/s5TwlgtfKNcG3EXJV0vJT8dgllC+c70AhYy7Sn8KM+6/wbpkVIc
Ed8WPXCZ8eXNKZdadifRL/dn+e9ePEeL9IZfBeIV4ajDsw1QwwsC86IVBs2PzbhFfH9VlJh3wg/N
EhmHX6tyQ0dy9u5PQ3qPh3AHrcosXXEzZJQ2vtwpG9zk9YDiWoTFoalVNTHnRMgaLiAKGXyF2JoM
KVOkddY6t5gsvdRpqy4ZW02+HUadAxlZx0StUdEAi+n3NCvNDynIMfFDyRVWCQ+m3RqE9LPlHxZ6
mZwcHSO3pmbwtMRhcv0d0H+WR1WlHomiCRlF7dW1HZQih4crMKNvDQieKKw5UjZQSFrcVCoZ6+BJ
OkWxpdWsIKJKWXcS57aM1pNmcTdrm9l0s3BUwnuz3qGueYLqgY4AnUcjwG7Oh9VC2b9XCnd643ug
0B3sRkj211p2wQSHbEcKk9MyXjN5VSC+5lgVpAbkPB0INcxG8emhMvwwqYkkBw8gR5jbuuJ/GSQo
LnfkQRdBK8xGPHT27v2a5y9VcLFYoiDgO6IddK/Ziq4J8WvVkEFQW1xdlkKZbd/YF5kc6mQ1PZ4N
yOykvfBKQezKsggVGTkYgeOezQUawx7e+y1AcQtp5Z5QUC+mT1PjRcQpZPR3IpXXXm06rzFOGaKd
YqhCYIdYuuW3waUKyHxgFbWy/z2NatPer/AtjiqEPLEqBQPG/essm0KOiR0YFr7qTX80bK+jpONV
I0ZX6dbf/agj0Qr/cLXM/S/U9Yfqda4nEvtL5DM0MMR1U5TKrGWCCuQkfS4b/ZUr4aKTRFYMOkKy
rvvQjlMOMTIm274wZ8J4yfsgV1j0XulAgtprflLCJNkMEwgcIG7icaBdZ6kAo8pi9XFBkdp7hV9X
aHL/aWhiadA61CkpkchXIoMscnAvzrVs7LJ+xHiIMbiofClt0b01vk1jm1TnHu+6t5pQU4447vpy
/z5zsw4XC2NB8zlj2kRHdaos6I0bkPUNm0KUTVnpWDcK+kkLX0pCD+xp+uKSsgslyp5V7wqun3gh
5XSrKOs0mLTi+j91AoTXjF4/pemkYe7Qi6M5l1n7oC2ZFTdz0picoBZrL79cmpf3yJ2ED5j8N+Qo
1dAtagn2ZMHiaizOpxknpx6J950kZMRjjnFvJx0iBninoVhEIsNLYx1uGqLpfYdZvWgkhRKnp9yq
Hvnl5fsQbS1boeadd/jOXKNAOnKBQEPtrcS7CTvAbiHxlugNmXJimQt0Hw9rbkzi3si/j5nFCR5R
r6d/DBZxMj8gifnNqDtW6b35svz1TBUPbLw3qv7afNOZF0O7cNP79MIIBO1yiyhjPy9TpYhobjRo
oRqwFmI+SeXZ1eh09ewOcKYlmu/0coIsVQiS7ZxUD/1H8HtuqSH4Jw+JnngLGcSlMTpEOLysPKiJ
JkDTI5HeMEWt3Mj8AnL8dQNc+IrT2Ibe7OpHLZ5T9Tp4NNfBNkZPxGQoZHsmGvk73NlHE/DGx+3T
BA4x9o9B3nDf4nBDXUUY1OHeksLU92aWVY3mC+bW3kdMBAMTt9IWftzdT2tgnq/XtQ0CO8QFyYVa
ms0D17ewqgah1y7+ndcuE47RwxB5rk7CnJ+IWO+zVWNbnue2A9XD8wqjqhOav1jynDF/JBEL6MZO
Y11DrjHsk6RkhjLn336taJt3qY25zOZwRkRBWLWvrGaAJpNuUSqK7zZkXIceBbM7zg/AdrK66DLv
8q1szsryrFl5JWhCcn1YKupThsnTraiFSCcdDzVUQyXelWCkwpcWIIJ35UkbPSlDpEqb8i/U940o
3v4x28aboP0UU6fK3IM9hkNz4XqmvfNqSGGuWpHFB0aSPr2TtK1Io2FOb9ifEs0kD0wO/bOHO0mp
qFRLy1rYO5g8xpCvtrfaBu7yxHHor0Uunr/+r/2vaMUzQcyLISlMp59gF2/PHMi1qwZSLDXFvEoW
rJGtjWNn7ON3IQgA7JVb34h0p65qPFxBiP9vC6q0DMIZKIT6cgO2b3WmDPBWrlfaxTf8Ex32kZSk
4xdDwEjgj1Jp3c2NzxUohJsntWfpVQp5P9oW7u/oJalL47Prv0PE+GXjCSpFAJgQI01onVD4fd5o
GULhGP4o41qeMoQTaDRV46WkuCH/pEnXbYDWIw2NNvqhgM0Tjyyn50xJlGoGosCEp3MpRiQaoKHV
Zj7PNU16fcEasM6X4efb0V9wb4zzppbrOVrxjYEr3vyCfSqgxcsAwcrDx09fIP82BmLRtjrbrlmw
tRRdhjeMF+FuclA1Gk07l4ou+LXOx0F0X+PIwmErEFkFML7OG3AqkTtsAH/H2Nnbbqz798sdKPFU
7H1h9teHDn6YZmDxEjTtBjgD52Wt0KSXLdifK1fMuVoOWBmaGIvsoNEKHUd03Q/9hd4+5yzoYtHV
CxAgo5Le/rdzKeXZxr+AGtlzq1xBK4ElLY1b5KVv3ZWYV/bZQaRL6mPYYpVBqGwXdE4eTIN266aX
bc4ED7h072NzuCNqiQVjI6TvtOw30r2TdLa0AGwnbE1K7Gq6iveoC/+PMVuWRRj6Df4KzkFZIu2h
pAHccrj+8In7uFAf/BlawtwtNgys2ArnY+wFVRLdM8AHtzXKBYqxX0Ll+wxed4iLrpNww0kFzVki
b28ndJoRlQL5TIsfaiilUPxABRpxO93frFsoflhjNvW5NZ/17wk2eQmgPDO/T2OZ6PANUeg77NUz
31atcgeXuKMU7o4WXu/K2ZU2QW9MPONpNzZ6XDAjjhpoY++SRmK01ZaAjnNymJ5Vx9VqyhgoulVD
cyBakepx8eubujVxc3HjzfHyZZZ7hCPNjedO0SDX67ajsXn7kStk2u498JGvUKUN7ew1f1ENbEJR
Y7unhmnb9Odn5CAQBMCmFJjAFEQRHXhBs/P1Px00M0J34A1XFBKUsCvSVkgiTr75VCt/lZ9i3+9l
VMRf7cFs+qjNbl7S6HfzAS7SGrq9+29mr/Xz8CzLP32OMMJaHiPUDmrQ8oWFqGQMRVUc7r03G3uz
4LSrfIhDErgD/ynjFNpdhyUcjfYRMDXJsMVVQolLQcOY3beoSEDmUyhqLJ/NF8djpPiJuZioPBQ6
RB055i9HkJAiYMOWsV2oKfVVsOQ0P5PAfTIw52uBhfdBmw+ZWZzCfS1LWHbZ7gUW2z3hED/SpJq2
g8pMrljbRsl9ZZEL/HzU8/GaWh7w6SW2kre73dwVBEuhBy8UNZ0gUJSzvSALaJSFPJpjjefQyrP5
ELWq3ui/Qq68musK+ikVHfs87b577dUnrHRyLdgONX4e0ivaGM/M1jYQ1xd+QP580QF38wiF+Upc
pDTeu6JqfMNpKd1yjqbCRv52Q+Xx7/n/bCc5YTQAcJ32Iu/pVME8hJcK91iKf9DqHI8p1HUoRDmr
EyqU/8a6KhZPOXN1li/BHzvjQMSMBuOb3F3QblEAHQ0YhS2wp4B22aak4et1k66HpKt5QVjp4g2U
M3Pu2/QcnbYHn50xvRBllvcOMVFQZkTZLb7nmrxfdQ4ha67MLXGRSfDCWflwI47cMxrOrTwt8IrN
jZy99lgf0acSaNUbD5YOql2Oo5kNORT/JNpMVeJYvxqGXee3C81xOLlqKHxo4FpthCaTSDOPfTif
yxcHdpD9a3e/mHHCUHoFOtJF+78J2Zd51oeTM44yt/q7iJDvW2dA0AzrLtTB35++IVUdgmZ1H9S/
UenhIZf4zrdsFKWWqXzR5fRfztNwyAAtbL/qnIMHyvWOeSpDaIrQovegifZAhTAczRMTF6SfwPt8
NEK1Qw2reyEhlFnwikMVZ05H9j55UDx8v/MBAgGX2jZrdgcVkhgtkhx4cE6O4qD655tLrT76elbn
c57lDFN5vrBXKNCDCyvoW52oo5xaGSNmiblBb0TTYwst/IZ/TV/OIiv6KNXMavgnzzzT3pVu6D91
X9S/afPoNSEmo1FeJSq2oGPxN72iX1KOuSmJoPzHLbyEZnP1MD5GPQF9aw2jo7HBsdUTVLAwhfLi
WVUUCuBr80Chg6zvJlH5Aw7jCeKod3TGn4MeJETzzmxeH8PeP+8VBGXQLmW/qt14ioiKKgXmOb0U
jLVjoGbFHN1hKtQ0PSLC2cdhl+1iIQlwhCn2qRidMwM4no+QbvXFGnUpOFnEn0zjYIe7JoV0FGKW
WLlLZqDM7kJPulxtmbiKC+eNwePPy9IEE9mUD03jG+O5EDzV9KPD1Jmaaw3KLsiwozBryJv00ZDV
1qiyqSTyjj2kwlXxV9iIlj6ZckRAxMTBBxc2sLXFnXQCEDUJSuU/Ssgv45IgGEa1rX3wE3B/GcTK
7NsUJhBVbzJOZ6pnFX6WJS+lq/Z5kTwnvySpdbPy4pzqszP1ijDSdZJoZFjQV6v+nlJkHB1rJRPb
kiMZqOkVQS5L1HbbnJaiud7PmctGmNn69KmpRdCxDzqU/aPsea1ipfkcJk9/vhXY7o15To31rY8Y
o6ivtGWK7a/kTMxCXe99UqdiMw4QiwmpMDMGy/MbwKKhxIMqP4IIJ6ro9XA4mEirqeufjeJKJJG9
Z16d3GjeI1gOgemqOFz9rmEI+7rbyu0TSQvW8J+BUndwTlEEVwSJ1lvQRbGQsDuF0ZXDZuaT0QUn
SDb0gISIU8jOL1x/VpfO6NaLtgDQl+IfpoN1WbQABD9DLauHxNwMSpf/of8ew30A/J4wS9PQgzzG
p7ZlvpA0t6FYQyoZi94Sx/6PjWZqHFFQdwZLNPCEp4iGqg1xkJsyA7w1BJTl8x5VYQi7FqEjzYqa
6i1eJRFN4WNDR8uHPAV8kGaHeZelZIHdGF5huftA7CFbaOwCITidvnzRk2pkfsiCb6x2XbC95ukX
ODlFjmTpnRgWXIpnUOK3lRZdlMdJIApwKl2BVBBTukBazMaOU8kz1qsl3BUprCiVHAdV3jhdplS2
MM5yxGjTX1byGdfkF+b0gFUcECKauJ4TaHxQgeQMV6tJcVC5ULW66aMCl0naFv2d8t//Ra2YQGrG
keoskRdHwK85Yb8OrYlanUG7JkKItjol4yfuDVelVxE4EFbWkQjdkEObo6wmu9P2vKmI8+sBjfdP
wM6lBM7jiFX9yy9C+9BYzn2tXlRvM4KE8MzGn7j3NqacvWrayb0MzQ6Ktey15oJMWRbxFxn2Se4n
bVni4hpyiF2iaYYyosWvpOgQ6EpUsuieUceE4MwUlYrIR/UWH45TLFC3mRMs9Oeq4KmSx0JbLWuH
CtH5turE/uiithXDHzWOys0mimZ81AmCXFMWUI7qdGZGv/5Tt5uXKWuof7kihM2ydb79cohwhqf4
m0Jh1bHLNp+o+TPGvMVtCnmUT/diJqqhFR76dPnWHT0uHT3fwOHRXHrsYhNJa2gJRmOLHqOF/qJu
rFR4kaP5HIPxhX+PdGP5gEYKXraKB31IUXiOZhDimE3ZP8FLAX249dUT2V3N6vVcNlgYSJwqAxkn
zDyxosG8lnf4ZQWrYNswxgsma76pfQeeufFKBTScq/DGtjZN+z4q/ykCoQDgMbIH1uHJAIJ+aPud
ZRXZOYh3xA5Yz/pJDnNaJ2N9kNJzx/bJ1BKselLgp53l040WwFF9n7Zcbxu1J79AaW61jux9sVxv
0XauYX7x8Y5hVYH5r2lj535/s4Jsl/zEhtyfNHa1KPYXs6GtRCNwdg+MeOElMOLvBKCCND/So9TQ
oqJPKC/YRfeo76u3Wf+HdHcWoYHREYwXAAnKAdtxQ1fdzWjXnn41AZdRuTpb4oe/2L+LYhcbYdl9
6I+nSIHwwHbwgvukhQmuQpOqsDHbb9rha5Oxdkp0MLQnlhg54kvMEl5PmJerSdPb5DmsTOEAdncD
DzWy+roqz67vDdQDmB7LmdevDLNue7y/xSWlUqSqOAbP/MBQ3j0WK9+gy7zpaS+s8/uXN0oiMxcX
7OocQD3scVHeFTY7rMDXjmYhvmBSY9O7erkzv7PF6mwNrA11RMKoK6pTpGbAbfbxmncB6WuDhivc
vRChEhLrp1ohdKv8OmRPv89b7Qokwllsd6QDPOdsA3bJCXUot1MtYOKSfsfFMS4Xnnao1L1WhiZv
tmpK9LKSSGvI2sn4Psm+i8vlzrAkhLI9aarNUxDS6IeLHTALilQJ5xKRTorvTaB7o4ce5f5iDW+y
oNP5A6Sve2GGJBFz8ue18mSK5vBiH8XvCqVUEZQWcedkFEssY0yWTln2DzrSakeOHKXh41ZsF6ZR
cUuQWKuFUJG+SrWmKpR2B//PSzpLVxr5ZdBcGD1VZfe3vi6KDF1p/MAwY50YfdL/+pKTDeJlwhwx
d7DUqe1YepWjSWrcP1MIIPuJ8F8hh7OiwmaYSmiDATUGAOsVJ4cvOdjCoHW5hLoiRXxthZMh1WfO
HPej8Z+zWbfD5rWk7NJLfB+xiFdkVpmyXtkK3pnlAOPrYzsuI0jVx8QslPIYIUe8SWyqYCczbKWy
nW2IDPrxd5jYGzKETdMgMbxzADnJkdiz7uMX5i6xhs1TE6F0GUKEbP+xRC8ZkV4AZG58UCXH3ymB
t8ukZCa5Xt4AzEspzJNI7HQNuZrH5pUZcL8pHmgQcOunARkznnVjhFp5f7DT0ZVpEPJ6+ujIa0rE
P+nJmATx5/Zdo+ICB1ErFmQARY7/qVb5Qx8SsxOgHI7K7NmDD1uJ9YII/D2yzY69ao3xEPC6uwP0
uW9bQJLmiJhMhmuTA5HOod3QL4lEPhwwU8zkkHWtMcMLcEkTCyRPrRE5s271hbvdmg6om7+S9oWr
gokfxe0AhHe9mOTUaVYb7aK0n+xyVVm3bx4qOVSfA1Hr9jnfPwLxM9vNclRusSdo6JSjCYEkA36W
RJ05eceblAHGOJXzXEtqq0Y0QeQIVWdOrvyoPNzx7ip2YD+e94yzmUteoOq70+mMwaGC5CbZpkLn
Nlen34dqOUhF8gpi0mcZES0cOFz9PRbm5Afd4uGIqo12SpjSk67Si6eDxb7Mfja28PO2J/KmiKrV
QoO1ZnldUra5Vl5bnzOC6Thyio81qFqk0h/baaf9KcZIW0j6ahQDFm+7gE5IQE+vsVL70sFgSLLI
Y8CzaaDW16BTCRYd/zLcvps1AZV/+hjMfA7fBQpv5CBmDUaelMJDHKDkBEU21iUGv0sjSRRSqJxF
fDG0fYkf17LVIlw0ScPpjFZ8ZlCEJe1kIhmxWIC+xaxvMWxUjVBrLpEKnxMy5miFbQYaF/OaJ5OZ
den+C1XfDT2BknYLcVsFtGR5mz6TZvSByySuaKIZq4yErODTpIAXbl3u2UXBSny7KhnVXnxH4tcb
BLEl3wCbPbV5WRGTHx93JMMeRbGuRB0I9vHetCBT0FURQBVnoPfTDsdiqj//ts0lVSacJhfU2KAp
cOxvMjoZoTPq8YlIA6IEw23VwlXzcFbx3nxqZCPXnMo7LRmEjIcD1khB5IXdy+A57ujBt9LpM7MR
+riXrtUCHg0H8dpgXL99CRMPL12XZOF9UYnJMqAZHkPk9ddFIV7CHq6MhQmWvwhyFh/Ww9yEdW85
sQUipBYl0InjCBgRpdlZvyt7RcjgXJ7yh6U+jkYnTSc5hqLhDnTjKzt9F23+NDoSG7FcKjD/74Ao
YxvaY/nNp6l0SH5/lBABQ8k5r763xK2gTEA47qQERrek7Q5bSAbQqMgJhRAXLckNaQA63c+SSjpB
OBv88OqhtmPIh1KhiHZgZKx3Pbb+AXOf/yvgiuL34/zgb1TTXo2Nb7s0gdbojzCJnqyzYbp7Hc27
k8ASaqoAW309fGDBamZaGdRx3kJrbsxPX9BzbU0Y1oW5eK5e7M3hcd4nZr7+oUsbR8uii/l+WPqk
iEscCA1L8W+mzcEm+3jrH6OxPF6afCpB9JLdM8XvKhMJOeaQTaz+1QXpintXb4j4Wu7BvtQdeaVw
qy8V/i44lwnGxJKA+DLiPvv6a0JkmGW4QIyen7Brtks0DY1AOt2JUF70CZEWhh7NrMUzrk/lHW0X
pJ5c4K32SmQIrFuwIKE7ean/+o9/6E+RNAdvCRWWWcYojsvS4n8i9SlypzLFSCAhUufl1wGLkXg8
Ukl1ph0ve4rD02vR+x/655vLijXjN/zYeb/rwM+1rp67l4LAr0QG2gIUu9ts5PDDyDpxjGPBEdIs
Dc6skcMk5oQIsI+II+++yyRUTmh5vpcTXY08cQ/ucieLtkyaE8GaHA2rrFeqgbsnifFgv10T6Iml
kPMmDJWifMFgQv1m20mCy5Fj8VgYunZwhdIeEarNmh9xp2zO0ufEuG7LvD4VlPPa6sYiXjHDygON
WoT1MifSiNCwE80oSA4f75gL5LPCbOGSIlXLNYp6Ft+Jc1qv6DsMyDMC2Np8w6nI6RQtNmbbZ4/0
PlTnKx3jC/X+y89A0OYIY04avY6OFlEXg8RFfSdV+srZyTfUtGaj/ankFAjVQ+PnIs0OsoB0M+AO
Qk6Vwp7ufiZr8ZGH4vT6gnOpHvFNJaOcxTwoHEGLGjEeAU3hIhcn90Tc7HTomWQBaeGZFka3AMY7
CUBRv5UTXUmD6S6Xo2ECzbGE17yZITwPPAIdJBbm+J7sjh3qUUXP27niiZwNnMN5DXnQ0KtH/bDI
brjpW/6ihO5E3rsOQx4Q402ZDcNkwb8y30AaGSMfzLmpmZdvXQKbuVIvIl++MgJM17pQYTvbftLj
2x/eUxrpMZ+kKF2XCuTW+5s9R65Cp6nGD8p0bHh8Frv+O9SePD1gAuzByjJ7ukGFxgc7w2c1jye3
bka7EceDD+n+67839gZwfjfXSRJrL76d5SoaEnTdaRMMlQ7AQ6olUSt4KaQOIk6JJOchDdReSicN
6YXRmzWQV18kg3OpQxQYG1rmz+e1o+cCiP2H7Hacr6xPL40jkIajO+1vgsOghTstayIP/uKNpOFW
CTWZBv0fWOP6GeO4zvdNhY3hkl/Cd3Y+Q3jJKgcxfyCemkPoAxq3OMIEUQ0oS3mR497xP2Aa0bsu
otAUUxQZw3aomr5GVkEK3hotcKaGbBvEb82n7NZdMgup9pjGE06K+O/XPAmBdA82tuVdsAiy64rk
PYQZJrEnQhOrs+v3swOtPk7nAUnSUa6m25LbNRYzmVfbCpRWMNsHHQ8hqa2+CG96dJPKWcjwFt6g
LtMJkkIVvJ1zfVnmUbolT/W9Hz3h+Eoc28ldMuO5tMqvZgRu7Oj5iZboUSjBr+D+9hrXFI7mzpc/
D95KYuWzdRyK6rnfXVhBy60ZxpEDdl/vPcDoORSVqhhKkcXYTihDnst0xvX1GC3vKKsGMmHTXDVx
0DBpOWNm8UORisqsPOp9h4nXAteL2vz2lAVA50c5DbSzmGuIbhqXVQn6raJdPYlpEAQLWs07U7dX
gy4jmztTPV5n2QsVySo+zZnreCXsaYGJUabfFEywk8wg7DFsylaM/XRMXpO28R+Dfaq6EZQy9BqK
JVgFdatuAtjP08yYzJlQXwEBUqET8jWD4JOwduySlAK2x5YWLqqEWdzclh+EsmT0EAl42rcBt+7H
VCa6zbLF/UFLSTzbTKrvs9k/RrV57rkLCLS0kgnOT9QupU8TrUL9dCfUiF9w/4tWsF4eX3wxCsiv
hQJiiuGh+igbnFQ00mut9gm+Fyvn92DdRg4Kja7bq2XJCUNLLb55M7FRYCMu1GRaWqN02Zsic2ZB
t3bO9XCW64X4oEtStgNzx6jBNlx47kFDhuVryn6sQM6zbogt9HEWdrhFYkQqYiY7MaFUJAEEEOIr
j9EuC1zockeR6+GV2JDUHiKcrgx3W2iA4ncguKbUxbNjlIcAzpPNYbtJV0BU40pn7iPSjySFiJ5Q
l9Lo0XRh+nYRPoYRb+Krcb6JZu4VJb9HMH/iF0QW81K5l9P5QGbpmg/K7NwrpyG50Z4nrbJyKd4b
+Gu4PAeiCBf/+A6PvKblOGC9hdseOl9qxgw0T7bKHT9m79gT18yAzoTpmBSi410gxI/0pDGMKyee
Um8v5AwObW5R52QjLxnllvhK15+LkU6Cv5imUhj7nrZAg+AnN+a1ifwchBEPAZOMn4Ukf4OE0qyN
88eb+jNzXzWoafp8nKNyiGMPpz3JYtV5kC1casstI61/1TTMhZ4smowR0Y50a4XSFH0Or487GdB0
amVu706UMZsd8uKCNMHBBrlF7XALmDj5LByOXTGy7VwvZkLR6/ArsDuYHtEQ7mxwW8rnq+CaPekD
y3is1TEkPtMDmpLFz2eFqPOStB0Clj3XazDT+FQo+q4txuzL/zUwl12vkuRxpgRi6pM3wBCDShYy
Pd0xz63dHwUcyzr+KQ+Yz2D0yDSkXfM1k71ZIINoYEZJikR8bWTOLjA1x9UR8RSwjfRGgzAc76Co
DftipYILkB9M52fjMqGGe0IX4qAghF1eRPlrcfyr6r/n3NppCeVSMONTChJjbAGe4MgVdKEV6UQO
Wp4cDf+qqLa0ks18SMUyDaRKz9iWbpvR9/J8mPILwhe9KK/SWj2GPO6cuW4vy/l2VbebaTQW1eoN
t+E7hSmJzKiJPF/PIRsQLJVmJwS0Fg88u2QZqIskBZDVYSN0eDM6O51DgfA7T0SiznbUZ4Nz1I2/
LlY1WtCPG7DXTjedSZw9XgWTJ8j1FBvqA+fzjD8Ao9k0CpZ1+RTcBYXyywvD4DKnaaDcp64/2Puw
p0JMiXnbV1/Kginnmd6J8hnd0htjqRrvZk3yiT+g3tVVzuh9wkrCeUQXXU4IK3+ABT8WW1ZgCVf7
paJKC5IIetZG2XZa2QDt8vNyPk8m9cBby5SeZ2furwmNOguPuywf5DHlCvWav9Wz+6vO4t6qS3Vt
qwml7hkQiEDk6RGgxAYyvPnWGrZMsJtwLgxtvxTV/RuHtPya4Wfzt3ac1PAOEKLkSnIFjiFtWV7U
7f5GZx8VIPPKBUvT4Fuw7nK467uY3n3n11YWu5u+1ZnaWpyRgJ3+1+K81LFOllJXutDT8LoNxLxz
RvPywh+wJA7Fxl1uxtBHxCSwfu+QgIKCDxoLcGAONJPlMj5vXVQfi1JVIcsAQQ7YRBEBzPPd6Uoz
scVOVDTKhF9AX9Bhp/t7qpzYwEZfT04rEcauEVbxE4cEVEe5xfT5p3RA07EGLv3Af56WKB9iUUPB
zbvz78gD9E0GSiACehQFxa3dEyQXfn+wasvQ9+GBdGDLIMJnBwsNOIM2944lV8K9ax8DIUqNuod2
j7akV8beAf1omlHLiCsn9vZDkV0xLXNpUUnhxmwlI79LOkH343mc8WokzqloG0V40PwhW5sMDoQ+
6t01fHWwuQudXSLGKscNpYxUZ6jJjLkEFAzj3UMGTpDVFWf3y32f9o/TkxhhiAH8R1EyCmpZOkMX
jRtCTWCHlPw4lfBoP4ZFftAtFIoiknu20srNfumr1chx/WPS554UWD8r4ZX8m2RbjL3sVH7jWDxk
Utt+2k9z6vClZp2jzYoo6VoP8vylcoEpcjtO+YwrokDTaFUhQQoIyLteOOKjG7yEZwarOB42XKuO
ANt+K6Q+bmyR1ZYrW0SSevoNUrr27of9Uz6YtmToJjgH00jd1of7P5xy+FNjkWVchVzpLk0bbdbo
9d1CwCXj5nbXlCAkTjI3lVXBWpSIlTMlG33964AyzM1qy6sAl5HlBhLhOIz3FL8oRHRHkWon0sOg
OMJhz8Fyec2USghN+iV4LaLuT9TeOat5Bb7sQ0WoSjJmrxroOjJioRm12gLevN//ly4CGSYZTfCf
h188dtcyvGbEzYWLO/a2Hrn/Xl0aA8cFfLqOaaxey976OOU8ByKNf37htFRUy2ITdCg9tCscZ/M5
gHkJcVtqXrkPPGQhtpHCm5z1r31pWXnO+DHik36UHr9fpVYJOJdVKf92ljYUyfoi+nfMmlk8vKU1
WzVvwcM5K1ncaGpCGyhL11qYmaON0xa0xTV02PEWXnBBjCmQ6gLlzCAtxCjvpb8nwFzVLF8xMrjh
ZJMqA8p5MPXTDUhJ5fCQfGeAvZYFBK5kGryud7gVERJ+euhpLA+5roHrb0ZldrhCZuS8kqklP2yJ
yooX9Yn65Fsky0bPkW452BOhwAIdMzD6mgqMACbyOlsMLdEvhV/IySP4F+nB759CCcYV12cv750G
K3z/wJENrD2Wg0h4C5pBAH5/PI/kYw7zeXZYCfPBNZOv1sZqgp3/7BHv7usXEKnUQFL0zfBYt1tU
1bHnhUXkX66m097iJQEkB+GPEWn7dgvfC0K6iOyiyci8WVpmbkFxR9+YD8FoQtfgoeJ6GWv+JGdX
p37t2cSW2SZGq7WGBMP9R+4QG5ilvJvXSBRLU9iCn9321GvPDFRQJRWKOiPUNjIulOQ+mzzqRLO1
qSfVncKm3cQtzpbvg4oW4++RZqVZc/RDjmPfIFbOfhJtkvIL9zSHZDcd8PObSpdNIyjMWmFsC5pk
P4ohNhtxVTxysxYevcayt+cpi0y29y2N9nipH64SuM2/RlxhSN3bIhCRxTQ578ZtZxqmAmCcLRln
cHxAra169OZ0JMwnnIckkEZ5+RU1ek9tUG3RyUBWITEG1HH52DZva9t7fsBiyPy5xRi+GnIGDQRL
AMjWs6CBv5lcSKFp071qX8t91efFgwAX0xkLk+Sya+fhav+kJqZwdeD0M8shEhdY8KGLSxMqR1I1
IKHkOfJe9tmFJ2zxkalplVttkgomU1szyJ3fkkOfUm++v2iwb/1Xg9Laui/St/Vh2u/aocOuM/UV
axUaFgWIs1f4GSIaJk0k7fLz+5Ync3Wruht1O3t8uE5YeydBB0oRQgXakQ9iyg4H4Kb94S9Vzr6K
qmmSg/gFQZYqmW1LxIpLOwEy/o3px7+onWgL5rR+RJ1ywXl3hHBsm3W7jqQ9anOy4LxyCavm2U1n
WhSPeZRjH24UQAM34teT5Y7cxt5aKuy9xOa7n1hTBMhCHOyooi6+K9oD6cKKo3Ync/kjFEzi0ABE
Vag6OwB4Ip84LQ4mhhLfS5rcKV4nlpq+Xf1xW6SN1Z054xKWNkJuxb9nTsz0nb3X4onRUhkao6RV
3gXJ4JiD7Il0kV/m1ISTW7k2ImtXu4rReRWQos/QgQBIIaj1wYCryc4ivzW5ANVj0zWF1kbP/o3x
jE996/O1x5LQH1vecvy4YNk/hkWPD1WQ/d7rjWOSac1q+tans4yrgcMcK8swOrDaQhSOaes5QAka
knGXEb07MEjlOqVjqr5XB8iaHnx0dSq3roMej720aweM49ZE+CTd25ZyfrI2IAXPNifsiCB6Zvpa
+nkfSJx7unt6sr1MtbEk+NqXflknlSFdkRm5WA85crXaUlvODRac5ZbPQ8PK3uWRzltvC8Kgd4od
bItK/vQeAcvlpeErJaZeE3eBqi409ZleaVc2fGSJKTJWP0XyiaN4+6Dc4fxWkYuCwGso7Xhu77Ly
YLnRQ8aco1gOuYTZaMpth4kAuQg7nfQiBxIY2szGrE5yXINPb24oFm8LRuO8SWa78na+f0U2evMu
wzV84hfjvHUSFpRmDdAlvs2cnkVdUKcmnuCWbhJVMG/Y92BUN5DMU9kAcZSZYxafgSMLpt3Xqu1M
1GpaiYsbpCn01BSAauQIIGnLuk/nJipN375AMnty+URi4bJAMgAMQCOR7XboQ07iecdI80UHuKVB
W09c+RCp7e70ghYLNy9hcOcjEx2jrfCeImm2LbSS3w1kT0IkeU1KsGUf5uftIH8/KdwzouXYQsth
GfulTGzMrUa0UnRXvq19+EuoNqfc4Sm2XztzfuLWzIOU4CEdYLAtyVr4fBqjpz92q3ttlIM1qPN4
nZFf5bUYoInZcyXRk/8K7LkI6WcQKKEF/l81KsIJBhpJ7Kxqij7HxRGzJvPDMzbLgjImhD0U1poR
dQAC/HdL0wiGu2GvsazQPvnwpgzi2n0xVkliPiWJJi6g30E9l9sne80LU0UaQgeFFXqhGlpKBnQP
igAOBGPTMSiTKnnPkEG2mvySEQV+uZ+cvWmHCpEy3NQfnkwlLqREXK3oPB6qTfxd/jUMz4/SvdhN
AV+DWdRJSWgMOTylxcRzXnsI+c9FmXgkuetyH0BPeImKYWZRE/4gZRpGyQsfoDDs+AEWNtOcO/TJ
goRv67k3+Oe/AQ8qOeXvEj9fqUmxRLrs9HD1BEAPKhBVaQCmlWZ6xJmXq055XKhykRkZLrl+eoii
oM0J5xPvxe93b01j0TbUcq5L3bJlnHrlTlW24o8Csed5n1Y1cQ/k+DIMEgYQIOY4+z/ipu17A6Fk
No0/W5md9y06K/0T3TZneXOP2eMq0oZa8XFsah/4/K8hro0WyjFB9pe8Jy6zvWkWfxw7BLZue+mz
DsSWsQaJeI8jN3deU2ZPWrdDwe1dUdYx2TZI9w/yEtJyWbHhaz/ZqcGoTEEyx/7zhLPzRIsWL2HY
B7foGYjurm/BL2OQtqdAeu/IIInUk9KKEpvcFOjnn6BkwPB/HIacQm4veFDBq09r8MIcU8gZYNHP
AjAKaCUr8hwNrc+7hV71CEg0CbPWUsVBjiqYYHsLOsuQsxF+bLTUNd6rd0ppLb/GV5M6wO5teN9S
VzalmjAZ9JHye4qbnBnLlpCRIEoC0blp3uHHfZ8T0QZC0mLhRb0raQkWce4tckPfR6dSY+JY5Fj3
TM9ahOuLiNDxPSWjjKYXnur/9oJUp/Df5EjCbhpaOeFgHGcEjozI57AoOisrNPlL77uNowH6wwX6
D/U5CEJD8FSR+TAniMB6nSgbWpJ/IyYMRwCGLmu2/DUD6aoZLnPj4xFazAw/RAvLBiYnpf9qbKco
5G/UQ1CVbC6ciuA1B1FBxgqVX9yfXLroZ5ItIydLr4tzA5+woM0fUvC37KF1vsYU2tyuIVc+JiV0
w21QfPs8TzpO+OR9lAbFc3xgJSY7fwgM/5zmz01L3vMRpeiwQn6oAJmcFn1Y4xCY6jzxJdr6U+1J
lQ6esEPrGne4dtXbDQM6/vgFbDuGLXcWHoUJ4Cp7A9UOm3Bb9I/V+/JbkeBCvqDHkdyYviJI5OmB
q/VJC8rUrRY2BVGsQITTZA9ZbmXu044cG7XPYievPyg/SFeieRsfcjRsBLZLJoax0iKwe/GjIuUN
5Jn8IdWv0IhO77cF4O1PRFRmLtO7omFzOb7QSk4Lf/v20uOWJynnRWzPyCTXUuC16HiXjLmIif9H
ynBOWZ8FWe5Si17ru9myJSBO8fE2oCp5wvUrwnzRezwsXr/g1hkqVLsrVx9lVl4uiYrNFag+7EDA
vqNUdDVjgDqqDulpCMkaokK4BCMnbkIB1aGBeB2eHeWJ7N39fouNKJahTqACwDx3q1fCupPPPDjk
rl1FWedtM5xxphRtPtALJRjspgK7eESSxfTO0hsvN7x2/diU4Tz+EHk4pdG1AM94FBtAV9+oUf/u
O/Jfj12O5KO8D7U78yKkm+0gGZxtGzYA+Tszlflj3c0kVSi7OyLwAWfgCXsgTzRH/TPIclGAOjND
5m+15vYbEJIxgMvsPBGLsNs6DHnQVcCsMqCDe1Q0+y9pcQsrcrO6zyUpWe2K4lUiX4ZvLHk6fxqa
H2YN0zr4inv1Q1pMxiC/S8HNhM9piXw+Jv8xMj4VacEM7+KL4A/Z8YZ3SB49gN7f9qhb3yz/+S++
5NVwhbCS6r8AtHHfmoCKZtRzE4Qksw3ywhe3RevaktSrSE6jKroJ9iQcITeH1to0aKs65BInrdSf
sF6sAiLDk9pAEKk1EEf5kimQRytTOOlM6Gx/OPkz1QL+QWzqsFMVj6m2aniXvLAxfI+K+s1JKT26
z6069vAp8Kohj868dJ+pvUJ8BSgywkBrL2fwONspHtDJO8Djqzowuu9bmy+w/6q6HUbVZ+lCmx2N
EYINW/qz5ZMZQdkcLlRCiMSyeLQqV92RW9mhKAjklmxQ5fSsmea+0YkVrZLU6Q0uTUIgQ2MqrrRk
7RHDfC9xjOELRGZUJYTAjzv3N7ZzvhJ80vZlZaE7rwVAFOkOINA5QWNSTez1qezs1F4U9H1bV7f2
Rjvf0rmQDqQG++aLm8gLQbc2jvXF08W5CSQUBwx7GHczmchFVWIy6AU3QGxiiUEqkGXJTFfwFuhp
9qmZDIqLRq6Yhlep/PQ8yzKsh3Io0bj6lavELDKElELQpEIxAKqKM1KXIz17w+1YJyKYv0Yf66MB
1ZydcKOpFu+SbudaBhoyt8xHWTLWXRs8xMy+AXA/WhL4a8/nc3YD6/LYNtL/rwX/ydVB2rT3KkS+
v0KjAtkLCzZUDzEesIz9o/dl8ELPsPz5qoymvMSiQtnxjbiV4hIWKMQQjeSGjRi8ZXEyZrGQFJO0
42x5sUktiDOV1N85ZCDRiVD8xynoLhpAfU5OBsaJKbkf4uCv6l3F8E2YHR86WrzbXb8AteSLmddN
32lO2UwfwM0Fxac6MxNhwh1FKjdmzpdvg40U+LFI1+JtGISki0XVXv23SHp0QQwlYiPHfBEwg8V+
XVGkYn/Ir7sGbLVSKUpunJI9cnUb19l0F50UrWwlIwhrYlOxPk95fZFxbj8sO+c6NHyZyWxnpry9
JVnGfPKl6/hT9ib8JN0SDgjEd25fJqESU9NaY8qyj9Xw9M3RPUkTijxpZ172DpD6iBRJSx7Zp2Ug
MCioLbdcRcM01CndzuQXoySUN+BgVJYUy+Ke6djWetMORzLf4MuQzZTgAkjvw7zRPUH6CX0OObDi
fkIdsD4mgOo1zGQT4kc5Zg6iauRtisQ8u1jfJArNLwrULpSjQZnPmnaZJ24HIgyf8P1Ig5IZkdXF
4+iISFQKX2rr+jYehKq2lbvq8v7O3MLez/aDWC+xtTytUXts9XMrFBJabouNDlMlgllLyMSf1IQ9
eWYofMtgb8NF9nLK4FY5Uo+fOqSP8Dq2hE/RGoJWSNzD7iCisYazUoTU9jHe2xsSpeTgk7bYK9y9
k0QQmc3XlXwdTp1eoZLTx6pEhzm4DvPAXMXwb8tyO9LpY2aWgrPYJfpqJ5GTxQeICW8NVu7DVsb7
xWe1hVCtdka4aBV1DKUVJiJMKLrKaE+OXqxxIMEKVuGup2imvPBs5V5quei44lxcSN3XqZeTeS53
e5R4wk9zdqK+gf7FHjvWc5DMhTLjIY6kJ0T90ezfBRYSRI5DdeCHU2VsVrusXf1QqUa1rHmg7qWl
J6J+q9dItK2icy3C0Tvpx0EPbGgYsqEZ1C3sIfEOfT2QkgU/YrFzIL4jnub912TUpjQrIA6+EHEN
VBs0SGd88A2T+3o8/WiK6FdlBsoptRAj4xDMWREK0iCMvDROv+O5ITDDLlR2DlCwCJ3P2BdhK4hs
NoxlOb9yQ54Fzgn3xdRB/LwezqoO/5cyHWmPw3EZAETNgYs/Vza7a3H5JdKSiNG4hUbJuOC3Vm/T
hosaBcbW2Mtt+I+uKfBhXInc7GKOhzITa8eaXTbnhc7TbOnIEBnxNm3Qw8vC9ipYrXYXmQNibiEo
0oVnnOngU+nLDkpRkdJXwuQUSjuXz4q0WXT1S6VquvGtzYlgwZKkGt1ECQIwfpWU+UNSFQHlXjrC
Aks66LDR0A8XD8e/5Df38KjWZGdR9HLEKoC3YbnJuq91xtTwDcEQt62LTfytmdQL8qoU79lMK2eK
/CTbVpWi1dCgftWHvpyipA85Xwd2UcoWXAVeMZ0dS5l5gHTyTkpafYfQWkS3PvneUMb0qgOE1tXL
cJbyAZrcOISM2SKquNsX/x68ZsFFfOHee0LvzvSjw/zLy/HGLu5JCMc2HiZYUbop8tM80vanoOE0
3L1agGwCR03uCYE2FtHO0sPXbLRtpkde+BeB2vTo8f0SZj6kj/JBQ5EqXgdRWJO7QwUttEd4oSw/
FWdf4hcm5jJuexp3E1gw8W20rlBT8VWibM/7ihuBK0algti8bJK2fcBI0/XkAsIIzyPGd3J0p/NQ
XCqlmXXGLhx8fg+ea5JLy2rGKe5aiWvU3QH+syEgqXRc/bqdwFW5JJbQjPGfODxaBVrx2kSVM9LJ
TsAB7S0EmEwexSteV3pgc4zqtXCu9mH5UJxZJjzQnvUI8Tlg80Rsdc/Nh6FaZUn3Rc9KUJ9MFstC
xZEclcy9Lmha2s5loWybDWB5JfWQQJO7UiPKOdT4Y4xE7rSF44m/B5bS8fCFGEyUwBNGUf04IcV8
HU3JBDVxvxttcKp9jCXk4eEUB8G2/eKMrW5k2c0cdGi0UkY0fmmH3TwVF/122DOQg+oL1SlRsAxG
zIPgfz6ECVNUT0hWMH1Y6l++M0kn+P6fsFAVpKIFz1ji5xUR9BQt3lcaZK6x8H5DGgvUk5QQ6Oye
t/2CdzATvotLhP8j3QeGg3EWJPXErgpteE+Biy9oqNSB5PiCm5G7b0SPRdRPm9Qv4PYiBP5DALkY
+9bSJ1QbWYwE9GJvFRboUOttUHE2gZIlO4xuRHe3IApkR2vSLrnitn7uUImBkKZqjr34uCGtvQ0T
VFDrzNCuq2z/Tqtnfh7qvq8e6YYW6H297cTwW8CbTdj8NTn5aVyrdzIHLvz/LRQj9dPgRgvE7ZcJ
BK8v2BLs5QajwJn/vXAT0UFrxdKINLJIoeg7tD442Z2LUjWiXDycJfO8BfwbYsYfBbVx9RL/pNva
Q67pB80iKONOUthTgyIpL1qTlXGuGc1VzAwB4LFLElXqPsYIvdfRvkz6WdLSPu2P7AbOR4ufHIr8
+Zg6pmsFq/ZY6pM9gLYIzi6rsUe5USpPFYHfK8TxXZA8LmXTVqGOaqHSCleM6j666/4B6C9Xgbk2
yrkbOVVfO4W0KOEjNP1ZBRG8eJI6OEiU55n6n85rKu0/tBhhx4ezXbkVS9YvWZXLmUHvmZWrBU3G
uO7ENaN0TGf6L8TEGkv2
`pragma protect end_protected
