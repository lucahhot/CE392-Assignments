��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{j�X.;߅ţ3n���/}T���. ��I���U1�B1�ͷ�I�i	sԯ�Ú-$H�0ߐ�5��o�4l�a-ޫ"���X4��錵;�ՏT���TnP,�"_��s-w=����V2,���R{��<�����_�ؾ1se���§��-������TW�ե�m��m�AP�3�Og�%��[T���9��_�?�&��,X�MSH��iR�6J�E��ă�c5�+u|B�lz��Ļ�"��������KnĿ�(��ނ�v�YS��������,סNO��.PU]����2TU��M	�yB�;y� �m�<��pT����X����3J�K~ڨX�M���2vS�-�!�1��$Q�Ϯ��Ǯ1 ��$#��si�����G��c^v:�F;ێ���к�Ftk+:%auJ��P���kѢ��� 2�ڒ��C����iI�j�����%��S�r�
ݥWƍ��O�q��l�u�znt���/Q �_���&\�꼔PFæ�S���7a�tr��Z�zu3P�����r����M�R*�j5¼k���&�C:�U��f�G(�����Z̊�I��/(���ߤ�k��>���E�b3����F��^Z��;�x�gi��M��>����m����!�@��'�>55�I4�~{l?O��
��B'�E�.ޣ��p�q�wm^���]�➲�񷀄zI
�"�j��jF�4��^I�p��}W�	��,��;�Y�OT�B�-���/�'�8 C�ÆbՖL��E��9�ڟ��>�r���JK�_���r��r��Ұ)o�ow��_V�z�X`��'��|p�3Q�º��RlFҘp�PU�x:��9�T^E����n�ff.�=ky���L1(e$;��`#ȑ�۳����jv�Tg��x�X^�l�p-ޥ��6�?y�<���U�I�o�O�l��:���c�_y�b4t��`����ORo �빜
��U�Z�a`
�_��i?J� ݥu;k��Z� ���6�P۟h{h ߿v�/�����R�~�k�暩��V}�ȦZܾ�-i����%|�70׸��<}z�<�I1����]�aN,g�X{����9��j�s��-�(�4Iߣ��$R�X=�N1�z�!�eB~�FL<�&��zI	%W>)J3�IG9�
7!|���>��I]��`֚b�뉱�zv?��H�>��+��� �J=�@�5=ۭ�L�+ۻ�ۭ���.�iW(�)�ЧK�
Jntv��s�ʸ��8T���"�w
��lX�� �@W�G��E/�W#:��h������Փ��p�3�f����u�M*�̴nH��E�Я�%x�p9��J"�E�Fb'�|�}O��2���(dj�G5=7�����d0.��N�w����+�Ŗ�=�P&J�2�>�K�U�B��DZ��z(䭊M�(.��DˠE�ʫ<�}/�;M�Ri�
!\�R�
���y,�jW����A�8��`�N�b�S����D�C�y�ؽ�y�'M[�T:)㮾+���GY��b�E�g��h~q��V�
��N�}�����W�iY��ZX��=���]7�L�&DL���z�5�a�a0x��Z�.6���J7%T4�^���-Nԏi���t�M�KGa����ڵ[���5`X=�1G���.ֽ�uv�8�aA���m՚�L�8q	�ⶇq��9�g�=��1��0D�M��uJ�6�6T��J��)C�ՕK�J&� ���K�g��nK�n�|]�~��A�������k�'����XҲR���R��[?5��զQ	%�pw�/z5�����/\-�뇼�U'u�v3S(�/�c�*h�Q�FBP�9>=���b���0�~Z0`/�<��3���*ׁ[�aG"��t��s�is��S�5N�l,�]���Q�)��j�An�.� quj���0�-�r��c+�G&��D˼�@��sh"�<T��툚:�9cEA��o��4o#�uR��yC7��}2�oWz_o�bqn0"�w�?Nf��ŧVT�UTK3�
���I�����G�a�@�|�[
�B�Δ�j�~�z���G��0�FU �{����:��ʩo{y��5
X��]:Z�`�u��:�.�{���vM�)�t쇗k+���{���6KL������^�ֹ������p�gG�C�~�y:]'��8m��!����%%��s��>��mJ 5J�[ST|�*�_ٷ��aT��C^���6�/����9��c��mM��E�<�'����~wp�i�A!���\ϣ'æN�v�d��i��?��ȋNp������=*�	�/�z�@s)B�fJ�H���1M��f��"��;��#:��Jq�=�YT�Y���%�����*�&(����;>��w������];���["�C�4 =_�.�l��u1�4p�:��Ra�Y��oې;�;�$l�Y�C;�+�#e��1*��s�nMm�<8a�����;�
�5���ƣ\آ]�`���8B%�4��"y/|�<������0�lFt~C��!���z�K��M�]�_�J �]��� I�},�Q�F�$����%�Z-Wa��'ƙ�����Ȝ�N�Ehfk}�0�Gk���\0�QI<�ד�ؕ�Pk������"n��Ǌ<*�Bg�U�#��3���{z.zC�câ�`X�u^�]�d���U�V�2�n�iFKu(�q'� 4q���.T^o�3�l���"�UI��+ˎ��T���f	+牨i�iu� ,R�c�\ą�SՅ?��q�������-�[1[t�ק���xw�E�ǻ�����;B���ל��������P��$��%�᪕s��}܇�F?K/���N> X���F���m��h��z)hhҋy�Ҳ�X9�}�pUt�P�b2���{U��J����[�f��M`+wm(wZ�+�u���3.��d�Ƶ�Ŀ{e��mF\]cU�Ҽ����[��<������]�"W'���\��^Ҧ�B��m�Ռ�Ц�����`���:�̠ws��yi��'�+�yi����TKC����"3"�9�"�y����R��HJ_���d�I?�������$�(�T���ZC�QcEz��k�HN���d�3O�S�o��I�Vv�jv���V��+9��Qk�ć��Q�:���2 �,)b���Ȗ�I�͕�ާ	^�_�P�5��˱��1|(�V�S^�a����ek�ۇ/ &Q)xMl(?y!DR��1��u�u}b���-���e��}��^�i{���j�4s���͗�29���s�.:0<�^ٝ<��͛5�@�g���*�3=g� �����J��=�Vէ[�?;�9~3u�����������t!��#�Xin�Uk����,\�awB�S�!'Fb�� �x�;�������xZzI��Zֺ�2VՔ�|��~�,b��gNaa�f�5<�z�6J	6�_[1�n�{C2T�"��c��q�r�!�-}}� �v�)o@�/S��x�LBc�����������7H���رK.C�I��'ƻ|�H,W\�gl2�4z���zj~�!j
6%�I6���]�����@�Ҿ�Q�:������õj���h�!�I�?.��YX�u�fH��t��eI����8�7Y}5��!!#�U���v>O�`��W
�U�}�=��+$���1Kr�ƈ�^O%E,]l�U�a�r�CF[� ��/ސ����Ln<���X�a9�����/��c�2]Ml	 _�MW����L�ߎ����d��KC����ߙ8PNhx�VXKQT�xX��$f�'���W��rc;��&��&�rw�nS�Ɂ�J����WBF�Z��D!]		hȱWn���zC�ט<x/�)?��F��R��~U>�:*n�8�K9�ڸ�06I���m�Ƙ�`�S�R���N�eB�_�W:�w��u܅�_5!_:��JՔZ` ��JiQ0H�g�%�vY&��+I��:�E:��{p��nWHH�Ѥ\i�������ƍe#]�r1�
�#���@4+S�j��C,D`w�ڬc\�?�`*trWR�@$�߲sf��{�^,R�6����S�h���\̉�|y�$z:���ij�hgo�TV�pX�$�����WTв�e�qNZ��=c��hʤcK}G�LڲmX%�}Tct��̠s�g����6�\�`�ĘQ�F���Ԟ�T�?�4��>��}���s$a����A�W�����y��M�(�����ٍ`/���E��cw��@ ��U[��)ԧL�3	����%�-V�;�������N��6��9g�S���N�P��{8y6p,;i,4}�$�Eg�{ߦ�};<���'&Ӻ���Lg������#�cסa��M��P�C���f�	��,Q�����7�gL���٨A������~_��;�^U��2j������<?�^�+�j�6�X�:6�bV�vg'c5�����5�\\��[�*�{W{� 2:Y���e��ˏ�F�xpʳ4o}��V,xQ��г��]m�y\^��ۦs꫽���l(�.*.r��UN�$�>���Mw$?�l�uP��uՑ^�K	m�H��i*T��yT~�<��"��TT��	(E잰;�A�@�
�'� J#.:�f�:��^f�2�t��-�j�~''���v�囊��]�Z��d�r7b>Au��W��=��W��4u���Y���#	��1~���c�d����ϒ�@S���1C��ճ&�@�S��6��L�sW�D��ҋ@��)P�;�*�˼+�s��4_�E�j��|I,��o{�����P��u�1��MTz��t�4�s��t��G��=�
�P�ј�����e/հ;Gĳ����v��"n)�w%�^���Y�fkǒ�����Ĳ����WW������t��ނ9Ž߂=6Jpg��	��?���Uڒ��U'�-h�u�v����`J�P_�9�U�w_gU���~1 ��.@���HE�_�ED���z%�Ž���9.���K�*H S�f�ξS���L��[��H�EF!��"]�JQ��� J��%}�m�(�O�WLY��<��e+bA����4#(gɥ`|���8"��B��=c���/��*���|�-���L\�G���Ʈx�=6�M�R%��n��J�)0?��W��vO��� �)��_)A�S}P�Obg�C�\�҂\_�klԙF/i����`qw�x9��/����<*�8����'���\C]n_FK�zG�
|��Dh��ҽ~�ZNt'NP�k^j"*m��L'�E���'-і�� �|1��X0{}��7�n���8$�*�f�?3�\5ҕ��bv��Z{��0���aq��w�K�{P�`�'�F��3�"Ֆ��]�smx?r$;���A{�)e�À�u4�c�Y�(_>o9����