`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lJmFCnt6FUmMcrR5Iymg5VL373rA/HPhGHXbxW1vGrj07cJOkv9KIfgcyhvq/uSI
ziFnGn8mIdAlPSP/gBANafuAIPdFpBGVkBOWM4AKO6q79YwKtWsFyAcenkzhIBvn
1WgnRFeAlMWKWJBsTQD4E2eBAHZ8ImtNTGCTKwFRCSc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8400)
O2DcwildLH3i+oXx/T/gy4S/vpkk5idfZFqnrrfh+hAodYvOvbWahJL4mSV7ZJZ6
YOs0wgO/ZVRj4CsYYla2v+DKGu7V/HeOQfGnPsnItaakiymJ9vYip1trLdI/jheF
3UtEhkNIqF1ZYGgiSp9vCbrs+NgPpo4671WAgYEbPHnYPlY2BHHUFtOtVPU8ydf7
4DgYJviVfIUWGcMvICIGrikU99M7wdcJ6wns9zOwiQ69fdNUtzYcF7p8omsuMc2h
+oQ2NJvkOXh/nVgDmPfWtOG1arxKlXumD5W7sVrMdGRk+TJ/w13S83bbnMupp803
xSuwAFm5cFYcN5YFm/mc3zdIRuwQE/EMD0Y6XtJtm0rXZNzSJ+9MHCXi3vnk31WC
KzPoE6Uou9mO1InUGHuejelUOkb4lcp8nx1gubn0WZHiNl996l4yyFy9WW73Gs3v
MTuTBeGo3k0+8spEohLFcEYg4qqgnbSid1Ikyct36KELimNFgzypDEmZKtufjIex
rn1Be7VUuOexqBB8u15spGGA5dQ6Vs8ar+pJzm11wfxL4xzEzrS5LeDt6cMgLQRB
J9Xl/zvSyl/KRaoE3Sib8SbWGtaQsmDJY9tvnBz1CuB3T4CNi4bRG+1lX5ej7oko
lCIkoazk4/zww8U4OZaJiPYB2l0dulmQTJMZ0F6g5r0iuuYi6fSumSCpwcqcVK/Q
ayhgYybl9iYZZUe67+vAKWyQMKk8n5AmvuC/vBRoTTOpJVMoYXbcFLh5CBlNMigX
CHgoxXqiQ5ur9sNna1MCuSC2ruGXWZKDjFGmPJQ3uWxph9HIydgTBLeoTYDTaJt9
tqL2RDYIVTxJKn/v8YkH/+Sv98sEwkCr3RwU83nFYEZpsl7cxrmEBONRUdPNqmQd
jgp58HcqMgJgawvDQpjysd7rN2CVlGcpQuMSyqP5ILBI/DjcTkisbAXRJoKLpk65
XOL1FClDWxrf3UPXeMoTjJmxjM/eHubTd3Rw+e8wEiIEjpYvLEbSrP0LtyKVJjcg
Wq7vXYdx2EiKCwEneyikuDonIDcHh9V4cJ3UUvVRU0Sz0xS8KnyrZ67FGy849NN3
4mi2VgYGQAbijS91yAvID0LHmtLPOOINZbqtL5cvn5jFspCXsfbQ716R/OXlE5Me
yrUf33F7Kw9pW1yBoPVRy92rw4YtW8qOihKropVI3ogULNtIzsIS8oKgM2BztNEM
IsHtHVOdw1TuWkj0ORpSoe5LTIHyTVnFG2QH/+tCcNHiTqNnyJctbFAOqH3szCG+
EEXkq5G7RQhf9Qtfdh+a3Y/Q5HojVc7+TDff3rvMhiGy2/3zkSh/0BVL3lWfQ10z
MmTjKQjHroYy0KCeVpPcF4JTyQ2ga/RTTGez8ZGiZrwAHEsyx31A473enRIVJvg4
cyRsRjZILyC6JpFrEvX3zJhv5+dMYZ+Icd7VcnL73336wABdPGCc+zUYvNJLZdqC
DG/drMvmBtLI/zUrCvKc/fIoZNg2dqs4tdHbJriJ3Onsq+uQ+dDuVFT1Mdva/Llm
3XzfPAlM2gevPdXwKa9f66909/9oMaQzEu6inREUSzEQ6sOK2MmRn61O1FZpG24g
JYKL0S9VP6mFEQW2DfIneTRb8FG+glLkoEqJDNmnqLoBoeawXmO5Tsp5DuDx3loo
l7wSivhv7Abpt9q42XXbrEaatK0jTJRRIgRttcsLs7qUdXBVZHsqjNX8nUWsMCpw
+E4YdVoP+0h1A4TDTeBHwYCLkoUifZ+B3HvMzi9O76QTLCe2YQPbajvA1/mJeiTI
kwuBZiyFEhnicotqvippblk9RbdykGkO2XQdHUyKj/KF6ZvbB5mqFXwM8gedaeGY
gAOTPomY3/Hm99yD/DlTtUYtqUPIB5vD2PB4rNHF2TX3hCqTSINHLG97Qse6Ry3q
6ImX2FIxD3AxMI8S+/B8q4ThSqCLbAgsX7Ow1Zstf3u8T9na7EeROZD9ndIP4D3l
/4M+YSOzN7x0vMnX1qxXmM9PFa7vpkbrbcrvYrZFiQLFgjf0FyF60WyEAyxamaXE
rvyRBXfMJRXcki/HoyDB6k15NXggBkdsWjo95s4Zb1OE/c0zZwCokdfXVQapVJeA
3qwGgg8xLCcKjlRrwAOIow1gLHMhcqCH54nC5j5zlsYf2ZMtoYgKPCEaThMW1aqz
Sa0vlh/iM/Xp4yx/twxSra/5sAVAx/AwwuDH0pxELCy+y8S1IlKpKDBNbhBYeicL
3ljDXHYfuhtOIQ3u3gSy+7AkhIZcbfw6zzR2erodJW9/L7IvjnvNifbST316yvl0
FTXvYVA3hvzJo1moto9ERtJe3vJVsKAKyw2N1WHlzqSai3gIjXct2ACSNvKL8o1q
LD5RLB0u8QjmvG3CBafkrWiQzu1q3PNpdopy0S+4tiMNY07II80pCerkVreAYntO
86C7kgmtARRyOewsRQ77VRc0UG2lVqc6aHewZiZNKWmxTAVP75fLZ5g9yWFmXq7v
SmpNuavsVvjQQ75dR2VKSslgyG0SHDE0JBxj03cUEd482t3Lmem3ZDbmRvL9n8bg
ay1gKyLOv/o8Es5z0prv+Aw+FFoekiLD5umneoJJ6gseiB3w07U/bUATCKYqLLPU
+SYVA5gYX8LlNFWRs8Ylnd4R7YBmzEp0knr1qMMR5+aGW3xo9UZ4Oiss1MbQ0VU8
yRcYGCzfFCLunCHZJaJ7Ms5gQu6Pb3k1FxvEG3DQ+Bt8xe81Vaf33q1V5983J0Wp
1dOYpj9KX6Eh2fUZzpmOk3S+0LM0pIQ/kdmb5nHselHE28DqhYyYo6ENDG/MRXuW
kaMjmSJudWOm1ptHHYHtrcr057hZutlbSxfl5TrG7JQNhuma2/l8d0e6kImZQXWM
SEexlOyTxyYDKETyra5VdmJhT2KqGveE78GBT8QX2985QOle/Mggnrgdl07qa2N4
CcI7I/8npi6VmJvxkLpdYvGfJNKwLt0Dn2X+UcS+1ei+/TYgtaEOKlnk0JQ595vb
MvZBMA9JjosSaQXAzmW3wO7xKshmz2XO1QB4CnCdauXEWSbjEMr0zIbT5Sp3L4Eq
BmSvq+LL5m26aa9qgHBMht2SWgLmlbKE8JNHiY+ICkSHzKdw5yHjKHJYmsQb3EJD
aSlEwul1JokuOm1I3xM1OIBGEURXOfJoMhzZy4SIKNaWYJhIWo2/s/2QWKXs3vua
eF+0GDcWt+PI4da1iTEyOK5j4Esu2GGlvdz37atIugbAECH1OvLyEDic0vOmr5Vv
AL6Ju+RaxcWBxOnqFuasRMZmli1Z8mJcHz1DKz7XXEbDBPsVJcbH07h9OfrbbyKv
6nS/Gts/az/C+GbHdmdQZkIqfcpbouJpuDHxEEhFn0LRJA7E8/7eb2jeKBVqNTDp
RkURTvn4A+afkq9wlGfODIYd4BuQno47zmaHqds670Llb2BCoZ1Wm8tkhoMRzUJ6
4yNPA7/M67OEfFSaRo5ej/TjtM56KrBtd1e23/68tdqe9ydrKBZ+1oT00J4MmzXM
QRbDDDr2g2r9BOdkxMvmelH7omumi96e8qwoFrkecUvPzfFqbSXLEf83osXWGbo5
X+r1g/aouCJ5QyapjasaN06gBBUnYoyNOZWwBmA0AQIPZBwbWsEYzi5YE6lSVTZS
NzLniGtbj2gowZNg0sQ5c17tvJIwtMRj3f+TjoGcRoVvatj2xNOJJqY7AqkXnk2B
tId6Dxfm++iz0giINi8m8gdjyNesBrcJS+Ai8ZNl3iOE6xghrtyv8uZ+fnVNq4/I
o6JXUuTkaFyoEZNhyamiUMdJw1vmQSwsgxwCcxLltyibZ4+pK+N/la3fxUaEqM0A
fzMUkzvUqlvSw+J6mx4AFyOBXVo1ZTHmb6TayAPUKzJ858rr85hELGPK8M1AkYe9
6zfFFgcKMwe+VNUcrHabeltKDfwK5CkNyvcwk69eLngmOkMHbPJRffO5LdmqJPmx
UgajWcXNulrfWF7MWqAbYkhiDv+ErPpROMJvGatKpb6fxzh2gRdxZSPnm2CHtshH
NxWG40SLzaodBaZiyv8VOsm8v7LYNr9D1zaMyvMrZ1mJNayFT7WK79Wn3npUD1Jr
M6zKecQ/VjTE6ELRpUvBgQpoLfk8BGUxaKn+UoKHCSfT4EYfv3RmmgIEpmXG57RV
QaW/i0HD2Q9w06C9r1EmtU387KJ74ErCkHByUtGi1+Nyj4UFpLpiI+2IMMdqo89v
4Q6hHqNFYxz6hkXqcve8Cn1v93+2Yv4TKf8sAq5va48N6zAwy0rtywUuKSv6IPKg
Fu5LTeYlQqqAvlbSsXtakq0ozqctQEsdZS9LuIO0zm+VLILgY+NlRlUPkKiNXKhx
j+lJas5z5DOJZeJ/x55Y9eV5SU/m9NkoqT4aqGzkb3tnqlCniJ51Xb0W+8ugMzpH
jzqRJ8oVl+O4BbP/eULqT0+TflwC320qUchoFfFCsT8fByk3mqJLSCASni2e69AD
yz5OJNnyrlNZRREAOH3DQpl6XRlkeuzdcCoAeJVgMr6e48MJ8zRH9P+O1A9I8mhk
f/busqBkK4HCL+7n5pEdKsZJVXezU2OrP7rYfo8c4Uve8DhdD84ycrKi8cR0mR+P
TfEYxZsh0tUON3obF12I8/JuNC8x0R1xd3I0VpbkbalXhm1D5zBFEyQc+skAktzX
YQoyeBj6kr/jq7kXdHAxUq2WnmghfnWaq5ZorPTgHz1YSqbVEVF+V4UFRoGeeg/4
Xppl7CPYKXMmwTfXMaIWyN/oaW1+5KQJ4A1EoXwYAxRQ43vww1Dan+gwQxzMqQjK
Ak0xxo8Iumu3+RQxp/9Xtx/LMs6BRVReK54VOWnBpcF0oTbMdCmpuBtiPtGIUwWj
h36vQfT1HJKB7EYz0Qkvl8eXVgTTOYMqmnLuFe7O7zXGO96XQZkFfsKeMjnawHhs
kGOFy/G+ny2lIgYhN8piKUweKkg+Qkt4SCxMfYcVJ3fg+k5lzKvx+yTgXPZLfL1m
ykU8MvchVduZ/P4HGj4ZQezPbEtTNdvC+3b87z4CBNW+iP4lpzEz2wPgpopYcPL+
ttl5ZhSakwlRLas4a5BY1OG56ubbbLCI476cJB0ZvISFuKwmXiMfM54E8ka3lWS/
+kcEvvBhS7GAiRMC0/qVjDV9ih1XSgop4En/9B/H4MwKc604UMbNguntIDhJbL2L
wfUf4YFmpIWqfzAdIuHRXMNOSwOlh7Rhndib8I466wzAreyB2Vmd33JdDNqgYDrh
fOVppjKrzbdG/FzVII+NfXojRPuN5Jr9t1JCUFOv1Qeji3PQNvdpwj9a8f8ztq2R
9Y12UzYIYLqqa07FoFgQ7N8diugIsOMeYsB9tXB33sy97Rbw4ATdLMzSdJc/5q85
yWsRl0F8ccswki1Duo1S75nDqje2ScPQjeavh0k6QwYuF4D9C8jw5SQjMyfVMNH/
WiE+b8+8D+PblzshHPJzZBY3r3GHFTe9NLL7LyywboJ2Tne+Z1E7VUntOCyn04ak
7LKxOTaXneo1P1sfNxZoejdmsDJJIobCV4hlheAZHj9KpMRqzo5+L24CJ5Wofmeb
rrh0qaeF4F7m9XxyecIjtCxuzgnCsin17j3XSr8cIGaqqp15lMQM/6o1Ab7JaSNY
0D0M8fKXydDeaaa26lAUsIBF2WmV3IMG4N9cy0ihmmPEEfWb8cKa5pHvTUQl/VWx
tkg9SdiLBNenTkA1Und5rYfJa91WWdrhzBA33MSURM9si3cJ8Xbqrjb5PuqFQYWM
6v1LLutLeDe2SwuxnQkzmDlVTN0xoIB/B6mGysiD3jXmoNXGOJ5WOhnngUYKnwUw
ZXMgA9ObJ7AkSsbrvw5ct23N+ZXeBF3/R/uNreDRyF7jO4xxJ1RROg9Y1p+gLVjn
5N/zj395EVXNbP4TIayy1jFV6aEEo0ZPP1BtS71+gddI2UurCE9ypTYb4HCgm3i+
90ISwzWoA9ghTqyO6sTxDHe2WKktFC0OxsZL9WOXa9cLB8+oThc2HkfhV+i/L0g5
tX7O9/cma152oOeVm/993UgaQUp24/hGm1zQShP9X8ja0zohRxahtQ/0bA+0GdMd
GK05/OBTK0FpWTmvs/FQxBgBBO7C0Y2tuBPJvz/xrquxr892mi4BNcP5lF8ihpSW
D0WYaZ/gg3iSnmkG++AXFYiIuY7W9sC0yItuxOSOgPtEGlj5X/9n/thbGLwRDaUe
eGXH8du3jxKY6jFQBTrBjqMKAt6Fgy8X5ylOEXVL4OwjkBOK0KQCSMDaM64Nipti
ByZcQ3afPNy/0ecVBNAhOU2T/QmB57OTqUXn0xrfSnxFKooGpMtd2WdAPYZlwVCp
88WuqmGfHkd2PtFfQn9D2w+Dn9tQPBn1wyZrGtrCXkFksXYnwmtwMFMNKA3pYK7r
GO34JC1gal+B5cqKKewHs5Eg790AKJTzF+zV+YAcqnuDPLxAFkKxYI+7PcyeiKLl
Op03EvPqdPoYJ/QmWWLopbG9seqnb6ABAMwyJXWMR5zrsPQwHWjOc0k8ujJlFFpR
DGxa1I6dmQSHnozi6prhViWg/wE5mmlKl9bzvj4HD48U0gyf//SYTfej0fom/smI
E3k+/V4CHWlAzfDY8k5NKes6MWzfAPCApif12eEAifHqCNkWyuDb8aoTmC7vKByB
1drsQvFDjXfQDHkqsJg12+0K3885OoCtI0gR9GwiSrx6d1+EmJhQH3NXiU0v+Dlj
dOX2scYXNzlyvZoXBMhcJ03arWTCimPPxtS7Bj03gIQJWYDlRfcar/ZFTpr1Gi2E
NUD0s7zcyNCQHw83Z8mjXobO1HteaXZYgayWDeFYEUaMFpPcv3v2wTjuaUKM/lgd
0IMvD5cPbhY1ieJiiW5bi59H5A43LmtQuOWl2H/68uHwjeaaGduKs5aUKTsxT6TV
Jj+1CCISYG7xXMVY+xSj6cXp80o6ntyPl+yisOw+p23eQHxwSIdvIfWt1YXp9Zxr
WsCWQWi5yCz1LzXC7HsKaCroERFAugb8lsYdaiDdZZKJRnmUFQGHa0nuM/UQYQza
5U+wzqfvqTx8kawuwgth1F7ySuzGCFJaEsc0LahQZtPjxp/3aAp/DusxSLfxskNZ
oeJxVzCkuB6589m/z6fG1YZh90EodedLgkfsOZMXfJSV+yAgnCvFFb/pTJs1/z2p
UlwvZnY+VQltPdmG8bU6a5AtEjhEtkchLfiAe8u536ihG19EM89mRC6qAiOnNhvm
Y/JVOnYUqQtfJmLuCAwc2IxJu61j8a1AB9NW6fQggqCEZ1JAyhBttHLiA2XP7tdQ
7xGWo0Lil3yLjptss6Mm76pB54HOAkJUAmfiT8zKFmh6KXlQIOhTcCCgYzWFyeJh
NVa5IwcQbqBn0VBu/CS/1YkhxGBJMTKL+jn7cAGcJy/NshW2WVpySsYv96mxhlC9
Kt/VnJOvf2FRb2XhVzzsYs0Hr+hcBYtbENPvYgEVje6UYdmC5cyBD4K8vKPLMw9C
v2acm/6j6vRU5A5Hp14m1c/qIDcPEubRUeV7zt/WPe5yjl2lJaqVkX0vudQFYKcU
sw9yTJNbMl7cW9ixhfIBZFWx+4yrgrrYKSYppnZrJSEqDgXHNNCpvBVFPausuLuR
b3Q9F7Lp7qxvjC9et6GoXpiVEXO717X59G49Ot5vdYyY8Um7igrvUGkoMfJG28jv
Gq/TvwzsDDmuEiOlirVlfcRbIki+sraPTMjnlToe/jgoFitgdULI+NJnXKlT+e57
NdesfGZHs3MygRarD7OGbx5D4RTeCV+1LZuWEXcPst1/r5lklf/UkflyOu3LaGs5
Rau4hLA68JOrNzPqjtAnmDpTRAHrvoMqk7aTLxCJUsIqM6IVAS16uYI2fshPqA9I
uKcg1Lim0rdGJ5RL1FBDXPLay2cVukBLWcBXXV5O+zdL4mmlHf4nsH+Wkwm8oTLV
et0UifbKJ/ht5Yh2EOBLgiu0F7lLuDGCHzc8LwClL87Pdtd5rV1JO1Tz3OpVc3UR
uVfaedZ4f5LS0YORshrFz15xVDdhzpvlgksSsMXr56OQ/WGRBffGKNaGt7EKmMsG
G2D0Fg0BGEwPgStgpcD35bm9JKR/NE0x8YE03zW0obTmRK1ZysKqNu7dUW+sBwGe
pxJpzGeNhj5IJgySiWL07N5wNfMcE2m5AEo6E4gARvjtvqEwtQPfyizfhgbWsLMJ
0xFj7czMEyFmvdfn18No7SYs0rjMTvAMXmKVuQ1Sw6XJTOah0sOMYX0mRcqDt92a
p+jvmt+eazxX246EkbZNYd/TwRbgh49xS9Y/elN9JC7uIY4PfgCrg/HkoQTJddT9
vHDnZacqOnPHlFoCyHyu4s4hiqg1Sww/E1LwKgwV8QZgTh3PerQiCNjBcmVUKkMD
yQx/TA+aTA5oIWksoLEsaRjIUiGxK1X7pXIw2KClOO737/bGRp9yzUzseDNTIxAW
NREmaI0BAQqAoE+jb5xtlNLdtYD9YnND586Y6lPr/Sy+8JQb2rAq9ld99e2lTigx
igAkCgkwN+0OJcrokuxc7htPoW5clocPuvg1YyuMJ+O/xrv/OkMU5Ta2RHdyRXqR
m/YuX3MEfdJgMvRbfcGddhKS8Xa3VvANHzN5trG1zi//3dgZaPwt4AnmdmuCq8CP
CvPu/ZM2cNqUo7INkJvehjpvAUXqysAdB2qtTjcS7Dw2UWmP5vk8hpjAOwVKhrU+
i0NXXpn0GcB/NYHWvK6IlvH8QDmf1ybeRJPZDxurx7LxEo9iEQPDqaDLcANUbYzL
SRJSM+NLmOkThHtYHZCqSFB5/7HBxggcFxLIxQ0AAB7cR0mrfxeVhrucrMJhptBy
cAnimowYjQXEJ/fUVko5t/S5g5SO+AyQ2XkWhSy2EIAuVVAdAteuAhw1g2ed5Cnu
iZpE/tttvII7nIepXg5X9GW0Xr6W+E3phGjXqA7vc6M7GZzYT8D+CgBF7UpGKD8d
PyS5fEWjojFV7UeRAyOr5cl1aCFGZJy0XzZ1fiDBdbg0rT4dmEZSX7gHEHhnqqZf
BaxQ3eLw4SAl8818ixTA9SaEjlxjDs2HZibbpul2tdZlllICXZcNNTnesCP8Zjiu
1jxktUjHaYCJ1z4pKeRap9l0W/Jrs+SZFB8aZJPDTrGmpnxl8mnniMJeWwlZtq2r
vmgCVTirf/7Jn1q14Dn3J3L3nG1oJFbG6qgwCvpfp/xrM8tyCugMl7WczePVoQhl
19bifoJTkR3vy5JapnDK/ANcSDrm1GShGNM6X8DLDEiDWMh6U4pBNqM6K52yqWrB
zC50L46H+D1blVi61LpwmQsKE3trVJPQ1w4DZgvu4AnVvUOAGoYA5+2GZHtQAZUl
MJswDZ+8wAggbnWzLWxtIh+ME6jX2TyQWAu0jYndS7n4R9bdKCp8RFjeMH85Ffck
eZAHo8Emxi2SV9vIxNAtd8nskhZeHwOWl36P3V1jCDjhXiq9ckusvmQEolX9LYZM
UDXdd8jt1rDYrlJbECvFCjkA3sityQ2NTv1BtK+Aq0aREdt51VkrcRd5bU7J4tjp
HKLqQ4dyP6/vQ54E+B8/77t+YgkqDhumGqoAlLWum2BHohVU2akK/RaWsvFy+W2n
uqoWg7GnRBWWzyhUFlFcPZiq3SFqxI5uKwK+2RlQVOpV6eFXBxIemXExn/0LU+8B
1LaOY5nQ24CWlaoyiFQxaI6mTCZCQrFmmi2eDIFgvsC+5/ibuhqw3UQNjQ07ErPG
+bEph/goGsqSIoToIG54CuZz9e+sa6s77PjkbFdGCZUamSLrhP2BVVfV6PAj8JEC
gELk0X0MfCcJ+MvrK+Z7qiMJR5mG6s/jRV9MKvZRvK/xLdzFmldsi/vOkAmj8j9d
NUXZNeIhzpxYhLlS1g0LDOL2tybIg9PN0tNUPjp7ygnWYQuIWVDX9S850g6Kzf4j
Jqaw2KnYSmQqyCgO2DqNEq9s6/qi8fZVolYmTOvBau33Ft/T1l4SF3BNDAGtfeWC
CT/Y0uoWmNO0DsHyXCFBbkNB3n1bmQY9YObQknxbD5g1uBhdpNl658qwiF5DAVfL
JYbeXox5HJTH5eVFWyNF+CETZzNuhxyCKAs4/UYfmxtVc41fr45oxYqbUKxG3F5B
hCBvY7V3rrdpspkqSeA9jqY/sVNfyN5y9hFqWpTZfJVVhfTNArXwYbhDwkWSvPeU
3BtqrjBNaRziT8PydGvhzx8rBt2yzWH10i6TuWVLqbMTbWbdMUw/TiqTtZU3in+i
uvxqKmtEldbhZ3KeWKadzTU4HqBlO2Ran6eVmzxUwnLj/Aty+WR63plrrb96Bn8C
eix1rB6szyxtsPkocbTRobqpkpujNufzrXJTbkl7V4/jttfSFbW902mxZqAQmM3C
kMJEQkz+UfOyyaSPvZfS4OQVDmOVgiCGy1SLpf6tqdVrErRVp77OnpYvhWFtmykQ
tIJVSSqiuUNvHgUg/xW85MQ37JjOTyh3TgVLmyetqRLC0Z6wYieUKjqy4BHFc6IR
x0R6JhK0lKnG1E+NSXCwacYU1e2x43VYGGBEu6N1dggY5dVh9cF14h5Uh5m1JXXa
7N+vWEQstr+zyKWVqgFkJQJDb7uwF6Ys8T571RE+PUK25Fx3Osazje19nu5PdHQK
E0Q0ev84eDtjBctKdIZvIfD4/Ci+B4OQoxr3dm2/sIMtTT/NMiqm4oSqnHQ9CZ63
KBqA0SDjmDwMrbb+Xamrtw/TPFGAWRMrv+M51ijGXDE0CTs/BGGFdqOMn+D1Hw04
44UAI7C8pt5q5SgMJdGcPO6jGe6cXH9kJe5odK5nMzibNM/lgiQHhcyW66m5+TMR
dCCwqSG8fWuCdRp2Xw9v/It8JaSWpz+Tfgeqmex9ieWAoPWl4qF+LsfgVVU0FaLS
wwIYomta7RfUhPNL1f4sAa3XzxVrNaza01g7MwSH+ZBxvN0KlfwGMVkchXaPs8/L
DRQVBgXaic/olkKeXeqggDCiGO5rjTEtGsR1kvDbpddEc8aGxNAaeD6Usbv+VR8v
rCcwkLwuDH2fNIOy8beDYyDNFrpU6gfiRu9I7tyMYjYhFJobytmcAMYTrlKTOob/
T/wnM9Z9zS0gYKQA4Cxty+PsLlr8KQu2espFxUwXBAePTlsqzm7movcnjCrnbets
5xDPa/ROLmPayDRmRlSzdoQ8oGTqHoPymtDmX6w6oVoNmh7Hkfg0Iiyx9pAxrkI2
`pragma protect end_protected
