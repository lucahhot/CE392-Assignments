// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
AZt+jK8o6r4CwLCXX+KnSI7NXHEJ11+Wy9lTQvAD7rhwFT6LuYXIxOx9117LtH7j
tqMTCMe7NGsWkFmtaccLaDDwnRagHT+7NW9Gslt9K9Tu2xH3O4nk1HXWdobXSInv
CHW3H51EBo/7gEl/Pm6Swz4gvhle0fcF3uu1D7VWw9o=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 79088 )
`pragma protect data_block
DShbWqbtSzPju+23yL1DVBhiUEYBPG/h38y9hb3kiixiiidfMsi0xod9nt7UJ9EC
WqxVNsD4yX6h3fFZ1xFoD+Ijq6r1WxcUY0SQRh0HT7di8Ijv3j1WEIgg0QKtsgQz
VSt4R/fVTt23W9dAo1UhYW5NBo72FJ7KcPCFjeCPxZ+vvg0oT4/LDyeWivfRj6U3
8A9P7Unlk3xLNXCa/sZT6JxSKccd0lrTr/C/I8YA0QdAaJrNhQXK0MzRzv0h1+h1
5DpE+yRucBZxAIp5/JX1Dz4arGF4evPUfY/rLRHU8MOfwHd8EQboqXp7mnYQAW3x
rqOSXr3GIM2WEbcKlD3mWGrrD/lRQcPBNWBP0A71x6HbQsTUvSfWflMhdch9wQ5H
B4f/cCiwz8DxSB7nphuIhCc6WC6x3WY0iPzPPisVUGjPHUOCahkeExtIT+EFyMUi
2ZWIhCht9nEMs+7tvKBL3j0FZ3o8/axlRimLiJ25M49lPniMe8HkW7qZZxGKapiW
DWcI5FNmI8Ki00eqgNBzIsg8qJAO1nzx3xlU//gsQeSx6udG5UYvvzPAmQXPU+Br
SAisIgTYvejqmnB/zkwe30ghlbkg8g5lJH1LWXxsSoKo1PrjMNlQzmX0SxIuXXoQ
lujYmS1Cz4kO9m8aj/JAEXi8LVtVKZCMHe7DyVuA5kW9O1lM0DmiPgpj1p8Wzztz
oAiqP3sHTyF1lUcqpRgR3ZqQwG/KSNcbpEqAIUfx8ogZy4IPpWeAyv1TVCnSoWDD
MU6b+dLzeXpvWwSek0lm1S8d8zLitUDGtfGSDwc6qzFdHaG36e0P0MP7jPNTNhiW
jWhGo3oEkx4Gm3LyJ0STrX8hHnJAOPqUDoRdMx4ZVnwdcZB9vAcCuFNjdFFt30tV
xaCjJdR4JKLzu4nZhmC8jjVn2zVpZ+77k5hFTiAztJMkcapNIMpSo4LU3J8NF8QJ
c9pOVJFRwu6g8Fxm/45xqNJnFDPSYlbPqoTm36x7CZYMeDjaj46D6IhCWODklaN8
3etfCE+ymP6ziRVYX7RFK8IDdDkH92k401yfNF5KiQ3+EwcHvjmOzBRtEi7R3yDi
ZMoHwWEEpwCodu6s4x+O1XvjqmBopIwAdgOO89hjUwEawhjCZltJnqKF6sQmVQgi
uEs30RWTw6gXZKXq26pvtoozyJnz/wDrJtSKo6kEtLxY8BqXxTV9K5cpXSOg/oFk
RE4oypbGqrNqC/0kGiCEv4Pumgxmf2bnLNFrsRHZr/MGJ7AHEDoiasGKUWEw6LdK
GnXObJEDVvk7X3VUkmV/oT3a96RLFvdlTe1Ze6Te5XOleSw8HMRyeJ76CnGrz3Sn
YUxjhAp2CGQCPF2McZzvCbKHO2QAjYqxPFM8pp93SoNGBFCB48fBWXEkmyoxj9AL
0FZ4fvza4Smn4jmumiazaxLASMMi25vdet5ZZi5mjRwuDPOtrUGuWRcmA5czi8K3
sX77u4LYaDP0p6R1iD52PQB+Wc6ZjMahyATFaxPnax0siv9BQ9M8guSZkBnUvomG
pv7IeGqclXfLmankWjFLFQM6aGSUZO/IYkljlFtQNcHQtfppEppju3NPL6HHVeqo
cD1doQ8gax52rY1Sv9s1EImerbj3w8zCpGj0c3KvCZ3QvB7AMsjp7AouNSRtoEhn
AJyoIUe3N0kyv3njMRJONraMf0YL5+fyXh9Ru1GYrCL0U7vnW1ub/lQNhrXIfXU/
qURTKGjpfW2juKjp318XaDL4FhxOcceucUcGRjJC2YVZFCzGRkf/OdTjB5SjppT5
Vm1QEIxUdgpRTr8KuaqMEtJlmjnvEKP8RfooYRKMWlcQwjqrujmJ2wAWEg6YMbQ4
jF+x/ozgHKnx7HcOrh26sgEgu43dEfPawwAcJayS2YP78hb0oTBK2xIXf67vXYpI
VlHx1rt9VZ55ZV4gtXJnOCmgAGoxKPf97xhsYnQyWGEZ16Gm63oH5vTz1UCopqN6
F6TWE9F0/uWxQAuuMmrwwPqF2vggYH87/rhoNm37rBzNBX8ghSnZTr7WeKJnMZJS
gUST2x2+xlB3O769QYpapR8fZVlUbi/amBtWhfKNMn88z/kYrxHNZzr+7gmjy0DN
TYveuqlUFD1oMLLlLtVqLsBAkMKsv8JP2/eDO1LoQ2KmszCUbljMgqo53CBTNpF4
isxKK484kCX075D7b6SZmiJn44PkLOq4JDMT1ZG20F2NTsZlDjlhwXy0uwtqh629
IcTkI6i4Q7igLYLR+fnEX+AbXUQOxxWA/05V8X6hKKZ1CtG0vs773wBrcQIQhbSA
w6wDLSxjwdRAG5MhwDaYYpl/duXV4mLeyc2nyijwyjct52MQ0AtFFnfbPBBlzYBr
oQg7lBlnewjQrPZM9hkBp7NBtR72G4cTcX6aAxvjKhPJe9WXZFThoQHS0quTTdZB
+YtDbZZujU2mcvE0GOAqKp75FgOI5OLd5DsMmSFmdsQ/jY7OMuDYe4nsJdF2Jvl5
AdC983yWq4TGQeZjpBqSpbdH28A5vFSOVLsBIadG4Un1blQpsSWmbhWZene48NLi
mZkZ1FigCEJFtwDV6VRnyKIOK4UxLtl/6OjXBf1U+tTntxcTDUJuPwT9b5CGMSMd
NqBPLhDP705fJB95zTEkv3n22ECYEJV/eam5AfACO1PywngcDDtin0l/7sJqv11f
//myoYCrmWlp9sGj9PAuApyo/z1lxU7aTGKG+Edx3vlB/GTyGI+zox0aRy1wfKUE
iwz3O5cgjybk/VTyzjsecR+rC+5rwHfGHvSKaL3gK1ryjZF2Gqq9xlPFua1Er7I5
0Lm1ILxQ2X1MBo96Mo09D5LE6QzuF0FpZefaMLRA6h8TkDwKNjT50EhUY7Qv9aSh
YOhZla+cOm6ITIPFBEHbc8LWpKiHK5x/PXUc8khz2BkW76YLuBgnRbIIx9ymu2J4
dab7cgqnMP0vOVKkd425fgaoH9GKTzvHPh1rYNO+PRBKkF2hoe5/aBkdaA3s2dnW
5daaHJUud4Xl4+F8QVIR8ylaOmM1aibHfOL3wlMVr8EVlM8vPziA16MN7KsMzCrt
wrwGeo8Gm8RJ+CkA64zOIBdxh5wQu3/ClGmwfm4qFgTIBvzq/6CBdhgwAKZTzMl/
a+w7udxtatdzUFeAEV91ROaeepO3UBE8ZxkSNQZz0h5i0rsRITqEB9Hig1/YXnc7
pwUvOwBO9a1XQE6fqrsLMYB7EJuvS6r327hpTkrgl9TuL8P0hMNkPAL3HRL6VEWS
QmeslSkI6vQMZlDptb9b6Jx5XOjeEQGYG8Ryyvenw47295yuJPPdWF7cbC6BoVai
LyD4sxYSrV5JfO+NBkwGIeWpGbAvEv4jtbDnXVSyz4Hwr99t0YEB1hqws7kEKpem
3JWrXH4lWkirkGX7m9aGe06aIx0WeD0Zvxygg64w2zGqIeBYKiXgIj71xmOLW5WD
WuaVksbMDMLd4q2UXg65L6lV8rN3jyGB7QMpcPt7hHgOxVPN0MScvHzJRBe3ysKl
sgkcx7AfcAiUpFSZFhOdnsLhkDg7iC3NA5WayYnLWIErD4Qz8sOb+lgxJ2AdYI9c
uqy8pzdn8aFXuaBYiKR29pXPk4OHxDsIojIONrOqx9ANQRNFMhqT0sLs7qTBXKQk
adrqnj6svZ5kPmC/7Cj7lO9DD+xBBOuF/uenTS5DnAnTjtT67HgSovqmAjTaDD0q
JFb85ESLU29uPyvXth3klJlk5iM8Yu5P1kH1ofcY0L3nVEAW3+jouCB3DiShPPwc
lnmbwtMrXFoSaM7ZYkmHPYQ8URkZWb+y/pB8iwhLEeoLVTupyJ8WZDIzLx8gGOrj
ndQka8LsZWlHceMbh4vxA/BtTXCmPlluLec01qKslYfrkOu+MY5YwW+kSMwWifjv
WFFshDdTiZaqbqdgpEYjxXrSQhz5brTaDH6nA7youMcQJJxAKcKRL7xCKgnygldd
mn2Nqy405D5u+WyQOLJlQ2/e8t96jZu/lJIKolo11F9mqEu0+RxXLgeBmlFHEZJH
9+Q+gGlF1SzvH/R64lpYsfPnj7EQe6/po146fZx58xDBfEiQ7+jV7oiAzW5RsZZG
CbwNOQAQMDLv1Y4jU4Jya0QYM8XFocIi5FioH8GhIS9kTKoccFuSMadyuhMTmP0e
Slnht9zZE0r+eyLqsMJEfzTxkf5xkafH0kS1gThVTGniRguXwlVcoZpssQ3agQGK
8586rfc1z0GeRTE8dt0aMUqOv1jDdSYZgsCfgA+l4Vk9Xwi+kiaiei6uiK9hjD0A
f8idCagrRpsGbWeUzQaBnXaUS/juk92d9+UfYApKfQGGXv45xAa58CyS99RQYvoJ
t61/ZvxNLS/mLiD4gei5L8VNQmfWcgainlqTcExPhtFuET9eLKhsG6ph56d50S3d
z1JSQHHMpM56bK4ZFylVb7u/aE+CJA50k5jNp0KNsku704X2t5abi1iA23dmQqOu
l03XHwCxm8Arn+hey8oFzd7fONmI35C75S0CCGwosCD5+usFXLxHO8hK9EuPB9ih
K2BqnYSIqzWH3gLHq5+FL7Q7b5FwbRN4uutaZx/eHtX7h5umteAFGR3JICCd/vFq
eMPq7cXRikFop0CpWcHO1stSd7SUYNf5UtJZH2d0oEp7U3mISZwbcCqxqcgawnsB
zAMwjqwn1ZWhlyix1p+lnDjUM0QvTIuYOx8yPqMajcAEMJfFdCossmS0CN42LTPt
YLsw3StfmSQSV1Qh+/SylYCQQ3uIaboMEaBP7KlNRy8WwoL8swTFD8gPJfICw85C
iZNCYoCLQ6ENDTHi90Wts+IZBcfE9NirSIlhbz8OB+RH6eO8errdQPYJFGLFfikq
0LHgZFiT2PFFGg1g5wVu0aVykh5X04Um5CepLjShklaEhizGV5UwW+QCJcAXrIoZ
ks+eiwL1TqMPQmxw5Avg9uUMY5S1fz5hGS+KjWRvZqLjSka5dhfgZCMp/gx850ue
NejUBTDQ6tDajrPfem+BTNOoBuqm3n39douv7wC140XF3AzKodRYJer6gfIF94C4
lkXU6D8JtGCZbWKCwtm/PHgE/s4K1UpgEinqrXcPVO+CI7NyAa1qPp2F7158o8UV
j0pOxEcH5jBJlSUdzh4lGaZRCKACDm5noWmuxx7bp3YTGkB3LPRu0psnBU2Udmkd
HddvemyfkElQv4IflIgJFTuCIsmZbpczIJ2krZHTc66Aovs89KNleMYfHDWgUnFa
CmlnaYBpM8Fc+EgUf+w8z8+jWpRQIk97VDH7Dk8iY4kIG8ukGJR8U1ijBCzG6EtD
LRJDr5uyUXuhsPsOeXl33cBOk4lgxew6GzF9mQs8I2UE/zpn2Zx7ncFP5OO7Ztbk
EA9bFTlAXkaN6Vr33WcmYKPA4hNGhjFCQPYuLyUHLD46KmgHVS9x9j2gIYUOre5y
DHX7abPs6yoW6QzRp69o9O25I9sOiZ/zr2SKGihWCCRESyTfhJ7M51DTKfR/T/vV
NiRsvai/VAHgXxtM7ZBepYBc2an4PdZe+mLvR/XxIJlKYy92f3NKgqDexgsSNIhK
xaHmdqTyxhRFjfOG179Lhu0EahTDzWOO1pnKG4Pz7UP5DLXAH4gn83RFQDhjgqDq
ptB9RIHTP7q9TyFexOyNfeA68XiPwGARiWGqaB9sdjqj/h/KczkmPrFru3AnMFNE
e0/vH/sNKMPJHDdBkMRml5N8tQBVOWxdbMx4OroTn8Yt0qeM0Jev/SAmtbow2sgg
W8s18mW5M2IbDRj7iroxdGEqV1Kz0Oo4FMEMUNBtHowRahz7brBBVGV8SWjZ30vU
cvZ8se58FUKJBwRp7A36Kx8yjKmNbYbQV3ybY/HI4fHarQX8Mvi0rHR/LGK9VQHB
SvN9yVCwxo6AT2KsGI51xRW51BOmHJ2fTsynys2yXmtS88a0WdrqMyA7DemrSK01
Nc5TA1q/DIeTkqFJUeCd+F2+/aHAdkdisjwRoNApzJ7fERoqb5xXqnn+or4lIn5s
rvMzs/ce4BkLhap0XwyGhJuMf+vMV438ZoScAebvx5Pw0bmRTaJRy6/THE+ZVJaf
MdAopWgpVFSFb1Bki6kkC/YT2vqZruFeyEIpFRAgvhBgeHK5oKTlw8EskfATZRPR
zjtuBqYYSEsz7PvesjJEuC1mIJfF4R67LA4XljqJeXG53S8UaQGvOBlYSgeTOWCZ
TdJe3BMER/0sw0hfgkjAEl27BFDbVsECx4S4SfG7hqeV2OGK36kOfA0aOLSYyDsT
x+Mgbb/YVdNaSXo43uhTkM2xVsjxvahYkh75W0hO8hxfKPmInH8+8tB20mC0J7GL
XcmM8cDeYrARmDxzpDi4NsKZd6IbCAJuqRsSISjcUjRmY0/L3gadJg3m0xKyK9qW
xBvEP3K1gl6Gq4WRmP22sjLIHdDQd1K9zMvfTeLONhJ+eSEcPmUqjWJ9sepcSaVP
lJbfnYCU0/nn0dnLVzysvKxhhvnFH1pdCGQaiqdma34lP1UzEga2k7yzikktmctI
02lhn3bigncFW7/n8tlWY3ze+cT5Jvap06DNp+a143n280udaDk4Gifx/0QP6IZ0
bEPdZgygSZQh8OOdm23l82IHWbbsr+QDmKCcWIn44ebcdUnaqIaDhbnmYLeFi/Bj
sivLUlDUXALZgDVpr9RI0KcsiJL2+FoTRYhwXtoRdy1yvr0ED4ANx9Rhz3ATN4cV
JMYycidF1Z2KU4C9a0xye9MfBCK3d1r5uNnAcSoQyNljAvTkEm+Pw/zgbWoPAXUZ
pjIB16KXg0Q4BM2eOz6urb/s6Ozu0bYM8e/twmHNBSkbdWXpLOpkJE448qUMQ4sJ
mdN5EAQiwJmSEsr7bfQZIL6J3s3wbr/nxEd110l+L7QQRsvK/S9JElJDt8ZRifMT
RMGFKUE1NnOJVql35+uKrMQYCEHEoK28I5LqV0aVX9aajXWG0bZ+4a/B/gRLbZta
oYBB90gGjp1yXsVl+gmtpFMJApbYR0eRxpboD2UhMKrY/d4ysrd6KUnBQUHM4n4D
OMAT/PZtN+6DBqwNZnTuuAE2Hb91pbVSQu+tSI2MTTxzkq2NnRXwX9k4qkKAWFvh
phl0HfZY0zdL45T9sT5EHgi1yFmtb2zbxRlFA//r2jXlulol0QcNjBQjcqjewmoT
aj0oJqAVgHX5A2wCXrEmEt/SwtH7eX1lgbr0vDHvQ/iR7qrnwt3ofnd2eYjQ6Anl
pMLJ+DxF0jCDPabvKAY0AtFB2l0eh06iGSeDRePScV8Mo1yUMFinhj51sZ4KSGFe
rrw3sbNNZn14K53oKQuQwCwHK8Nrahnb7q85cVmeiUlUKZ1IVbg1UZUQbxvRVn3D
dAlVOgb/9s2W4Z6Cj2wH+6vERYuZwwYq5pzBnMnSASbQyY7Jx1Hi20J1KOhCYpVg
gxxtVm2HmBuHblMrGZiexgBYKojOb+b3ejIvmtrXfV2fk3EN9mQTDRgnorb2rUCQ
ry3qWRCiu/injWmM4G9U0i2Wt1vtMSlFhvsmi+OCwLaqcch88tAB+7dZQry76+AU
un9EpxusvhJZtRyKNwLeXvf4yspViTfW5uOtxyXSwH+xuAYsvPdkdquatBXvpq5L
Fao3qmDrgFHW6YrAykwH7JsxhgXlxtsvx8hvad6QCFjeGrTDQAcMXpC2Sw/H9xGg
s2GUpAT5Y6u61tj19skNdcOrmLq1xCVv9fr6m9jrrBO1InU53eqEg6UzqI35mo/W
TdDAGeLxyGAumtHd2H43KUgBwOXlYYbETTAI3fT546ixPKoPIf0ahwJhBD1X3XT8
reinmHAgoKJK1o8iTrY5ixh1rs9GQ9PDjZggHa6k+G7tRXYN0aYfFnXeb5eXUlS1
dRtPIW1Dd5GcjfVrGYQ8cQwF+PZEa/BBmA97W05GHoT1hg3WvximPaSl+W4pgBPH
xUpJZ9ynrzVWhEmZgENLCP8wCyZXeMIzBDZYoMQkFBMp7XBCVACksYaRVXnFumzY
gE3bnDsnqK7ehRk1SBmF0A4Ysv8ScV8ybMwEe+AJlx39HWyWHjqJJnoZ881YGCiQ
kd+rHbOoYGH0Re7PBcYJai8+m+Ig16ey9N/lRaRZnFb3KRE0CcHoBjQdrsXxc6a6
MTOROKsoFctnz16EgfGGF2kj0L98c0KKJgxPxbo4bg2X+Iyor5qvWOddoe4cl9fU
em4D+hU2L7sOXO6DIMGsfQkfUhfHeblR5W94t9YvP9FBzkjnUaunC+faXmfyYtHM
a7+FZF/xvwuwWLq9ZPk//0iwNLoIzyOk9deIwaMK+UlORHGV3KzD2wW36MM/hMVZ
DW+uzq47okXUcp+RCHehf1bvf6u8IzNg6jbOWL8cJB9gHqyEiZNmwDdNFr+9ACb4
KMvvNq27lmjcyabqH4+2Q35OWzvyUlUAv7tFyOnQQel6gsZjvXWK+R2J+710CPcf
hI4eDTQOCh9hISFhYCqnF4QW02gtPj9YQiF6RhxA8X9bNwGoLKApKUVTOkG+kPu7
e9xETYRRmMcXy+KILOoHDpwFsUSUwQ5lUGsOFW0dFdP5loz76/gJQk1DFe4DU9g6
pEA3i8+w6sCVzvct2eYYc2RVcXkkBVAfD6ddtQ3D0F7YZt9krIbxGipNBlBr3kvW
NKcVbPrsMYXYMWNiU8n2R2ddZ1ZnXV6iK90d+IglGq3zJgw49m8zUAGLSJml0vwa
jwYe6R+NRlIQHM2CPVfkVdc+RpAx1xfajtUX/diDN0nRxl/wK3WQsDGxRsMcr2L6
8xTFWVQs5hIEWF88ZXo7cLitRWC7asBahRM3eKmcY6wFpDd1xbYZv56nO8FxjHnX
EYvYxx+pErZyPExQSMvrazxlaYyIJSsppXZQ0Gc8AiFH0YV9v9gIs9adoB696o4J
rVu8MURHtP258TizUbRI3W8PL9yX6Il/JhJvgqZjHXWrNW14pMlDPmR/h64+7zop
84f08cZ73r8pU6HAp12fKzNni8RS6ejBJfTZmlaFpvYgxywhCFgUKJ4YyTlNO9mA
zKDS9MSBW4Gmg5YboQd8kKWqvZGJc+n+VfYl+2HHEywNFobjG8W2yCJAXFuVtvVg
hcwEIQQet2tBy9TOINp1XfiIGBKQmnCb6ZtvxNn0lNItW8ySeitMLmP1iFNIJ9+x
xP/WZ3zKl8qylE9SRbRqZ/emtadxvbDBj1WkJALIq3iDOc5YGMMBBkh1nEzk+K5l
Kq5CCJhUBP4iXhFbQcvY5WvuDJzMLjyu9zJ07xoawnoaikEcrUq9lPCVFK86vrSi
ZFpwuZfSPuFUAe0lhZHwbE+Q3fxAIyOXe/2SpTZ08SsQwYp6flVZSVn9wkBm7BB8
+Ajb+85UQXE1SfYpbfu/LiqN1b2QU4oiSs6nrzRZ4gupLQysbzvCOQc3zuW8pmiQ
khCv5fB3lGu7/Kx5ez+lyF8J6VvhswViXh4p55TgjhNLHJlx1W+G2FSFP/tAHuZk
khI6PgWtGHAUFvVl5yo6xNoJXh5hL8uxDwk7MxIjfEi1s/AjtOEsnJ0+PdO58+vK
okZrSom8fcFT7y+q26/IZuRGH8EdIXhq70aEYHVy2B+CXFvK4MqveBqMsa6qvpuH
c3H3Umqu/ZUxeCLeI56k2IdQBFyHw5xaJrf0Lc+9n1v97iyoVe/wehfddk6Cvend
K/e4RMPogu/ysrQYmcwrN2XoqYLzNSH1VD7fGvuiJRAORWnuGYRtxvCtxshFUaJc
6TRuQNvMvBvbimE1LdAiAqUnNxsb0GgTGiLQm9+FziG+RKn4ifrmChJhmpIKtULG
oDY1s3aSdccfLdeF349tkuRYdJhe8nmhbINtJ8V4QR9S8IsxI1XBOYtc231/mlvQ
dSUYm/ssIuXqyyajU7tgOrwmWUROTFQ+UHW5N0YofgNplZHbaeshrCnclFG0+h4r
0aaHP2Ne4HX3bZjZZl/TLN6U7Rz9TgQi06Rnh7bOOZ0RD+z697XOShL9SIBeQq1N
aucJ2gkeq018ZpGooPMP0o4PlBeilzQNM1MwXIvNLn+JUY8nMp6jy3fEZHdoXgVC
+qmJjXPrekjzekYoHndjXmZwJ/g48LKw0kMu8y2rjBV1W1JLlaRLxLYWRfgl94Fl
LTPWuNPJ4x92ly+YSpNaWUtGVyDanu1C8raE3e0vdm/d7+WO9svdOet6QCdBmTMt
cWPyJhEx5ftb68zlM5CVTs9g79QRa0UnYaaKKk0RwjyscKjPE8r8Id0YMt2kwUkg
WdXub6N4lRYROC6BIyAkQ4mxN9iDJ7xphS3SCn/LgvW3V2T3SxeMrxkcNft1kLVO
pjew63WpkBON6lc3cmQcGOEVEQbkoM4vBgyB5yWnRYO3zpWLs6ZBa8LElRfC85xQ
uG1Cr6Lk8/Pe+6uoRj7/dhLgL2LLW8DlmfaHK1CV/uqZRTLeHOYZiIH8S7CyG/U3
2P3weoZ1JnmtKDbH0BpQyCknyKau68Dbcsj1b22XrUMM2KaYUgWleLcl6StlU2aE
Rw39F8LIoHVlHttc49JlQ5a+8/LaPzNGru+pB9YLaHyXZ0HILhi3njQ07LKVyvf9
h8R3hCdSnp484y7t5TAuVD9PrAa5R2MpUEeCKbG9th/zp7v3jZ/x/nxwl+lfaa1Z
Ld7W9MsV3/Hm40pA8lw2a5rv72chKzFss50Y67YiLFFfGsYEOKBXnGeeyQU1V8kO
kd3Fd6idR72gGcqDFD3JjLHrNl3yrdRHjnsbqetEcvSj3cXcb9TJcyCOd6CezfEp
bwFOMcQsUN4Wm4Fz7zos1tkEvxyHCVqo1I2x513jtvOkr3SLELeB5TGu8Zx0uQcQ
yn2cH9qDlB70U6KNjvfJ4dIOS2AT8AiwcD2dynezemqeBpJR1YE3GWxZdbWqrc/W
+IhZggOG2wvZ4om3CX+eg0hN/EzBNSaaT2w6y3sjl8E4qfRU9NqaduFXLEKJEjvf
ZyIh/7kJtvcXHpt7ZbJKnpWdKhlAb7sbOqEQiyaCioZq28d77L37v8q0Fe56luFV
090HeOPxkC2UBEliYD8+O/IJbUlNFW/8bj9MwHC/IvYzfkuAFpPD5OEoo5f66mQz
vz78vPI65o/ORXdRT4xytBD7CPrtXRXxPNk1rSi8sLc/La3hTqB7YVoWP+j10X0W
1I9mV+yuJy/koXhNRRrrV41rpK6nIfi9xiLd7tharQMzVt5v96YmOt1XYNHCuYnc
DE0rfJp6j3dTx/RsnBGALZYXyW24bFYuYt6YP0aldT3ophQd8sMctqHhZwuIghdL
ie6wYxav140u4uQz7gFoHanfA8swnPRJSsZ0K+Qjsn8UeZqX18zsbNNFgw2vpoOE
wF9qS3r/pOA34tRnwdKi2L2AzVPqwMozCJTjWzNaq3gv9dU9qyIBc3hqzHu/V7FA
R00je9mL/MG1EUlQbkg5eBxryrIztHL3EjhfCFdvODx1NipO5I0qdt882UdKUA2Y
6W4BLESNwV5FuYkZE5LvXJk+mLRdLL2c3eAO2e1hi+AW/0LPAzYVQFc5hzoDsfRW
ObDNgT9WOZ3acOY9f5KErsRovs0vJmnAQgRmagSWSK5fR5hqgXJEacj/V/u5LL7J
+K+FmHxYM922yhuwOstj8FH5FdJSQGBrkN533KRlYQaN2jr/i1A7TZ+aGAfI9Jiq
tzaGJQws8Z75a3O9LaypgJtyWk/M8xtRzFVd4rR4qS0Sk6RY1FePfBi2IFUO3Cjh
aZpVFtUHT0hehC+xV51ctCh8tJ7/todZYg54jmC3NV0KG5bhMvGGA0DHbNfmPPfx
Bqs4LDyvU2Su1OXquS1+d3spU1bvosktb7BY1b2bE6nYQinTVZrlNgUs9uXLPFiS
n3ew1sLrWD+jI3Dc3/bBhKA4X8VIN+ytXmHTKkcnh5JJ4ZFtjOTvZ+QmPlSfoIhW
MiqLbTDq7p4aG8rUqcapGcY5AxT0oqBKCQSRei3Us6iX8GepT8FEH4q5yuYLmvrW
IW5qkVuQcd24W7lNJJBAK/Lbkpyh6bi+X+iAjGxf90uiRuCQiOQU482wH7ZhMg7j
/0rG1Qi88lgpG5YU7u5dwm9VGZA8DwKbybJnZgSxPBADqxX6Z2mB03q1wdb0dNr6
kLZed0Ai/M2StL+RXI1BNqCbM7UQvFxFpDldXhXvXqySXs4dcRo9DB4YObfHgtth
VNV5mSM19qsJnK3UZTBNup6LAaSeewuILBb9UP8tpM5H+GMQCEQiBZmZbGaTUmMd
04Doh3UeFvaNUajn9OVD+7P7tYYX1d7V+cAu+KvLsWzgiBvzd1Vyin3S5xDkeBHW
m1Z/VxkfFyW8wNbZ3PfUjmrA3pGl9aHD2RvSQGzAM9uu/w7bxcqKn/Bj+UV0MiKZ
L+5Ot1g0ynx+gjCUxuzNvaghepjKoJLkada0KG8+zb2TZ+LGcfdBD6UNddmKoTeB
TeUeDAiNKQge1unb9cgdWF20nv//oi98fMFyTrdX/336wgzEHEsBAK6bgAwuwqfB
vftAxjPniObHsH4TglW2JGb6Xypifpgl7FdNyNiq+Vtk0c2n3F9rtTuIWrtZY4tx
1a0o17KLlmLuqgXBcQzziizF4Mg3oqFNjQXwAwtTVxIICq33NHe63ZQvqQABqoZZ
55K3I2HkK7JRd5D9/oshVvUH6d5Vj+MyPt73eEdNuEDPhAuDu9820ItmB/zczm2J
kHwHVlNGrUiHhUAHuyJRgBBnbH/ymVzRmE2lB90Y8rCaSCHz11Dg3S//nQ8rDhyV
8BMRvY3jQ5nplLctaH61xhaHr5S6X0vgLsOZfZCroB7rWoGsnrhv+waCLmq6m6NT
77xiB+46CLLz0fPvhvRxzSTi0OAO8N+4umZy9uDVYJuneW/zsL/XXDXITFUbp6tc
OLkHVxB6MmDPyon5yU0bjf4pJCK0CQPPRNfl4oyC+MbKEDBJ3w7p1Ltt/YBIwuGR
nfgYPiSjnpr9zy6VsG6e2gKpsLkYu09uiHF5QIRpWu1YLWWpYToCI9OIUnXct81l
uImpjiGtA95jFKIekKNTdn6iZXy/S2IbX5rCjWY52449h6SgkDxa3iyQPHGiikGu
OZa7pAHB/VVnb/kHm7+DQCuleUWxsAj5Rs9xRRnNkOble74YR84VmyiT3IMf9oTq
Gyk2glgcGt66MDJaAWRl4E3kDhFJMOXDTED1OuVXZ2HdoFs83UaGA6lyMj1tQU4c
0fgWmktl9BwUpnmyJxpd8J5DLWXEpite4N0//uRt+uW0JT23NVLmz+bVGNKf9HFp
ho9zFDQE1AdLCXifdD2o1Neqio7lFenNZjVDB5EOGKPB/O3JtB4edhxDM9m7Bt+s
8qHqhnk1on8vqcs555/a6Gf2CG0PyJcjwOHDviO9+Qqyp71brKfBD6+xPP17ZQX/
9azXR5FydtQ2zRJUsIPyAKl50vdOvFR5BV1MsBrdsVR5qsPW9nNVfo+Rhf2qU0ZP
AjQ5+Au7gL8Ly53xVe89JKLqha9szNry5XM9ZV2UhGwsOfxEwClEHK6M/nW/blpp
7bq2sw2BmjYP2jyNZ0OH8WNZ14fOxTMwUJN+yItC6wypdtCsK4xCk5w9IBx4e5Y0
MzZ7/zFAqct1+JnxzUxM+nd0SXk8SlILBn9Lp7hFshZdY08C/YmYw5ho7vIyUflN
8uhcumgD/uX/eXcNCtxk858mvGukJ5bTdUSaGpQ7FBkYLl3bVUaJV9twZyhm7RoV
THg1eLkFfM+MchF7c+22oji13uN+v9ZyNpgrc3o32SLRm1MexI+JkeiIN8PGdLLQ
vE1kiRyqHF6/LuahH4jLjCVkdxLxnNc01HvemsLQGsv0pS72+DGdPMgPEqvAW6dK
Xpw94DlW3NgizWCJFf56qJtbrZUZZFGq5iwP2KR9oVa5sJlu0gvErai2lGIz77MR
T4usz2ckAhFXwpnKY9ym4lnWcFgtbDmVSeGvwbx3bi0q60n75vH1Rd4RhsK0Ev6X
mFgLcgvrFwfT57wOU35ke4CMJEzYBodTIvlrT9Rda2HmEaodIbUGlRf6KdpcO0TT
RPXedqWX9AfeEBlTZJlSVjztoZA0zyNPethi9SZgMFYyrhSbqAgSmHaXPKNmZ31n
KErGn/2J5mSC7tI84gKW58thiJW0FRZXcQAelckjoeaIPuUm4Jph1ewdAciz/S75
/TWx8yyXSAVKDufU4F4vPa+9m5Bx+K7/wWOnhf7GFR5Czf1/nEAz123fNAbNk9HN
Uem/GZMQZoWPkpOrEALuUlXOL3jHPhbCB2Bry4/kweiebkYNn99f08G+QhQzHjSV
ty4yoZMaR/5FllqH0BeJZ3qqaBC4pSrApus8896P8/mI0L/IIsfAug3FBCpzl9Fb
7gwhZ7+OcDpAO5s4daZDxQ5n4vn1wjbxswCigVWY6qOfGevy9OTKHuNZ4bKsTOVb
a7enY6CxG32OG/41cEj8HPytUtV1lmSWfFFQINtKfYja3v1fszgRVbKTjqt3E+JV
2ez0MpK6x1Qqs1o5I2vf9oNViDRJzKOk1QWLe0Bj9WrLDRqj9vrhpRcVAoF1u2Iz
q4WtKZyjTbQajUfH2dL36Byy+CLzUdddof4FT6BQM6BuT6iMpN+2AYRq4fydHxpL
xlEIuhsYDwUWpkerM9P3hVCi6sn46jBLD/CzoE8xSbQiflAAmfL4L2lD3Z3UCUsy
8bP7qtG+XHOjoIV1tT7Sdys5Vj0Ng2XBu0BhrzhyhioZbOpSUhjdN5drbwlrzwFB
bM5kRcIlo9vkKLObG9Y6EoS+Y3MTD3XLqs5C2N4PHyZkyW0x9FSEBtUKvbN0/8N9
zaa33NuLsZ+s8ubH/ZJQbnVG98u2hiPF8MH089alPurbPuYp1dVc85zSHBZ9MJS9
xyxl3o3CO3bLB2ExCp35QEkR3SQfiXSVmbZ93mtytShdYjx3RKOFX8j34LWpgoXe
VQpe6bDnIHCcOMQtLFmYYcHjJ73b0tyO2+4KCDhQqDjigk+x1QYrcM/jih7hvoQY
vuX4eVvufwsSKCHktqX2X25lVVBYpsS2gPSD6DplnivFqw7ITpjSO4W6xEzqqWHJ
A3a6wrD4rIuNWlxzZkzNErDs9GtVPLbOLpzMcq/4lprzvEk0m5aSnWiIETqXx1xq
oM5gIlO4omV7rKpTyc/3d6uCluYs96JlHRxiE9PcVWrTbFXhDMSFRGv6wgw5BERr
bmaq1IiwEf957ZQvZ6Ap0VbQf1MGgrQ6dOj21i9BjgIwslpB5OxOK4j6j+ij6RZw
RonNwY2ihFPz9sSyhRLVLvEMrj5kHAsn1auDysHtMvhUeEPSzDLJQJmt+TXNuELf
XK3SgugSFD206gge7z+vlly9+dPQjnNID3RqKg8LsIRANiUFHGBMvKj4ZhkyxqPK
gD9eY9UoqUpTvtNYXnu96K825eTmD+0tHAjX+yV7TyyN0jAQWWaSK1pXQ2PgbLl8
ZDXbA3IKHzJhmczl2fjR41yE1bWgJsGK3S8+W0Vv4bXGpHCXZiJh9eJOFfahfdzV
CjP5G7lCFPdvSym3V40uKNBODzDg4ed9+7i2+b2oIF/K2Kjz7GYtYWEwpZiDuvoB
B93SD5bf7TE99LrJVO9QN2iRwxT9flGuKnFJbm66cMuTUBX5VkpYFA/ACBfoO7Pp
fMfL3djy01ct7CUEu52aPMnvqnAE7DaUtT/+A1gE4OrzW2sBixi+S1FoZ2uNPxmQ
nvkYdvBrYhBLRp9PNr/8xwPLkGwZp0SlPNe1LtmEGmkrr7d7vJKJjnQ7oIkfYmWi
5cP4/4uzxG7LOiDHRUmAYNANywksLnATu+JRaMaf+ZXGTIIh9gFhmI2B/HLqSPpz
7i3UFi+4UMI/NMJ9TZcZJ3vifs+qXROHiaNau7UHI7TAoym8IE+gD13z3jjcLr6P
S1fz+J0dbq4aWYQX/Ku05wrpOP4Qjz8zAlRBfG9XqB4YavKiO9Fm2ELGoVFdExDJ
YHJDlV3+xz/Uq7iCefVASUFj2vJFn57b/AGwbTzlvtgxDrqijL+FCM0pnLwwrvU+
cK8dHLEERQSQresJpGU4wXL5Ve6hveSORTW+RtVsKGR8dUj/CDmR/rAXH5oBTOR7
jiLbfgTnb3wa+4AoTExCB3ssbLEqDhcz4GSVQrBbA3lRKXbQbZ1k5TtCapyBPShX
YjaLwfJuAJknc4TUjkymmr7zKj13j1Exgf08csp5jfpN8VHmV4kDDxd4Hq309gCR
sp721daYA1prVrlBUSxSvfVwK58VE72rvl1mk5fqimDV8Vlvfvu7S3feOug8KO3+
nQ/kACwHbuOI19B+Ps8hWbmC0Iip/nQpDKp/9Pm6nOwJQizR9N+UVSuivL9RofXb
OZwiDIc3++e004fS5dsPyAgSKOy4PtmV1kx5NHRgL1kV+X2UJAVdDtqjVzXXybLG
zz+jOIticImoBdtTokz6dYizJ8oZOcWy0uPxIY44NF+ZCZX2VZcQUsrQw5Rlt0Ex
VB8T0DuF84RPCgpRusjIiWCctyC0kQkcMBEOESuCyTV9DhhR98mjVez/N7Taok2f
teG4FuPF0hK3mi+vHbfcnuCp30Eg7RfyTdqoNXhRilyfGnfYQcUaanv5GjGQpwjw
JhgP2MbXhP5tA2MAMkGdkY6Zg0o6KFNCyOTIHkMq8NH+MIIxheLEuoFVuC9WuSsF
UzU2vFA3OvLfUxHYiQVC3+kAL5rDBqdR8HqQExI1v08HKPRQ+oaWcD2rzd1nHoX2
ExulWutooTugf9m1olJLsQwRc+3x4+y4qRWRGpEN8DGt/pBdZ433ohrCQd37uMJd
gCty1O4ksoH+nTwRA0P0+Xk4VITUQE31/yPToZt9LkeGPLRCzOIQLfWH0T+Z0iWf
cfU9egApnRN04VOcUiH1HQ5XziwizTcbXLqF4lQyXPbfdaNV4ZnVJd4c9W9FUDkm
sSOZITxstbNfuxqI5Wyxj2tw5YUR10kHF97jLb/1eOm0+ABnnKgWhKO5Ik5KVEcD
okte+lCQaHIorUusWgRdaMtv3X/6yYZiNnd8SfWkZbHYsg3UhiRh8opbfeg9rSpI
CBv0aODdsNVxqLAJ08P81sMG7uCXqh4yqF0XiBhFleQxdqgxjnswP69R7gnWZSND
vhBk4j6hgbnFPkJyqTAvRJDO8aOHvlxVraaSEv471LrPe/1XxbP4LTdmW+pXnRb3
uVzfTvyVDHOWWrrPKQ1fvK4U9pTM8mQU5Bnb0LZVNYqXMxLJfBSDPjSb+5KltTg8
aPchyDAX8ZPQ7OftphQM9pjXzN0Jw6cchy/VysgH0ubkLwWdxAiAIm7GdMtCJpjo
08XnTfAOS2n1muH5LP2hthXMMR61BPvPSwWxlzT+99PdwED61Eq9pY/y57z8FeI3
sgQgW+tiO8A2oYsinTyyyIqE3HXDZ7CJwHN558qtkbxPMxkDTUE/kVdmfRsChJrx
wPuKk5vxdB/Vl3DP+s4kbHB2jdc8hJZs8r+A799MQCeiZR+Z+l7c/+Fg6TVm2Xns
tZn8R87y7yfi9iciSeNeic7hikM5g13RYlWgW/XFoHwn8rMEqd/S5JX/nu5qaqDR
oN0uxvNSONBFd7K9lVvhZhnBVDp4+83yDqRHUegawhMSPy4YV1hQsQnb1QbK+lYE
KXKKDoN4q8NZkmIgZApZk76VNYn/YAA+e2PjHek/kBXYKNhtE06ftR0aPSyFk/vs
937jhASa2l0eCvxi7iqH7QJ6LiEbTWVOJUj217uFnbZUklFr9m4vVuGJnT30z+/C
3E/VEM82fPdJ7/1dJw87DeXzb6/jb+nB5iWEtT0BAZuPA4ELdyvbvxALfNvikrSg
NERj6PdvUQPtbIB5yfAqoK3jGUsawiZU3y26BxVqnfe3ZN8QRujMY7e3Gp/dJ0Oa
YnioHMpBUVGaGzGUCI8vlJVxondbBhRcNwbyaVGMXVLC6bnN2qqhASatRbp+IywD
QgziNQCPzPqEaUy1CdswfYa4ktNLqRhN6JOgnqQ10+ei850zXj/KnMhDginRqTmV
frBS05t9cxSyQJcYqDUdwCS6PZZ8j0TNLRxFSEkNAlRe6ZeniKtzesWbJC4ui+Gv
BVFkfzJN8ziLZ2G1jA7E3URe7kBwVid3ydfeSr5NRlOF4imAFeEwW79cj8FNy/mq
X7HxM4wukWdQIkHO3qAdVnuPmCzm7fmoNVHoKVOA01FKIoPj3z3qSKMarVH8+otl
eOckTg4jjYpkQK/Am+M6zNzBu3sNTeklyhvR2MW96Ho5i0Z9EMexlafPxmzz+CVU
UaWHpUeB3dLhdEl0GPRJidRrNPn2L5TOYn9AT4n/pq0ocYstZzQE84p+Wz44/fio
lner2E43z3JTNwOdoe1o7hPFcquPSTR2dp7JBuRmfty1fTg7Og721vv6ol5QJuNM
NTOs+xK1CAGFmz7FsSdQz2SPr4Dm3sbIpAkNErO3ER0RIlFYh5LHltMG/4NOfCCx
c9hXttZnH56xA1gIy8xHPgUj8zd4W4B6i5xY5sLPuEfmvyEBGOFTLyBSVjpx+qzS
R0KAsDU4OzY2AuBbs7xuvRxNOKFtvWIa/EytsCABZ6+XIyy+wQqCIKn5JCPcPCsf
Y7W8SU2sPTfWelJ+jwbAM3sI10F3kG1RMrwvljX+e+ZThXbbsUwlWqvMvPwv7Z9c
dv8WAwe3gOZ6OC+WczZY7ttnyhIZ0gUS5b0+SvwWJgCLmBC2WLIk0OLfSKsmzkwf
gxCLPLMJYkjThpU+RkNyOHP5eQY+XglR2IkbjnnBkMHI0CIwrq+l3iiInrPOsvM1
x6JY5JJDKd1PtVwqUGjCOzxtTumKaSu6B1X+0W7S+crT1czpvlIAh2oaG5S4JzjA
Jip1rHm6GjUnR6j0vk/Ovspq5ZlQHQVJHC6xVqPBLjzMIU1GJTp5vjhLPlipb4E2
vA8VSiiKL357mLh/wtQMyx5hH7LuFNUiRAn3wT9QukJn2gUSrBEALgGvaUYl5T9u
MrzIv0WyEelRNK33vC//ofikqqLMSXnxx9ayB3QBSitJFM6o+3BSuwRuKbHcyhMY
5ry/XacxLQrtK7STJoXAYr5Ao0B0co9kLt/ty1y8XxRiKDuBT5QbScbRfbHePY3W
FV1ZDs9WBi0acp8TbSSVZUWiKr6fjbUGSzWtb6/iwY8luGh+xyFXhu6hY47v/euy
A0xG/ynFH+7EoXbPNB+xrbdfNiTVn1xC2mwriW+dihGDKXLh1Je+hOh8zxdjoo57
AmTeOYrG+rbMa2xLklQQ1qm4Re6l/zd7G2w43amxM3kjSk7xdHqbSor+XHpeOjak
kImbqR98kmW++s1Okkij0GQmgcH4bZeLgqIdPqolkM/0zGF7XCLpR9tstXGjSGoy
BFso5WYL5P6mXbr6flwr8WDlpL4upBIRhYElExzxNNaRulcd5tN13W0ez3EqtYjC
gvUeY/OueLVSDwYfTHXOTceFFE9RJdJPueMR405P9r4HhG9t2MAGx407ZRdG6lhq
35TL1rieUx9inEfq1qpRRcx5D9s1DrdUUvU+fQfpRFCHoDAUJv/EeID7vuOVmxzn
C4+/vrPAm7wytCfbRCQgsCRUUxecdWXtkFr0SzDF8gNyHycEe4pbNTCKlO7Ipff2
TK9zSdy2TwsGL6+apk0+DYKuhIE9zevAmmcVTC3RkTnVTV3nXFLXgtDUgwZ61Kcj
87YSYoY3pf/che2ySn6GK9alssJJc4l9My4pNRad5/qmxXnj1pB/xfqPQ14lEJAW
eqUGDaFYbyWr89wpMqriKvwrvG3BkyV2iyYOC8viOFO9IDT38A0dL1ZQtMZSlVWU
9G0rVc7p9MRclLkjNTgnZo+cjrSBLutQpPgJAwaawN0AxLD62bwUJCweSleM30wK
+qXw7GJjmcimu5TU+sE8wmP1Zysk1/hvYgZUpR8HHlLBexy3CfMexx9ergWrzZjR
hdwsg4RO1ivv/GPSAbq0O2PrkXRWE3Zn0ZdIqIHBnIR3BmxLZ6r4zvjCVqcavsWI
tJ/k3JDlnIMODRMeLydR+J84jEdBOwIUPOftBev4b1PoKFmJo+AXB6nrDlixHN8f
Pt1dmwUs8WRaF2lYBXVPIH5kzXr8H/fpggKfV3pYbEQ6zoEC5dJHoRMHNay2mimq
79e7IcXzKfdZjaCj0hgCBD91OlmeVn+bmfdlzcRL4EcT3B9W1dMSHrZBsQXZhiH/
LyO+JpMpxB405TB8gFyMXVuip855bt7y2rRhmmEhd4j+6PA14yuLse8AekLYF5hu
u+oHLMQ2tgZvpsxnzdwSx98xI4u36Y5sgsR+MrxEGwRewKe7UhGkyA5VVBfFT+GA
blD/PuUeuddPAHiufmwh6xMmEm3bI3nB6SeDWzdHTqCy2sksViPNU3ztVi5Yod1M
XfF2dW/MGfOmr8u0QiHczW14os0T4Z3d6TWCLl7wHN73cxPpKc06DfA8bSP1NaIl
5v/iZyciBFmpy6bCc9i3qSfPp65sOLxUB/1lDfFBsWTlr2eioWcW130kBGOqNwkq
swbXGZI8lupXGjGAEEIBklhP2tVePIaZvhltUW3wz8aPCj/IA5ILfgXvHarWfjD5
Ms1VYEgHly9YJts5iQPmCK4Mhx6oKGEk86FBUl+bpiMvOpvAsm/+u/JQUaPeVF3u
QQvZoH20vfHhu4WnLBqP2FBjB/c0SAWTlLix4lCimpGq2esOMCY/Q1cB9X9Ia1T6
52Aev0ezynXabQ8gqGTBG5JjXEnuXNqLt7Irr3lnEuscuJnZddK6eg0RjBd5Kof4
l3iqO08xpKDzurWI17mwlk+fsCe6Aj9Xld7eM9MBUu04YKxLgNhp0c1908TXiPDf
3P7mevOehCVoyuGIKAaD4VS0jFfZjnC5GDAUYYjY0AgrIf8mCtOdV6NdLYN5v12i
K31yDazxGubaAr8pzB4QTPl0yLRnSY9A9zkF89vS82Zl68KIBNXJrECChNeEjsgV
bZ995Pe3pm7T03+rQKKllLHzob3GfzK/0k2PZ9TVyVszZKEPi+Xzzws+KYzwfFNP
PL6PwXk0MBW8jj+q1BZGCmk+Q/ftKoT4nnIHmjcLYQ78TI9CLMB50bKL2PjahBQH
vz6p0CvAbVUBwXebjU0fAo241511JGJ5BGlOP70jFDkq1VV0Ef4rkATIO9mJ5g8S
69wR9GHiT4JcwIO9+q0mpbI+Q5Gj+2Uyth3aWPunpJNXylu6TsrZSy3b9DvPLls0
qPRLfmQfXNQlfq3MSZ6qoP2+Ggsl1Wg5Va9Is5eHwDNVQO6zqMhNKp7EwE5xCGbh
BFw1659hP++VuXGDLDwxm29osN2KvUmIJcYIPGdpnbvZWGLnqPm9qk/vaNTq+5po
91uYtz/fNqvgFmgD+MXAjGSHKSouwtGGw/hf6tIhg9Zt1qlueZbBSFUWI+VgeAZ3
7Dl27ZdqPtVdZMWjxmrNd/wRcZVnI/tyqHCjzlTAFiQpRvsdLmq4NYdL58Q0fCuV
CdrI0L43pzt4s+pg6LiFwg8mi9UZZpCId6NNrj9+3Qu1Js4UXC8b77dBSlR8HVP+
B/zC0bPNe4RHfgQHnZ5GAsw+8ugmuiwQ9smCDQ665ptT5IEUbVwXIQpDJ78NQDcw
ZVpGKJfZhRdlmqalBSyBkaDnMowkmmElb4HqeqeLkWoFwN5p/HdOTlrACsnP2o4Q
zT+fF+UPNuUuXHDrxj8uFxoSz5p5qO7uiDYaJKzaHwuZD2KfmH7CNWCyNwpDaJiD
+2/lxCLosVaPi3yGvDiUydcScRqAnX8k+XSbqhGmZXkjS+IeBDc++1K3eRPj+Ems
HDSIzb3Bp3U33fw6md46vjnhk9xtE6uB+FarWG4b6hmbQredtByqgztMmrXvgs0N
u3YOBxtqOxiE9bIRl2nZxjy+dfaeymjCZaLcUdmBoVzX4vVaCYNBMyW2AxxJUHqV
liv/6IDm4Gl7NG6DlZgtX78SAnCeJjMeIslHi4IUKA0V3M6bhl18c0MPl1KhyN0s
uM3Zyc6tzkwQPOwBIxeQLYf0fmlXxBIAVZ4uC+aA/AAkW701+D46/vrsTHppeOyO
NfrgWvf3LpSPkaVhUxEhus8dD8703nobLpK8Qob0MbQ4dBoRVV0dKL8UlwRqGAUc
rOrcOhMrZAGcFhj0Q42UTXPiyKPThbvVcfha+fWjw9S0uEYL6Ib970nxCN+Ww0zW
OfM+une5DieBlRxJ6I+tlbiRE/VxS8o5U8uqZmv7AcDZXz5/EXZh89+fnXIqFCga
4rrp3Fqme6X5CWP3CLgf0z674mzdxOBM5/LPaXU5hwfWDykfvgRD74HBpgzbCyJX
mCdp+H7KMHVGnauGRQomhoSLhbbIC5uWTZfWcis66aQ4Pfr9HYlA95a3X5jg8ePR
HYUpWkSCDKQYi25O8ffcy929iad/254MB4vHFCeLApKkefvG+P8SNipC+sM3amQi
4PRHNC2isKjtjJf7/cJzRdRHuuiceQnmN6nzK5L+DU0cgrwmeHglG0uRVxSaVlSf
s2gCRxpBv4lDUPg6FH0KsPrJMzPMJcLqBR3k9VmLfI67Dm39Z2LaoNHE/mnz3mg/
3E4Pcw5Tx7Gt68VUTw/4Ji04UCSzDu35hBnjGKP8w2YbHa1ofwK1nZ1ziNcmoa2Y
cU2/JT4DobIJoT0UdnQYLCOBtLTVfMUefReoFSvjmhePom0sxxDZLscxM/XJwOJ9
Pe5SmuTYqpMNfqoa6sO37jYiCoe8LGRXZ6b6FvIMcPx7jhtjLE5Jg2SAlH59s1JU
lY+ro+bFIw28HVJU4+rDZckhqaWxDvHwfNUXy5+ZoVSsUX9L7G5KPph3AlghcIFd
WFs8+xxwz4FI98XQYCyc/ifzx38utq2scRo4yv2DiSCIOlV6M/kPPkU0KvrfUysa
PnrG1RnrwsO6bnLp+YZfKW4tuOBrWQIjKKcBFzBH1AXh9vIDcecPCmDT0RxFX0IQ
3X05ZGEyy97HQ20yJ0QdB4GAmeMVFlJiq28+l/iLHXmd/9GMIIg4Kz2u72nCn6Xc
ZNfP8KmKIOZb5mN/IGv/51UgJVrOWb5qq5z4NGwWVeLpTXylITqPVSu2lmon5/rE
ndCCQDDht20/6e1Z7hkTeueaWilo16cOZifsS+SBKmaWsokeik2LyG9DaihJReJw
qB6XEJPHqqg8/76WfpnpdixelHleUh9/Hj2QfVYq98f+UwjINKQnAWOpB4b3OkJp
KhezziHzlF1Rp1XlQk5kCmt3LokPGG/SlPyGL1Hnq/Iw1PA83DssiT2wnwHZvoKw
oZhhOmtGN5K8f9G6tSSXxYJ0JFJuQ4YpR2TsF3g37ih8/kGBZIiscyG440UUX//+
TelRIUHXRZvxaoJ/MaFoCRmu9qpwhhRNOfRL8ecF8uzgzoVBmkAPqEGY681cNc8o
L000sR8VA+hQu6himH/rUYWUXDL0OfwKm6mFEYa+tdQad5R+eUA3lzOWSC5CvE++
wkgnKgrxE3ORwDjEmw6a22++H95WHeyJv2aw5itRrKwPx2gXqt4Grt5reP1UHY7e
TjtdZpNDZJ9TkhXfIcNkRm4px7b6FlsNvo8zrlPCrkFbsnDhTHuum5nBIAXQpyIV
YRnTWPU87gZo1gxVVA5A6oGGKbmCWVuUmBIX6Ks7xHkkvy8u//arnYj8N8aqGs58
ZavgTBNgjBFGuxcBM432MuDlOL7BsicnuLDMlSlYAn47h8aImWIC6vADEfRwHfS5
6SSkNjnB2wqQkvZjyK0I+fWPgjpncO7fZiyaWhxu6T8pbF9673G1TVZClrXmikU9
KRicRP0aB8798d8fS4/2tGo2not0mGZac9DHZlOjZr51VKeiDLIj7N9QqZod761/
Z/AvFYYdsxa4GRq2uDHxcna+jhVjq/1K4+oHV2ELFOB/xXBFEAixX0AL0J0kICTe
0RlFI7UcgbzZQUYxMSr54EGFqCN0IntOVpSh0cTTuVJ+PhXFtL359H2psgO7mwia
K49POw2Inodm1n6XJbJ80obV9dZX/f0PDOzV1NCLhMXhEyK4ETNopbPuALntA1X9
2z+x8ifJ8w66h0qEb3YqZb6I8u1LNSWiaktAv/fLi1FAZPFxk/aDXRVeWe0tRgxP
KUH0NMgJ6WvBpSjqTwbPG6y57/PD9ayzqBNpaXdfrY5NNK9iZQqtguulJmQi1R3E
l3I/jRNxpxMcud0bAoLP2aOjwLymDghwUvUafSdSURznTpd0x79OjQfKsseZip3F
a/cbm/Bi6iuB9bJCdH+1JVH8kuxD2XHmb1m7gNUnGUVfhEzo1K1OOZCyMlDIiy6y
R5qtu1LdnQeC/XWpR0fBuIAmb31tU8b9IGH2ydOxmdMTPpwui8G0aeDf1LGhQVQ/
T6TtNxwM5h+e/R2b5QualyuPysah6WoYrU71NwBQ09cYsz39Z3HCww5RbC/0KByu
Dp75SxDpqa9AyR+2npYCTVicodL6Y2Pw2sNvqz0xawEjjolPDO4iIm6fAPAH5SY1
k9GYTXXHXpyOmnHwIOS+F0LnNlgci/CpFSFRyPnXufI8cVIyCSj3CTyf/Kl7s725
e/LtN+93rjXDMHlCnlvNQq4QLJ0bLQWe5ypCEOuiLFtILy5ihCE8JFZf1wuLDrAW
6DXHH+XScajzbFxFf+yJPReszLac7m75fY9bMhnwq691T9XlJrVI+2FAe+pF/R75
XcWIb00ZIjfe8N1yE2K7JsdMZcZFecyMJyqnmfRJFNtg6DrTmFcgFgJTr/sWuzh0
JRpmhQqBeBCbVb7Uzt2hEnkpXnekW3SDcTPziTJkvPJvXOQxpNQS5PbaT3gFyi66
jNhG+zSLsEnXEgRjHL61oQ+ePEh/B9aMy6aRJd7os4/eIWsYYi1nYKpyai+VGdj4
22uCrF685IbR99fZFTzt7cJK0n1totpagfSWXaCH0GV+JXkFsh1TcdcnomljMTTp
28mgn9oKM1J1UWQqIBaqezKpCNr81p6itIL1cIwrNfOT9g7xvuY4v8WWrYBlFnFt
R+oSMjg9gYYaLtl+ZfnABrMv1TytTisiy01EAqgCXFodUFuayRajCrdXCWoS+ZMB
U2br4KMTaH7yujsEqyKzBorXTRMYSKjIU7uorkVx6n5z5HhgNbPc5JTVDw5hcEzs
nk12AjGJGsxS9dqVAfBDlLCJTffj6WJcNpIb835HsWtT6hVG/Bcb5iCoir4nwvhW
loJvLgOSbiln0V5orvXsmtHS0UACLwrD6G2FXB2DKjWvOFYpLyhEqF8lngTio4ik
3FvOPZEhoyeAPaZzeqBnLJx493gFNmKXTRHxjAHdo82UG+Zzuy8Ekxhv5UAMSI0r
OEj6KeZYAKQk1/L5G4tiFloICPjWkw7ncROQB7N+uTxEAGhvj/o+vV8D3Shqtd3G
6u6zJ37towclrE4Z1YZfHFORqXW9BSAm/nrklQK/ja/sqqmcpvOaq/gnKOH2Atg2
nF4Kt4jS+T3olXDZ8hJAWB04RkIqlQGdzmYQmU8dRZOxD5M5RKvMnUg6IL81y/VV
H4W0ghTE72j8RppK05gJNxfx2g5rvi2N7zILL5JP1dXLiCz/FhiUas5078ImUfwR
lcrExAeb3TKiFdbd7YZ8X5PnSndBBO8IcITXVI5E/qwm/recEM1EwuMq8sHpYwX5
GDMVJRnpRp73RheZ6riyi+dbOpdZUz68VZoUxdN3isQEUj0qMEmwRvIQSlajLrOg
q/Oq+jEVXMf4HrWeNEBh+G/pTAk1BflfKuxEE9Y0Ad9ri5JYH6uAgv+QKUF7BfiW
vz9eiq5AjSFxwTtZbefXVUx61x3sKBRycL2qYFDHqAlcFmWqON8syv3r0tuq5oa/
2NfiFfTndFK73uZhGVAhZ0kxasILIL+5HTQwNazJMhY1pstqFBKoC6o48D5zRLh9
rGy01xs/AsRKhGgfcMSQkKqiGi7brS+Nh+gG62O6x2HKkmPQ2jmXy9MLHXqrey9f
RBqoBt17v1Snoqnm0SW1M9lsjOk+Gia0shzQEbpkVqo8Bc5AQGZmXO5MH6SDeifj
Rlw7FVV/3OWnwSlhtoVf+P+YsKHgt6jjPIf2X7llOVa8hy8HWLmFsdDfxSHDJA83
6W9DPiAGVFmxc4AK37rexi26UQ5Z+ZJn9RpfcczKbeSVz2H01mHuDxHd1ZjKZav8
Mo9bm6f1YaP6IvdATvREE0kTvLMb0inbs7boTNmZv3PfVWvF0tH+wxWTmL6ypSf/
YUf6me2JhcfJAHE4SpL9A+C4wOvTZLlvo4IbY57fwtgQXwdleLAQZMqTRwaCPIxe
okFZbWDN6B6uCHzUAg10/NnuUfPr8VHMFrEkb5efpBtNXLPwjrRn58vgEr83W5Od
br6uaFpPHAM88SofsNYZNICZjYdh9GPNpXgrhWoAjIgm4HPWRoe02P0YOzz2LFrX
SimoX7o4d7oT/wu0XGagtedl285yBtQOuZnfwaJV7X1aSvaMhA0LPM2Djo78H99A
nuOB9WpmtdlGz6cmemxwIU+tM5vCUX9z7QaHeMi0XE7IqREz4NB1E7A3wylLW9/V
kXb3oHk8GhgDqyZP9S8ZuQX5m03A+dHgDd0Fdzx3MCFs6Rq9ubtKq0yn//H3X6/V
v4zHgySd5CDUnmMhMMoL5FJJLJakDxwnLGa6fBguZj71Fs9r0A6sgGjIkyQypd/0
j9zRRNMh1ToiHrALnCwlw4iNmDmpD9U/N7K2OwvkavuKryqrz4hyuoS4zM6ggKJS
Rr97ZwkonMSqkVvJwxfcZ05PxrBMnAN2ztTPvhrVnO7a+zQqrMohv5SafbivP3/d
wKom9f2OeKYTDoIRNQWS0i+mV9PpavNi8KjMQaUvuAwtSOrjAaJJXxZkij1uPwWu
qA7nvGuTsBNJ3JRqz+Y3zEw2xhNi8Wt88lr6v25u54w6ltaWtXXNjgF5AE6cZS4x
Lt5TLZqsUwujrYVz96/AxbxnNlOf0f2tyD42/1WYrpY1ACbUkhhtOhyxWSic9urs
vBPpRLizKPbeGUljWnZyFM5MZapSFCBWU4NvnDcOrmtdypZZaEmUSjqG5UaKRwEl
jW0t2/W3fiVwLd0LWxm9sAqq602Nq2Lf/PP2qYyep0qGmBfSbwLE+bIp5GMQDa7v
MZbW3ockIxvubCEXnV2NSN3m68xicuuG14SkLuYlv7Zwylt5D9pEuOnB9ouHUDDO
3jVGb4zRTW2eRXeAKdOpiDsuYMihqEm/JovMYEQnYXweYbcgDYAZjGa1WvzaOWga
8owuJkxyWxivCOQjfjTNknqyW3xkYlE24niTQAuWFLe8Hv+M8p53RI2yV+XYXRm/
2rci3WftN1m1Qn/Y0jr2PV+weyVs44qKi/gTbzpi/vCE+gd86EbepQ/BgdsLKAal
ZoCxQzkWb4mYRMmgOqTwsBvvQL5SrHCXf7tYVJKQe0WHxc01w/c43Oc7vF5eyGvN
hf9va2A1OHtI5MRqbO04pul7cajkSuBOJt7tOrzwF3yF6BgQwF4pWrWpn7Wj+u6A
XGxgmSUXbI4K5TaxbtR7VcTBrrfTP5vrlaxDbIMXi4bLR4q34wHqtpD1q7xwYJN6
1JCP18gfpYe2x37MvopNAOo1Bh5Egu+uYF7pqGQn//0D4TfQWNNvwl5n1JShtMl0
7XOmrrH2+aHIBFnQbzhoDglv/f11ByGAalpYIOjQ1IADGy2V34JmPqSVrBiuXTVn
eOlUPRO/qBB6T3Ej3Ze7GtxMLU102208HPX64/7R6QbKty3eWHHWL+7+HWvEz32H
G9HxRtGaNZFRwn9m0Qj0W5i1vkakvymw/QHmfVEIJV9KTk4hor+UkBFO0bdBMifi
gCL8u3iqBcfKDoABuwJFK4+OCdvwXry79fLHhyBcMS6Po93tQoOLqrk4VtjKSkxI
7fWFy4JbMYizWqroixDEuutVznZSkFegq1ydZO8rIeZRcWA565+vrlz5+KN9UmL4
sz1PQcp7m9U848fnuJYsRbgFB31ZWwlVmehg7eJyO6EZvkrU/Q72M19oSd7LRfv2
QyG37344ApfmxE0YEZ5Vdhoby34CVHMdXLq5xrTZayXySxU/sUU8yPG65NiM3R5Q
WjsmBNkZLIqVnt5dDWcLL545FpA/BNzPaSRvm0V7/zaMZHU2XCXJ0JbFtrdJ71rI
TI6uiv/JJRMSFp+NZpgj3O7TC9PrK61ECPSHByg9k8PCqdnBphPog17jGVqirHbW
Vcwjxs8z6I79lMZ3Gw1fmGC/CsO/sWhPTO+tj0dczMVmQbhl6sKK1WRUdbY5RO0n
OUeo4TLmr5i5l/WJNBJyu+Xq2/32HNzzCulaDhDr5kdmseQeWgBhf4bcNWiLoppf
uyeB4FhTBYMu0nHiAdVI/H8fBZqWbOsVndayegrA0vQUC/7jLxD4k5+5SSQDIJm5
KCBND+vV6uee402fu+6WDr2n1yUgQZI62liHBA851YtU6zzfhSzAppQo99EFbMXL
4XEhE9LQ35AWr5jBtaoYS2/MhXRlYxRcTXNK9/otWJrdgYmcL2Ewodw3zjqAUQhU
JCQD2f++R6z/rOqn65t1Qw9in2odsQbqZuFcdu81o9SNH9CxqybdUjPOapQk/UpE
rBh2yqUPVBnqEUMClGUehrLn1fbsq3htOR/ruH8oDFmE2e88mENLa39llj8YCn02
q2ekdGPo7Oxui4cfQha/k49M3CHWrsHuKX9zfwGZSEYYPW/Mw/uajX15yTeAfKd1
fcjxSUHCokoUp3ZGW8alU2TTEVohIJGUu96bsplcjpIW+RAugX+pEKCF0+hs6fNu
9IwHsgp69qIblOfQ0ggAJGtZp1v7ecrvFuhpK4RlK4qe2qmIAzdz50gwbunPi+da
WzbZN+MKo00ynEJf79vzuYy1NS4dJqmmQmQFhSjsLau6Pv0+RseV6NiK2Dzh8p6f
eulr9zUELP1MVFONfStEDMZ76+hZyR4carVC1VWLSbExkOpLENNwGfD450WuflY9
YGDKpWy3DpE2NsPaWR2+bVC5vvfGRheYD7FkTT4Z+BdBga8rhpl3dix+5qFSIOkc
rfVFHM5b7H11GwYjACXV1M9ownzTyHL6A3kp1mLi+h4W0CGA2wCqRKTbUi7T3es9
Wi+sNdh4ql1NbazYYsv+KRtDuHagRXRA27M2YcwkS48Eup60zPBlpzHKkKRy/eVa
Rjt6waQKH8U1Elhe8emCUtRETJxCSggp4fbt0fF+e8IC69T8d+hvEaJYQCvpWZ6z
7W5sZpwyWnqKav9aAcC4wOmnkpSxxaJ7K/Tc57sTUJo/jR4rJHNWlYbvktnTFLAp
LjStrEtuZtemfluxyXo1/SSiB5bUEIC0SV/d5Kee4Vim43kEdoQcjWLPtfE0Kadz
IgaTOoaPSL+WiKVPYwSC53DMp5Dki1ANZYergQCdgMUOigiF8jPjVeR1+TmqBi+B
NOsCNpCaPc/wrireLfnyiX03n1lqWvOTrOckj0bHwsaSiBW+tfe3MzxDw74Pbt8Q
sZgZk9eXF72UCBidm3kO9wfyFXnQyKswlAhh4dxge69Uxclv5A9idfcXM0RatgD7
t4FSKMkjtDVsv5R0wCSHRIulfN/+sr/A1ADyaDzQMwSZL3D9aY6Qm9B0T4u4lIpp
G0DGQ8F2+5KhCoCXMNIu9UMFSbzlqjsDznSTRjeDYDSt6jcQ55z8/Q9Z0w1+Trk1
iUh06ivDR3YkK8Wc/VnGmCPqTazk7KVv1doJaac7AI7++WiwtP5l34RGOmoGtkoQ
IuUzw4MR7rQjzuVJR6NDewLGxWmwd5w3DNtYlD5N8VVZRRbTJzTumT3ubsVnG9gM
4upnbimmb6trpWhDllclxME+4Yl1Z8UU/MuOQGwAe+ggISD5L2zGvTaIGSmW0LSx
c3rvZOv6IxtZUnvZvBxDsqlDqJuZ41gIWoVuW4s+9z8Dw8FE/C1Z/ZtXE5IowidH
M8HO/q8u9DOvKHZ10SGLI3E0a3n4VBs2/Fc2HEqy4WGK2dpPfiklrvdwhm6DhRH+
g5xIXGVcfiKVVwj/xgnWJAR5zss2qq0BHPdmaH45uSJLi062DL8TuUvHTDkqCmXV
K7OATV2qrnv/BygwW+ubdo3INapLeIs3h+ecfIAvHTUBxDznGcyU3ZiLgLMbZhbo
rqMzgNV+zlU/x6graqV9JuCIj0mMuFwFJEuCLBYctBBDnCy+KYGebF0Kof5V/GJL
jbZFA0ekFDPi0fz5iaya9G2hrnOY1fTp/8bMv6fepwG3icRB4+k6qsAIodnsmlgI
VlBn0lq2bgcXa8l74A+aAlrU6EFcICgtBOxy8qg56X8u12Bk1pjR8ajYRqbUpvl+
5FalXAKwTsSEGKvzLBhlLm8BXR/fF+UdUIXzXMae8US2SYSr4n8D7tOgjJb9LoAP
h1tRxlglJjAlHENSDEQ4uChw3U9vEt9C0YpFFoApOoISQIv3IzS64hU+9LViKSZy
+xJLxZQLCybi9kEULQ1V43yLC3Z2WBu17YvPATCw2xh69eWzEMZx4s/emNiuTJIC
5Bz5g64jgNhMlHo9lxxqhOA5wRVP2rLvsC60L4GZRw+k7X4v+cSTIPs1GO5HrlLL
Lg6sZY/LmVC/gHvKBRdkQvCgGraWU+zCLcXutg0lkf0QlIdIYobBNHW7PX+qqYW2
6i7FVUJFL+zvxs/0wIJhCFXZICCrqmSS+F8BvBEl78NMn77vCo+IxZj++ZBjs3uS
uWTliWveAyFzaOpQLdG/cl55NhsQxHEt8JAxzwRfj25a1M5L9J3qtS0y9TpRicOV
CXOMs93sZG1lktFYUhCN1twwc3XbW/Zg/guumTJ2vwuboB4MZYNakOPQB7SeArm3
AzJ1vE3mp2kXRJK2e2qApwL9bqBjKm4pjusCoueiCAFla5btd588hTB6Mph7MsE8
pg1jQDX7pXS+iI8MrVR6n0o44phJqu+e7SRks9fZAstgg/vm32QtC7sNkfw27ySz
ld78UJf4bNAY3BE2Ss4pYF0x3BQtoMXtyVRfwwkWdzz+fXlT+Ynq7fY8PHGzuTvE
6FJXiddBun5oq1OP1M44m5kJbRpKVLX+9xCMrIbsq3qygpb4oy8aq0yoJt1oSUqO
adDWvpgB9TlqNsRtIt5KG2B8vUiR0fFa7ttCHfg42na2Il6GJVYIjCPHKqrgZzzc
5rnONVGdxsHSF0MEuaZPUURdGhLX/M8Hxz4yUzJIaI7RKKgCC1//6JJiSUUtNtB2
sW7GSU6biFTCzXySYU8oYPn0pGmgnbnkNU4GTCOTziSTLEGlSWII94zwVwB4bWcu
5wVpJXHTszi9pqx0FyzhO+phYcgltBoUUjF+5PYSvOAoW3n1mypTr3qGu1IfOBiC
/NxZvMu3IhrUpaltz4z53N8ZAT8PChO3gloxCSdDpnAexGOLvNzYdvLUP9fW7khi
A3yhQzmshAYzvc2vLEtjc3KdH8cUtD7H5rCVg/DyQVmONmoW5409XDtVmt13pr/p
bycrt5UzkkCCaSIgnqUZ0lUqe3+ORHuPTZPIezV/OmKaQcJaTCZYxUhe2KQB4uV5
JilFqVUH2/Zsl5bF/vvhzyBZQ6ZNegw/o+jGS8n4Xp2MeHpn08m/g7Jii3Dc3Umt
j6qkDx7N6jwn1LPwo7rfG53rjJIWbwpPpTm+XlRUkHIZbmLai63CmmgAHM46sqXq
S/IBRxNlo1phA1xyEbBX9wUFbRHqB8TN/0RDzoUMw7PdUbxz6yxvobv4sHq0WN63
KSzdy5XgDQaG0fimBobBBAJuZEsO+KZtNwhS9uvIgj6ijKHAZmxwCp7gmFXCSkdy
BjcWth9teKDqSj/dftqR2/yyHQU7bpCTHRPuXBgrZsKJENy6uP1DpDwxUDRzAvO6
mVgdc2Fc3Yi0GkMcPXpni6Giqf8s63Ti5JC+VDgIwIbE/r3aaz2lPaVC5awMLext
Q2t61t9LKzJBmZ7p441AmQmV9s1GxDqbJqNrRExt8uvFasXwz/TfRe9qCEJ8IIwr
HjclTV9/QxQD/v0+31mzUFv+l4Fidd5n5c4y/f7xViiGdL3gtgd3NuMfipXD/5O5
RPARaNQPSeJh2VXgT3dth50gcysaMCXFTujan9mGmKdaByw3oB31pdhLE/99zMQh
Tk0R48zq+UA5fpznJQiH3ReXvxZcLzajrabuNMpbWA5GQRDvCU8Vpcwnt9ssJM9W
ZgMGwgioEVMSkBDPvcnsVBlNgVYr2Z9Xr8OZx+0TpjX3GDelIZmHjWUM5x2XvadN
BKsyZBKbMLG6EPGGXCx/jp1tECoN69b3fKIp9CrgG0FYBOOtz2rY1UySMXAdj4vk
LgqS1FRicy7j69ycBFzd1erliyn2E7RtKgE46515fwSZ8DmDA1QXqthz/iR4rySm
UNS6Ina7yY8TxXr5THAPysc6HqEdSEoyxHH6/Q3pQ2a5sooXR+KG1/O6f21DzFnT
ebVVeHyyo27Xn0Z4BPDuhHnMuUaiyaNkvanXOn6YOwzmn4sjFcNOat0u49T+uJ9P
hfM5d+6O5eYqJCItzNIykkDerNzbNy+cm1VnYpQzbJ9vVz5vDSF8a3aMTay3R1HB
zqQo2phF8jFe4QZve+HD6zRLwivI7i/gH5wRcxFMQ/eMqYBgGaZAMhshP0kIA/qy
PvBP9QgfKUgCAAu8uz2LMg7YaylAZcAEZET9ViKUdDYFu4ZOgtBKBinHJIM7wmFf
SF4bw1F/48fAQyirOGo3uuXt65MZ+Jy3QGyGs2pO2Qf+FpMhyMw14zPdll9r9nHX
mVb6qq7qnH3F9LYpDGXK7moocRK2GcVDbaQ5CEUpNJQE3m7bKEfD8XdjO7MD46bG
lLyHEBy5taQUnX7GC8bO2t+j3yhtmpo8PXfRGQHXFrHTE6AtM49Qf819YRAgCFMJ
5SDJc5ubfHX21PkSTucuppr9sA4+cjedo2qVT/w7eWV7uDqKnqDiJub9tTqlWIb7
WRquZhecZ4CXTCG45OK/h0s9NYlzUZPE3ZRzxH4L04929u4+9qYUauNgbtOy+a2a
UAALsjWAPyF1YYJD+w/cf7j7sLdfptn2NXeb9qnBrCzV8lS+EpydEmd1Iu8zrjG9
ZjLEpNYOh+DatwlWwfcHat5SrJ1SAZBsxNkJd+Q7amLGWs0YLvPZ8JZeNRPQY/Z9
OREYBW+xdeVg+10R+ncNR9BD6g4xKAM0TwIoeedVdO1glAtsmH1712zPYyPxsllc
Be0Qkl6qjLqt9pcB2BZZDsvpmkOetcvq2smHvWjQk6Sx6dxLcuaNsLRU0Dws5bha
9mg8L2mvnAZAJufHTci1SFSIvZMxm/TwbPCJGTvEU3ODZ+dGR6sQ27gmmNK0WBGW
paTE3cwVO0VGw428EJtQ240ublmN3+p/UVQCIiAOPxzbqref/cEPRIEZ4d61lh2N
SnhBE+Nj0VgLmnvJgxeCVkcXu9fWGNpxV/9R5dQ4xoqbQupbRUOaChppJAYvaY+K
VydJ+3TL4VoOk2d1NDylc+z9Hlvudlejxs724BXCu0Puo4L+wwJAkqoEN3g1ALuX
ugx2dwCV/OG9TGUVY6vRTxeaGeeyOh2pZv/EImDn8bPZK2nFy65FSdY3mWrX7igj
WMbRBk8tEc4WIPUvQ90iKToz/mAWUxx3wF2n/KPgN0AFIshkWCs0PLtMuShgO+ee
dd+5k/92XGwMfrE6NmqPtMBaKRHa7O9fvMDrXsObrG4Q8+u11bWSPSYvzDOFEwrk
ZmnQl2AX98Ob0veQ5MK9cEazmN9B2mEV6Mx3gzx+c38rNGOHFJREPL1ywRaeoAT8
94dsG0Vj7S7xSls1zBjzx4TqKML7J+9ILMBVSVi9zg7+UEc5DFjdy/qEedOLqQXB
U+Zv4p2RbBnMfyNaSVHPdnlUWEBiCY14OEnT1S3GF2kBYLiRYHX45bZGjosv9snG
3pFg2KzhY9hDacHUIqlgghVeVTU0aplFspvY7HST6ZuMfNPeqZyd9lucaPQRjl4I
rmoTz77lDmpNZl1eequNQlNJI7bUFNrnSoSFCg0EpjjteYXo6/Mxi/UXULlG48df
Hp5vi4MSLHyo+1myUAdXhnWMs6ER1EkNHienW7nj4RsGlU+DJBzRIxTckjctbVf/
18inSQ+StplK9tggDE7H7t7As1MBSiTuiBbF3Pc/k5BDMizS0zrXXzM2v6NSR8F1
O9KAMt5VUPv0qYK76xAqqLZ0JadtV63fDHZL3xHaef6YrThbH9lFgNuwEoLcm/V5
R+g6xHoaJO4MLF+H5VO9k8UtkRm9VtoyXjhq9g4qi/fbgH6qnIKhkkuoczXVOvhD
S70oaO0aaXtFuAWvDMgyB1cb/YanDCp34NGc5JnapMesEH2ssYeYECqZJDCEPb2w
4Oc7Ne/CIQth6FyuKFzbONLi/mGQaruS5m3xNtgJ+/EusL5yn3Gc5u9H69JX+jYR
nwbW5UtAQjIMJLtBallTeruzvkCI93EYbIuXAjtmWj3I3Jb31lCfz/P/AzuraH3L
yiL/9va5lpGYbiijxR28vZxOBH6cUO7TI4MlE1XWGyGmPHBua/BI4gWGL1YZWxW5
gh9RMnCTNUmZcoThY6tBQH7F7ER2+fi6anVcfRiIxiv5/FeDOHt+Eum2IKWIqPBG
shlJjUoQTlLQOxaxubPT848vxW9RAogIMAusmZIz9qFCNXIBbFh34XvpcXpIGh7d
PZNHlbkH+rt4Fsbo2r/91ZjJaVjxTho04TyzHSkdkPnJ4oqd45hTjXrslq3u9X4V
k6PB6nRsvCsM5uXntyO369MAjZVNMSFO8eP4DDr2EKr5kbR8zaSPzLFkXJZmhees
idOvveiNQqYj3Am42kzKFQRwUCIhMtYrMJpxYFvFowxXEUwczgCAF7Ve3nlwvC3m
S9b+7t36GI85OAfcnamndfVJfzki8QczZbuCA3NFUTrmo9jVbL5uzp25ZWFMMCJA
zaFpRxoqkEKJowwBHICp2Hf/zysGggylHYqjp5VXDuycqEVATLQin2nNZ+GWcY++
Kb2u0ZxOCRtnltfrVg0UPnV4GBeFRcw25jfm5pmgFu5tQ+mJU3nbUK6/XOBdbggB
b8d95xzaqjX654bLETtkf0hWl8ofz/yPVfHZ6o4GUDCXeDQUgzFxpiUZcV9ZPuS2
qAkFS3S9aPOHjW5+GCwe4sO0fHQAxtkOdXBcEn6DiEi0CATqmnxM2Z0RoggjGswx
DwLEqopNa3iXqcMB/4wQ4JQRPzw5CKdSvj2+6ruKC6GCQQVRco/TZ9SNBPnAqA7I
lXFxThNUl7a9/qYV4hv1Srx58EzqW817SFvFT+USlc2l6ZN4Kv6vOoeUu+Eg328n
L2krPA4HY36HxR8RqjehZaQnWK01IBeaR2KWTa0792beNbrvrmjebkOoAExloEuV
laVgvQbOGrgpIAvmg0B/wkutIQDayAed5zoPx6dJtwy+dsbWd3jN/UReuwUzMuhE
Bkm7X+1AdHcoScUVZiyPof/XfLmZnq5KPkW6DPkskSjULl9w9sp7fkslbNn94mm1
zQM4kglSCr2IyfbZNH7YQfcANVPTic+G/61gPOb3VgWLJ9JogJS7JkT5AoSuay0/
Kp9Ab/j82lLC2nYEr25slfQFD9AYIbt9a0gF8rYJ3vFgVFH6uP/yOkn9WZ1S275V
2zCRccL45yG35Hot0giH2QQNkvFnutE9pSreEzxQARxg+BFBj7OC93hFeeRpNnK/
bzTQe4mz0J1kezj8lWjob8f5F5DL3NKsObcdutAOlbUBS5g9zgiw6LOd7yZSNUST
M2x9YZ8LTWP+evaQHgGOz+Rvyp7NVg8lVa4L2TQfrO49lOKcmmO1d+ofUk9DGfwN
ZgxtXAM93VdFOrfUvwe36CZ1WrW5XzgBzH4Pt8hwq9q1B/14/2AzxH4+EOh0RGIs
b99TFBbfAPrvJIobc6+FO2M2uHY73cks9/T2UOYah0DDUBTlQlYMkLiTQ3FDPfMi
jNf/ekJrvtCJczWBqUpML7K6ZFnA4px20pUOF218NfCo4BhGZcRXXlGJgI13BGv2
3CfwdMve6RHAPBfMnK20VvacC234e6HvRyBX32iQaFJJ8UfX4X2fxCiuglPzqNQM
66frao2kp6xOSIvQiMQIUqxhXr8M85vVFQntcaUvv2ZCLmecV3A6a4BijP9+frGu
hvhTz/EX/vVJWnZnSRd3EI7L3yZmqfokMKPEXLKNMCkIWLFrC6iTmp6MgtMJJ6so
vv7TBS6MkQ9LIoaQBOAZoei7kVnfdBS1ZSBXvk2fHqda6bZWv6FpYy11XIAmSzf7
wtBunVA+HL52hy7ZP7GJAM709Y91/nm14F+WiskNFfroanQHfyuEjwmb+yf+tXKe
UY+rIZ4Vykfwo1bL4NfNuTGKBwMvOL/Qle4RRfr69Tg85coxDfcIEV2tWdfWdGGF
iE7tBsvhVg0hN7wurakXKp01sWIVV/qrJLUsz1xgPociITUI8ZVzdNjy7hxojB6T
L2iBalx2XmESkL/r2dvJBj/H+ewD7KenVSFKkIZhzTCmlK0S9XQcpCLEFbeE6Bdb
y+df3El6C/Lp79O+LWpRQN8CtjUTxtoi98Fid1noRxbXgsziY8BPf77qUJGvHX4+
c5ndOJ7GbjktM84jJ+2oC6WCiuF4kBI5sDkf4RaKp3GKt/c4uE61adC6iqWthUg2
hvtrhccNp2OPckjqJpRNOB02tOB/3l2Rv8Zs6iIRTSgQmityR+L60wDC9z+OjfJZ
But/mlY7PUwCR2nfocmXJNhD//ecUeGqmkDxfRPX1I9DXAO7klDzkyv5T7Ap9ygn
j6SaLh8qFetFj3tYodavswOb6Okg5PbWFQU/3DB9qgziSojbec3mg6WaarQYc1sg
b69svcaDfNqUAC/+RW1kvjAn3yOpIUiScahxU0T7+VKeiOWsOSFvYY8N9eN/N3v3
ZfpztpkRoaU70D1ekKkukFlozJtF0JTD+WwvvkM0wGvS4x8ndIIfqw4NBlSqwur6
PJpo7byT7ht+BkkD6S2q+rlG2QeqiUyiZo6+uYDerYxLQVFy20c/KiuTGiyEXg14
IKzxWVTy9SkI+N9HWeqjWazkQxlFvDsR6/cdinusmp00kRAiJYDsYChmnfp5Xo7Q
zTxn/+oc2ZO3AFc4W6PNFuyC1I5AEO5TcoVTHze1u8EixnYvGqf4MHpGjUdKSVgw
q63aHQ4FL39tJaT0ZhoLpAuMRxmnbqXZL4Yde2MqBKZUZgYa5oqI/UHQf2YSB7Bm
GX6brVQbojtshlvauQQ1r6CS+lecjbk/IOMzJZEwCXwx1UM79hUMHJZX/tqn/cPX
5KdqMekmHE5MJkYuvsxPlWRr01ImjfOaODR/c0KN1+wbzuzfzu16MHUJT/ZOytaX
LCVKu17FTCySbanzKkwln26mdKliLNkYXfTDHAWZ8sN62l29pLDZaIPupDQdRSIL
fj1pl/kDRXaAT4EHOZGYyoGC1Z5fHF3UXeaMM/IQUw25wzbQJjQnZVILe2xjbtEi
PqZy0LFZ7dmwC/zwLAi+LPPw24nDx3T66+sKXXBXhRW2Ca7TshA4NoNeA643YdhE
j4hrAUA/j9QdAaq0MylngYG/uNRg6GcR8dnOvE/JeI6GxhxV5MFcU1pzzZHYUsIM
GLNFlumD97EogFafe3Sg4x2y0mHCZCkb6xsCwWz4LCSUeXDDvCshlUsIGHdXlA0S
wzvKMOqpthxA3CkYoZJ0bOjMM8CmdfM/Zb4kLyquo+cvZERvY57hE6ip2JLGEmWl
5YsUBdyNr887ohVCPppAKZwVNQNSmRd67GxumupEgr8V8xaodkdGTFAdePAS5xIA
Oi5s/u6Kzma0P8J8EK0kcNK2OQ/u7APbYxXgN8xRofCIiMNmNT2FDfYtlcqBiR83
wS8dJYcHAAi8QZkZDXeRWgVYTny4tp18WmjNzd8RO4fmMuIZgic2sZb8x+/KdQkF
Xy0BBZ9RHWmGEH87jrEEkOzdWld6KqeJi9qsgn1XztvlMeKcTE9mdHK83X/+AzsL
Ztx4pgPZFVwzCO+eRddQ4clhNqOiQc+vNo0mbKOwI2HvAidYNnaqLnAUkFyw00RD
XyXFI3gi0Qt3sbAVBWy/LXE+fBAQ7YMMfMM+L2JlRBGC+cFPpQFH8tJSYPVq8dJJ
tC/3eiE2a3TTBXirsgvPEl7Zd9x+psmRQ4pexZltd9ZU39BxrU/GTwCWi+vzO4e1
xCBXaufGa32ZFTyhowVmRgZoJ/G2KsZN2Vu3pnob23mhdw2eSIa+9fqtIRKJJhFH
xSXZR1gn71K4KJkGJ21iLJrY/JVbO1QlmOwswInigru2ZaCXHzCtQzwlQPtH7cXY
AO08Bj96MUtOoEf0ObVq4ace6QKZMMN6gz2QKbsEEeMFEE3Vcrp/jnBGZHufh/PB
XBUA4yubOI2nMBWclX+0sZMHoW1bL3uZdC5n9WLiZxV4r9PMNIvGAtllwSr+lDhc
29IZ7JUb2Ihmi3no8/QYFOAwpAI42XgDWe5+MZq1hl5hC8ZOmauFM+b095GLYrfR
BcmDdD+GSNwM4SnuYr+TZ6ShNsxToKkQCyfaPGmKuJEC6W2DlUwq67y1U4PG6O1I
fWk/QYXMngCoyTrPk4FQBjukcHn8QCTQlKGVEvWwyPAe1kY2FjhvW30tBBAth5UO
yf2CQ8wRa2Fg9nFITNNqVlG/nUEHAqMADG9snWRgjg0dV87cbGmsuxVK3D9Z/sP3
XQdLmOYaOdTW0WcntEgNh324AnwGBVf0Fkp8+oKXGblzDNPPHunD6HB9D+zp/HUi
S8KLDfn0EP/CFP6KvEN+6lzrOF9RVQPRvLZ4Yox46gkhAcWDnb2ggSfos031RhsU
EHvDp/tVRpxirYkX41a04rwbVaBLUxyYO8ABfVzEVmkpG6+d0jZKD+DGU8IGiVuX
5uspLS6d0PAXOhhyLUzgSIBLC7hRybZeh6bjkogXIajBapuOBN/Q2jOmKytOEnTC
0uEHKbV9eML9XcZUVCOcML0s1i1JLwUdwY6UBM1muPwT5uJqXgkzhiUYq8SK/Hww
Wr13bs3GUq8awsOncMO+mibsmCeSayJuF3hr7o7G1quY/EsF6fKUxHtkathqGWYW
AEdf2a0FkTeY2AEC/pRJ/elf0dUakAFReuDyu73dbSOmBSSW/a3yDvv1vqf1N6e2
xhSYiSL+nhU7UlWhjMysUhKyHVbaOWtpInSWvqQY/yIi/sQlEa0DvrVc/OgQdU7z
NBPCeLktjw2+/N6HlmJPWASqBueKomBT0JUoRtbhdob2aaM5brX9bdsb34D575cR
/rG/kBydeQUbj1RNbxaQWrePL/3d0q7Noiye+TZ/qfo75bOmyhXJ9z677472kl8U
B0bQVnlIMxXHdosflFDassNB5Jj6iLdXaiQojGjsLJJzvmPmTRAfWmkf4S6nsVhN
pDNUIK2ERylPG9YZmMW9BWINU/TSDLSP2MVJrv62pz0wV7Z14GUE0VBan9NQmj4u
+9dZJp9nR4AfhcfLh8xA47vHEKVHEYlODtL2OaQKXZs8ZvBAVKVJVAgW34nA+sEm
kPaxLAwM84C5bVtXk5TzeLJUZNJn+U/AtbrnUWdutC/3pBDzyIXobOn5mKEi6VHL
cSqJI1DQStLA2Lfnb977f8yQyUkQG05qHD1P22QdgAkJ0Ktob9CqZyiMZNTUH5sh
XVRuQ6yoCBKkyPFPpCWwG0eFrxS1VOZr6eQ3KwK9IQIOYL4PU7B9m5TksrPTz4YS
RPaYtttRSu5jT/tylew9ZXbXvGCpboKtvfKyVa9uy2WmNn5eVCTgQ5jCu6tV+xn+
C+g18VYydUk4aVJPG8Ljf70t4Gl4j57+6P2z8IQUpeFg9dafucDALbkPLRgjmfQw
oLQJathZmhLtmGfoc1krkw/sJAgplPD7JNAbmgecEsWyAVTCCUztO8DI29nIzC3b
ZvVicHbIbCrvVspDiaoyA5e882p/r76DNxoMdu8in1NqS/jYCVbygMVe9dVS34EX
vErImY3Uk9yQwCIj7SZLjeRr85jDQjSqFk3DmY4TtRNxdYe28cP1toDxOnFy/ell
C+8y465zVvMBi6iLAOQ2zy84UqOK3x9qsH5ohUYqoXtTgxonf1MrXVrUClwTi0O2
/oqAvK0F4b70ik0jbvlv6ZU4tKs6Y4Md3yarEkL/m5I/XufQ6et/s0t4ZLNyTuIk
IPpLCRCeZINvw+pqtuDeuiaAqOCsoJuXenA34maXfpGdwMUQLeqT4H64lnw6EpiC
jwsk1QC9BY/2G4ekrAgZbPU5I6wRYu2CnlPlVg9uLqU6pt/zDyTaw1P/59VEycTP
NE4XT5K/8zzXSLTJjyTqOKa0+YBtJeCQ+0KACF0MNlaYLa+klOVwxdAoYFEVxWuz
wVX6MFPiIwWi7qwxMkm4Ycac5016GlYZ3FT3HkuaiJAYdN15UnWZNWCzy3H6Y7Pp
c3TeQ1X+j9cUlFNGaWzXRsYzDsVt4cYRfajOMYmKIFo77TDDkdoQw+Tm9NWjf9Za
bjjHzafFRprb+3M1YvNFClZtDqCQH6kzmDFXIe0Jrh9JepufSyaVN0VCntzcety1
SvPEOJC7fN5plwF6hgfWArHo3gSMMRBPsVb68rzzrrFV7Qhmcm7my4urEc1l9ccC
YGS31vYR2PwnFZjGAX3W2zTdMMRSJtrzrhW+oh7Xa9jIz/0QqObDFoUAqgW3Q/fK
HBRz/OyMcjIu4oU3uS0A+WHEz3ot8iNOQcowIgGPEpOPiyBKmanip4mC/S+MRlT9
cqJYvnMucLvE2/1G2VRdF3k+MprV+eazU2DMW21fFcDeGCZ5MFWL7IJ4dsQhum22
hYlCXrhrZC6V8YKbhBRfc8QtWWz9tqoUhXOvg+nxeK+zt47EVWyn95wvQi+mmBsG
UWXbA9jXb19QXdwUgHgjdJXugC2E/AVVpnRXhx9gq5/h68TaXiQiUNmUwJhmK2S8
18LlbLENKAnfleel0Slp9dWhl8+boMMTY0Ub+WSYpMKIbNug4D2KW20vJN8e80kP
/LqsSGD9Lm9u9hDEZDXfOvoq13C1Ehbo+U7PB9J0Nx1PMRKoZZY1gkvkTImB0YGa
0BN65kug4CVHB4PxalNeJsJk0VU4k4yjwCf6fTDNUgJWu0DP1P7z5Z5YDsOylRs9
ZIPGRlRSutiTtzC+RocKr1CTyYN6mrjMpHmwNYd55ws0kjNvpu4+MBf+UVtH4KYH
ddJ5lIXT06x/TGzbxeGHFMWyZecJLxWuIWi9gAVfUNMtm0QCMdS7PVx6TZzOblv8
sgdVl1/P4X31ixlw7d+Q+TDU9j5lnB3pCBWiw9J4jEEnElBXxJ5VHYB8Jr9//JXl
nV0Dk48NVNzaVdc5F9GP4jyqkHYMZl1bZ1/mPq6xD5K4R1OhWxaT6EGpYBdWOo0/
0GzM2G7HV26hR9L4Ufj1Sr6DVXsP6CdDhIaOzNHQi5Kn+6QSDI4g81lG7yTmwXRb
bsz4f9sfP5zFslUju8DNSXwM2MExYbUrGkrPEEJfJnzKfxkngP3R8OkRXUmQyfLU
JtNOT1XyNGZ6EtOLHJLIHWmqkgAlqZGY9eH8VHdEBxzDHwq9UDURvgGL64JfC1u6
yUZ50n/asrPh4y8rFc6pBV6Z7P/889OH1DPnNhTIJHa7sgEXP/+AdsvL1qaJKvlO
Z4RrT/S56WRoIKsx3ktPzbHk69ELq82/wQ9ZKT3aOEJJ23gFfZ0V/9gca3C0PIA7
V8m939ULf6psILgzRxKmMeFQ2nELMRlDJCIEkVyC3H7lMoXhCgyvoY8q/7VD5b4f
S/Po9rNaPOZxXqKABYF/+tX4HoDp9Il/2D7RhggyKjhAShCvN6+tScq5CsAvJq/2
92RZPwdNwx7tpKjWJ1+wGYNrKYk178+9XSHS8RiMxA+wz6EoY9zVRKCTgDK7Dtf+
/kdO5IBqZBPHGMRTlM/WWSLmfD4wLIqQtDNui72vhI1OXurOmdhtQA045Yqig+0J
+CrEyhFZhH/SXiUy+itp2Iy6vNFpviQXTwoIsGCCuKBWeQy5xmqB9FJwFBukQ1FE
jifcxEjL+IrDUGDjqexuRsKXvE85fOO+4vaNcO+nTRbEnlWh7jiH/6ZsIafgm27J
znbpFt7C+X7bQ9od/iVyzO6mH9m+pKJ337DeGKaH0WWkvgjUaIq9IcxflqJT2DAz
T75TDSIGOsEcKhkBCnMUpwIt18qYuJ7gqRoAAf5CAomoHb4dtQgYuqk/dEkYQtnc
HW0HnS4Swo8/l2DNp1VquQEgPAsiz3tX0V8pBdvQEEwqIyPftMkVLECnGPvyzoL/
HTVNf+jjlwJUrEWylomfzkFQdabSJVa1+/PjHgE6U2hYtcq9k9mx6n9vFmeJ0z31
dBhgkqzh2FxxC4Sc7ei2Tyuny0zwVKha1OBCSdAplbs5TKZB+o50seMgW0AwQ8FH
end3A9Kxuy3hfQUuarKIG8LMdc02yY7JwUjzqtjiPoqUX9wPL/wZMo8oDFAMugs2
v1Rs1KJXmX4MHbWi8ThawIH0G3WjWGogDVMJS/lPI6dquVNtULJqXC/1Ux2qs6DJ
MM18f+FZFL17gxp7h1K2zdSOwst2YOfK2Bzl3TohAXgj5u4RW1PJA1I/aNGTtXNG
Xk9jwC1VGNyrOErUzG9IEns5+K3LLGv7YAYTKu9W39oZPZH0l1+pppjLUqf7L4bF
IbiEpXMUk75ESCGCCSh1B+jDFBVpTONGJZDuQDXR2ocu5TQnjIbJls5H1I03IylG
OTMbpNSNlMJ/HCOshUqh9e+1brN6fZjvlgohcdS5GfAOONZnnXahdsThDEczYrRd
kG1Bn5BJYH1G+XL2/bVt4RvRvcyGEwsUL0rfjVVb39ye82EwhL6+KyJzayK1ArjG
xTeVp6taxqoy06VOUXFMSwDIw4Nv1zf1lg+FA/mhJ7RDhaY59w1uL3l7wK6nnUG5
skelY/7AKv+4/sfGKsTLII8Iq+n0VLCdhdB82YBQxJjEiya9lXD8nu8Sh9iNPIgm
dbj4oDfnvcs9JxMWxIYQJIqF4t7tECmf+xf2L0/TlC4KWXCCQViy0b4UOMl/QbvK
oT1ZyXaEA5xTNbGbTuIgnciufzMxF0ykB9r3eqAay0FzlDllKN9i79MbpUC6UQcV
Wjufy9CPMiRQ0dxwvdrdLHBu3w2+PaNkLsDahpIM4xoh8KWyalbYhVEJFWty53gS
9gMCRIWirMmNg7V3lLoLebAvw2kF0iWNk3s84rF+o8JsT/tUa1xfrS/z/+wxFpMN
qoUE3dxcT9ZmfM3s+9/7qN6YJsEt2ahES4DKgMgMPkM0BfklSV6yHu5CttCob+qK
8orSXjfE7kJzDYa8GF/Lby7HgWSqOFkMD1AgbSHy1bJVvEemxEn9bvR+ngVDw25p
YyQ9uBFm35LklVh0R+jGe/7t0M/ZKU6wIqiuX398fh2mgQ5bZxvMFzxrebP/O+Nn
WYa4A45znMyiH/xn/Aaq/XeRN46cWoNlDMOamQusEd96isE5t6Cqj1u8DC4/CHmc
wUdficnBjOnUoBwiB1nVpXbpChR0Q8Hxoxf1GXVEb72elDq6lyVt6YDKgumiWMqz
9t/+WefWfIYdPxFdsvkMhNz9Yhoq6rViC6nAo5pLE3VEbofKfHCpe/Kw3PT9uEOs
tNx40ViLoebVsrOxWDFQkq9MozuTnxqjTudGT/DVwrXWVvZDP5fOwrKIU82VB+p5
wvkvsFDBo7XDiBrtLtPAspQ8fKQMy9NjUilC7vj4hjkGOoo4sdp2oFt/5deLIx7Q
pNYqYLegdljveylWNeJ/iUC0oviuwD51hjJsqbLoYmIIjBwOQIrsz77Fwz5ibXwm
+5Hmyo8wS9oG3vJ+DlaT5YxkZznlAFZBjSC/Fv02t8ftxsQhMAAi+/1Jl7fybHVj
ETBehyvRMkEO6Wj6PRcW8Xee+rnHVfk3L8B06fAKRGQXPKsBMfOAQnMkxWcjviXh
tw66e8n5dSMJcvezXb7kkn3Vl4hsH/kRdTJo0EzWJH3aoaG4CzsIMd9TylTg4eyi
20/f6herwpYsvA4/+kxJgyBdjNR15rvZvBA1Y2asZxSZlVktVEmlTGRlZTKQt8EL
1IkwfqArjuOzeWjN5ClHPOxwb8UG8DpAqsz9YnPWQfeVo5URO3gu16lEUIvekfH3
1utb5G+9RzSr6bO9t1v0GB6/Il8Jhx8DkYNJYDfQpl3q3aNyY1/buWl9F4FZsB4D
Uzyd7WtBdoKBV89xo52/ufUlijGsK0nTiRDQjDymjp3y8ykvB1xBMgEXNOZUD2/D
jQiIO3/FIUzE46PQtjvz1KPnVgeReEjwr0NG5kPUblBfG/C0JYBZXUswYJQvzJGv
ru8Wi0BCCYtvrG5iG0b1kwIREODWa3ZbdBrhWDakjlwHthbK48UZf5Ad1GmJ40+N
H6N1fcY1MyXK0N0vtqQ9/T5N80dY1CpFNPob9RdiesRYKVjuWZxINdDIBIYy8gkU
ObxUHOos9e5gSsJe3fOff5JShxBppwtkD8VVQpXmdp0Zew/XXeGDOxI2TMW6vcwC
hUw13KVcFaDUqcAfZCq3A9KqX9V83qX8MLLA6ikPCmDJ4jol8UiIjjPOq/dGiqeA
GV73gsHDmA3QP5DiE39oE9Hl8w+EZBoiNkq7rkLuBfOV/38Kt5mSNEsU/DCp7gL/
DiUlUkmFUfSsrRVF4waPUTT1w89ACOurf2+4PCcN911MStoZ95gDq4MGSuxv/Laq
NiGJFzVqOrzjG5Ww2QhDsbceWMfNrZIvbbDZCLOct0pUSk4SxFTWM5EEgSNhVu65
mh7Et7wtIV5w36paipW4xJeu8E+LvAsec7nWczsjKgjTasTniFR/d3jcvooGTEew
jtOyd4wHH93M4WwgedvB5QV9J5sg0A0bMsuxI784K3lPy1Bi/gcU33xhQJ/htjC9
orTJHDoPmIzf5sJEuDgZEFo1fktEXG8bpvKNd8DKKXPkGTVTFP3VZXPXEV6bUGRT
rpRU87r7kYpUxkN+z9PsED7DiLh3OtOnPs9I2J/tAlRy0t/GWEtn/DIAFkdBLTeX
QgWxzufF3P+frCNWHHtMfZaLac+ZOZPWONEFKJsOZpxnQL1tJH0kSu8Ii9HbRFh0
amRDabVfWJLVOAjDEHxp9emUcV0peyH/qK7StSilmONQiGSK3Xwwmk7UVwj0oO6f
A6tlDPlEZe1mWFVijLdELaGycei5okmQzXpzafPlfhtAYIN6+1c6SWKlFyXBJtOF
oPqA/0h4xKuS8RjGpRqtdFuBVdO9ktKC1AaeQbm8KtwNy3TWo8RY6hEchENglacF
Yph6qTOF3cNpI1O9FnslPiimb4jDUsOQwyJQhE/yKytv3RKDy7sGMQS9+xr27bWQ
exP6wp6fUNzR/NEVfsy16y4TXpnzKrRyJ9M68juS2+vfGSP9s2DxXiq3x3fGffD9
qJ768tcCJ8YeMuOHvKXcmS7wtTU5+PldYNZ1DnQZs2RrUp5JANTLmLCn+dMRgMhG
2Q/5/NlxD0nBWG8bqfFrV1ABDSutreFEfQ1omVtni1iKyS+DR7A2TInVRIvRhmXZ
yrUfRrXmCVNCrpxClLlurR37c4CLdPXXUNYTMNicZrjWbZpV72mM+ksLkMAukVU8
g5ROumLo74+GT9UCgbhfjt8E4+pnM4txwNESRMbP3WwCuiXPuZM6llIabs5A/Gkt
LjhXLOXQGg5GIV0g+FuchshJTp88EiJYfkiVvsE+3mAs0GAgEMTck5QjfYizo9f1
bh5qb+WIXPSmDJWuPYY3ugMN5FyJk9SX6M3/IPD/YvjM4alu0Jk7QEJO8SfAT/sE
leu6DxxYpBp7JJ1Tgw7vYeLZCkI6MXD0p6/WlH9z3TrDINpv26YkRnapeL2hldVa
O3t3zb5jt4J1L9zdZDR99qK+wsr/LdkUEM1tR5s5PmegT4OOArvan2QzSqxkIGGS
RsXCJga+YQovNamOkUmLGv6EfVjVy4QKF4egjCuorXY31aiEytpRKklIHVuOQgkR
4hXyz0k+3s2qog5n8wv9E5QDUtTSXjtzVk5gM3R7kSlCKdN59NDlkbgh3g6pIvZW
M4UQ6oImFkEyzB7J0Hcg7vabfMIw3DohW61GEKlqebePLpgKrzXZGL8uPUh+ZhFG
LW1jAfA3KihxvWiAtxJN+5lNRcF10bobXUl8FiIK4dz0tmT3s7cCkwOtUZCG6kNb
JPh1sLaPMnizfIfFUOJdXQDTZqAevRSMH0WjS+GhhYac5GEeL5i3Ln40nnMsMqg9
w5NwaCgLwwPZSoEGNhJuQ5eskNt/YnOy+eh1EaIHOzOcw++oVghxwbXB2KctOuJy
7xso3eqAQvBcukF9QdlLitGlnKkdi6fTrA9I3ii8b7LbwT088SSSHpq3ybWlOvVE
WoCedZxwJ9UPcecBgvLpN4uSFA+seEtSrWFkssJnASi91httRkkrX1STYdBMB6Uc
R4didJoVv+1fuQ/6FsbAGoCX6DsHBhQ55/BRZYnlHerW0twl+822dn5efDRwCy2m
O0dR2auAVyAz4N8gxkUWxZMzs2eSoDiqC154kV0wWKobDgZmzBLRmkSztCJ+j6Bs
6Vm6k8fx7elaETb+ID4ezlUsGrzI6H+xJhvZcw90OdZzNAiR+HiDZGhe27sZRAAa
hQbUnSu5OzoGJwwxeCvFiz9ZGZ4/5ez3KmpTpTESwVJ0kO342FIgrTKjGpfV9b1G
21/Vw67U2O1MIzpjsUGzcF+fQc+5RnGHX7uV36TJc7dlcpj1BTRJhOFizbj4DkFt
Mt/MGy4c+fPIUcP3l0RNTWxw4vfZWZjzZHELcWw6jItDjmNWyCtCAUAMzYLc4ixh
NrwW06yPKwwutiugDMqaP4u3/IWQ5tCduwgpuqEMzR3KCW/B4xhyUN+iZCUGtvak
tY7AjwLjhB2t0L/AtCyCnS9EAIU4FWIakTJJt/ZKrT/LzKUUsh33aLrrqzzBO2qc
IqmqPr7uCxAryOhKDiGwTviGVqJStUCNIKQ3aTShSnbeshh1pwW1DVz1zSmECgKh
82s6egwICsMd53ovui5RiRSiDjR/klRQWd7zPkyBho0u6+GvI+nYCiJNCTl88yRv
axmIs7ZyQAZFpJ5MWmh0frOaqaBDHf7y9dyJSXaVhuRV8HY3osvjV5aGhbUPeYf1
TAVA2oL7PccNDD+7GxBpxBU8fapRyyfvV9Ak9ytSNAiHGSknabTqWJLaupfuLQMn
MYv6VUtJlABapLYQdN4M9Xrgq6xEc96upuDfzUeWWuqj78ExYTzXD3Bdhw9GJZXt
C5Ls6+VtjNTU1lSViFelnKGG0SbVUggvJXFnHS6W3BPOmmKvIe+P7zT9rMURL6FO
+uCqBoRqYxC6hUx1HCfjb+J7sIIAZSddHp0tFhaQ2cuzCfThYEf0hedPVxFFKf33
z47RF+17SEALC9LCBLXPJdJAFwoPsPGLriOiL9gXd6S/00tkjPyWlKqqAdzbSJKp
/0FLJ9svjKaNn8bOnMHAP0yIBidHyW0Cr6fnQFpAGcLjsz4cBSe6QRjXCXwVplFm
3Vtqe79Nk6hzdA4UpL5Lilr9YkuBFYzFAbcWhXnHkdhFcvHVspiIH0W8JHgqJD0A
2QvaOJJ+gIlLvVoAHfy/0h/vd7O3iFUZEv8tltiOpV+KBIhs3CgkCZ5xXp7rUWho
HKhy4Exb+oqBMV2dua1hV7lZXxuzoiUIrMKUHvFkx+HKyQVPOEhUU3TnrWm6sbi0
XEV2NfSxtdhgZzYP9EfUK5+oxFDs1MdvHhjaM+frwZFEycmxJO3W2iUn5rpC9M+u
u9hgTvBrI+N0gX79bfrUMMpF9tmVo42hDtzt2+pf/g9vrF5EsRLht2i2Qs4TYz0k
JgCu/cjgGIqO+5FkzwB26qeMCB5uXTZcgh+3JbQQVsvdWBgi2ehubZgYcZW+b0gX
+qGuAuFNjFOu9jZ4QYXCIKV3cIjDRkh9BcUsjQEbIn/NWC8xuMjvGBT5uwwz0uUO
xeBXlqdIDaUuCNr6pHJyVVsZ1PCji4uBFo9Ch7JWSY4JlAJuIrayuPesXDlJZGZP
/meNIvZ5WDtQpmAtyfEJ7kXhNY56OY4c6k8+Vz/uoLwLgCVZxgblhn+vWICjQkA1
Kn+twv8jDsVs/+CCv8XApMrqEb1odDvXZ/Vvw+ZpVXxB/Ge5zeP7XPm18vxJg7po
nFoCZGNxpfXWzcFl4Eu5Y4KL/WHCjmovw9kRGkBN7MgeOrtXoB+E7axBUZyfEGOK
3zRkm7DdWNQ8uqK18BMSDfAr97AaEZYCp3XzQ3rC4Ab4wx0iVcWqfWgG5J4g9rqn
1QfCqwiH2yMgR9efPI62UklTMMT+OuFhUUkqOK3W6VkRjAZZruJaZSg+UaeeP+Ip
dhjzlA6QLFqnsN/uYZ8XvS4evRHk4vJHSOwK6WfQa/nCp0guw/dWlfdF9E8dbJ1O
bRgEDW0Wd0aK5ERZPpko30mIMHg39jSwN7stYo022uz0kkdvtaVuzn0V4Fheo7z5
Ak8bKCiG52eiPPXo20Wj3H1zNOV9tUukyKgio1w1lsZ5UdRuenT82BNPBhTjBnVH
iyEKvxZWjbISQ1zxo2ih310OAVjsO36KaN089sHEf1lD+rzfWBRLg68xJxXgSCQw
2MwC2FLPtqTHTItq4HcG0GbovBny3dIQ/QRTYpbXSWQuTYYeXXEzwr/B+6AlASgc
ygUMNSrlhzGVpzEumOlxjgXzP60aIiHxmmGQUASrUyepCeO0E2BdKdyQq37kTWTl
CLZLvYIyyxyHP0V4DzmsrnpvX2GMXSHCoZmiRbY17qLdg2YBKhTkgLQjLE38zFyq
dvtgl79CnChcVxLc3NOAQ1odDmGicUzO19hepcpkPrg1BL/8U4jHLW+WThJCs5uK
37BjHCn+zHTyqsN8u5+qMy4Vz51iWdiHQ2KdDRiUGIYLhLeR8cqYC/CVnds+Zh++
fClHlY+cn/hXes4yUYpCTQLX3v9vgeM3Zf2F4a5xhRaCJZS+FzJ4lY38CYK7dK/3
F0hTJK1wIniciDclpjLwPWvBJJlkvCfesnJdhREBXKYO5UReiydevjZbNLWqJyRd
kwXQAmVXus9QgGRjKs4uvTfEqRdSbWwEQtGFZCVv9bEfPZ+jc+tyNIE+c+PnIDuh
kVwdZIYj5sOAOALwo3RqOHHngQJl6KDhrj2VHPzO+W07OhDZDhcotAbgIccBiX/k
q180sN6amzm69/lpYJB27+tq8bazHICPNsnL2x2adkqGktuTxALtLG1qpb4lQdxn
n1UL2UmfFD3z8rTe/TRc3NCxYtq/XF28cwAybeBX0/MbnxUTag3sAYmi+6fB0MEn
K5k76XsC1F7lHUrerByRdJ48qtPzcWVGWurXHbkNDtmKZMZrLRSt8cj120A65OO+
v9kZ3QNOlldIqV2rZTYwM1BpXE6Fv8kwgIueTuu0N8kccczaQv14Z3mwPRGL/BgT
omue24+4yGcislTJJxNshL+gdUYcUg6uqVjthoS2GHKLfmhxv0VUY1EL3Bxy2pJP
3AlmJiW2gAwkE4QPQ4vCmHBOK52Trx2n+4EGHt53aVL4wjK0CcfnYICOgSo/KMYP
Kb9SU6QQefv7Ok18LQeVUn8nJldUBPYizwnMmym0zAOsLB8j34bkDS3gy4I4L7NG
qz0M4QLNVsev0vfPxGJjF+u1o9a0rYq7R/uzXXx/+Rfjxk2T3IxzDncb7coSqIso
huLPuz6yjHDcD9hgnlKLZ6VBLPVcJVK933B3z4QOE8ZZXpD8FjOuhUAXH4Uzu1oC
2mGmXdM9oPOjj3WCsb56IxH07oQcwN/ZHkC9rKgvSS82esWFuykTky0+9AAPYyhe
KuMDxkRWtHpGt12EUY0cYg9dgkG25VwLGNF9ild/l5ZAQoIRxsMxMRlKMzjvGItF
pMWpN8UHRFAu7kdPdOv7h3oNCoF3coXYrlaHm47FTST7F6ZgPXcBN9u9lLpQBgq1
5xh/+qnknGuWb3exzN0BRcN3HYnEsew03+m6fncWbFlwHxKcz1fwJQUINQY63TiF
oQAqlt2saI9Y6Gx6V6xe0Xu66G+AVjdwkwAuZCwcTx3bCMyE9XerDWvEqmRSaH42
eJvNgbp3RGMBqChSgS+OS3Z1QMUXAXZRR9D+ijWNrDb1a8UpoukDASbyNzvDnwGm
n4AjOpcG7DvMT8uyLaKQmgz0s6qhD1bsW2j1SdTu3UoZhih8Ut3uw8y/rUJ032u2
kqTp46iSMcOO54JXxJooyJs01JLL3wDNVMV2j74yTYawgZ37FMH8NnVMYKZK+a2y
RAj85ECI+tejF7t6RdaSHkzYRsZtmMCNrH9FTPbSTGSZzV8wXrt/4Ucf4lX/eCGX
50Tb1wQxLUa3ILXv1N8gxJlMK1TSqxeqYlsoTjZPPxAkHyL/Xm/wvDs/RktQ7zsa
ZS2BTnnr1wwvWVwn+xjCWra/zW1unYi7os9f9Dg0I8FobtNfmtL24IcRK9Ks54Wh
QPcBEab+VwZ7eZrK3CHy8SE45G1rfKZo63OgsLVIT7WY5GRuJ4aj2Iv2lZjOuQSC
Ng+3M6WoT0O6ksOszo7oxjxDdLGw2B9rAFpyLBlDr7O9wEwX0yQ88hFu8Rlm+vno
+oYBwQiTKMoU2+9nVVUDsRMrG9YdJqf/V0Vvimq5rwByulWLKwzg1hkbxZklWow4
lIIVy6VbyF9Hfx6490oXWngi6ws3DxRSk1nAKaUn1cdzpFAjJhmLvAqe3NglvwOE
tkVnd20s8SuJzJkPp0UJ+UGYrRzW1h/BNDYZUcZBuBQpEWsQHKTL4PIXkJ803WEI
MTC6OHdlChz2c+Vgt8sWJF2bmh4riZAu8fHe70qc5CzsYE31yJN91FzP7V6G97S/
QOF2ux830X3Y1pVc/tWgvqXM5JDGouGD6hQ0pL1n8JqUN1qqDEfigeBKuwR5TEd0
sTdTUUvEkUYpdW3EJ+tMnDx9mktEm8wTL6N+OMudO/yWWeWPKhI+aiEFt9lX4D43
mGKTfciDpRKEg8ys/WG7bIo5lwfHimx4wwXXE3BytmLGFqSXzeUIisytm2MvDZTZ
NawuUsVYIIuhqtx00szPBVCZitWKzPnSoRn1TKkXV7NfzPOCPrItS6Ayj8tB6oTu
otckcRPdv0oUc8lZDrhuzZr+3TEguRF8rKxTAa3t3oCcgtzwUAuwbK5ZBHiE4qdB
9TPTPkUAHfE16h4c6E6h/OELlEXEuxQlAUysCYMF83lLXueFGH2WM3SkzMJ2tScG
bpt0pjk1sJ8ZfxO9oqp5sqYH1Da6ZJLjT0U7mr9FdIhb2sYXVYcImjWiUR565IpP
eCP8O+5O+ZkziaJ74lY1S17THWLP261R2r8M+f3dO75x0jGfQBFmx0CIKWKXXUmB
Q7vPJA0Va4rORGr15jr88nOhoNzZ8KUBH0nxmjNYiLN6f8728d3dDiYY7+72G80O
LLDOI2bsLYMbmOZnF4W29DJvC3+OIx6LYMdkiuXpXIhDqAlQUFknKS2BQCtgK73b
cHvrg92/asgkdrRu3LlXU/C++7zPNX8znXXZJUktXNgAImQGw+GqHroJAMqsESCp
839s4zcKVGNMW7LnztxzzOf6XdyDsPf4kNQWvvsSGlhJy8gKR6aE5eC6kxieDFgA
ulcCCz6jHtJjIgneI3MYXL4OrcnCHLG1ImzqEbO46KEAGkAu/+VEODuKqKdIKUnY
DzqyB0/dL3uNOY9qnZUuuVPt2WVh2dbt5GDjlSrW9NhO79QVUGZeoRzDWQpqgTlW
l8u/DcylKaPftTYJjw3ngMTm3en/Oruy6xhHLD0LYk/3hBaEmy9/kYDy5nVBdR6D
w1T/nG96Is2ULocRhIkqDhEoQXI3iNmtuVAQIMnq03LwDZOEppOhg7o0k7MNQ4FE
0npHk2iEjP3evn82iSeJtMaC5JfA5uWf/VwcENzUGeeYCIlcCwoEgtGNurOi2Wi8
2uK+MGhewbYZfw6CfeYRj1qgnvlQX+Vx/4w5voQ6NSjYeg2Jiv2C8asPiQSX2cG3
JgyNq+a7CV6+GqY+Ct5/SEN5aJiyVDA4Dn3dYbq14cMlpfWaJ/JhT8Yp2P7U7ocb
5/NUpETM3cAoOp67hOCu3toR8fRg6AGyP8ixZACVmj/kkduMgbw8eGal8YnP7ru3
gQ9XytEpGoBu7EKEU9sdfLRcYr8rKbS820RGXXFcLMZF9AjQKqKA6aqGAyXiPSrq
4OXvXro5VPIfmvNgY7zV+H9KCqeSbnX0xMI/vy7n5GJU4q45F5AzKzHIyTaaFw+I
C0YSyaNTpAxpoWot0hZhpyYN5w/EqlEG0k4xzG98Ja1V2Z1zTETzJ3tSoY3Av1BV
ywvg+5r805S+WPoMp1vq1T7lrvw6fm1Rm/UrfHuyw1QDIABRczwmuULKFN77IieM
Kt2mGePDKPJR2qB+HbZodLmzJ3TJEF8hbcngqYHx47+aDyCXbS6UalqS9QuGKDRW
Rksw270JE340J//6+qBP/6X7i4W8oDNL7CIgQM6LszXKul3b2yj0EpUqXcYKPwgp
ew/RwCXnNcWBy+2ZL0E5VkASZ6+gv3ZJL9zoPyHI3UrVsa4j2eNF0LeWftNO8pBt
kPphNpVaixlKWjvw3/B8BwHyAcQ2WLtIrrFqNbgm9c6MiCJ/Ry5vVvi6DD26Ylzj
zu/0vWr/y0O+D/niAJv5qjV0bDUPmga1TEMVwck5rQVsRQpmLplWGAqwEWNdELKJ
78N0m5IyJyxD6PbJTWEJJs/dYKtTNOI5s5lS7bMa4z18reUE04UojE4/O432UOJq
qXRipetJ/dllIpj2UMdzUzzlkDLZ5OkvSPcVdJi7K2U6HbrxhjmlUeBSp24fuF6G
gNe6fXkD7z/lhevNvR5hOYjAvIR/N4IqsBrhBr/DJT8YC0iKgq+KyM3VG1LGptQa
PVraasAjyeq4l8u2whg93K80DS4ZHLXoE0oAO8ZZXJItLodEXASLVX6yok++MrQ5
8YH+BmENvLNZ7rlivZZ+viHg6h9UTwN/Uw4lyVzEBVAbJGJIWEDR40219d7zKSI1
/+rNzHox3YYvHpfAQfLlYXZCFgy7T0rFYzlZpZgHtUVme498kOjwjzj9k8U8pppD
3zK8re0zjN7DYwRe5eOheMIuR8DrSc1EjKwGQD6su/uHkGzm1ok8Da2FmDlD/Kn4
lLJgYkl9vF75uJr7XnImoYgaUldGdZLCq7w1gZOVVyYnXseq6uWAHw5jSeHADRjg
ZRKliDfg6H5fN10Zd40BVYgZ02HmurGSIBc3XvkDTDQ+238V7KFRPwIgn4b58IA/
iPVo6HU2aZgcAzCH8mkpujSsxmcOasb0SrvDk2OjtX8j6TeT1e+vOuGgtfk9oeh4
4r+PZxrgI3muyqock+swzQvw9DbUlYcFefyXnZE7KCv64roILTqizTNC7bMlsLJA
Qq3/WEzkiykA9DGuec6QMdLzJqhPqBTOvjaXqEPYGZGjSFWGmmv2Y3Z38Qf46ygy
DJXUZfPezBZxUv41kB7grgCNHPRn4KTYQNw5djyoU8xXX3fo7zLwpwS2zBsEtFv/
bvyMux9+iFOaiEXx3dpghaP/CpY+jHFgQWmvLh59EoQFpU3HrEJnIumjnp8T3osa
xSVo06sXaG6FYLAT2zeAuy/EGcM4mlLIXlZnHhpVXSOz+odrBZrpSWG7X5sjBKoH
trFBKaRmADojVHS9a6rMHeCYW5uLizrqBRNh+1fU5bhU5GiarS0VGJLNG/8dd4bp
dqKh7wEoB/Fv9ddqKqL4f6zLso5GuIZJS6zg7dlB1XzrfaK+Ht8Qe4spwwcRs5BW
Wd3nr7MXN4N4UPMN0M8W32VzYpvxZ82pG3WhdLk5t4iRBOqciX1AvZp1iO95eMYQ
9luvhLzj+qYM4yMbqIerAS7bAe2KcC/xWHPi5B9hWoRnREEFn3HIuAWkMDQhtPj6
iiyI9Qvj4otRfX+XCA+S8qYVXLB9kg9CUVnQ5SQycZDpkvypK5acu5AuB572Smn7
bcM3XtDUZvVTCLaCvZkuINPdbfatD9cfj+ld3IEEy6K6KYavJNgdwixGTSd7V9WB
nyQtYfnNCsJuLx2E8R+9l/4uTQ90yCAzf08cGD5HMjs18j69N55UIimBj8jAr25E
t2esHCzu0rvJcJDQE/oiupRwkwFgB/7n625Z9xaZcYDNORDf7j4xleL+Z08z+Lbv
CklPQpJQB926t8g3IrGFAC7qVrM4yvoWcNF10OUFkmWrgEf5d31uUxqsCQV6zrC0
mBjkM6d9zSELiB07sVPhRf2/bzWBhi84sonc2VHkonjQBjb6tZhqsxUMIau3Knek
2JhKrN2Pn9kevQTmhCu3tc+Y4qyknVCeguUNmDXFQI7mG4zch6WzIsUCx45n1Z7S
fAw9QGlVITVKv4eGqx5s/n+/gOyuHRso9ah1/C/WhbNFmhTYBRMwnfm4KLHgiw7n
HWz3YSMyiDwBzolsad0cNaYHITZnG39OzrXDRrYoAnIGoYbi1uEHmBAjnN4PC90h
lkZfdBgmPWkDrjZjQswXNVexSeM4D8sHC/QmIOQ8SKxYuR0yFCo2tYiwqcRuSDz2
hSxkaaR3opTpIaSmu0vFfc1lo+fMZSQGIYtEVqLIzthcb4Sygw9gyEurgkIyFArn
SdfNsemChFoPlLtLbhifp0ruBIIL6X0+ksAcLpT0p2c+arwAuFzonSY4lDCYQoAD
IqUGuIifqz5hJJ2h/+BdGMqF68158R7cEPxkUIhh1d3vdf1JioS7bJMTrMV+Lxgf
qQz4e5hTY+/4kNurHUB+7VQMzrwDDbFV3g641KnCUsAJUaQLwDU15ZBPzPF6ZGoZ
Uz3Z8mDYVAjOKOIL5MOkRZeHR3/Zf72f3C3gUPJMce4BfHr1dyyHhNJdodZbrw7f
WeT3YW9Tc8kv/K7kjXvnnphP+mw3E9GwMHSsVgg7oPA78rroqQ+rhNTNzc1ZFAf5
OZWwHTdvNwopfSsqr2ZaZyJvZ/dlQ2j8c0Kk45/aC3e5rXNhB6FD+LgrJs2Pmb6d
cb9NFjJVzWiygIyLdhGkvs+LxJ55BT5qBTRWyeYSM4ROVae1OCyzJx095TumsDbp
p98w0+3VnyjnOkPe8nj5JNqfM1zXRJzyN0We/eJ1Cg076mExr+g3kQ6oyfvaNpqa
Puo3zfDsK1A7v9YNIKCBvM6OjkOTjWjroRGYQV/Gijmm57eTAeOyCOccJr/F5T7l
d4eDywuPkl1k/4L4R+usxMCvFJDQtyWPTuqqCNT5E2BCzmoI2Tu/nVMRoJ0ctV02
ABjahwU6HFsYqYrnpkqH8Os1D9SEHLv2n3qDhX04934nxu6WPbkBP9NZTMjMIMPn
jcI0moFrQyF5LKEy+rjKDnrGMPAcNlSu4yt5WyfLhKIwquTgJc+gd/i335Lm61Dk
OaHUx6dg0/0m8hOEQiVXWJynPcJKovVy1ON053pNsxbfSsyXmMchTqrtNo80udgJ
CWUa91mwKlf4qRCPAQg76sLFKp3o8t9phN9d5lz3AeTCUKqj8pZ9EgmQSV2sfffx
qX+rACVcpQCRsPPLi/173APA1Sh43qRyXVQDFN7wh6eVmy/ST88GtmKc9bg9aIML
h3WxcK+2pRPnWZ+FPP0I0/eLgGZfgW7CSPJnuP4HQP+Rv/ygJhrOtwo8mC4Jz8mL
tFtXWBRGo9ad9w1oHKkhdjwBvSXSUrxtS59rKnWwElxkZqI31u31auVBELD9l/u4
yN2B4fUKPzl+bteCQD+wAprQOodLk+oiLti/0RBc9Qruc8uCZZsQlX4gYFPb+g6W
thlMOARfFIfPp1garvHWhxfi4XprXul8B7X7VvZSHlUFAN3cKonZsOvgwGvgZefz
SNmHTTiZtXFsCfcVA8Wro/EBwarStQUwE4erRTQ7JhbJkVUKv3C5hy9Z10JoL4Hb
ax0RSO+iRwsFlbd4fFUGyhWJKn7MBWHP9MZ9LkxIbYgZRJMHYCB3KbgQ+0eVOzGm
wg7nOlCeDXHtQ11eDaCEgWOa3khpgeStxV6t5P/0QBaCaOweX5qf5oVTy+JHk0pK
D8eCRXpVLuLVe9tjDOOA9YwmNU/rsal/+H9rGNpIqFnHJ39gWurEaqbHSv9uPqMY
n0/SNtvDA7SU9gCYgAIw7J/yxG8NT+4v/7+Ldvs0O9Nlxe0IMu6LI7d3i1hn1msk
trA0WHawGTsEFphTyBi7bigj4v7Pi0osK8GixhDr3RXqiJFqNJHXK54oHlD/1MeL
LX9+tU4rLzmkDTx8sipDrW36FZZ/a5jscQeoTkpimFaMAFoEXXzJC8JXY5DNfYcb
LH1t91pHSpzASO86m25gSHwQDU3Z4n4grkC510ooWqIZy99RkmlXFPRsdryuCAkW
Ylb3EdHQpsRMzeDu2GCFpHxjGVUUZeWSBncXxOn5vu8mqD0ZbfOGFANaQGV/cnkx
71R5L438XBV6r+tN1lhdNtdsiIstz8rj92+gCOyIWr8tynCgQ3J9COD9Rr8ZjPWp
HBAs+EfLOncjbPlg5ljlXcf/LDu/RK3z0AlVGe7GZ9iEQUTiLjtgvQuQ5JdxhRIH
pa8P74jxByihFhohvkUU3xuZZN4btZraQk6TGhqItbL+qHMaBaCRhc2wlIwL65h6
+8DeV/yb6uQ48is4ezAW5qjRG4X/wVQRTuSb4COtBjWv+jVxe1s6SaNELG/LqUnw
qiKuoBByEZBEnoP3/mb1gZhsDyWTOWLAYvS9j7ZPcrjSwoW/PKRk2GkkeLpdcX7u
MzwTPTQTjDb6ei977Xs33YIcMtOYaFS1NBBM+cLlSCaT1uXb0C99IOasijD6Uppa
GE/ue25fnThzAsTJTcQNpyPra5GdHxuVBFb21+JwIHuPFhzQj+m+IyESwrdPM/eF
5Zolj1aoe1buVKsqp3SewC6q04PFHOm0KFsDA/VYprjpF1r180DQFM0d6wb+ojFJ
Xe8tcEE2aXofi7+zNXnzCDgLwuAjkLiWXmBRmudqIG+45gDp3SB+s8cMkvoDuDnv
U/7ZkLia/KbSkz6hR5lfbIrPHL7xlIgJ1p5CLxS3evLXHVUDMN2KHWrEIFCc6eb5
Ox7a5uXgEhRqv0U9en/rhLNzyA0BlTV5oXQuf7hEDn/XXBdeZkHL1U12/m0smwVC
Jo/NJtOp7e+mlEhr2uGg0R6jJi8BriUWBu4Tw9ZC9ltxKrEbWqnjmZIVE4sUL57U
0vruUxYU+9oNfYh+oRItrsH/vKZN2+vR9O+wOq/4A5igrTr5D+QSwsFtiVhbgled
l2UH3mOd20c5tqrM93pji8JPeOsWGplOIqAPGQSr6mHTjtWcvCn0eJSccCBKWg/g
U1iLIB4RoWyqXbyLWWtnjcOL3TCDPJNENrJY1L+ZHnvgRaoihEVlpx+znbp+mUS3
RffZf6EdZSCySkbunn7XIF9XqxrN7F863g9w0mSEFwMEA08HVRs0d/emWZ2zoB+k
wrqIoZLR2Vg4m3TASfzHkEjstC6ho7WWAN6rkgtdFM34rNmGZaYMhK4rV7rRlLzm
UtPz2AsgLPs1pyufjs8coKQOIAWqNWJL/skiJgoFr0XyM45l6ba8cF3zQ1FJv1CA
NfjkN3Dea42Fg2XUODKayeAjNJx2NIW3TTLN2tkMExJHZTe5HN7b4Gm0BKkGJK1S
aVUBZo5LeBGAiF1S38Qebn7d7ONiSQtDJ37Ilq4ZYV11mrtP5lLc9ESMnY97s6dk
JbFbXjT1eMx+xrYGf0dHuJm9vwFd15nCctEZCv9oztLv1Qibz+SLx82PcsjSZhL4
FxUrvMmedGm5yyIml44U+9pl/iwR//XLiGDdARSwcC+sgvj8z54ITlHs02ISNAA4
6gXu6y2KNq76lihAvqpfx3KSJfYqdhPzAESeVTATKLMIDhglX+NTYmbPsoHVTjg1
c768hZMLAjxDRAy/tPvykwIPcL3EHTgLZsqXcydh+6ZfpSn6ul5I7GPXhujw9wIP
PQDVM15chaZ1RciSIBtjEoHuIv/pMV8mJ5yv/RX2AO1DufT78p6vZivoxKM3ikfO
SpD9LGiji6kwYcsg9H1B+584ElPLYcHwhVKZDz0PelNOUPKmKfcQLXVmb4Uf8EwV
aADnkBbggQdl2XBYLASy6GXwjGXJ7P5FPJI+DGLpSn0YUeTLK7WgUznBvlxVDJrY
7MYXfnw9pPyqnE8NFtb6ZtbVvDkAvjAsWZZo3/h25SyDSwdtc9WiLL16RW/EP8jC
gSaRsbwIa+LkpKhJ6kxv/bhXIYY/jEsDcD2ULYmx98dBS8MzmloK76Oq+r7p5B4Z
Ruo2b8zZ/V5LjC+VQ66WCS0l0Oi5mBFgjiDZJonFZfHd8q9ZZac6tH/xSWERAuYN
1+owRrhHcaecRg6seeH4oTPqZPwm72QKduVLAwHxD94Y/coqxAiFvZcydx+gHUdd
4xLDATWf4TeD0lo6mskA7cby8sKkFMVJrhcYmr9SyVdq8AzTEDssePQvG3MVwgIR
EI1U2NwZj2rfP9e6XcQpWuyAgb2pFnrPez4g+9nuaoTqdabL20tczAAJnd7Uir0X
rPT09efbXE4QdlqExPX0ht9U8hlPsewq8xfA8h7zKmfxqHO5bCr0pZBWOgtlwnmc
vwaq1t92kYmX4eY8Da9ZA0WGB+yB6YE7HlWVyDvgrGrCqaS3OIMDOXyph5DX6r38
5S8vPuw0yPRhS9GAQJQiihKW0gYOlLFgrp88hx6hAj4VmeUWF3Ohw/4EFkNSFZ1/
UuSrRq+vM9Zlvk7GHg3f57f14ETEpLM3THYxtY+KjB5CPIXO+1tYMgH9ruu5WvGr
CFesYO259UB2WaY31h1bMl8YobVId9hMgS+mitg+bDZ5y0o55sZLDl+1AcyU/fuz
fw1sKDCsA8k7FDYQkbmsUbPjc/z3W54AanHtcL/rkWU9JKA+lCT98dWvLqWyNSdE
M7tWQHTK8XjjXJ30Oaw90smb+1GOzUH+V/VaU7YQ7I2yZPt8p9CDfMND53jJ4UNR
UdFWexPW/fuzT0gPmg5bTsxHvhfRsRqN8JNpWDdvo4sllgAlhAtsTT7YJExpMOjd
63fl/g+lRrfC8fAcD9XKsle8hA1cV+qkWbIzARdkdFW8rfx/Ei+sR0cl67QuZDx0
M4U2kQ/pAATYwrj9yCBjjaI1j3a5GJMZ1OMiPMTNeoG1VgID/QF4tpbQLjQWXRrj
izgU/7ixofvNnOYgFehwnayVL8+0oWouCoQj803McqYHpCMAUV463UtArdu0CDDU
2A0Oq8u4/GrUq4HO3P+mj4H5kYVDM9vIK3of6Wezknyp/YOyIRgvXB5X7nj/LAv1
R1/Nk4OAWCLkE/0jPTKJtB9dcdEsOoEPrQWDN6A7uSj871l5w315YTITqbNcSsx/
Ij29aMk5YJPeFP+XBcN2Cuj6h5a3sHW8t1Hubx5CbQHLlu2qBqIw/TgpXJPZpXK1
7SLMwtCFGHXGSgp72/fiXO5uqQM4UoZEnepF57PXwt9fYTBEmsO+J1Ps88i0AOtq
dxqLKJ97AGpjqomib2Ad3J8WeU/ER2hzn7y3ZlCEv7XTZcHParIrSj1FNUwsxB8m
xxLJIu2+9aLQy/3QAJ5sTJvmMDXs54sjrVqEhwjpcPMoyV2ZgR3qGdNZU11YcV5H
lZEWZuXhN9n96bFMtDs08td5RzHOfgM0Hl+gP5qgtkclpeaVKldhl5nZ5b7pQwyd
B+ZVhBdQYtSLRzK2tLB2xqLggGO2iYzAjwRObv268rrkJlVN/T29XDakUAfhLpyD
T9J4FDI4QO1IQMbmheFHfXVKG8sGW/qJ7uioYOMcW38gEjvNXxTEX1fwTQXDVxhb
VYe0LzGKSDsn9o2X9ycKKDKvkY0nuwDkXy4OonOQ7kKeDId7LX0ucQF54rEpfJQy
1XnocndeXlhYAGgX6H9ZCiPVhLuSBGXVVu8zhE68svb+VveX/QtlLE8QatlEtgKg
PX7sN60aj89LQlkHkKRWCClg7+phwENDi0wREB5S0e479VoKUFBu+xK8UGPMEt59
zNtxEnM6ogWaSwNX5JfgTDUMkUKS1pN4DSxTACkW/dtAomLuIai9kQu1UsJTCG04
wttHCteh/KEa3hY15bWMKbErkVI/OVYOcAZbI5dWNZBCVQCEiRpCRGyhBKNmxzFB
/5lpeDNtI2IMOyPjYkKV6lelUdUQXTSYkaFvfEroYIMudPFj+2nmtkkqik8IZvXZ
o9mWED7easN7tYm5xCTfZvQ2W5XZbvs0saktAZPxVnCsXNTgX6f5XjENPx4pNNWJ
KRe8S4ltG0y19UV/kcz2Zr8lxiQMJcW/XbwOSR+m/qQ8a2idknoANmd/IxqEwAHb
RLFGSpvWlxjY5t8ktjTYNypgC/zKgwmWmSvX9n1jxbyevsFFhl8vAgjryyDMZXOk
Tn3Vfu7ka4ihY1xr7rcSqDhZIi9J4VnPgA6xwzc33bliPqN17Ma9uLlUEqNUf0ui
K0XL5S3Ss+Urk/jmNhP02Mg/W5N+F2CcnmkTILpUYGt8CE2V3vddYqkJBQVGa2WU
/B/qD6/n+OQO2R34hOsy6UotSMtek9CUXfW3gfPNU4N9L2M3eYlrvxnCjorslueD
hcuJJah2LApFla2I+f92QkC4YlpZPdXuTVS5HKYPNlwEdC5KJrgvJ4V5WGejXAUW
arE17mYYlGDDpNyXGuM33sotr98tZOBWCVbQuPtSMwqm7hpaEoKR9O0Zsmqak5yP
SZ5P8F7iP1H2d5G9qbo0QZS6bN1kW13dnjORWHjtDlduCTYQ9qoxalPZ/HiFGQno
U5Y/wdW1BuCTDv6AnuqlMx2qN44pnYnJ1/d5LqXTiUdgMqSZUat/tZ98cAwC4ka+
lxtjg9q1lfMRXuZPQ0Q9YViTO5vUwlx4PL4zA9SVcxrluZOY98L1oNaweRZnX6bV
+N3X1tBSB8+fBMEolYe0g9qd+mq1CvJ5aOEeuUzfa/GmpQIweQkOMPS10ZJkqxcE
GKrmmAKoz+jHhP7s6MzLUSDBHHfjv01Nv1GfxqFa8iHQuMUO5odV/oAL8RCbXK1t
Y0YyRdrgk3IwenKHffIVdBiu/JTsekQZiqq0uHLIJf/2eqtZA0Iyvzw/8CJwM05F
i0lvN9k/7h2xmyexXWtWwoHOIm3PxPTh6LcbfLvJNhEvWM6jthewMacxzhXtuwwU
cLtQCVMMZ2Ddkn3YcxlQrR86cHwQL5gtz6B3q/fXNl2My+Q4FvhlHp00jLVE2GDF
79U9wkjN1lt4h2V38i8n+pw+rvwPmyStSKXQJE1RzJmY+5r8iu27nIuESeF0Wzp5
5HIJ703qeMqxQUIbYb+9f0gTEh+arupAshrZUitdWq+G2Jv3wrEVkKVZOaY768bf
B7sVhFUCSsnx7XdEVDwWh2dPXSdl4cCOl1UmlBaoI4v8FQChabYw/KkeHPyI6Urp
b0JVkWGLLFDaip/woLdLsLSAm8Wzp8OFLj4/db6kx5VkcCDyiofz+Yi/8FGc+S6u
u3EYE8zylrbjsSgPwjJM0ZlsOdvFimQF4cVTV0Pc6VpheNN/qc5fmk/OSFnviWG8
1FtXH6C7OS70eyTjEHqYE7VtrBF2WSvD4EgDdioM5+aj7f79C/rfGf7xwIEkDnhz
IX0NhlFgkKCJSgj306Iz5fjzXFmShyO7IqErCoL58ifoUeqXVtS573oh0QvBSIsW
Zr6nRm4mNvAjiyx9d2HcZZbHMqVJ/FVhfoczvPG57wQJ+0ziuU48FYbwQFqLOQsS
zvB6bpLC6QwWsawXVsCLT6B2QMREYWU9pjcSe585GNXzVcWnKq6jUyKVB79nEiqo
2C60ARdC1QopewwwIxHg9/h/SSrxrbsDkc6RSBIKeLSJv+AWkw9JVDtl6Ma4Idew
/FMwm1SC4zfslQldAlTn8uwvQhf/utbt81eZzHiCMD4ucBo5/ezRguTvEUQzm2uC
9Bs5t50pQk/CLtX+IwxW1cO4DDes8vmC7K6zUgYRPWwt2J4hv4V+ipcYw/tVAP/m
CeK+5PLAtSPPC0pFT2ZYGv7NxA4ADFAIt3e+CtUshPeXJgCoICgAe0w17udSh58T
y68XEwMhkMbkaCrBHrbMDmOOXm8Da0z0kzMVwmJrmq2p4Q3w4jl+LMNbXKHqXFpc
EgDe2VZTUKbYBtHEXjW+Miou2p75j+3ARHW5mgaODYNEqn48ha0pDnx3pb4g+uXf
tC97mAbqc87Zmx0O7LF3VGFHKtt3CLzgbhe5kDUc3cR8MeXtEQP1Hh8ii67P2eEQ
NGp9UzeEy9UDPTuZAP1gpEYcTwepQ1i56QFLAPDJwqEuw1eZhuvWyKoazg5Zrw/G
NDo4mFGUIuHWVzlnzUpJOMIHwX7cIY8BMeXHZQrfggjQJyAkIk9Q/T8DBnZPCmeP
V+r7lkWl06ARtBEg6h2Ay5GZ07m4ExnYZ4zEWhR+Pv8GI1spnve4EqKYaMFGfpSu
abOzhb90zAs52apIcdwvVVgh3GgfbhOy9u0eMshfItOWX/2plcWhPhoci4XXpliJ
j/gZ5y6KkEG6FaRW8cmFI0KQYvYJbLbJ3ayt2uHBpw4KaO83qUhbgb6gcjbE2ZHN
EKBFNfs/L12T6ei5x7Va8TcG2KH31XiVoYINtL+KnIIoTc7BkQRc2NvCvHP3cyOs
AbFE+TznQOmW3vQNI//nvV7xCUCogbCuvdi/12N2EZ8JRd0Vrru/fzeFfnt5rT7+
6DiFBYbl0lcaRXDkCZ35FDneQuacOEWwz2P8weEyo70H/iRglQm9btixpKuEedrL
c0wLdoOuL9h0ssNYfwHpaz4eE6GMlAAc/AKYkmJ7VSySSliq8E++IKKFr09ZIoiN
ZXKWlCoPGJYzOCyX5+hy61I8DgCAURAwe+OvFcJ7uwzV0v8GoyqLRqi1ArlYvSWb
tNZiKmpdp9p5dW2rwlB9O5uZ5JFIue9NHhF2wRPSAPChgFXUYkI2WLSWNnXojolO
1rNBTAH5E1kzigTD8RH5CH/lWMukPCUcDRsIfDGJtPzJ9/6SM5BQZZZmDJS+J6Lp
ShVWPYV1T7wM5DBnp5p+nJazmZ20Ig4JjNKN/qkbn7reJf6b7Zb+zT4ghJo9Iygp
aW/w9+C0rbu4bLZYEGt31zfgRWqed5sNLcqyZk/Pp7tWjnCdCX7/nowe2/6NGL7l
AYb3tzarUG3eG3pgS7yEkZDCAOj26TrQU3Ky8Q77OQ4rQIZDbnmC1Kt9L7TX1Rpd
H8a82SWJgK+vG3Kw1X11znxpPwizVJ/2jqEVvNz4grbgSyJlByain2KuuCi81o7d
/ePhPtaGYYWYV7kwnEf9oFf2NKTg4ldPiW4yDlst73QR7GNRSOCPuvZY4fgV0nsZ
ebuxQFrvsycaV06Z/ZDQghO8KhZqjVI96xuXKxotrS4QxThdx1nkBrMux0C7KBL4
0zUNDVqbYFABMHgEp40bPY7sOspAuBvte6qecSsHH8p9JnzPJe0HcsPwvSSFmgj5
L2GK9dmFb9hQw+/+GKZbIsmfiPzAH3eTPmyQoGZaaMH5dc6lvI+NgqPItZku3vrM
cCLpOMD2gpcbXkEu20NQm8IZTWpqFW/WqnY3qZig3gHvVGgn9Ffm2ks0qSQHAXSa
ULge+BeW8IzHyKxAL+W+Y3JyDt4+OxfZ3Xc6jzNu3GQ5O1UF7VUNN1DiO9wFI+Ex
Z9LKTGDzeJv/EC7wqPHciH8Tl3IJ+foZLeEzwPzh5j6XAzYps7ihQaeIafC2OlIl
M4mwNeaCPPyc720sq8a/J/Nl1syUEc0yu9IaHvRF1dXqqS5kNRIHYPHxy6fkXKK+
s9uAJlYJ7vJS7V0hMuiOwnKd46BXQX2IorjIlTl+DUML9LgpDnUuAX6cLCvoEJTs
3BQRkvZlmqm3doZb3YGvKIikJKYLCq8yGcvM+U+bBfhMxT/xWMjPE27CDhLO1QD6
qOZyneoxIgJVoUjWqNz0ZSTVQUsp6DSvO/zmQK9jdfsmrhOrAUfMWuq17RNrSLks
8oklclZTqUsmzU94FeRhCrkBtQ97rhSaeoPjpUWd6/DZF6kMsuHpumm/e1dn+Ivn
4ULyyhAZixYkY/dIapJrC0wkCieDwKUkwLEK9mUAaJUgOW/GN3E72CDnGhTCj7T8
oHAbuIVx2JeRtMkPwUo7DWIFe5YdNjx62QsJKFjV7z0nLC0Utmo3PoBdIQkcrqdT
EEm/pUUwFnLeQ0m5k8YSxTV6ANQCN8LxOTjqRUK5f9Nsr/KtZgvkNt4DwX5IYW+J
yZgghZ/xukkEjoio3ygodp6KTievoGbB+3cCqZzyC7rxJn19WMyGnz8eXKVX32MZ
iEZTnT7uXpCpXHuvqCoqalwLTcM9prSd6TNneJm6iH9Fcl5w3locguwLMcTjfCRw
toIpPKE/WWBPS8UQLQTF6tSNn9UOfd/XH3+HQ5kOdmD39fX0LSTtkBjREz35IeF4
evSXcAmfyRbY5UQVjEVVdNgGix0y/OVtIlPwwmQrpBtGoIQE1hd/2HmPvHKRoPPE
O/h/DrP4b39Pss2d4/0mRx9m2uJL3DtD3+T6u9tXD12+Oaty4tZPUFyIY8wxaV/f
aFXqZKY/YmwmOOnKEkAJcgjEzpOhg08TMNJ4+xuwYFugQag0ai+wEAdlGvGt7Qst
8FAfyHkigPiskjwlKywboNt8a2FMRFFvSZrhB34OZ0RmrADcWvXbjfaE7pijTJqI
S9Se+fvVK1MHmEM74ZACb1wVHtFjy51tDqOBlFwBi3m5f/oEKH5NmkJuH4T7FhAA
pD3Rt266sckQ6EZ5K8Cjuq/vHHgLmIrOyeomtyQRWK6vgUiUmm067l2zi1avtVCX
W2I8DspM2IHiDl2w7rfEVWhLr+ea72czg9YjDWCA+7azl2nqsjKlP/WrCIrKYa2B
h523KJRRezSYjbP4bgFJ71duRm4hqVVkc/gcaNnZquCGCCmibfBQOcR6ksK9T3dj
wYGK3LTUU74bfDEG+AJsvjCgxfRXBLjNP+VfdkPR7XGbjBxVP541hdT1GUtypRho
+4JyAeWINB56L1TVPcrR5iKhg6zQSxeaRJNy0KRAF76hO2PRvbKASnZ27wCiVysq
TXZ3QNvYtf2kKACTR0zT5fApgV6+TSXTLXvguPm8pt5kKWjB6ePpwz3TCuh37d1+
NVWWGickl416fhRkMw6iPy20H2TswkTzoKxPikq3vC1Mo3EikPkVQK0zAVqRgrJS
lYpt2SUysotB5h0Crnt1zYq3rYYeeFvoK1vhlHEwdDxpUwlYNVwTjdUiiY1NrZui
IpA/5iOAw0qNvQay+jtDZZNeDx3GVC7CAP0XF1tYGLiVmr5SxjXMUmHxOPa0tSMY
IWp5zofwiwBclbsWy6a+xh4jeE8FyGUhydcmClknpK06mAmknJIvk+eItNcYXDoK
1eQqyzj5hEFpXClSJAeZSUhSn8ZKPSYwzGo5Jml3EuHUJcIbbRPWbDwDki5uZWdK
f0BfHTEcv2fH/k2JyN5pDzDRno+yr07k2+hd1ECpaFuEfwc7rW9nfN/DfBuE0hox
Ofn+1frq+wmehvsZMvpm7T4RRWaJ7LHBOflX4QL4nzjoVsVKXOkVdk0uky/5ntS1
ICzvsRKJ0AVHxxNNvDY+j8ah7BbrKX+HNny4NEZWbFkxK0Wt7YCk3xGEM6nWSP1/
0Osqd3fZ4x/KlLlJW0gST34xHxHsUpVOpBLiivzvclsgsvF2l9iqcVxFPou+1LJv
2LgaPsZ5OMZ/Dm/ZRzdxjQg45wOSn1bm6lTx9o7Y/vVIU68q/Md8o71giDTzE3Zo
Z3oklQoHY3p63kdg9Y+rFJTGcflOo50G1LSF2QaTaUyivM6mRwXbD9Du9JkPZNtt
4KnjyiJUvh8hiw4viI+TjcN1mrT/csYdYQxIROlzVI1sih1q7kGji1YbcPyBgcBn
d8cQMHREY27yqo/OInP5KnLa5jH8P9hwCX+gLaENdkP+w+YtEKBvBltTYVHzFf+N
EKTLRBR596XKrHojdutSc2h9EOF7ZoBeOgws7sEigf7chWf+IaKUNDfzCjrx5cL/
Ow+ZvhIm1kq17X/8vQaMyBrW/KtumwKHhJ+SMYKdstdBiyTmZZu+rFdWsnbgGHjt
o2f1hUttfWvO32tWpYLH+FSlvoEOVNNVT3mzBoBY9ucwAhoBiYoHQKtz/OAEsNDo
PyZt784v7D7BOvkfHylgKqx0utItxsn6LFDCbAWN0AtCi2FnjpO5ft5qL8Nv9GQ1
fde0BGftZ5+GBasdan4ZtolrWbGGfbHtj9wUg04j2kSnmmvIBGIDXrKF89oqDkjw
QOdHhGmmz7Avliswn90BASdoEJd+ISkmdo5hx8UsAVnrl0w2I9Xjgm8W9HCTh3Vc
HqjwuoYiB8tNJPsLVGP1gb46ctcOYCDJY/aonaX+07+9P+RSCoOWsuGdH65UGYPs
up1ZMitQFxQVJVUsi/1tmOsxGoMpIFBx/njLtJR8YCg16dCSHP+DDnwp282QRaRF
U/PFvYzm+8d9aAqVyBdyvZmZIxdwc9J+w22Anct1b3rVW4b89/az0IjYFZ7yIFaq
8Ahe5xcvGh6+OwtqtO1CD4OHCf33/FiIX67twC0G6pSAhScUrIUiDtiOn/GeN/4r
DutWeb/h9C66NXRhFe2/6ir1pF0ZB/fFnfjzYHzX7/wXkAUZeH03m2iTv7UZ6aZk
hUgYXCSJavoVssWVeWDc60t1isfiSnOMWSWjaRZnmyGs8ueyDIOEnUCdG0tkP53W
KoWpe4l/y9bKfuUuXkUoflUx3aEodyULgGdGtJK+xDfxJ59i+YFyEy1UYn/K/JVZ
+P8X+RDrfvRjOOBmykqTPOU7uATI91CKwoQ1BbLd/MAP0pm3wjis88jv44iQwwW3
L8SJK+UXaej0uK6IAfFcUI7bOIiplB5LLDPWdSeG0b6gHAOqNdnxCyS94M+PKGPE
wwunxZ7KWaDTu+ePWzXIy+WLLZQ1YNkJ578cCT2bEJo6rRw8xWBkXcZOmDv1MghX
GRKUqujY3WqMTk2M0ITzabDaV++b9eH9u0s3OByBAtatRposZVW3Uh+ZsCGlU8Xx
sEG59JUQLnh5bGPymTPQGm6mCJ3pcShAwyyiWRjp19FiU7O3hTe/xM3Q4MVqwot/
ioEhYo9EdLS7onmzIYF3dWurnF8fAmrfSRyOcv6rmK004woqSWSuL7qQOl/AQoww
ei3R8K+AJBcDrFkdT4MDXpx+cTeZd4BImcLUJdmFF9YN3m69f6lQ9LVGbqxx4yO7
pWi4TgsGW0/5ED3hHfpPmk4TLwoCtXO5Wq79EX7zgzk44SxqPyIBCpWssExEhW7W
5kmke/cAW6ocfHpg/t039cL4DlLbZ6SuEwu8XvXnxTgRULHu7feawKB3CKbiJlpV
ZPoc160XP7dWkZAjd+Az4D0DVXpghF8aLGPZUphfBA7C5VeyPKGlS3DxmBSMn99d
Tfan0DKiSkvs8ZJJ4h6Ur2hfdDdegYfaJGHTyelwyF0dIIY4LxkRHIXqLgHvLq1P
ztd7iLrsswiggL2R8rThi6yM7Fm4lZUTi3c23w2WpY4WiraX7f3T4YHjpvbxZyUQ
VXkv5qrNovJGcjir1p2oOE6rjUkuQuQCQ9f2EPcL1YVeelXj7HZ23AzOt0dxTN91
VOQSjRLgoJyJmP1e5RJeeJUo+EpX2SOqEwQR5MvxgnKohOjJPM4PqEtrGF0ygRC9
jZCKNRx3nMa1D8g9VecLlvN5IWgiibW1Q4zgWmFYWAIOnWTYkzFZtIsJn1yTr2Gz
QME8nBOVS0evCEFX9XwvnLz+F0IQWqkR1BdMuLenumNlBeTQiJF+V9kJEmJkz1Ij
T2QXpJj2auxNsR7MaAE0eM7/KL7DmyXH81hPtBDyjsOba/CckbMNeH2O4J7BjxFK
hpvp/XYkSrh2qr3Q97FbpDjl8iroDKLE7V0SLB3s17lfki9YocWrVGF/Ga7YENHd
yjiRgjGzRJxcgiA3Xt9x+ag9l5PfjiY00ZVN7S6u47WgJedWCg78Zm19euVvvxPC
DZ5JbBwiJNvgEUGYLDRAIkwRbcvsS31X6MJLxmYo5eThhy7hQ/+/t+4rmNNYAoFs
vogUmbfJlR+0r8ghpAPnNcnz/ae8oHYTO1gmds+YtLCvXqFtGzhkdO9JSWddov91
kzPA1Lq4cTD7WAu4VmKtIyB8enoywUhYt0R48iQ399FdonqSVVo6oS0Hq1lD4lug
99/GKItPUg1t8knCKE4qDU7zc0ccvaYU3k4MxIblg8saing4C11WPzHueoUTVZZT
6bCDEVjv7D4yuJWk00HJ31S8UICoCsydYYeso39iOs5z+tjSnwO7C03+IkCEmygO
G0JTfBmJTk/tGjheec4puMnotn819O/KqXuI/WPwbzou6WhIhygZ5EOjGwHxnrHo
7E74W4AetgcHK8eZX/k1bSVq+qA5jW5sTDcbJJ5ajHVOb0utStSmCA1Ea1/nY+Ym
uGj45/xHwmK1NMSm7YY8ChCKV4Aby9p3jbjIJ38eGiij/SC0Z1H3gYI1FOy03VPF
PUYvC6/LViIgSow8jkXJTB0A6VSb25x6ei0ebTtZ/l8V8w5HopX/c/MMEifDsTcy
n57mZVdHRXHmHDyoo+kNT8wRKuqupzvqWMJZWULj16TEA64VZpXP/yC4a9+24Np/
Rl696ErHHK4gE4uwYiIkMjDF/dIMQVgmIaJ+1rV1J+3UBPD/Fdh927nlfjZ+CQ/W
ejL58zKM4OIwRgDNFQGYr1D6h1YYOGA4CXEfFQ+Rpx1dqnuFt/TGrtEKXiFem2N8
GhFuAqtc7YpKeYnK5r0fBWE42w2vUf8mYHbEpj8PsecfJSt/R0h/mQdc/Eulkg30
vm5ePqCdF5ra/qSCSNt0+CDGmZjqLPNLP63psVJyEwIE8pWW2uMhBg65uv7evHBA
xPLFLkqk4+RfyAxHhkEOzGzqZXWN5dT3h9ZtQTrrArcG9GQeTF1gVW6W7dYN4m6W
xlRpcbiyp6IVn/sYssUkaelbjeoL3y6Unp3E8Ji3LDFy+AUNGE0DtQl0hlM05OPg
P0gXJEs3Bb2ViNzitwbhFtibS2JDAgQbPMeyMQzH6ntJVccEsBzpym2tmPW++ahD
/TILGsVD/d7oYpInNrSJlP2FQmUxRDBKMt08tbGYSMRRZZ9zB01xNUYG5CnPm2U1
HCJLtrzR7+qMIzyhZHW1PLuusXMKdehISmG3NpVCICYAx4zx3J7W6V+F1NGsJVKP
bfTPkq+0Xt7+X1ugB3fkRyiUenxrURUfjs9VyUEVHAGL7wC63LeBrT313pQjodhU
FaifoXUHWM67Kfks3dKNE6tn9/cbvWwtdsSLP0M+wkn4Wq6KEdTBDC1FukYCANZ6
mhHGgeHT2T9nLtv05lK2EMTKDDEa4d1oN7aFQkfPKRd4SWQ0qiWN1QI4lLP/B13E
encfxEP4qys5jv36wR9vLPZwc0wY+eQch5OfATrkGKI9HL1dzkjJj9J88c/JrKBo
FP2kVlC7N3U+aT8pLsZVqW1ZEWmSEYEkLZI8Lc7PcL8r87zL8wDxGI8fTghCQFor
Jz1N6kDkr/tRLpW7CoqCBOnp1LWux2Eb3BI8ljG8XPGRoYKcovHDzXGABahf3bBW
HDFiFIy3U/hdspz5kK/wMcNbFvSLRuwHXOLWQcOzD8tbWoxcInrtJXsfRJ0OkdQo
Df+lS5JEqfEHqJz4J56v/N3RYreaMLcBU9VlmddHS4p5Yp4XbEZ0Gbu3Wq8vvLYw
YCy0ZeXVRLvAr6uyu/zFvRuFgrK/9VeYPAH2le3bbo6a9foLO81Cru7Ley8hS2KX
qPlvurO2eZ8m3lU/1QYU8mzL/qAIICTHV4cE2wjKKGzMjp9jco0FvH2AQ39bZ6EI
x1BY5V1d/9lUKlHxHkLHMbKp3OExrBNuRZRoJluOhLsAOJSdqC9e1WYZuaifQBIY
IWIFqHaYJ6+P9E8UtZeu/l3p2mo7RSQbQeUg3txlc3CylqYOj9Oa61xe8owXqW1t
3ap1k57AcpcapnfdmEK7nS2453RahomDfegeS3/mIcuC6s5b6TZsSvSP1a39JFYT
S8198Y8w582BJ9QN7cdZynL70XfASq5bi1rYQUWXSyhqDP3r27VwDfJXoRtB8v8D
N/f4o5I8izCIvSC7myag2mdi4PUNlOR7+hvtF/jvVlLymoC0Ed7o1Nlh+BMOGXCh
WEqsATulH88K5h5czahPwVHjexrON9T2tLoIcFQbJtpreWT+c+Un6WvBysw9JFys
ygE0yooGdZVg9WyqzXcz7WPQBdiXT9F5zsjG18fhiR3MnKWiYKWttobn7dbfbpKh
pdLezprwWR93zPia3MTpfX3HAQgg6SprbAWvpIhwmrOeikGiRibWUtDoYDSk7f7q
KEzv7fU1GcCy/EjMokH4rY0toXxU4aAzvU8cW6za/CMkkX5oSlJba2j78tmN1BFo
OQAhb0ngwQExX+Azwk6isbdxMTrzVVPFyXjtA+PiRlIRUVqU6Az5VXDQ41MDoV2+
0HVsEQ2I68j9oHVrcLHrdts7VQ+yeRWpuiXYsi8kBNLWg4P8beo0VZKelr2zSDDC
PsnHgKhdZCDcJpjItFhjpBQFEx3EVCcGwM75yNJtSdv/fFL23R9jfVh4OlESg7N8
6tD3AqDM6fCfc66Rozmqu1NKjW0NMp8TUxrTookbGJqLMew4kveRfdtK36siwxE9
hmdbStvqkPekbKi3cPNE3ka19RWM+yBebVMITICoWT0OnsGRJaGghsTWhEMYSWsu
zsjndyrbcnaLQy+xsm0qKpX0H6JUmrmN65MPjZdqYCVlS11uuAldGZKGl0jcerdP
iw2Bd8mGDSOsWTgd9+CsKr12V/3Acwzns0T/jnbL3vUot+UZeDGfhYtNiL0KbbXP
qmsjPF2POoLza6chqXeZ/1W97rue2AUb7QiKyP6lKvJ5asmXiOU9apySCRhIVU9l
5cc1s3CGZAp980VGp+XAm6QtDeFZAJlphKbwR3kJyzT7x5pJDsk9GFL2SrKAwsCj
jZjqldAswmoz+bR2xI3GWTP2oksD/nb4HT8KJErHSJ0eH6krUuPfct0G7kTOjrsq
ojxDhfelX9N51/tWExKvfvkji9gz0Q1rbV0KVeSeiwWzjwuw3+XCix3beDWThGR8
q5puaANPY+yjTkIWp9Z2dmdcd8Agrspj5ASn8fJtJXFbgYVrDdNB3MVLniRIDPWo
f/a9s+jNT/jaEWoEwkWTwbKDrAhp1XIFQidKAWpKN3Y4jJHXCTu6gg4rfACnSoVc
/mqVaZ2m3MYSkkitYMc9hdYX6GbjKrbV9O2mA9XaZgHMhR/1FqCwyUL1CbgIZGrT
YD8Nt5mqaT3bHBNQQ4a4LlX3iONJGdbDxVIHjnDxyrGzrUeLSB4RyQ5yhVB6G7a/
gNE0teOqenADgPoWFmYV2IIUxd9qTPXaVlvculrR/QnLkD7SHd5EJfeY0fnrvKKb
P62WBM9wymXo4CHuJC4Iq7Jk2OknNvouKp708acrkE4Qh584eHaqQPIUCUdKY+29
Dt9kYl1OAz3AjkCU3V1lV3QqCBJPHasuj0AL8f/NVsC88ChJ+OCN4PQyNNAJoHOu
MnhT2p0kUQcVRvaqYMLxW54KqmOL6fllLstjdSRiMKFLXp5haof4E6bOGVZmVDVD
8aNMv/Is2IkQmia+McRAIh57OhTVspFajYBdPqdJBQmcjGpYzO8U+w44ihh4utTj
SBmDBbMZLJo1LPVvFMGwiEJ95NVp9z6hN3vRaESNKG+oaDcks2M8A5ypaKMEOV3G
rREY2RlFmEfn7X52i0ZT4cXKw799rHObbR5Tcq2xfgEfKzhh5Eq37uF8/7Xo84rT
xGvQPqhHcrR1TdIYvPWiEcafk0IS07zuDLgwvrrmYRxj/nxB21aJAFKlN0fBzCtc
4ip1Nrkq6ew9JGB7uObRxskMqtnrnyAvC5MTkVgnGqw/QO5PQO+Yw3owPALaH0Au
GZP7zr6M+hS5NACffFL56fT9LhedysTnn0Mm5/KWd03T1h1LLbmAtMjqFB7nTj4S
AC84n02YL7s0qx2ulEpqZ1z10+Es0oJk+1rJ9tpdVc4IGuh2wml9lw2kQvtbIGil
JpX9tdR0zrynNIb0OnnLYdyLleRHZG8+wVTAM/Fjz5GLw3Ec/bqoaokP6MGzH1Ci
j219yzvynpTEnVEfmnXeCWuICaVUVRdg5s6HdKPw4QxXeQiMovPigGu0PWWtgaWw
aQDr3Frk0gadAIVjZhJQB5+IWV7SYVxyAWzf4a8kxlCkEu/egy1r4aHpcKleapBZ
skbjEm3gaitq5uOaMD0QA1fRpm32HUMf2zI7OrcEUEXCK5VneLGyev4p2vCGdI1z
shywKFmqVEORWoNGLW3x+NR4a5FOzqCU1pWETUcsUqWKc5XI8ZJJiRJZU2oN88p6
JJrRNEkXnknLgIZ2mEsJnp/VazyNZmN2QlxmsWuczPXv4JpT96K3Fez8jwcBQ0+U
/3dIJzjbnsUZqZjnkRjldK3/Z+gt/xFL1VKD4iGfmubqvxW2e0cj5hOeK9ceMH42
G/q+D04Uebmt7xWd80Pb15DRLIKHhl6jvRBYmBLo2Vj4GnL0DBbDqzgM/9R0sXN7
m2KqPAPd8uVfg8HEwi6RdQgLWbgFo+XyOVIh4Dw3wfO0f3ZvefYKtDIR1tV83jIX
Bmm0idWLKWR6tNRuN1ex7g8O7oO3e3GTjDkhnnq7Bhx2MNwBoJAoltR6NByhnUuf
JXejbx5G+kFtPXzn4uN89T2JyXgkg3ULWkkrb8tCr83+bZMmFbz/LkTCPWoDFl0l
x2dZLudi/LmlW19uRS2NAa3X4OTJ1Ec10VSC4S5MgktiC0U/eVDnzYEHNUO6ifQk
yoCn3AeEe4tMhHJoepMcwyNQbSTXvgdlRv63XI2g/oKCt5TNUBVPal8kZYpV71qY
cqZf3mpouEJlrfNLw//YkRwXx5LRHqo3HPY2oUkztTvumJdXcnPya/SALvJEXTIP
jx2Wx5JRSXg9NhqDUZljZWFqy3OddvxJPaa/WZTI/9sFXKp3sfvAYGUJ+ziHyF0v
W+/s/C8YQ7toLV8HhKoa7Zu0ZlHODDq+ejjab5W70ZZnFqn8497Npt1ktqzJbQ5D
sVQpuP8z+FhDhAhnqJlX3sA/edTosn0eANBlL678aj0x0K5CWwAtum2oXkmQNIQg
6IlJ6JT/xVRD9ZC7ApSXZEKyTj8MUBz9rYJMi6H/GfCC0iuDIi3iW+0opQv5IllJ
KjOijpQJQ5lebtLX1hE4mXmAlyF8yG69XsuKrhtEZ4N2bOJSZAmEh0XkTRSliuts
FxG7Owzd+NEViF04aB2O8dtgGkFd8VBAGk4n4gPgPJJ3jQW0yGx8m/aiULpEjThn
DWdrxrCnsO9WBo2mvKkwMPMhgL1XLUz5jaIHHbT829iiHmEUKng024/OEt5bZ+LF
7iQ33drDJqdGkBy6U6fbkSGX6nZgICXupqkPWxN29HQRvHAvhRXXM9sJP2pgMUkD
RK0obWXArr5sKpvTguu6bOeZy1XN4xbmk4crSqir6iwZkUCqf1rjQOumcpkJIf6E
oVLfQ6OGW8RiKI3QcSbWlYSIPMx8Ivw/jvukyfvJ4fvYtcGjuJwZGgbpIiyY/Y0G
/yeDCUPc9iidzt+VXBsDo3eJT41tZUij8WKbI9lmUhOp2FSfxN/kcs8SKx4cKL8p
2yRtuDMF1C9XuhyNNBtCdAAZGnkFL2uhq01CatKEzRZQRA+UwN7bw4+dGnNIxnGe
4r7+KyY9vsKGxi1lX3l5TP8N/9uWWqA7TonHXwEq3vSx4h2vbTA+hWSNy+o2D0Y8
OSMnihUlN0BPNWa//gITVGj9u/RRGSyVoHQH6ZuZfa3IS7kKTyVIa3sEEg5IXLDY
146pfbbBEUDsdeUh2z8A6pjh+ldM3QgxE7Z4XZQtPgHMLku1La1OHnKW+1fet7Pb
obcXoq3jxd+eHJlKfubECXT3lJjZPD6UN4HLfRfjBVafoLIGlKIpSRFkFCsMoK8o
Nb9LMN9N9DhNNzcpRZ1LldlkKLj2bzbkv2rPp4AoYdcPaxT11/8EVlNqYAx5EhPA
DZ8DHHFUkNTyayXOB0ibtAlgNlcNWMAfchlsTwXrQ3oxwWDz+sfbt4EKCcsFuI5b
CD+4WhELCRF0N3UD6K51GyazlcAgSe5BXzlJIDIXqUfL6sp0CQ6bnoPILa5niBJ3
9ALFSwnHjgNF0WuI/ljB1kFGHacmhUm8GM0hmRuzY9o41DqR2/o3ZFKTZQ8KXmlN
dQPPWz25f8wL+x0Ccm3JmWU3LeCKQphjDYIGrvSCgrloYL9DeM16Z5b2DbvdFcMW
p9QI4yILm2jklmpdRspWyr/iVoieNeeMtRxgWSffUBQcUl4a1dr/5VX9Ab3Docy/
ct1+t8IciFNS1qXtsL0pQSeBdNEWOJQ8LDNF/hyVVw8LmMaorg6QCtteKebYlOBB
KmVhcemufurnH+en35ZxBsXduCbsYLh7lBQ/eqJBR9vKp/hwBYtN2qTizPk6SxJ5
sykTpYvmYXS30tJSi/5gKojO6DdyFA1nMy4RcxXOf9Zbm3p3KXvvi7aZNjYbXOy4
imLqNT0j4/4WJbkoR1JHCl0UvqDd7esG6KBOCKsP3SpPM1OZ2XaIIcgmRx/sAY5D
QUE2n0FeEtstEXyxD4gFL4OY1hW1JwGf1E1pNOTB2TRmpS9LHlj9dIdUMhmTKrqC
3cmYn1USINZUC/JoXTDoX3DsriBIc1+16pzbfUnwoQquY76skraZx6Kya8MKMIZX
VOzkL0Pwcl+KZ2MsM1kcBUL4Z8H1l7L040AsZL8LHlf0gLJTAorEvv7fyh5Kyrrq
29TjAH9p9frzx/lqY0sFkNAVcx221RQBc2DoQf8o+eknXHrvcdAyO3wT5w4iFXtR
0JZsWrYPernLJf3jY//1jjaj/A+r06cP/IpGnJG087syrqWWWyU3jXOFHPu4ZTkv
SzFn6t4ExXS3FbI+O+Q1o62+T2CmZ7jF6kyJYUhYgKUIR9gre1GKc2p1X7ewW6BF
8jRSUPr8KMgF+gBx7lvbqSRKOqMTS0/qnn4cyxCGZngm1axZymG9TmBTifdw3KaJ
2wydZUgHiXyF4duVyLitN4iBvoyxz1qQp5kL3y0FqWKqaDEg7iz6ahsiwa8HeQ7q
g1xYnpa6+x7WWQluVemj9Zdky87lRkOCkV6ORyozbrr755PkTz8/mttNsoKCKpYV
Ez95zQmwQuTmrvhFkhSX+2TY0TxuF7siqoGpwlmtjmMVBwfFwrXAxMbhZVdXu2qs
mtpUCbs85m6V5xQgBUEp8sy3iEUGr34UYr8h6VPeyYk79b5eGJR6Un2y4yPePyBJ
kEg2cyNNVWfOjQQOywOuEiYEHdybjforhCLWQAHj39Y/L2/zb1cNch/lmxxxPD+3
4Xx1ErNgCxqraNfsBGmvs2FE2hFFOm87HVMoSjsZltc1Ea1d1/Xapq70zch4Hc/S
9yk1MRted1fle3abBnTyqaCLo2IANpQ3gVU5b2zIbUaKLuzZ05tpQiTmSHNX2HjF
BiVNJ3R3RXRawuVrfMQlpfrqw5WtDvUmrI0emo1eZKAoThOqEYl2A1t8RXf18M03
0VwHwejeBdgHSQm/lUNMD/hACUVvfMLYb3RTcwrFJboRwU3QebwIfmLgRyw8P9OQ
/rypZB1uL4li5cx1C70Vq2g5Of8uA3VmO+Q3zHos2Jo+rN+Uq7pbRhzfPqY8d2SR
gzKfPXANm8KqZIfDQXygPyODXrYvclRy4Ex7+xha6Sl4xanLWCXUc0wXzgbFZSLi
8fdELFzz8dPLovv2g8+2Fu4p2H01zNzXQt6ptNggrb8h1u6QOH4bvKmX1SjYfuW2
FhEEbyV9NyOrVv1JY8hk97pgrwJoXQ1PHjQ8N+BxMGo26htG7yXVeeVYx5DbYCUn
UB4G8JLRPTXvgJTvogLZKif4D8fYXaxN5+PZ9uWjyu6t/RgjZZH1sqBz4NgnEFCy
bBUgiKvtdQJznpY5Zg1ufPOgeDINJh/cVVoGeaHAIMJ4M18mB40bK5wTJ932kKrT
1Snw/mfcMtbXoz4LYCzWlnqanbmpj+pzgM4LDPLviFOq8J+9PkA4oorg34oy3hCx
Xb8gvgm3ESVhnZ002OiTPzaid6yOy5QApyhCFBtrqHdjlGVIOZspMXBzlWBl01Vl
TRtoaP6hxQZwKZbrrI1r7xHZBAq5s8Bd63LGbDzBqzmPZmNvBuSws0vbctFH+MWq
X3ZHkVUgddb8hGudCpoJuPVrjdCLTjQx/nC/H/tJFx8GyQFavH4rvpCBht2OJjIS
se7lMgtHGOcdxqqfDUwDPbWEL7+/d6M8DG/3bMWIKYGPLfGl7X02iiBCSaM2cB6w
O6da9VsuzsDsH13upLhvNqtSe/Z+xgpjYBZeaefFR8TNF52NljqzlUbJXBNDZW81
EJtnVMi+prERv78jyqQzhfmT8DsSMH72HrFlCPiIedJzS5fZ5FlZVwcHzjqzmr+v
bVZ+3HP+3XIEH51kthdNLqggxtK2IbEqBObxyFmgevcLH1gkHfWe6VSCuXP/PTYv
37lVqGvTo8iik5SWO13SxrylKF/IkANMOkXMPkLK5ZxEnQCbBGjz/X4OehTSafM7
katFYNAcZB09rLn3XzZmuu1JtY40/i/SRZ1E6cLjQQqeompy6M6HabW8R6AO2aSg
N25XLsnMYu19bWilN47hiKbUNGKBLRYTwfRkX3iH2/Fnho+gH18heLq/ua43zFpQ
YYGKcUW71gUcrFFk1QutA1WD6y0OnFHFxlPb2UDTg1kdX4aj7PiHMtT1JY3QrD4G
OPxcpwAiOSt0k/4dJq0EV1pP16oJIhFDm7srnh9dR67BXu9dMIwrxdxrqNnYNYJg
3y2BdjS0gzkkFhKcutbcwvjmQLGYYsPyL36GV5r2oZYWCg8sIIQs+OvkRdC5Ezz9
P9RMSB2ZDINbJ5uYwQEdywwvDW5fiFizmVHqVNYBiBJNAmr/JzcBeyi3C/tnmizh
NvC26Ii+u+C4F5gG0enDwCRAH3NkcLlttqZTKESQZuv2AYk7GUlWN3YaAmYM11IE
aKXIPkpJNbfIv66csPF1KOfbYHPjq/QoWHRJl6ZTAtV8yIMxrw1cXar7PHLy5al7
5CM2GGYw+tCpdfnhlDoWMIJ56KWE3CVCVYWmS1j6kZtzooKhv7+3dzpVFAFY11UD
JYyQnj8UvlYK3FFiW/b/HWMLRSzOQguDiUZ94FXKe5/LioY8lagAiv/FeVAPN19s
2mWF/CJLQs/80sTicO/0h7iq/f/m+q9iiyICP5JBBTY2Jxlz56QMpPHGjbeo83+z
JNc1HQExuvaFwwhDK4WwhwcP9Jd3XAmvDe9zsXFpaqFZGXPyQIxtvihLkbRqI+Jl
n801aRBX/YgiDgtmvmOi5x3KJ14ENS+eyo8amyADkjUCQMSjAQAhMDUbG41he0sN
+zazi/+yWvv9oNS31+dnbZatZMH/wy99qJ2iI3y3Rjg4K+VTyp0hx2XW/cLrNIiI
NvTsDkW7+OStK1a9ZQm6QbqOX2IhCESlG7m5Ax5aJLGoTq+drfVflKBTZ2zNwXXo
sb0tvRtT9Cn6/66jIcCLfyk54lWBjaKLSX3mn6lQrdPKCkxvCbWs8xXwqAe28bCR
+srSw8HXOQYzqpqUXCgnfOtDCYr56BQ3riQagxJpsTH0SOda4vCbqmlzp4UWOynf
sartw0fuFeJimNkD1GrAXftK3rkj+cK9MgzHN73OuBntg8R7L0bGsNgFIwNiXIEI
+qgzAMUUnOiLpiNUnybHZT82djbl7UCGj5nkS9AaeZQIFrFSXA51Yq54m1QscFKo
mdFvjdvkgqxRYm9QN54lu0ttY4mKu5SP9MrTppTeHgHCVO9uj4P2HG2+d/epy+1A
BibjYCp+kY531rZGvpowfLuZbEBcp1RVS9ZURJDIrjzKszUKGjHr2IEO+JK8yG28
C/LjpSXXt+7+rm9Vq6zsAS9p/ZnBHzV+JiSM+Lvu3If+cPwyF92Tsg13QSKo0vzU
wWD2xBQfqblzZrBLBsZebf9b7YjzX7tPrMpkQwYZQjtRMR/ZTRHVc1VJGPC0ifHr
/w9nbMtwBCwpz0N+fPmOBt+VHJvrRl31dIoT/2wHXiza2Lc7qAgYGC5uuuGiiyQi
A7lVNJ79mnM7QZd3GiFDJvnOMWEcZDx5R1R6OVQgiuRQumlhuwCjs/DH1x8RDltf
3zKTEkAN4hwkgIZYNmD9DCMoHh308k8Nn9Y79RZ8zves8HFjX0AiJYSOz93Epy5p
73fSoytWoZSrSVvkypHk3zP79j5mkonDzYXMRCI8wEfiriy236GCUVD9ot9aqtVR
5co4qP3Kik3Blq30Xv2+1nmRdCdf/npFqeMN/mCLUITA3qtQg8ecH7oh3hGe2vCH
hCQOI/sgQthUABfshQcCMmryurymjFNTVw5Sh1RSfR7YrblfZi5q74w4SVJoOlW1
2341DPkoMU1SgzwoGov2useQNrEQAt3+DMX86GEhhuvqR+RfFQl1JBBnWmZ1bLaT
7hy/Hzm+MUxjgJuLftN9ZyT/PNyWuL2P8ZLAm+LQDp/G80sR0WUzDGdefbL17XuA
rrpWNYgdn5EnB6hoYpyA3HqGECw5M20WyDciUuisfWEkTQWn9dHSZy0+knMp5S/0
KwGHlzvd5aMK77ILV7VRH8qYTf36Ka0zobvbvqOyPhnPFwmgEvTD4LKMyth5hgT8
fxiRuhZYA5Ln78IB0fAtmrJsVbNFxhoO2NdOWwaoiveGxGs7UQZ/7IMI57xyu5Jp
UOIRnaEqCw8/WQ3KbpL4tJm9YGCnaOp08GRAGwi/rVmrJh0j8PesIN0P0bIy566M
hr6rYON+nQlEYXcAoW/SpfwfuaK4fduoaZBUXy/gn8kfEhnJsUNFAQbKg+Fetxo1
OO9drbOtat5/mrZwgeiLHlViP29XBRsI9umEm+Su5Q0A7PDluL072IltwVX16BlC
uAxNNHTEvczwp6VHaF+ncU7lE/LtLlCX1WlEgwwjA58OgVLA6eYc++1YXfeslbl2
Dq3kPc3vbfPGviqu4XKbrg7uJotma/IdbRMvZeDpWQUTBCsbqLYod1zg5mSOv/Id
AVUS05JL0ECbtGYF2o9B6yyOu5RiEQ2pQjHBsIE/5gfEI/Txl1/vKJx9BB6yaTY4
B/y58YpmqerUTsMVQBedICPLT5Ms0eJQyI3ypM3vjLzMdJe7MRlJIWuXhxiq8c7w
h1QbHTjxvh+2JUfuX0e42qfAqGWf/1BA+Rcm+kPgVfT4jcVNI2K+p/iir7Tj3xh+
CY9fYoPijrJRwePF/sWoHUfau/Z7LJU8ZGHh9S+Yr/PxiE47WpDC7UCjfEHjV4AV
dnBkWUaXdUyuaIFnjpdNu6tN/+7+cg+5hJCILpl7N7/Ah2CI/BfTovZ8wOXOyybh
blSxy9qKhX5lWbAQwZjJt+qCWtHqS5uEpp+7yfOHAegTQwKGCx3jPXbXXOTlSF/s
iVNBSbfvxHZHx0oEJlVLU35617K64iRCJ7+QX8oftrgA1FyAUgxjxoOTm7qTuwJj
/bJojmx/nFi4ZE0n7Oww1q97k7qqs4irJMYv9J4Azqy/gnN0+fM6R4soO3GSBnOI
QbGmSkeKvWi0v6qUg4EHVnl7ElXYXJ36DqNVqA4T2YmUy+1Q/jfvXTL6Vyicghb/
QExhyyhVrRhkqNFYBtp+/VPdX71GZgfiMBgd3iXorVQDow7ZDAeu96SB5bef/f/U
TtfV53/TiylB1dYe5UIGloIYA+GxOCa9IyGVHK4G6VfOkH6vT8EukbGpfk1LDron
JYnzEssZnxmhb7bh/HNnKAyi88TjT4mC4rQTcR3aMtnrI6jL5rbvH79VuGkdOyIC
0EyHAg3rhrgfF61Kf+TzD9xazWdM20VYjROea0WwWxhXcL0s4eitsfgRGosAcXCP
DamwAHhwxGFme6ccc90gNl35ln6Jh8CXlK/cCg7/6DyGpRcK+j3U03eLLZgzZ/IE
7EoryFCMsKe/xJD6S5UbXu6R1JP3PZmulgimd+5HBeG+X9g1Eyl9ZiepmYDgAllv
9U6mqvcUD6vTM2d3PEtOt+BVb9qFN0Rg6k89YgbLRB9uvx3H8mM9MGQy7uoPY+Wu
wSEcXA9GR+5k+kiArsy8O20KN8mrLZTh66MVpSN81pN7edmv6+stCzCPeS0r6VnF
uoLy7ORk66qCKA7pelkrBvTtYPpW0rt1QyuYLei+nOiXJKw9Lz7UtGNWMkes/coa
H1gQwbCK54k3qGQX8joH0iepn7mmAucCZmc5Uvsyy80FK6VIOmyl293pbdU/HSRh
XnybYyFsGI5ovZ8zNwAmVUH5xEgGcggCAGMyjIt2Qlbtx/3GZIPUuaznb241AKqq
EN/gVjuF0n+IV5femzENAGiWphUDSWlOqJmFD2NjMpZKuj3piVQTDW9HUZuo25HA
EK1bF+oHqWrQpLgJJnvWY2IIn3eCVFb69uDLytdWuErgY0WmY4O3JDg1pqFYifti
bIbU1zZ1GFvKrEpQHK5UHDxAuUdaDh8p6FibQNfxjLi039owklKWutAZ47qftguA
Jkg6z4Cd9/oPZxoZWdQ4TTBa1GgPQL5zKHdnK9kpe0aMzH0SpI8E+mlljoUs8o2k
oYXeNTsMdUYwpj+RJ//dsYdqnz0MwnMx6XKCXyWxo67MTtkAqUgD9DRpmXhzaPNI
tAEBh7s+XyleYYSpts9SrodhM35oU1SKmrcbUk+cZTLOTx755AKRp0hnIiMBZvUd
JRGITarzHmRPtYg/KavZGfc6NwsSojwSDlcP2KDPi7D9AiGzXgZLzNDPXb+Ugsl+
jLBCx1Zh9iTzhgJ5q2L7sd2c9Gz8AduXQL3V+exoS5dM3g/O0dLfiC6Ux3ElpYjE
z2h6pBkEl0gecW3UwlGCRJ2rKPEHspXotebVl4YaGCBglEbTLUS4m02ZTDGrRzvR
YR+wdODTz+OraehuJTvdXbnVkRfY7quRTqheXuE+hlEbuvW49Slb1W4lz+M9Z7A6
ZTin+xbQbwq5S5bqoMvgDPqKr1c6qnUS9ACbwSPKU49T3963UHH0FKE9ksfNh/EL
kH5Ab6lBXOIlNMHwlLS9xHWaV55Yt4jf80lbT0gyTWyUPRVlX7DPgZ/3stwHbZrP
IYpDLyA6yhidz+xO459frA6gm886i9B/GDQOKl0IySfHKpbs9TjZ426yQP6dlO4f
NF71x2R8doSZq4dRIW9nefWgF12LtoQfsOXQWGpzsUDk4Nk7ClT/kSHNUlpwD6A2
2ctEBLl4Xw2tH6TCbN9BA6DD7YdHgS1c1/4Hh/PWTBUcAODNGIwuAOCpQRAgnbuq
8B9AV6WN9R/RPmi6vLBOteGOfLAUqQYD7eRKhHQEPvnQDhDpifBACi5g5Ns8m5ML
uztbOQbAaC//ry5IhFVo5EXcFK9GbZCdRTuD5Abn0GoLM8Zpv0HHR6vt3eTNlfHW
Fdm3fS3DtvD2Z6GsfA64vnyEe4X+DI9BHSszVEMAMa7k7LxWNF6/mfs/NgjRscRk
e27bpnJqhskNrd5pugpJy9g/l3Di7U0R4FUBQxYDqutsjYPg+RYkqOPDMdMwWSku
DLH8l59buTDGRvtM5hv7zaq4EGOjw+eA/IGwvMWNgpbHBr3PvrkFK4lqYgFMQUg7
dpMVWJcD6M79n3rLUt968Jqy+x/bDTqpp7GgXr8spp87mBNFbdCOsERMmM9TrAwb
f8C5bfEdB7DRN2bpJUpg95XwYQ8VE6cQDgWP/rQHo+ecYrhFewbgduCBjkzTtqej
hx/D0FXBr280fic6TEZmwH557z5yWgt5I86Hbc1b+2Vfy9iEbu12A13yylvWwtTh
htASPAhfqBWysF+nOpRHJxdSU5zc4/5nE9ih91HdLUP9YLwgboH1uxwaXwmuE/Zy
kYY1jVqNvMiEjfiyC51/FKfawEk0SpujyKNzlZfXvSLCijUAWcx9DJjOU1gDYQBU
K1UKXnyLzkCXHll5XJ6Ze4VY6jmGr+47YS+BbdHV0aonoQ/fZhYG/qPyjh2lcLpF
ay33zmJceRMJqeeHzQI7DLifoqp/nUvdUk926EujoMPQaoF2AhwdI1EnZfCw+3bE
6b6n03tNLsiB52a0KMj6bsxLUl5MOD4930befXnSyLohOikdICH2bWjUodtO47Aa
hmIQw/VfR9q72pdGkLs5CE/HdgrMhXDjpHR/7goGCDHuCBOMTm4bmQr2EV77xDJt
UXyremNn87tn1W7q9dBlkBnnRfHUr/0T8RKs3Jujx/dK4U/o5yxHlXvIREIk+IFE
X92sb4i2/M1TKbFjmnAKs0XpGVz506bmvYMskM49pKZamCcrjPie/sL6+Rd6qBvF
3rfbK09Ht0xV8yMDwhnrX1bh9JK8aiYR4BM6X3h3vr/hthZWU6GURFVpGMK0m4Am
ULgknWS9C7kAD0fr68EeMmCWBVDqUZA4+Nt0TXyviQ5ZV2Wi01ixg0RiX6Kzmyky
3YGMRnQTYfopRFI3w9bYBnyoTvwBzF4+fO6PHVZLIkWNMkpRhVX2S0AUqF81Za86
CfbNjha1dZ0NDExBd3kSbSQ22IqEVfedQIsycHosJNiOKszMLr7zopZ21ssZYHiT
xnh8YnG2t5NUpd7saZzLXITjpYB/pZ/1gnpwZQ2CJRFEeYAs9waz35KcBwIBc1+k
EsMmE+FqM3MN2yB0/58ZGLi/y8WkCXa3yhmfupHuVPojAbuVkkG5tfzD/bLkRKaG
EG1B0mgXOoJ4Tn6Kc7JFWk7L9Pzkr9zvx1Ne5JIq5U5ZcF01mh12IEVYev6qK8z5
IEZGovTA6/RxumcK5g/maHqN1T58kpkzvv1c+bZTm1KJN9FO02N3CjxPq8Umv8s8
e6jKeJvyel7pRdMc2fP9F3UDMlz7wCZkRa0qNhLrKYiaoJiszjyt2x9V4ellRfXJ
wDs7J4rH96Ut6bhHxd3nYLNWDR93WigLwQG9VcqpZDT417AJ/aeYDJmQd83W0rh5
oECj38poOGxQBHJjmgu6/UlXN3Xf8XY03XxuwtAeICh1Gj9ELIS0zvR00Ai51c2a
LOrTQBmmGAnU5skve0WmI1UM2Zu2WP0DrlARLhWxdPO6ay/rT/lE9BJQtWP+oyJQ
0n6KRz+NYNyB6G9FTk9haMEYq/IzVC7fCVkgGSYyS7lI69RrpJcjk7VNexaunz2b
x5UTN4Yx96eFTNP41PXjLXcC4Ur6rssTCwW6xCkjrdNbEkXWlwFbSyobHm1pd8oQ
LXmC/BWCsu/KHGEiEI1ZFea6ZjmX78GKFh6nN1H1/POQOxhUfOYjsLbyW/R6roJ5
zib/Yb4lrUrqlSuP+yTKsWbHXhUT7/vOv8O6TNsVWniaR8emV8omI/+L3xMwrv+i
DUyEol4HyeaCFhstWWtlVpTHFn1g6o/VxG3gTIkqi3frgtnwmZs0yXvCB7N3H44d
YL6Amv9uvRYJoJi1ZHo9W7fIUyPLGTpXeSO6zpzQ2SiHpcOSZ4IJn5gy1O69kDdq
HPTW1Rat5gyIUhN930VQk0t3OcFZ8M2ImTcCq0wfK8vof00eJngqS8nhqvAqMjcm
8nxy1wl5L8ZVIzVtq0mSdIJ55jIr7ZkDmqBfe9+UwrYCdUsqfOjWALOa+H6GC3Cq
47dxOp8/3CQUhVA0l3kDcOZTlmTHd3PGTBXR/8ML6JrhgZfO+ive+Ao2aTlXjFZ3
78ZILVYUJFASC+oW0GUMNg87QVw2tW7VsJx4OjQuuoEgj/6nl1N0EuHdbFhOTrmT
1vsmJa7h/RlcCu1Jn79dQOfl4Nr3ZiAUI3kGe0q08Md3QEyMZRyNVOAMywmNxwev
W26L3H7rIlkV71YtTnvhEyCwam+fO3ei2NJAa9MyAq7+lJ1H3J7WhKtl6QTcGBk6
YFng/kSoQtuXYLMyZrKDlEsOxYumXClgbffhZitebX8ds2IuIC3czoV93Ewj//NL
K9RduCwsug+v5VinCsrtwU6r8z+gLlOMkEXz8tlb5KkDGjvRiC6o188VR0ngDvXJ
kAJhejKQizVgvdUNpa2Ri6Y/T9k0uBYXfrW9PCN78vJifTNgeKpApmSDk3HvSrXP
R1xacB+Cnl4ohgW4BfW22DAkEsSUn4ehu9X0ShQkyN1eJnYf87HOhP5DevyIeVu8
vEz/fccFtJWYekamOydXTsF4ynFSYzAc3Ke2dLh4VW4ATxXjBKfaCH45QZQrvK09
dV9yMxUW+qD5SCTVpJh3cXipocjPWrH/xjBayQ1fPYYiG6hYvNokm6JHQdvAAXqT
DpFlEmdMmYEWiJy5a8nhNHKs4i3KpgQ0uaqtXcl0BqZ7hO8/wAovg9YXi0Y+++K3
tEvfDpAafeAzssy1yNhozoX2sGH5x1lJYgWzSg8R510y6p909/vrqpapcaFu7LzT
z07u8h80PhKFqX4SRZhJGTXsYBLUqjfPFzKWo46rwjPfXkmBROdV0f7NaQE7war4
x0w54i0IVxL22fFbfoDDviAVYmrqTVyJ0WtzNf4GbuzgciHsrTonfI2YOKappsj2
au/fmdUN9GUPEirZEbe2iPQXsJEDpApn6HRYfyTGKQMyCMGoeZlD0TBNEmWj7qO4
hyvZjoeYZjeV+y7a0QSBufg79Pkc1SZQjTMWJKU/X1Dl9FRS0kgH2boBEel0TfIp
RHsAOcxWBxgM1RQY8Ct5W2RFBdRbQcnomVPSWr70H0oxLsv98ZHxuUiZN9QGxQiU
jX6J5sKTqhyM56NH/EBvepEYCSVyY8F6MAOBxIzuYfmhUHQpErMqW5XS+tIjl1Bl
9jxEZqdCUMgDTEGXIx5vygvkvOQBJrrdOWhhTp0CQKY3VsnlHrGx72F0mI4jjZki
H/CLQH7iU0auCZ43+hI4wxt8aElXseWVVvFU23aInif5Tu0rAPIGDW/5U+pWa00R
tnbreI8wnOzQNlA2Es1nbUxMX89O+q4K4q7CanI95hXF5eC/vnfThE/bfmcOhCDg
JcVo7+YetZcBrNTjqBkErCNF4oNUiN3imrFTSVBt5r8BpFuhyQA1JAzNhZn6Bdbg
A5MoWB2CVlfWIzE0ihSDkZgvgwV7EmLC2q1jrPcl5bXSM4yasafQnVWhKcG+NL5L
yA2SIyhqrzCXCQ6c+MqvPT69jlMI96Y7WG7oGKoNP3rNw4bk1wiMV6h/UIGtZGbv
iGzNVaExCfsLKFUupSgKe3wTJG4ZLbsXn36nKrNsrSx/DBuRGKZis5n6iUfX79JF
85/u4udPqtUgZfPphRrklpHIiz/gkYL8+mjvyDjQdT2P4YBduW6TRdq/a0/3w0Jz
V7phpLXTLuBANJI/2iylhO3ZbbKSPD5U5uB5H19c9ubZQEwUsKTPFAqTroZulI3l
W530YOcIr3md/94ke2B4DKN/CGPOAG8inh4I6byEx+0Yv6frwRNASMjBGFlRhp2j
M/QfjvZ68BS/LRmgwtrqQyDFs5Q6aN0tHn9jdZ9fOalMqyUr6ltiUIhgCHbY3vfE
FWlpTIKoqHGgMH4H8g4Veciph5QX2dVlse6FIVU+SJjiGvvV8Z7stUUvxwRxEfm7
RNlTBpf6PepCuifmdp7iMBbV8Li3m/eWRGzpOHtwcmE7plk6Ypv+J3NpCJ4LFOxI
tHH2BGyFqcBVHLS43E/oHlJIvRasB6Vba5L+TA3+4voLuYe4U4BXu4VqizYEzw6H
KtU9FK6OHsA+P029FNP3ZEdGI9Zz2IxkS3AkvnCmEx+Dolw7s3MPpXBXniZ2lI+6
KE4zWktla/nbOEomlLng1EPXjoaNw6Ld1DZXpSCVe0TR0kBJbmQf+462Ih2KTBBZ
8Q8MANfFrip8qw6Rh1VfTNatpWWVK3bfezSDIU6cjkwzGrmTQcysWo1/ohdIRX4M
5WhjDBIGO4BlRQkgL2IVvuMRs6yGSsjyLJwDrkMwROL89wCj2A0/URTKY9tCsryg
nhA4QTXxLQzGZIWrd1Tj+4WxXq+a7AQ6pgrDPXoSwXDdArf73fT11i8rKn40PwDq
R/wovy34XoL0l5el45QJdpsZ7US7M+tFrX+gf2MvUyjt07lXbKgCS398pUgPHDtY
7ZGeEr7xBK4DoLcdxPccKKVWySZiALD2zXG7D+dwYuMlqeMP18VhWgTj5aaC72wN
dEU50INGrM6xVULtBuPOs+Uu88DNUOuszZtXQe/RhHDsp5FZAqgVOQV/v/a8ijnd
MxX1dIJ2KJr9BpWiunXWEziW4kE3s9y0jtZR6ePGbTpqxKGW7WdfffoqTA3WPWyK
9CtSK8K8k6NF3g8v695J6vwn+QtCbKaratfoiH79nQH+2LqN82Gx7hI+ONAd6Cu+
INNoZGIybduiWaQndb0tMNfE6dkzpicIvMla9Hfhu1EwapGY5xyoi9WR3GNFFAzH
h8zayhetPq4WuriABG3DeKHinqcj4p7axca3Pr1RjV2nusiPIP3r9noylzzMy3/L
hrz0mfziKIByrYlQprRhU4iJJdKapAESRACaaTbwalL1kQ9TN44HCfcYvg7yBjcg
/gnBy40MpxFbPiF5jgJwbiYH7QJOWRu2PvQjLmxUNZkohlwXdcQJM7meJZYQkZ3u
GcS/DzI6kE+CJZe4C31IfDZZNPM5VsIem4FktnhzCsUTc06VNUu1P+f+9zK0O+Si
HrZFBq2p5icrj8AfTem8NeGIyF4TV+tJX1wtAYatibsqHE2d81FmBEeckutjvC+2
2N0WefhI6YJBg4aNbZWG1i36+A/0n0yVKtbWjqCfYJ8d/iSwsPU1api5H0a3Jrg7
AXtf2l2b2PVRhnoQ+Nz3BtO4DOZgOc3M6EgxliP5gZmetM2z4IKZ+OLptg97fF8q
KvRzTbyZjUgSq1T1AsxDEE5laBOqNFJj496GeDOzgTiHae+RRTOuwF3zvlN+qsdb
2Bj5RUzJCps3lyaob57pmwZAmVtXSwyWWcpTT/yCOh8SJcEX2AztAWRs3SgTXr6P
Mexo1VZu0CoCZdw99HMY35UDrnWgQb3gMpdg7P74zA7A0II/HQg89BTyEUC12r3J
8YwHQ80fpPgwOjajub1BTBOoTuFupY2TZE3MIsLga7S8+X76kGQViCrm7/+DugC0
m4ic5bwgdEIv0/neBPnRO6EyuyXDmsCiW8AV5bXAmk5m9dHZz5f9JtbcEsXs3AjZ
HHmieIsfLDjjhgQi6TRMmgdOOZpWzqnxQjM7ZUtsVCdr0VRLn0l01Pa663K4MF83
IlriCNY9gw0jhC2shgNDdFQ509uD+uQDn0kCDCfwjxPecr+DgifdTXobwQWi4Csx
profvj71+e+9/ckgu7rS82cXBENX0aA4QjKUVQcDCue23LT9tBqai6PqK/m8kepy
vVWwjbZRNQl7aRWRe3m/tbL/cb5JnC65ovhFeh0lnFBXcpBDumMRrotBi+C9Dtfh
TouobLwC8bpvn1KV+sPEKlFS4NQUMVbSbGCZrRdA/JnM3CPumjCUB1hzFKtjDF9o
/XSPT0QcAWadLKQHiENfGvsDvgo5gMzyHv31yF4rfF4QX02NnMEsNPlXmS2CAyYj
EKRN/NIribQwjMxBfFphwm38MCIMifVRhVZZyVISf1fUiPs86eJVEygb1fSVUAtI
eBof9rPJrZSTRGmkq0qajw5/7dGBMhuKO/Qe5WX/vT0pBVolxr1eUyETDbhCiz0b
NO63hCnkn9FX5ZBbrdMi57mowS5lLuhGyfys5rud/ub6GM54Ah6Lutn2+Ub1NTXZ
ONLpAGBnQI+LsEx3knV7yc01gllssL8ZuXNblxjsVYPHxHCH2rl87zlQN6pQn+ZJ
6wjpszRzdWwvcOg04rIlUO5gvyesR5/Zd5oHliiFqB+3BvhHK7llNmQ2aIIZG6xl
1atNZg2ocT+ex4YRMjYtlLSz3HedudQ/bQmD9ETLrYa1CNzZ4QItkzgnujf93GBz
8z8kjrdejvey0Oo3xUAK1KNTZyfO50wAbiRGUVyycbPvDeG43eUyL6q5HhlABWdh
LCMc0Fe0DI168DeYAKBZ5Jj37tNSQdEkJSjuQA4do/VPzMLdPaE1wMrzmr7GtjaE
7RKE22AqQ7cNmoH7S3h/GujBWIddV+GbqwcWpXWBaMzmrfT7pbjj/OaFQh+bMUL6
KfTo7yjmwKD01QLLohpIGAa8HWHGGW7tiJx/FvJWHPLIVCsnQvKTpDxiihjwTGM3
7dhtj0mg77urH3X8x/PkZcg1g+ggcdCfslZ6oXssV56BemaPwD8i9nN1tNLe8KSl
vcr4YqEGwUydWJPSmBQER1dGJRpyVrY+MZUo/pXseAB+Ohr0NGdmLGcwNcwImFLL
IlGFg/Owzxv2v+/v5l1JzgQnj3vtJFCLFdSEiKKPKGldFc0Ap/IqgvilDGjsmznA
ef2hQpRmjB4wG3Xh98KjUSOrtOXnpWrw0JVVQ1QN1KHizwrh0ngVXseMdwJFDu+N
++qwg/S+2e5cHy/uhZEs7sTbz7+/vJBkuF64OTICCz94JSFbuURQE3QVWCMMV/zd
GP+FWIa4f5LzUaTJixYPNAjyKdfrIeqgeawlheafoqsRsQwpNyL5IU4GdunqXbAc
GPiDt9PnNsLFsm6XICkUT50e3OJQjUautzSeE5lXMnJDVM1cX2GOY5LlBP7xesVH
2SmUcL6U71pk/cFXUddwJw08JXJrh+FC9/O0AQBbc5lMfCmP1BBc5GyNaM8uiJgf
m2OwATof91Zs2aePn9k0KIPwKgklQyl7Wfj7gPwkkWNfqBbpSliav4mo7kX3fqR/
uVTwpRIMZQTlI8QPOICwdRboTZFeB/r9OERKEOW9gk/Rohl+da4ZKt/d0KquGjWd
xICEXWOt6p15GoH20r/Be11ZsAqRTE4d8sx9iYZ5+pKHpj9Ig5DP7uRFHBMSjTB/
/RsD6iUIVFz7Zu+r0V7XQ6sNnNIZUxzjYlJBUcqyTDknjkAXCeZhPmwLHhLVMDRN
bu0/+Uixl8plf6nOVh05T8K+1Ee9qEn28ZZe9p++Y3QSG5lZWqScbMG5Y1Gb9HJZ
8o0LZxClCdqaVvhmzUEltG6m5XQcq2W4s97hie9qtVdJKse588atATJ1ey/xl7bf
X4wf8Rq3rimlfrDaNgLJcDYDn5aEPzrlrBu0bWy5z8GSFOj5a43xYmI4Hlye4L9M
WkbkHl5c6QLE+XIvFK0SHO1BbmjeVDshZUr6sNyDxmwiKAncEpp4aO3JhXZfkABG
8ZAUkEHs+16k1a0O9ma59doqCzfiL31TGe1xji8Pkbo66auXVESmtFlmIXNY1U3i
nkwaSEqJK+eDVrxrv13EYj75ZGq6m9BhuZkNz+NgxCnD2GAjkzk5pt/1n0nxFKcT
XFeRwJKkkgssm/zlTf+bALZsEQOBJgSbqediXbE7CeLrhxYZYM5tiX+eMeJjbrHv
Zxf1HHNLwq/jiThOE6t88w7kBZgfBkqxRyA0nk67nJ94URtvG6JeGo+pGbCW0Fsv
AGKS0guCfu1u043gAMNjnrAXHEQlcVAj7NlYR6lVDHLmazvqCJuBy+xXyHl2tvxO
i2NbrOOEJwhTEFiBpYSi7Jar+wa7OC9z+j6JA0ZOna+3VXvth3vxAwJ09p2pZyPr
daHSfS2SLFCY59F0H1g4I/IDr4JNlBHTGszT4EnEW9VRHQVU+u0j7Hbz5AJKEnBx
G9/H+RZ3dTOsKxwBZ04gPVFxnUzRyQCP/QHUxfV6l3RH+T9UFaKNo6oPCdbtZsYr
HEXNVWC5XowKUqUyBgwn1wYrntMrIDuVd3JZ4axgA4FcGGTbzOrP5M6Smpse32Qr
HMbRr+PigfuKjYuH+SvyNhxDLREmrDoF++ODnD6JLyQ6vIQhHHOtmC8Yh9cYJo4u
+BLXkDArOC2hbPD3zL/fEMC6ezK4ig6SCFYt+zbDqUhVpdrA7lKmhFuQJ7cPgtqr
uX4eEjQp2wOJLsGPtJ73+To+//KocnI2nroMwCCDOByHwh/3JOYs0XSHyZhd5zGi
GCaQvwlRUH7qzTIoViVyWpuBvzWCdYjKx6xBk8exukYFyi5fD1zYi39wzowNW7J7
I/asNosROM5vWzgOouEDw39iS7ZhVpwPwkJX54lvUvK8IEHH/P5TCq37HSMStwoy
fyQbRiKSkDqZobILROdhInmf3pF2DsqrgBEMe26V1wUT4vym0Sl/pVv1DHIuuKzs
asKKydAvuLeGrzBW876GQWbwEke/uiSVXoXc28Afn+pnitceh343KtQrDy+nRtQU
TRQ6k7qITP9FEkr6got8pMuw18DvAr4hvUxIoNoPqAEa1uvbGb8v2L/uLm61LgL/
uM5H+XualqBYph+LoHIiVaWeRBbc2F4DkQwfr8IsM3Ml+Wd3MEt0yPHUaFXASZIv
wLVgVUIBV+BCRAnwrGatNvbBl0vA5tDhxzX11njR8+fP1AkLx5wJGIGCjzFc92q+
fvFQaaQvCOhW3gRtTTAZxsjJCzGCg9gk4/KJA4wKF1mdIuUvdWEz+moqH7tpwBj/
3zvdkz8ATkwldFzrha2+0mhqwzCsH+7/7AS2ZliO92Hhh1rIadK1ETjwXudytFbO
JXLHAl7aXQziObDV5qQideYUH5JgFxyRAH1baHWJVUTGUDTd6hzvuSihH1O7M+wj
j7380/9l4GdHC5w4bXI6c0UlvUs2pVjkNoGBE2adq7NNMe3WniQlduxt16YbDvuy
9aUOp3jP+TUG0rgB8JU4LZMQ0TuMLz0BqPVHtW2JoleeQQI0JueBg0UpxyOOzb6a
sQ1E7pO20OdjqhHjlKUDhHOKrnEo70Jfqek5ZgX76NXzbqhfVA/2C0iiW49bc4Lv
tx+sKEirgVXLvQEYyONF3aACTTa0SnkIg72QVxhZLaIZ/NGxeTlN6iPK2xSOsYrt
biBLEs0bssjFfl2ioxc5RZmg4iUUci8XpoA82UgKA2sO8ebNt4Cddxfdwxq5BGdI
dKu3AwK4FDON+ziVTnYtAOXlJaG6JPAobv0cd8+34KTUXaxN6GuayueydBrjOeMT
30hnt3cko4hIVLDf99hpEfnluNC5A1VCTMLbB8z1mQNk6dcZr8PE7KvQ6x4FnQMu
yQDvcJIFvVma8WR1edmqJ9VhZJmzQvraQPiNw71DdHRsMxD5WQ8x7UUmMSrYtpSs
1TRxPFc5mkmJUt1E6sAxGoykkKHxJ0g0X81T9Bf3Hl1X84MIc5rDbp6sWZRROreV
lfqsYVSlq0XgYzJQ8zfXPSlpeQM+POC+dGF3FGUHX8r4R1J186ukagZZOhRNXkbV
wWuZhyhp8gLRhgYyqOEWwqRt6ZgLdzYW4q1djRuEKCL4IhW0FMa6bWHecUodj0yY
vC84LjNM8k1mpJ4UI0i04jC+uo6REAPj7Syka3DADfNM4t6xPWoZUpXHL8fpdEl8
xaMm0FOcvQLBJ2I53TS6eUSh/qpwjt/eNYpR3He3cgNowaBeWEsFHRIPpPnsuML4
u/PNfX6hRs4K5eBTQLt+CVdgMYaEpv335SJ9ZmE7GNgOKlnGSuN4BZamH/X8qNt9
4UDiZYMriO6QWVHJgKHfs3N0u4NNK6VtaHDjteQ8MycaivxeLCVR5KKjmnh0CvNt
d4a5l6uPFjp0X6KYdd8Tl2hmSM+G+8+8mP6c3mqFXJfeL8dNcNGFiqP5KO72bhTN
LBuPXSIeBaNvQ7irKdowWenksBYL2/BjBzYL9kR3axhMG7upd22qu2H1xFnwP4YP
sMnQhF5sbsQ/F+oBhX+PQuXuWB/225do/Y6xUU7X35F1iT/Pv1TNJwobuflXih/9
OugoWnZFGxdfnWOXEjdtgdP8fJeRJ279vvqfKZwI4Swf3xuaZbOjXZVt5pHVH2QT
j7cDsawlpeaPiR9p3ZddYyGScAYY3eeoaFyGFfRi2yuJTUq14SMh4a/xSbteVh7g
QS5If82OlOnaN8FQQKOGLbKKh29tCV3lgZqhURAGvenWG6NjGd0nkMlnQdNAfycR
rcvqV/IAN5awYs5T1uksRLVGT78EnqFN2bNQBz+jHicYYVDIzpyVNTB0YZUqAYj6
UpssELe8h0K+4sCBYZ7wWfq7gWGBF+783tlSI3O4gBNR5Biwe2zRXAlsINWyerWe
JjZ6O+b10Dv+0zvhkjvVO2Svp6xMStBoPqoTMFXiRAJCHthT7S0ZEHC4HIK9oMtF
3TDZTTCLExFFKWBfMtGrw+W+xDRSbJrPLfGE4YjxWFncpwQZWUGM7/ctiXTvpsK2
zcbu5UUAlWODfaPBeOEcj3tE6Yt8uBQWwhL2iysLwWHQsLAMYLTcnDUBVv9KClB0
KVewC1dPIvw7T+wEZ+KPL9loy51x2sEEkJQhRi7DMBh5XOOpgJhTV3SP0GPisb6U
URJ1zwxdLDpUUeasFQgW8y9gXJzX+WbHShOOo5yvruFSUXyxuJuas2ozdjL+r4Ni
eL314iMTCR+akfGJdoYhpT9YRUhUU8rnfcjiwFNqvGVzuiliVosndOvDN+GKfLC/
LGP7gm75EYoJDSacLTLgXcI2jKjYSbbmNuMWNj/nU+zqHJ7kE+FtBaD6rPmMQP5x
eiyprkb1mZQTU6vRUy2nc54UlzHEP06VvLBks6c/LiSnUNS9Zwq9ZAS+E8R4u8mF
baqMMzMfsdjIJmZc6YTiWi6424aw1d+6rFo3txBNZxkepvZPJXNEWpfBILjEouTJ
BPd6EFbe3fQt2+7e6TJaMQnNzMEDYcmT/KybVerGtwDmwTMQGMEnK+8+bcqu2q/O
ks2KAqpEAaoLd8osqJr04xFA4Fvye91sSkN65p+Kz7uWOg21c5yQzSEWPJHCgel5
WT8oTZp3NI/c14qiSeGPSHulV33tF2tW+f19CrfB3YQHJVqSytnmuZbQ/pmjQDY9
e8i5OmycimkBEGFxYP9AzoW15J0ThEss5DsB2lanHZEnckRmJp6VB+TJpripNB/y
Rh+VMduxuNzH9+sPErLuBRDwAwQIAcc4yx0snkDe3LCW90zbJYxWnkin8MuUL6a9
guSqW4yTbq10L4lrS1xjW5vFNZSFltC9mSoA8bvwz6xZO/oqD+8bb3PQBJKci6NQ
WxHBwF2Xb80Iw6ki+ekCyvJgMcNsQPHSsB49Stj2QzMn1D2umIg1uxYdU6FGKNLF
UkeKY8Ysz5Zg0tiBrt+5AP3NoFOYbkNObGz4H/eK8JziYeiBmzBrPXU2Xh78l/n8
j6bWGxsSMxhu3hxnSTWQVnV+Oii+cVb1S7ppumYUfG+Oo4QAiOhj+dvHXy/cUQ8L
e/cDKs8BMHo+ar4UwwRurBAs7VoUB6iJ48Zk80lF3hYxy0jGahF2rRuPumiqeMzE
3W0BbhboeCDq5aPKpHexWGtDGQ4Wv1kxTN21PDFfhv+JzVepWDdiJ8cp/M1ihbIk
3sEuJdGlXRivcwEnhpDNFe9HGqa9PsQoFDcnI7gJNDCN1Vk6lr4jooHj117XMxC/
nqVstI5wugk2Yf+AH0NpkbbcM6riMky0eOn/oIP7FdtgmY0JSsRwUPlgfrXOgKts
LSFXJHtsvbaY9VeJwSFqicrIhsrONk/lnD1bkWQ8wE42sPi2n+t0PJ3FtX1AAgRR
nPPfaqrmUVYWUAvZmHb84VBrdfgech/elnRPqhLlWGvGLcWgVqjU+rPy0abL3wC/
UeYyWjLvVy4u/5p6wxGtlUGOXS4IbRCJ6vfnT1SvkNo/HM93s42Qx79NF9WXeWPI
N02nbruevTEjFnMSQHDvfCO9gjCQiBMSZbGowhL6MTlu03gAhlasdsI+CwnQQRvq
+Zr3dkTjAf0Uq3t5U4XB+HYpUoLGK/vgstuZqaqfN0vh9OFuLVTy2T2qfmgKYHZz
8KK9JJHhJiu/Td+UGoby2YmOZMbP/QMxGFazmq1Ou3KiQ/kcbJnhe9nBFXTBrM/u
RVp3iV0uj9wpOnHkFu9TGng8CcuCbG7Zkoi8LOUZX18uwvODCrOfSYivXKn4wklN
cIS7dnR49sHR7XeJjdGumrSD/NZtLsGLrAktxFRn+aeRPKObxPysDCzyNq77jmAR
uB/LFo1nWjh4wZ+DixpCbiq80vL5gyflwowrg2eB37KF2Y2W0f1wI4/hiLjxZ6+h
i2IfvOL2i0gwGrDI/zeRdhGVKEwVV35xBtvfAAbystNbKLzAbKv3p22yRb3YwMpA
qZFxd5zhOW3E3ai+bJjrlKrA+z66MewS8mmywtUKjFS//qjEpgaC9EwAp/aYvgLa
YX7EUDOQFOjvcKO0fI6zjOCmybhV8dHRFqAqQjEjy91l4k9uJNYksj51PDtUA7wT
bLkRg+6M2iqTQ+7+g6Hnq36Yabw0wXWqVOk4ade+xftqptcBve78zEJ+gUohsdDC
fdBfrvkBEwLx+Rsl8x8XK4QP7ACf4qSfpzYCPVmSixDKoYwfS0rlU/gFuhih4p6x
HRF/i34skr/JryfImP7Zp8U162tIPWsDOCwZcVVvv4vpgrnVWu80DGCWppJvm9qY
IZEToNZ8icjtwgg9SNkWxH6ZdY1mzDdwBW2v7ToDPHDRuYNRseteQ1+vFE4AwoJ8
xFN9clds8gS6xQWZtdkClQB48uTFuwyvXndjWPhLgCWNhOur6zd4FEEO/O1BvMp3
XJ0wN1zJ+DWGKHXZ3ccKXUsvW+7mIBa9oltmJk6QLHcjhz+O6rR5tfdaxl/Wflhp
8G7VT2MIWU01jg9K0tPLGGU9H7RLc9RvoqIU6MXWztoLc5Dhn9/xOA2fYZUtFJVe
RgvRYfwBa7J1OVF6v/ggYWtF+5GRx+b90kWFZG9AlwrRLKJkxccs7hp6Q4impV6G
qW4P4dFFQg3REAbRJFWj5mVT3wNrcwsg9O1ekifM6cwdB/Z7cBRf+QKVTfeoagNj
g36ZZnIENOZxlfZWBuq8pA2YpPKzgqWaqeyLyvDmxz7+LIfmg9xazCvy6sSeG+Hp
XKDoZG1/WN4M/bgM3wz22CWVnDv/H9fnc/sBEzr526jkEnDIUGMDGPz/MTOSmPgh
BRdhnvrVjoWsdGqRh0NxHW388OMKUW9eMWv7kFD+v0khJbktouEG3FcveTHjn/tH
C/rZF5YfXRJKEG8nACWv3mJ/6i8xXk+i8BbFhOBBTred6nzZAViLZRywjzRLdV1q
GXicTKKe2sc35x6e/AYNynqZMeEnfqb+gq4El2PKmnkOzGHD/kPcKtyw3qPLNavA
esl2jbq1vtQh9Ni/CotpxS2/qG90R61x3RX8mYL6RH2ovo3ijeuKr2IP4zhGdUP1
6soKEjz2tVtPtCS4geqGm0IZ2siH2QkGGDQyvTu7jh+QdcyrhQ7MztHHssN+5ZbW
AYR4Ze/tmvYr79cajrtWzSMvEq/JLu6X5KIKtdaUKgoTwlpeXwz30VnYaznMuFaQ
A75C7uiyI/wv2LTJ8gNMcpt7XGLPzCSEi202NAVYuiXvle+DhujgcBJbdPh3nQ+3
T8lNpKsEd+WntidY44KJnSYmW+Ke+LrFDgDlZ8/Q8+wkadMxndfpwAEfO2uzXzAF
B90wktCDDe4/t3sMOkiHqdCr2MdSSOMz35hC+Y2i61OljzPPxL35xYB2CZ4McrYY
Uq0DAF1qpgoNohaLdIuxJZCw6OYX6QIzdiQO53LruL14BM+U+KL4129qjamZ5WsV
8uPbhfgTwkw/1Amytm/CiMmVq5AFKPk2pdH9l6e4dtM1X4sZn/trH8HwjxXi8kNz
q/uiri9kgLKiey+wznl7Pki5+0fgm0r8cckUJns7Yyqv4KZ+JhXMD0gkskUGbtzq
83QDG6v+gr020HN43oteepe7k4pGpk/ixdZNr3hpl/ptQ/py8phAvHHH+jDqIxBc
wzuphRs850yTvi6r1ZwVwDTyvUD6TP6s/C+arkZRO53qe80ta8YlJD5h2xCMDz5Z
TFj9ijV9+xXqBP/FFEEczrybiuFPBqOH0nFtEGQeaF62ookC8LqQtlNt8qSNWs8D
TxGMpOs9u1VMzx9xm5B8N9pWi4XBnxtJ9pXGAqwESfrSNn50W4wunhCaEAuJeEhw
sB8GT7kv+m/8wX2hHKBZLV+u4dNIJnitvSAMmW3rvDCfkOh48db9AgfGEWTOJVs9
cBH2juO/UQpSmyyz5pLoU6w3uiED7Ovd5Ep1pvL4bLLfNvHUm8lb7bH0l4KyZct4
b+cq9ijnNmMku78h067FHqBjDjJoMXGH7K8QmvGXXoHyX++IYkZy02m7PbA5ZnHQ
xEA2KMN30sUI0AAdapX2o/qe7qh5shq7hd/bRxmpa3aL2WU8vqk7mlhOxYFGp6kO
XSJKQ7CZdozs2l7vCQmDtg0qDbGZYuvkFjVQKcyc8p4yol0rXnihVvG2DjlFmPO7
XMKd4mGBAZk61GVFNdq4KkBCUX2TE3wFVQMLIJ8GewBmuHKqDUvQ9NhBiOEIxXVz
ExNc9T7rhUe9HJY9PTXm1Y7f+74sTIy+6QmZuHHz6eRJ1iU4F18/lfW3Vh8Ygwbk
Vt695mY1dIyZArFIO0DyK47G37tJIaE4Adp56wamQdYAJJB0yT9JUf0h7wYzkuJZ
4CpGQPVorIoqRmN27bpS7h7p2GX/JNK118JB3p6wkNe30hnPN9jXSTvLMfTsgipa
IOmi7d+jCLEzd4e6wXUqlQfMI6gPKC5VuwvdA5yHTUcrVGYxQeoGj73uREuVIs6M
wwvlw30aVC+OcYzK4i81iHaWS8lh9i/6mOpLHk5hyVYzH3YLyjPpxG3OvBNn+y/8
ISPkeHhDOHtqumSiAIqK0TME5hMrNU1scliD9iVtumbgF+6eteWp9KZbx6ZsSO/7
gWIEvjPSX7JIOJfTbRTT8B/cgqX7hemYRxgaXkP7gHvXRlN5FV6EaBQLSvEI1YyN
UoQDhC5ePGHBp54uZNi2lZWSRpBn/SSFbcE4ClIQiT17Io/0j3SwNMnT08yJfNmM
zhtgb5cLF9NofzenIfRVY7F0C86TrBZ8lI+1e81Ij2x76QmNoIQVqvqC4X4R8+5y
ImZ0jzrx9o9L8MdpFkQ7KUnNusWjuKZ7wS2JC39lspxhQw/KTNT/Lb8MzFNxzw7D
RYc61h2fLdDDF6KVysQgixTnph4Xs3UTr2DFPCOg4z+jyOQftzvNE+5OL6FmvrQ1
dUFmZWREvuYmynLl9+3QYZrSvYzk3zowGjEMPIO4u0zLrjHnwdZqx2dvguLg0911
PkQcKrT5thvGW/z47czTr9Zvzj8zUok65f1GUO7GRXkdYDIwtEVylArlw75SO8bj
KVz2RjKfQgWXrb0n+hyhcfsI5xRZgCfuC6efk+guTZbcvbU3T+zIXQei0QAf8aZ5
xAairaEbaGw3+5U44Uo5fT7VWG8F/+FBLiUwks9DVVD9PPSksxcXkOu4cPyriPE7
O6yc1PfdjFnT5U2xxnnW9bG8aYh7yGxXaRxdQcLycExMo3MVltD0Qx7bOMDgTl4I
d/WFPn1ryq2h7/0gcN1IxDNDtaQ0NQko3UKL2kywl+1+xHkp1KURt7e7DKiKli/Y
gcfrTLYZ/PnlKvlxBl+egU0FveAvOKADo1OpQan9r7bZMPA9WdiYMv/JNYby9yV1
uzIEeZmmaBVNqlRkEPon4YdQXk7uU5UkNkfLlUIgTj4pCnrKUEovGrmcYBPob5ia
CsPNMYB6x6O4u8noCfa/cjqAfC2EdiVUpPJZTnh/SmAKqt37RB28/K9ObkVJUNMl
KVTWJGuRCXX8gv95tfbCqyao4vB4AoInA0ddG0+ZkE183Edepctv3t30u8LDC2jX
JpUARGzOQHakEGqeBB5g92ayRAa2Kf4M9XCgi60hj/pHyoCq+Ua+5U9z76C/Y1AR
WB1GhJI1HeJfgIeJrxiG5yELFIFdfkciv5zsJZkdF6JlR7//DI0kaX0nesjPxL8t
6A7WA5pWPZd4JPpkupzv2n0Fx51D/8rwTelJzPoDuKHGdojmlkq2rgG4TPvhy4k7
z4nedPY3Y24rYitRVME6eTTX9gU6oVyPBQJf1eUK3KDFQmyRNJunnfiQbrEr423Q
REsSi/ePJyYm4oB32VNlVo7Cqs92672RueyoBko90yZha87v6rBd1dDDX0xzvEpj
96+Bv4GiDISdCXJkOkbxyebA5VNggi1dHDd3rRuvf9ScFmyNh8BKf2bZSkdxRXzf
de2HwLBxPam9crqRQnvR+yFpSmfCIXa5zyswobIwSjTiSJG6DZvGNWh5YFjDB9j2
lUk+MYmrz83rnM4orhaNmg2rzUoxPF6+6VCSQelDESaeCngqrYGOO5P7YEVi7i4J
V/stiClW+jhU+aM6H3aAnLk1MHyD9Dd8Acp5IHBjmR2sAdulOavHvlHV70zGCtbr
UnHDdgYoLwkSzboasvZ3PFk9Ffk388GBKrnXYnjfLZ3u6rqAc4sMtq0/bu4cK5tv
rN491SkdgQdIYmo/Nt5AbYjQw0L0vb1vVx1eVO/ZBk1cROZvzCQX7rRfChTbEsPb
5TuhrGrbFwP+fI/N1fJ5eKKo0eYn3hE16XX0PM67larOndGr/TAcSFKUCZqmyEdX
uCtjw0CSrhYtSncJqnCTSo7Yidr+kR3S1A4G+S3fW3cik8t8smoyrtIvgP02xNFn
S4L6A425W6UdokuEJ4qyNVtFSsiW+CMd3dpx/6cmrWfV6m+vXP+rtyzUVezgK2tH
nHqvD3bPsxvLhz6AboaPzMV4OQRvFL68KpPAlL+hlc3M74lWOThVbFAVfg9J92JR
801CL2j3UHA5OYPDpotKsXNQfX64WcakVqvanP2vgEh2AU1806HjTHxlx89Zp/YL
YylCUo+BpXh1qCOTz2OArzhP4NcU0yDQpBRMVABbNKy/2M4FH8pm3GxL4gc4zA9z
dTGy/fhgDibdVQLoBPC6EFXYNAQOqgx57SR88qGyUYOuaWDheVnKLPwITa75kZ5p
RKctMESHXn9VMdy9/EwnTpa/lFJe+OtBF6l6MregWYF3FAREkRoPFySKQEqip3Pb
tz2An8tybn+Y+IeaM2nciq6OiFiwk9H9u7KtyMEUdGxLsiWkKn1DRRmUT/mijb+3
ZK170/ZZLCaxjkWbL0tLAawS6ql/bQtT4pSbnLcPoiFi4a4Cz3clXgGKF4n3CFv3
Q+P38PmqdML1umFmsMxVwFI8KgMEX48TGErkI84VZdwBVVNgY6e8w3jXUiJYgctY
rxoRUwt9IAjHZS/2l+8d74X+oFflTN8mFPguSmlWRI7rIswgAMMlKRclMeDUTujN
yWKOm1LfGUejaL9KtY6vRrzJepVMRIV+8HXUaQVg/nx92YBxkl8DBKxKR7miLqF2
t6nsGv9DaKCye7JdCMygU2VRCIjZc6lsZQ29VLqbuhfDz+VhBO2BMldwcbj4BgF9
A/CYwuY2H+Ye9DNPg7e9pAVgMaz69JNBzv8dDVO3dJhPhjaMoJnakhif3DBxyk96
fPFlupWDvnto8WG7pAsAgWBjBcK9YkFF1h3KnegbfqDOESBlCRLY9Jjg24Hcxq+9
U38rYKPvTcbjTphSQi35RBwPkvoIrD9Mb+bInF+ISW7tPWNtb8togWJ+dYxsMhRN
ZUBpqU6eGVaVtKI2ii+ISNfN2+HXctbhTrCZBCR8F6O+fhRjyIuPVg8RNnEw+4PL
80zpmj9GfDiCxdqCZa/o1+bvOUo8Q8ya66euu6OzmVhOUGqLE/iXPiHqqKl0XsS8
8C34bWl1GsqvLl2P/fQ8Gz8CJtpZzir8wfOUz8C9Ony8AiBmjvxmkLeJqKP81aHP
FTelxeCIIfFCqOUEciU31oJs4eg2LWj2KW/4e8KOR40lNX0iqrMR/eDx8GTCz0N2
1lSNhzK1ZOS672+tC+v0n3NyldZQj3u5W2oGOMsJf+4dBDukn0Kzc4TFtb4RED1d
I9E8c5B20VKoHcMi3oLRptSl5qT/rt1FOzd7q8C8+Pncy7U09MAlcF8myrFnKcSY
dFZ4p/hP0FX/+sLfr26V1fuJsM6bvzRGmgQEzK/nlkFv4WChYJS46eDV2Dtf0D9e
aEZJxRo4h77YuxU3pvMdfgmebOLSCKXd38m0DPEaQ+Dq/evfc4ZS6I5Tpj60BjRx
3H0dboOMBPBdL6cHPE3IQ6Vo2AsBchYzPELB12G4GecMmDCEK2Z3Lzq7Bf+mcmtY
2JUha+d0RgRzBIRBOQS7lKNr5ab5y0HCDgmTcCQlAHKtnFZpCKK3ACXsAkk1Ydyc
z41yWC6FGsdCyN7Q4zWMdPiLL5rab+7Z16jZb7bzVo60BUKo+FyEEfrDT6hH4AvM
oLbI7ZJVpZLeoxJylywbJz/WTm+5tIZxaJc8cxjjbXajJxex7Grp1o06USTbJrYx
AL2K3hhBV+f6P1wVUraisak2+W2qNOq/y6BtC820juAlbvyyl5tJ050FQZeNRNJc
AWWao2a7m1fuLzdWO0CIKpaAGIx43V1lL7wOUxys+Q9MrWZNB3y6bcrQTqZqIIak
xvcyr4Q+t7ztDN3XzTvysIeuC/8By63h0MZOGwwlu9Mf21b6/QxJOh3D6tH+LkYk
UAmzVNCsLjnFm8Clqt77UheZH6ryh5305bMr8ZVnhyeabXspU+atkVIUmMKC337I
luwsljYwXkEfeuVUSO2uzIcLE8pK3Dq9TcQ2MRLgsUh3tiQppWOOL+Z0pheVUDLP
XDO/LdRquCkiJgYmpjcv9xibSeilY+1m/YbKvNfLfzMDaCsGYzMguANLXaN/K6ms
W89u+HJ7NY2UvFXuQlHscNb0YaV4vWJv4t2Uf+esf7pycJAUBaZPstkHUu4TsPZX
dZxQ41Js2U40rx8rRJUtERPVW2nhkeFXfqPocndZ1y8j7nx6mDh5AYmj4ppbnZX9
qvNi0Wwlx9jqiOM2N6nE7ixpM8ziTumafP+lW+ZD7sZegeHb4dpFTGMbeiQnEJ1K
cfJ17INW9FweaOS9e6GZ5LSU6chU4qaqjnliz5LJ4SI9PuLOzEFNFaWxKBqzWd09
yMWP+K5odCEba5o3jkU2L4ybmAmVzZBf9hx5NQ3LYvfI9wN5hkod4B5lq7Ck9rio
efrPCrC2gG/nAOGuwXGZGQHL9T0/7DEAM0tgmVnJMPknQdfTjmp4qUQB7HMlr2AQ
/iDrDyC02xbBNVeXYKAK6DDJV29dLz0RuUcC1MMegMyExSCq0aNXuLKquEx7RCnm
aGvdC/9JemkG09B9jxAilE1EUHeWV8b0YXwI9TmCYK18TcAHgIL4tM/QnOK/0m62
WorA+8FpoFjEjuXGl1XcnECBaQk+6+ruXGp1LtJBQYyuebRT3BOXLoqvANV8FtCp
xLlZ3gEZYROJjyjiDSqAQN5Vr52DIz5ya9eSHaR2LpDckV2zyr8GtR3rNz8asPKD
bo6OnUq24+08bfVONlHYTlU9AX1ZgGWzRZt4OCNXpkY9SYAovEzQXGCZqBP9d1Vv
7oFJfxyJWb9PXONdcb+Ox+doVV6F0N+50bA12ZeeIfP/03KmrMKuRLZtu9h5PfYa
W3iI55OiyAI+AVc9VIRkMBYLXK/bl7JHI7c6ExPtD2ebPxsPGI2Jl/7sHvjGcr01
sn2IPfxVB1CuY/zuWIRB5vvoE0Y8CBk+TOiqrSAYX5s6GMmWa+AZberkkyLUO6TH
awmppYVjOd+6wHLS7ZvsC9Lyy9z/pLogzh993hKHezPdswh6p7UDlSOywloAl1V8
Ob+Jdekbv/CxuCLx5MQRHACtkGHrdrUc5t3p3KdDR/q5wWMl+Nuq6OAsNVCI9UQg
vDYLIm09JR8v06cUteYL/e6MyMpbR4KEgocXaQgkc//1D1dcn7v1naeN4fMiKyYr
39swrYwATC9B7uqbu4o9eL9ZVhIOmh3hFGmjt+qvppdO8yh+TnBpQ54B0K/+uv/R
vgz8xqKvCoyZ4pZ1LgTDHyu42wdBLVwR194DPjIIHgs7RL7WE2xO+nPSZ9JGVViB
aLdYZgBNmT2TyUtV/UhzpOxWdneEe451LTgshKJBhmp4n2HALeGYToyUoSa9EVxP
fukUPvU2pfs/dFQobRbq1QrwMqQbK/jhvwxtkWcBqULUcoJhfrHmFfSI8qar8/Tb
YnaTScER8cBGSKirdeuG77T0p+sbkOqMXx1oecqVKyKbRmn7g/PFpz3d3Y7BSSfq
8q0PHIEPCrrDphS8K9xf4aQ02Or7D0Sahfgr2E5N774WYLbrOWU3sJZWoSzzs01q
GUsnjJjB3dUlS5Myzuns6I7APEwAzy8fnfbb1yBWjjeshZ4QxecjkEBm3y2IJwlx
qhrFUjsSWFD9R4ZZAQ+PEdaeSjWFCTthkVRyT6iEdeE8ddYYzeLptwMlngfa0vc/
/uLpb8eVjqMjmGiPa5MQ9Bj9RM9+NmcdRRnsjUF5gtqoJjutTopuWEubM/f8436e
oiq+csnLD6GMgqlUCb37aX6sLNZS3rl9joSgoxzbGTF9XMOdiNav24pS/Anhg/Q6
a7M0jqXbuEKbkRxNPSiyr3SvySib9M5l1RK4nzgL+e2bI60mDjulvK7xWB58I8fK
YbKgGo9+yTt30YrqttJYH9CxItMbT3I4FfqBCFUJsBhOCDX6B1xTVwuMP/1cU115
gSwXz6RWG4ecQ6WxzNNPccqM1iBk7dcYdpQ9nxLGtSd7oKeTwgup0nW4kKxAp9+C
4ZS+oNZ661qCdTb0TRE2D8fhj2sNS8XpbNSXT9GTTxHmQwJdSdilLYK4XbvE7aov
6IKvDz1rOswQuwlCpJNq7u0jibh7qTUVBHaQLSTU6YRU4tg0ht6xwgz3TE/nR2GP
Vb1C3hjxSHFHLmiPc9cVNcDWWwix3fA066lGobzX1sXMoTHWaVr2wi4Zh7pfzOcq
10fFzW4JAlUJQbIubraPmcYZjnk/3FzRzX7QfrCBHpzcINjCU3wT1mLSuF4x2lDc
rj6XvynBgo3I4TRSjQTragAMiquwGGaVHMO6IkW5kkxdKNI+72mgc+ipmQSIxf/F
WiNLpFDZJvKQXW7KJc2NjAYwvqgXMqCdG/jlEpmYzssCWgOmc9XhfEEt70/ocPTe
IHQw64/8FNT5E2eF2O1UuziamKHgh6roWTxuBr2RPjD59JGRthgitct3DW1v6Nwa
ZqwA9ITEX1f105hHgZs6zrS9uP7QSdcojLS9hIojQl29zIqXAfrq9Jvz4uqiKuFf
cJCzJeLU9t88se0axNjZUw78xGXG7D7saGlVl7wKa+jvXhgb5wCnVQE0Pc20ZSWA
r/7gzMEzG+IMiDCF6p8jcR7NMW9IaoCq4NzU2bWrVgRCHS28rdbQ4Lm/hgENWyww
Ivk9er+5RWbBMaOHPzgK5ym2Ne616EaVpBOwBl45UZnt8rfhFOv+hplile5D8EG3
vt/GeHfEyVRqprG5WUsZitfjr4GUd8M2pGOwQnULXrw/Hr7mmmeTxp2dFGojgT43
TssM3viOVpgsrDcBhwqfganNyDAPsXY9FqWU6X70cjZ6JJJrndLeVZ3aF8DD/bZ2
33/SCfTVAiHam93ofP3VFafjIIJYtMzwON1Hq3OMPDf/QpZ5Wt0EYl7IiibjuAXK
ndTOjHn0xI0B9ekYA/N+KDPXH3sDTn337jeyyEZLDJG7CbdEdVgK1sp4Nwnql5SQ
d5v/9yCbyTG3ykpYBdsdWgK1Tv1Xk1LFw/iiL0HLscXD2AprvDPOVg+eZLdIMTNJ
QTfPqCIQXZfbw+RDOe14SPKSAtwfJXai8IGHI6HTtDYvQGjy+nrreJWtDqAo0488
XTe3iA52l7f8CCMO4YzlNM6unha9crGzco1N2GuJSCxLnNgOD91Y6c6Ad8sq6fYZ
JOQA06U9gBVQdg00oMxY7CgEG3RG5kA9g+fOlh0RPE5YJtUP+rUHL9MuvxBaKFVt
/DpYASOmJRHBy6vffJV5EBDqWnqW3ljCXW0ZVgw5KZsNLDa8QuI0bvz6/Gj6WwPr
aWMFJ7NIe54I+1Equ6r2RNRdzUqtdbOIeMyQxp34cAVqpcQ7MyI55aYoOqgMIF/M
WVyh2vC5UbqYFPZmKWTNixZvJ4iV2z+xKQUvhFFhQScZQHEUhShaRV6EK/mCcbgP
6hrT/6m57LJWgrr1Z072UZ7JkkDqTT0AdzrabQkpBBWA9fVmoiC+wS9bKLyAjgqn
9AqrZD4faD6ZJbpjN1yQPIFR/TkGJ91CNwSj3L+zl6kPRzMRbhFUlkLb2YUL7I2m
BfA0Lve5JXRPy1PG4sSDjH7GxqrSVE0+EtSYMgKhSoOvxn9IbXBneakr13Hcu53A
W1bDv5bsrCcYgOZCicszMpAV5zfsVv1hgZ+mpgG39Je+9QK0aNQc+Sh1oucJMDvO
7oemi6e7uhBe35fUoDkP7mcZhkHkyHEQ+HRrdvYcxP9HhKrxlT4CVrlAbA5S9F9m
IJ1VnD5uN9SY8COYSbNGwHqyYsmb8dJkIT5F5hJSRQe1pv7f4eZ5Pz8Zs23j+Y7b
kVCmRG3qVOMHtOWNfGgR0wq9sd5H1Uyr9kuqx1vA6h7K+VHpA/iTzUTXn5fTgGPl
qjH39o3q7NcrQZlVYQjo8mbpWmtNy9PyjUoo5/kPDHJu4l364+S6yIBm3IiinHyB
UxtmRgj7ht/hESqJ5Vfvy5APQofFCJEJUTo/VxrDe+Q34p7OJ1S/j/zPnN4nSURb
MbaIjFbwTMiyhfU1uwKBv/aGKvUnY5hvIYrOa3SRZGh6Y5MOo49xkMNBPt0GLKOB
UsHmCl6pNVPBvU0QKO5PVIrgNbvtNpUTl03EoxO8/Qn3o927eQQvyXuPNIhc28mv
u1m3S2vSZCOkQGqceNjyjS+ny2HfvDpqvlaPhGqKOsY0m6HJOWSrA6rWfsel6hta
bHf2HzOs3w6mEydaD8LlQq7xOZZzdL+nURg/OnJgw8rt4BHdfx2Ys6hcpoS68Zo/
mB6VmfzvJV7BZz8JrinRAYyd/RXx02ZVrS1pn/ynrXnttgvEb/DdWNFt9w8d51Uv
/rl8jvcEbj7UtZ2pmb5M77yD0HYgwbQv5wwBm8uX/u7c6GOwGLnPFxsWVC0M9xGo
DhP/jmuBbXCxvEhAjvmIpGsEqyBHKyPtL2ronA5MG29lgsUJLj/KnQiXiIRD1Qrw
nBnXXi/L8lwyniVHEXMItWO5/o/Dv7fXq69ox7GRh2R1i4ZEwpaz6pXdPidaax7Q
DUlnC6osoQRrKKI9Wga2B/axucLmrJ3q7s925W5+kwwl3tqOkfWJPuKIODdUQkix
ualWXMiK30Umz5nkmIQ6UEVKtINdMF76j3w2/7Se5mX4UDFQmqrsSs0WolMSX7tl
WU5CzDbHgdiZ7SQn/dkyHPK2obhG70Orm6LpGGAOKnuE4LSWzvsmZlhlcwJJkXv1
PI5FwQl37FbGqFwG7qniCOsrHbFdPN2jioqvyNHFt3NNRTVqEf/TNqz3vVj/eVQ+
vryG0uND1lN5WM/Jx2i56xkKZU0pWpEOAJFiaZ2JI091UBolkeD6dqlmeG7GHRYV
U6M78WvJpJoPeG7d5uLHeELktGt+wa2EbIVwWAtaLqc=

`pragma protect end_protected
