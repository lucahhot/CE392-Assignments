`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lHcAHQV/7WANURqaubpJpQZxLPYl6QkW+HoxiYdQK1YbJCnXrFPpbIpbBKp17VFJ
Gl54Y0RumW6M0khNV7aLe1sRDNOs/sD6Bi0EuICHCckxmNd+F7XC8QElEGYQQgDG
dNqXYYcUm5E6r0gGfSQ84fKxE06mb1I89Ik0ncXDpuM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6960)
vjOrR4pPDdSA/TbhdCLL2tmPTAqZl3CajaXQOmwYtAUuAUfGHxbcbbl+/YSG7ZWg
G+hr5UFd6U95BILxzpVajGjS7a3oJYfjD2vpWH7PzkBDErvHAwkbu8mo3QBenOVs
UyX74F1jOXTYKAP2fLthpbqvZhVJqBvpXMLsMseRzUo6T5m/94f+pmJ7u6nK6vzf
CGJno6yoQjI21PxiBnsQf7wMOthA+5WESe5FaXL5ABUysS1j8rbmHaVn0PJLTQjO
Wutvew6sMPF0jceAEXxOBU35nI41XHMhXBapkN3Po+oVPGM1zE0y7xV1jivaL3PA
pJ4BxSf9pVVee4Jiif7t/iwyRnILP0LEcKoaPdt5zLXcKAlIOkAjKvukSahi6jtw
JSr8aEcfJ0L/NWjdFDmkvbhlCm0b7XQUkK6KZ3WgTQLxdOjybMzqO0VaGN+rUV41
5M7AyFZ1dhbOToALqZ93RLfoEuJGb+hFAh1k7ZltmEdn6P8BiriLeUP0Tu/jGHa5
tgu1H+Q0WU34liJLsj0EwY2Wgm8TUtlg9HdYgt43vqIFmJW0j/f2eA3MLLb9bReq
TJ0LoA7f85XP106rEsbHCs9MFXOIG6qHcFkCShzbCLaFioEU0D/ACNwFHejXst3W
NG4CVVueX1qW5vkLmJEHL7Sa4OEjbXcvw0djGJM+OqqFffj5BAxLwXfD5OU+ApYA
q4j7frRNhATirSxwkGeGjbQuEZAimnZ337Iw9YhmbCDSCSi4SEAkigS+aejKRLGK
NJjjAjmJUQIzvFPijcS3j0LZuX5nQI/HmPS/d5WQ2V9nlNaqyuqlL5Dk1PJVXwog
IOyZ/bXJK2WG7yEqJAFEgQR2tfubTKIqjzSwa2aVDMbK8rmNtTcRzPwoTsS4rq4a
pSt92pi/jHewbe84lOpOgMD9E78AWW+Beqd23x67AlkY2fdSkSQNndGnRekCsa4T
5jDmDzUVyAGO9wv6gUlWDR1ZfmIx87I6AYtPbnHPyAiqLS9U57wtLHK2T0FV6nt9
QKaHExI5HVR/BkKc7xguw1yKdCI683M2MKGlOIvXwXvUt3JHgP6CP5Rj72u7Skgh
JkFW0QaMegTWfZ0PIoQHc3op7GznexFLkH9zMcbs+dXLTWDK6b0Lw3GHQaSPQS9I
rYZbKAvf2WtcLdt8kzfh7VQNZOhGtRYXKq7CnhdXDt8MT3FqizPzk9OiPj337VG/
Mnt+xjeiG+gPxPggM60pWsKj/zV6+/dPhc9cyaNY7kfsROeNPftZzkkNWvflPWzD
zEWpe57akBf1iokR7lfwAkXJ2Hf1ONJpBDEcSZyGoE7h9slWlci/HuD51CcWfI0A
UJMOmBqCnW2DysPIBJ0DXUXn18+pP6vigJ1AVVzKzbV/invIrBHT+3Med/rSmrWu
0jSobgsD0Vy5R8ikNvnTY5PT6jTGC5+Ph9N0qWGggu7d5KHz4avyoKyELWO576Yv
lZqyR8i09DJZQAcaQHqoO6f+1Lr+IiaY3AocH/AcIJojbpHiTzbZdWxdXuX6dBwH
YUJEWKKVLZq2rIqMEBWKGe6f/iW3Wcp4VhHgHnUsCl4CYnHRjG12yJL+lTB8F1T/
hXipd+cF7/SeJZSTMBCN2O+orwmHwgj+oTwqJa70QdNf6knWxMLFrJd/PsS4dXhX
gSQ13nWiMQG73u50tvtBxRpyrY4K/wITpCsQyCrlE597vTuHF2RiwS6ZQCtf87z2
mkNtjaYT3/ePT+tfrWY5/HrxlILVGhkBoPX8oBfINTFEHHFVne++eoF6oVGdmaJS
V5wjNuFeUi6S+/M0zGu93/Xus4pNGiGedWlsW3U+uXk8dO37DNkkpSLbMp94RjBb
+MBL3j2jgidL/izlXKldG8EWhCGrWTEeh28TOJ16NOxU1YnHDrQOuNidVzqag+VM
GaoeC7WCaE7OjG7zdZWSUi0pyV/1oMfG7j9xSKNudWep3hcx3iEbGptnm6EyG5Hx
gL/NduWKLYChYLe4m6s5j4Rvl2mIhq4i2B+HNCKBZTKwyp+KuAk821PgcqInrFHp
P/D93sQOn5fS4oiaWSxWPIL6B+qhWznoGKFEDbQZpE6ayqg3ykYOdesh/7nyVb6t
HCPKo62Nq5K5i49mX9dGe23Ix3Myg7e1A1Ln5BphTNoXTlshCTM/1lBNivCMq0lt
ZTDDj9EdhepG+ehRism+vZU0Rdn89c85FIWU3Oy0ucvIkQUBdEEyZlewKYgZkgXu
CjqADAKRrMXtmMyx/sQixnTsnavd2uXhCrfvnMhIosqySy0kjOQhlj/pHjHjvuk8
9n6vC0dYuJE5s/kMPughAyXQz7kL54Dfumi++pzXSOe5E7I751YomeWoq5VnEKeC
pjtDFpx12CD9H6GJwYJ5sfycJE/YOesnQxLPepGxtNgJHX5jCDPninElqjm456AZ
ydn8UzPW5c4reJHEZeAsXMESxkCcBV3OJ8OWYbuWkt2XqBqEFdvt44hHfLNtcMnD
q1N96j3c8OGMl4j4qcehqKYTj4n7TI7NrZot9eKhAeVqN863scv8wVyN60p3Rr4q
uPy+/EiWt3HhSzQaZgWJlpqsDgGGwF+u9ud8FwzM78dlvkH7CWZd+he4ma7R/t4D
BtzMsQVym96pTlp64HgZzNMvDwDVx3zq0V5sVkaH11qiERFoj0lvWp0I9guYge2u
bXUc7/ECYFwlbWJYYDmH9Bt3TN9QHYvg4fRxCHO1VDxtmlZ49V1VV3nyp4stomRR
mgas8wCynhf/vqGkss9IG4nFI0F69NFqvephEt91JUpx6VNU6QqQpF1SBjvUnMBR
o4WnJMcodYKMNMHGz6uCYeXU2/YGGZcM87e0aZpBopASWq15kKijMgWrUXRL6F+P
MWwEHP3L5yEDIeE8zi1q19WoJqehDG18djP8DvJ5XZxAYT8aEjOXDzrOgYX7P6G1
6m3uKKrDk3Qk7scNxqzbBrOjeH4CS+RHEGyxkRZc4Ap+iC1mB546ZqaTfKVcHyE3
J/SwPIpZukBYa4dtKMDao+ybUKR4jDF2DSBTBMgCAPNfqXHfGsJvdY6tx7l1Jmu1
ANnI7MrCOdz4EqcDE7fzJaBBfskNZRiSiT49EGnFDBttuUy32yqA8Hre2OxuAlmv
U2phoklgxmlpTtCBCnRLSH+vu7GuPsPNdi+QLcAumfCeb23nHlO7aQWQj1XyWFIO
BlY5Lf519+tSe2jlmZzKNK8VYAB9ri1WBZklon2Dr+Zp8SLyXzC4lHLuKcSZcUdM
H1M5TuT8U/K7QBAO03I6M5sjSmUqoLBl88EPMLHf9I9pHE27aIQisiW5kEUgO+iM
27Ww7Lw1srUUwXytCXYKoRwCX4h6hh5IZGMOsmHa6cMUJQxIkeiyNUgq2nZDEAAz
f5aIHCVZOyEVnlFwsOI9ZvZDhqehsuhqio/Yx+yp8pFJ61YP9oyzu3sG5YN70Eh2
ulydrLABQsiI/psXMwYrcyOY/BUN7GdHBe8CH2ENjVbGq8JHrta3Z4CT/byfXMtc
w0dDCEyiElUItOT+7QjfecWmvVBvt2Xe06csbTYz2+A4HkWB67RGKE2aOfOVwVII
FasYvdzjYfVNOIbmMQiCbMEjKSSwfSTEu7ihI1SPP5vJKjzaHiAUODMzRhLa2nGU
S2HFkjoibQAI92fh3hF+MeHnFRb7PXAWPDB+/2c2V/2+yqirg5Sp8iM+jFSqcVj6
omkUQDSsL7hw4A19mjxXQX9B6GdUgWcim6Inh92ow+wPKIqwbitS5K9NIRi2lbOS
JqOjTKdGjyglx4Cn3+rzth44CH8f4UJimYl6jP0Ju4jWGs3aQ/WETafI2HxA6AwN
DBAs4b1+i3KSKImjP/9SKanjEAcajup5KytPGV+HxnibCAs5Yl+LejK+G7C4JZ/G
WrL6nkBy7pr2JCw4K1UXWAk0/9dzZqZmWUGGdSdpEIQU6oX5NAdrfnEXcoOhU7rZ
8sVPQqFjxFwmVhZVamCkymLDo8mc3tdt3+5Wqfbgwa8X6MyDzOmLAIhSe5JGBneE
N/gTR9CcImk7xApfwEb6yJRP67QwBiLNHaF9H/qsy9U9VQtlzjL+wfnnwiN8ecM1
zO2MlAtOfVrmF2ML6+jQPaai7tyZp7GDPwwcujOZNKaDz24uBUxhEmfh3cVgY0Hw
gE2H76ef6DQo7NjncPGgFSVSCOPFOubQm8UUcTCAg92YExpRKw1zQfMghUIIfAWB
l/r9/1Re4E+dTF6upZu4Ow3Ds11CPoiT7fz8l6eUTEJHoADFiunObov5yddnvElX
RZvrIU+Cdw05ihd06k8jsk2HOmSe2jDZiCBVT6Ut2V8CjyOdz60VO6tdSV1wVV6y
7R0d/5jPHnT7RFnNn3nqHrEdO4hIDqnsXL1rNYkujmgrcNRn2CbTqD3x+qRABee6
eHEJB0nFEXdlQh01t/yNfiUO/ZzmhAXfyuP0SWohD/VNMrw4smB94959fUJnRuef
qOdyoK6yJiOla5LN0kEszhBLi2WjzpIyv3QWt+7Y6dpSstkk1WQMh/lXR0fwM9Uy
Da5BTYJEllZjzPNI99Pal5fyc3Qe3JAi8Wln9QHHHgonHwIA5C51eYLP/pEbIPv1
+eeqAwTJiy3G6KMDiSNMvJG1YmMUbAYiRIXGpHZJd25dms1H1MK+itrfT1cR2TQG
aAPHNGdrwXPH/3U6pb6k31WNchVfUhjPDDo64Gu1QdYfldga+/xiTdNVM32SqqIN
TgmD7XoaYmjcGa3yHEQS1ZNaeL7ZUdyuFEIDECfS34weyF5NTVogbhbr6SlvVD/9
iB8+OZKed5lz1fuPPknyzi/1Qcxn8qfxsYPHnALlCo9+bhmtNRDW2mj+2bfrrHus
7qk9TxtIAeZE9FHWi4xUUzMI6g/Ga0gZZfcMQxG6owTyxT+xdg5nrAPuby72QZ6z
vQ3iZaEs8oe0OU7cszZQT1h8pX9m9PUg4XMPOaqgOkcqoUyqMliOsgvuJZWjiOt8
y/mTsDx1m/D3pqzgpN4shRbLkygazfWFbIPYECQn6/CtFuaxTgBW3EpOI+vY7UxC
LdZfgsaHTXXI7hWLm4OVno8yFM8cThmb/2mafZQ3NRKQQS4yz5QSOThD5TU/q3nQ
ghXjLnQll0NC7EJLzEdT7y1IFD0fPXFWw7oqFwl24HTolEXwpm4SuU5WrACbPRVd
ihVPqQAftfxAelQkpoSWyBpUvI737E4U/oZAPCB5RpyIhhx6xYy+/sslzLhs1WXM
IFI/xWlxpym8bFy0jL5tbtvvc4DcnwKHE/GvRf7xpJxRx7D7ScDVGmnv5do6/YGf
q2jh/Imq4R+9PY+9uyBQyjAjtxj9/r0OCo37erI/O8Z99gK/3t/RHbMeXPvA8nRK
bql0eYgAkpqHhkbJcYaAYaAOX5R42NJYWINcHnoGN9xmt9GsjKLOgnLA7107kJM4
gsiWuPveEzxkMM2IhG57GWcOwhqMPAkkFZlBE5tx1fSGPUYv7BB1iyUut/Wbr/rj
GvxApBVvTTs7RZHaz1+7i7J2HIQvdOiwTSQdIdUG5FzYFRYahv1DKe1EzzR2d75Z
2J1UcQ1bMd5Ba8+z++WfPGPiFCE6yrLWypB0eesvf8EeVlmx17muAyB6f28sL1om
lHK+rAwyU7yWl8kCwwhTCZtsKEyzIeF2VJdobQaPFz9HuFxtMwHAaHuTqEjBRTjl
kEEMwDxUVXjeTV93AVpP5KkxZ4TiBnMMJQO0Fe6e7lzLKBrHoST6A7PaMUhnnqCw
IMU+SnbksUJ+sa69VXMlE5izP7C765RPtz+g+W2C3rk0YN7YmBsKnUq6309Ad9Qf
dBFjW/lQpDLrgdFzcXqn1MoRCBYAT8b0+SgE9NU2f1YBsh8GcUEUCi77MlMYy911
eGyRIE1BGAThcaP7d3HyfOuPewR/NmFNU/5k6OTYkX3DDy15rFtO601FlAAo42Bc
JDHX/DimWHkZ5aVhai98FmMGxQiMHO0dQIu24HNXlsS5nt8esj84qCxOJOjLwiAI
jByaGG3XvVvJPXzVvIwVWUBGSRnmOyiB1ZziMRANLOs6Xqrbjj30UubTiFkvEuCz
0lHBz5k5wjt6C1gUU95tQhE+xwZlLNWqI4wQ//IayEKQCtD/yWUiyHIV4zVdFDkk
Rrzi847dg3l7nWEzIRAg1JBqWIg6OKcbHi6yAAxA7Y/bz5/bVlMbFbxoLn1EM0Hu
k5ZfQraxgExk5Ab8UYUh813EMId4v3ToPVoEYhZmCn6EaIlyR4PeNH6Rt0ioKR1T
5Erg2y1uP0kvR3TE5BYv7Gl1n/NyaZyRtnYIMVZXwj/ffC0yyerNEefBdBXPKUtR
dxeoAZP+PNNvZ8RnLIiciHpDJv+A7fKJ36+oh0BgJJSCMQ78jVer56xj40xailDq
L6rY5JIaCUmDMAb1pnMvekMGgp7JpxTuN6YZ3gsClXRhU8UWOTCqIkUGvmr+Lt9O
p0vYyOedjccdNgDm/jAwayAD67FyTWXAkBdH9Ex/VzQU6PLO3Zqq64uw5QPLsj8/
1hmDRrHkYSIuiciCJHDebqk/xVTktbOyfZJU5dq7d+kOwzL10cekmsQXG6mR2xZb
duMLNfuZpY9RfLgoBikoagUc67QEl2I2sVHFZ9ViWwJ9CuBe23w/Udli4EFxqeGO
lliRzeo6mdfYjW19oV7IGlB6EFAdr1sU2XkZI9NknF3uyfk/bFBk6OiGLI1MtqG/
8Ljnlz4eQ551ySUBWcl4X+UnPwLMx0KDz39j0sWK5zh3MMpArf68gDTNub+6wy3O
wlwqY5eA6UKFC5ZqFB9GZn/hC20AMuXrTs0oxAKOHYJiwtPxCuyL8rVxFN9l9JAL
O5Tfwyy+XAYLQkvnTMddUmkZ5xQtLvD1c8e60iUIK4VSnPDPgNYvY3s82PsOMwr/
A3YjtgiOKGdgr6h+lVtorO/ecBgXfU2+L3HYUteirDKXtQ4bA+heizyp4AcyJRVE
LXyFhXjYTzG/I8irnLIqsxF3ddJDrzhusKw1m3RwM72LLEhZRQJoYRPL3GMlTHnd
/rvzl0fPEoZGKZ/K9A/KfwmM7ToknZ7rby3NZGZ9DMXOFCOqb3m5VVZM0JTDGvZl
n+SgLIP82BtXHOvQQLO0z9Z0Nba5QC3T90T5o40ctMsixT3X7qGBnPJvfKSax7J8
1F/ppHAA+dtUHehJ2d3oZfAFpdy0h3TcnLs8KkbIqhGCKk/2Jiz3F1NqFbdFbN6W
7ZMszDCxvBElGbpX+xBwOmXd8JJWXKSlkN03x2po3kWU2mdcdxcWELFfOzMhz6EH
AB60KNPMVnbMAiZ8DkCtDbbDvmtq0WBO132Bl5VLfUkPH0/z2s3LmCy9JhROELiF
23dH5+0Y/wcxp/pYrsLEC7RcPYLcFpLOYCWOkhZxWgUUWIf1R4W5JfRAHsaVk/Nf
H9XQkNKTIfpLylbwTBf+bP3RdAI/gI57jZJbXjY/A8qqIYFR2TgJKKKFppA90MG0
Wj3oWkFVpdM8ZMmy53hf2NV51Zrc+Wv28wffSS18/JcNM2ykVt0DAmowNEzRFNw2
aFKPONDhTjhgAvsflAqTi92kIW+C6pFP8EyojfbYLUrb9lEmz6ZZzdFoqOOsF5sX
BeJcbd1smzsjkYbZSmWqPy1EADkzpne9ZJJH3kfowiJjdHW22lXd5LLYqtu4ET5T
bPwWS8VD2KWM1BngwEiKWcxwq6YyuaC5JK+rulvTjPtI/+hBLoVie9UgTmJYS5Sv
NoBGa8Tpnmr3mgvIsFN2CYYUW/MjJ0dRLoZE/2g2M4GCr9kYjZTRIFuiOLJiIvos
OMo1cMCTSVqWS8ts8zpcDndwIR4vsjM1YHQVkOFiGmFZJLpGrw8roFkYXdcmcMd+
4eGmwcJ5Dzv0dCjvtp0Us3pImR3+R9EsSOQNjVKbny4xzXG2xmxSDCiIbgNDVGME
63t/V4KAX85j6zKCddYnFMkVAQpKMfsfx8kd8WP5F3yNvi3POknCgZ7FVbW72WRT
rBEbU271Yl35mSMzX/vT7vwb/OEVzwXsr1TylRB024MuvuOLRUv6k9Gpd9QEplZL
jRnnoGG92tXrM3PFGJrHnCUQtntuuqnEcABfkF5V0DmYbN8N0hmlCEXtsR3nJW4q
eOtvIyEGiQpJ3PXbKzaIp0/q89BUOH98GABVOfMHfr+R3ahF+FrfDnFC3P58mFir
jnTOvC/RO4LUa65IMC0fEsDQgL5Hb9jmoOI85rLqxk+l8iV7XGWHu1cdQEH0JPD/
5qr/qRQJCRj1nw9DpNXInbr9hm3nF5KQDsq0dXleK9D3VLrB8hMh5XmIzPxPJvc9
VYm9VBopjq+p87gN1ByHxuL7c75UrYS8KHRhPuDY8CvyjIjbZMP9onBsOzSb7a2j
tpm2oujzhdTWRWrd5dUANYtvJQ4ZPPJak60QPC/AcIU788lsATMnB65i/0UyB+iz
IVYm4ochLJgFibZrUL6q5Uneqa8FXPhK/7PEvx2VPKasK4ZFAKCIb0d0TayiLQMM
WHk6/wNgpL8gt1eW1CiEvX/2tsxgzGhe6eZsJiKHkE8+FxnMOuXRtBK8VyGBZAP+
uanxRcNj6ZxfhMfrqduBDVoxX6SRwGLno5PzyIPW3EiVbiwY3flqoCLsZo14ZT94
LCLroOym3dv+0on6ILW044/EwSfdJDfYb1ABwNUe6FBzeM0h9UUFGYLr+vk60Zse
Ox+32vvyuPy52plfcephxPcIPxsD9358i6GkitTRQYwFwWHQ0DecpQo3mtEu/20Z
TDvpzjDYkcoME1QjO/eb/3oyVlUNBRxg84q4WVpACZV5NB+7jQgAHOoIBiEK9TmK
6nSCtuNnn4+cGCLd4nTIapmeIr7DYv7ALdaLvZGF3vDoCRNNazwOUltsHX84k9ew
4LE2VT00Nh456rDejCigRClCvJhhc1dkvvWznS1ag5LWoH68FuTJv8i+4BHjxFzp
tYekdhriP6dECblz57G6vmKVf+tB4ma8T6RQUrIZPJn+mygbksRFEgSMyK+zY1BP
+S+Awwng92ci9eVkiNzo+7wSFaDLkUT5kCQ+p+sMBe0Hf32Gntd0iFHeP/fn0fFh
gSC6J8gZTgpep4Aheov6La9Bz1UjsEw7uRw4ZbQyZCAGWL5Vam8w2+3IqDeBQE3n
qLstD70c6VjTC7pN0UHcl+QChCG7n0tkIbEHIFHmezwPChJAw6f4VeY9qA7PG12/
zTR26iY0U5H2Ec3CF0e3fMs0walfRC6T0OHZOsSXEBdFO5phChtu5005fFdCaVS3
`pragma protect end_protected
