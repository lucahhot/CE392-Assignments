��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�a�ȝ똞ݪDQ�Y�I>F��Ѕl��=���v�	՟�l�(u8������O�Y|'䰪W�b�c�2��/k���� ����s�����k{��]��2+%	�sR�����<�r&L[����9���i=!���	E�(����<X��S�"bQ�L2�� ��{�G��C��7׺:*?�(fX�2�fL�ˠn.�m�^3���î��oP����_��A��G�� �����c-p�!�h�=�I9Cǚ�o0���	�
L0"���aL,xE|�0�S�^'�lE����
�7\����nD�2ǎMm��v,���>�!�������Dg���$(�Af���ַU�Ir�d1P�tա{��~L �]P��<y�+fk��]�_�I�d*��KS���ޏ����8Q=+�2�v��2�G��v����_��dԓm�Ѿh������ p�佛O�}�l��EPp�+�U���eM�'��(��u`
��^��}�<�C6��&��q��'4X����ޓ�/6�%�\��g ƣg�D}{r��I�T�t�G��!7s�Z��;���FM�e�/��Rc)��OlXPe C�"�$�K �Ә�+�v�<�Y�_��@Nh���;��e�I�.��jfo��RS��& zH��x4+|��d�Q���30g��Շ?&�\C%���W�za�Lul�{�ѿ�GI͎��W}�zƺ�g��K��P��#$/���~�ƚ�>mCܞA�+���0i/ny/�n�03�x�U���a�|6���rI����3]卡���~�F �:�����׹�n�*g��1�o�����&5�ɶ�yVy�����z�Z�&n��,&�%��{�HeӨ�؃r�p�ߪH���@���lo+c�&���2ʩ��N�Ή�ki*)*�ɔ-�=�E�f1SUd�V��٤���~h��v�6�P	+�Q��4�"��C���O��N��2�qE�"�^k����N�1�a~���x���R"eS���)̔:�����PJQ�Ĩ��P���?ON@a�� ��f��?De�Q��}��؎���,�R��ʖ���`e#�ۻ��!�ʐ��ǃm�W~*��\58�����:�C��Z(0�1ވsA�O8�Zݯ:�b̐D��F��\?EGҲ�$K���O��W�5|`�0%�ޙvaB{q�|�]���f���R����F���ǂ�-&����~D1?����q{�Ѫ{�C���a�ߪ���+Ӳ`�t���pjJx�YP?����⤾z�r[�H�B�Q,�%���^�h����`�Y��l8}9�n�JVT��9�A\4��$|��?��Է1`~��1[pd+&
���㠋�����p_�M떽=�\�>k�ɚ�e��ױ�`�gm
Cz���d-[p����Gޒ��w�^oL2~�c����'춿��Нgt��KG�������}�W$�#��� Ny��e�bD�S�'�N���%��Ȑf6���,�r쌔��a����e`m�|�j�s��L��7O����N�8�JV0ɟ[ن@W���K��k�&����F�`��ku�ݖ���w�F6��
g�܌3!� 2�C"�~�q؄��9�x�����"�����x�~���>��wv�U��jO��m�L��@������W�(0iȚ!e ;�?��C����
3�V[*���. :mR��:=}��� ���|sf�֚����|��+��c�a���P1F�(3��K֤T�>M�w,��鯯'��=���r��� ��+� ���'�s���x���/��jƌ*"��`��|�E}���П..Nm�ͺ9u�Z���׹�O�8�lg�}h�6e�'q-���[�ߓ��y��dPر_���wy,�FA���8�|��=rp��۵|]ّ���]Wr�K`Y�^te��X�a�VnY���2�T���1��Q��Lu�Ӿf�]����K�{�ǯ3�]蕡���^�#?�.|"r���>tOn01!
��%͊��R�ɇ�s.R�ֲh�z���ec�A�.X���A-���X&��Nr٤sP�S��x�ޗa]�whQ�#�����E#'%��1c�G��j�N���V����Υ�IO��4��N 1��
�=�Ga��_�v��XLj���l_G�9�w����{����jP[�]��md�$a���p��ӱd���8[�Y+,�j���'�����L(d�E�ov�&���1WC\eڠ1