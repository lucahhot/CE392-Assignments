// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
PXkqLE9AyKJ3DhTpe2PhXaWgUj15iQxsc3yzTG3EwY+JUEPTzE3xmyXoGSZWSK6SAVgvSpMsgY2s
/S9GeHEwWd2wwEaROxIWjOxJ7wPjDdMbcR7y2g1nFjE7gQ5wHx8aRuXgkNacmK1/odESi+PqKvNT
Xgv7l2pcu+2ySMQlGPlm+LC9ghAa/W8z+4PYvaR2yaZlmKsgdcFzaHh6JpGFHQGIuJAIeas4goV7
KFkedUta1jIv6kKTFgtmZijtdMxt3y7353ltXV3ooyGkqSfzseKrU3qz/bSrQJuLAmtFK73ZqJRg
u/Xce7xNPA75GA0Ud4tl2GxJ6jcPBnwvXx0QQg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 35408)
cDz1zXTDtiBVknBdi8t024zUBHX6YeynXomZeWZxt07QJHspBZ8t5QNaUDNMIrV7NE3YIAY6EeeL
I2MeADR4WqvXibKkEZkBCW+iNE/T9amcNnJcs54UKrjvAcoqbF3HJVCMnv0MQwfS0k6G5caSD6uw
7M0Pyh4vFJVJjvu9u7fOxOYS9t/64yzfSgiYmka9XqG5fN/DJVSO5G1VISsRznLXD6kvE8JGs0pF
aEPHA5C1vHFbMmu4lL20G6sdjHdhShKV2aimj0w2ktASsH9ZYDAs1DYO+cUjOx51AJEBRwKhafh/
VC56d0rxoJffRcz+ufE8Ez9OsPj+YcXru9Fq4/aegENdO+11aCKLExfplQGT5jKPlozItSUWVmAS
dfo9pcZh1zDnVRfl2zeWj3PNwIKo/jnG2Yl946JH4qC8CSa3Ez8LNyBZhVyU401ObDb5NmAzvSwv
MD47SjjQmDZSdejXQ0jOx9DuuJMWuXI3+9rjuEQrZBXVZcePUWDyUa0VIqCihH4pPLc5NNl2dT7Y
O2AsQpkZnhp/Vx7UEKz3LDqEnGvO+VhVcA97pONLLNEQihKLCoWE05fYRt1e2hNp7UqN3W147IX3
CmXbfQk3kLgvlf5y3VPVSetGJjhRfC1f2SPLTKI13Cu2xJyLEz6nXHkJUw8sqzYB/DAyWcv5QI7m
/B81pm+dlBmbF3RrVsm1kaCGqA74Pnr1wNG9gTc0ZawpckfZwdkVSFZvNRq1tw6j0jKuh67x3bAi
T9IZ+IeswRf9azOaiqdu0Ac2JAmeadB6extzujk+srtteP6rE2SxbVly6wlB2UA8ssrELiymoAqM
C5cNhkAXEwcpJGetrHhvS50fvg4tFZqm1+l+HAma/wuJLODVJv012LWO5BHyQw+7wUGBmZmIrcx4
IeBRaypu8Q34m3hUqDzp8Ue3bNheNbjjzbQfYobYaUpE0arPdRIebU667UghEgTby+geV7tYiEEK
ex1jWdhFaUz233MThKYJZwM1AKJnqfDd9MXTTpai49ZAJJsPfRoD6tP8yOEGZT5lI8UijKDm0M4p
9GKq9JaQDq1BuEivn4LU0t+S658E1ZgYikqzbqiUi0FUdy+W02CAjnEqbL4USlcd7tULTz4SBj8J
rva0pcl2RY0Rw+QX5UL1IhRSgjXE2AdLU2y5cqpxFPNcIDfVMU+jkz2wqiKJzidaZ5uOV4W/efuD
4zXYyxafDCIAH4kx2r+wSCyiTzj1zmefT5VpGy9B8g5Ni1YTj4H5z6Mi0ztLxlr1QIYV2+GnHA7z
sJDUocxyJUiHLtoQf1YcVrTjKLlQi/ibfN1jQXCfskDzeGwQIAxHkfRv+cexfL9ptjgC2ZxsrAST
v12dreQRxaZQclxu28Av7J/yrMz7DMwQa50djwB78VViu/Oj3Fp3KMPWtamG2PhQ451rKGA1gN3B
prLKjjFNsJiqb5M/aqCRob9lO6V3xiJrKzWx8JpHtEWeQe3+ddg8jOGZ6c8HtQ74PQUKY/bfGSkU
1TdcrnuN0Rn0VjT4swOcDhY11zeSRiyDCpy7t85CrDLy6d0kJlNssosX6qaLtsfasNYtMFgHyvPc
SB87XUaf+eZmPnGMHVNJfb+Jq9IC3tGPmQgrVym743jq5B0tVzZUizVixwL/paaqwOVPKKOdTroG
mJQojItzVFN/p0hqopxOadiCoGDJ1bgrpfU+NmEI+RuXXaTrIDhYbzJyCBMEYUsMR+27p4Y+bQXb
zdYZnsPaINtDihF+Sk3alZyhAszWbRI5Vb6QTskt+H4AVKBXWk3Nzz2QXTb7+nXLraVs4CuU0mYS
twIhLsudxBR7YUNgilwJB17wrIheQigBpM8Z1sLKznKiaPMGtN8o/4egUk4nfBPigWa3MP5RnJwf
SPrVAtk90uFeB+FXjAj1daO1m6FF1+5xDDk/SZ4KPSdPKH6nKNkkYqQOdADb3heoS1vu7bwStaZU
STSvADEOEfinDf1wtSA9wtRKuRsRpCDKHwfPlaGQreXGaLAA4Ji3/+qYnwO3qIC596/ixk5iBVsM
etDS/n9jHjmuhrXKEd4h98ceHQa3C/dzZmmY8g+2mV5A44CrAmAOdu/8nj4lEIDAsqxnuuVE6ctL
W9B8C0ebMWDRq5iMqXfeydgcAuZtmKU7JUPMUfyWT6NlgkbXZeVWupsRZI7gDzSwDsHEfafl68je
456zWNcB9Di5bAjgPEOOxynvOqhIBdS+II+sw5qpydrDKrWGQmxG3Q8sW9osRWImzvz4v1fT6FM6
aHsEWBZ8MjWEa1M21vv34Z75plgaynP2PW1bkHHgzdqds3WpVUH8tTcLRFY+b9fB3r3thCiVLnwF
6hljP/2xq2uai+ANrS9V36nU5qVQ6vFvz7lPl2M4NrozwM/rnruf2GeuVSYFNSXqRi/X96CuLG81
geQ1HBGfy3+sMjhoDxPjM1tDo84AhmYlaLWIjHFKzyo71iNRmxaDfC/3YsD5klNFBpzBV1Ugd4OH
eJtXnW41DRA9GuKzlIJUJvssuGuc6uwUjmT/I4hi03Y8zsdj10TD+3Y8Wx3ntaC1uyhEfgAAudlP
nxPYHOE85IvjveoaXf7FwEwMZwJN/AlmBvlFOZCUwl3ixwTfriAqqufvHiqIEwv890bpwhmSU1zC
gpNj3lNNsDVjThXRP+lA7Hd4C9x15/bkAIA0aveIHDKDV8dd24PVi/ks/VEoBOlAD6UtxBlTHb9m
OHLx+THnACu6r1VQhlflg72IT6GDq+XvCjhr0R332RcsEBX5JlpvXrJTN6i57cfTvPm3OQptitRZ
O3sGrPEqA6hCWhe5liBRNWLvaJbVFHHLoU+Q2T8rc/5B/WM9ILRLMwsrtelAiFIQnIa6ukzwTEzO
o9BnjriB2XZ1wx6X9H/7VCM71ZxK5R77EoIo62b2btbMT2sTdyWXghFi7gMshkTHonsZm6gAYkGk
Yx7Zx5f8nN/D3eUqilDfW5xaw1WnQ1+11UbmfwQex410LKS+YNlu7rLn1j0frHJwau4oGJ4dqUN1
h/qpErgnhe0/qhtbBzdZgf3+u8szt4nfMveNM7TtgpQvZONLN3h7wbxbKttsWYah2bCjZX7ODs6k
tptK7DvodNK3RjG5HVHIK9dlqgj/yOnf/598WmAAQyoXmeha0uZxnjlexTe3vQ7v6n/UyCLzne7D
+dc2idrL0r3plNKGnssANEhj09xUC0B3PI6lh4WlTpuR8YqnViaChTMSU7SK0yWWbP1z/28QpSNh
pGYpFZAOPjfPNyhcKZN8ghEdARjbaJbnXlDwD3QLUK2Rn+K3VygGjRTAmzxLqC8Ix9YTBybAaAP4
echZrAuOcus2uefV+a5xgKvIcj94YvdIMRwsrXyDaknGQNXvtHnDYEbF0a96oqAZ9iiwNiwPm/F4
EUUMsKw9GfUp1gIPam6CNNrZ8kuu+sCYhfNyMfLUdtYTAjtocxaMOPly0oUDQHWyzgAsYfmgHo5W
f1OO7qCpMp8cLFbOT3XINqzWS5/UIC+1CVFKBpKVwbvJeIOEohtOiEkv9DDLgSA0Y7s9PbWfCrwh
OjVY6l7MnGMWDiuGSY8wOSUpmY0puEEZRdxhLM0EwfPs+/5BXCd0sHPtDys2Jab4eLlFd8tKNr1S
/H7W9lCXH6fXfaomYdMErQHyYmvOYveED0XQDot0lRBR+wafKOid3Egrq8loT/TFs4q5GslqdR0h
Hzb6LnaFCjGG1rvZhvFIovRwBXlo4fFPJbfQNSOa56ayl0flvQj4NzSiQzJTUYuYhMwq2xZ4UUBL
lLhRJhW8iQuVE+xvrdCTxZ/clQtbZ6G1KbN6pZLlH/GymIklZGPa610zhroZ2BcwVmClRHux40Ot
/GRFe38LYWk9l8RnSU59IVp41Ww6S9BFCH0l1k+qfdQheM9ZCjc2VyySeoodfvMKs3dWLc0zjoQE
/2bafGkr8w7z0Pvqh3nVckKnYG37tM0kJsTBo2oyOAW9VZCRkCIEzdImDWjchY9uVb4uzJIjZCBp
mvEQYp6aY06ZvH1HUwaHyNPHPlxfsIBWlJtUX0e3v/jS6YvlC0bTwMojlkHLRsIBDKie3vk1CkQd
n0IuaujQYFku3JSZiBiKqY92wVJGHZfj19TbuQIKkylNI2+WYLQ6aDfDNWtTioBMdyreg9F0eQU7
pY6LQF58kY2rtr6DYl3qvuu94VwhhE0D9JeE+3mZ6ZGQQKf3PFf01XhvHxNnHR6KETSO56PxrwiZ
nTEi4aKLzU+FR/vST4nwtDAd4N3KxUO6g16x8rVP06cyrlNEX7eJVv5c/+d9USm67DRnugUnmB4B
oyKxK48W2aMLsVkf319/v9YvdA5BLrcKUFNIqOGheVKbe7O9D8H987njZln5qYu3p2EWZLoaf2yj
bHNygJ+IgPF+3Z0qoNB5i2RbnwaMdLGC8D70veL3utWFYPWXCUjSB95TwEf2/KP3J5aErzjb0Uup
CUN4ap12630Qs3Del/gZR6uT5EMjV+o/8rjyYPRvOFJUET6q8VfzPvtuVJIvG2IlQwygB7HHMfG4
F5+oVj6xU8zTOX/EYUlrB6dwYX+h0sioQadrlEs/6MWeK9THNihHvYCWUCWojpRMrTPjqkLps8os
j9jKQsMlCNihZxlDWztVYQG0NCEL+MFGj9cF0JSGwKR1+fSvMpP/OEXqSihTjCUPzkuZ8hisNNdG
Ipq9XBZ/az3oC5BOX8Z0SWvxWT3Jkt6DgCdYvTTaGf1j8L+Es/5elAhuguXYyBX7gt0BDSpSTlS8
IFAQUzR/fzohkD5t+MMh3otDJ4HeOWI07m7VZCjhBEq1gXSw9fYkIh4/FGzjgsHkZ7ZwTupLhvZ+
OaLWGtRy4k6+aRN4sVuAOMhjWJve0FPYrIpKaZMdS6Ted1CVwwBjUbIRWYYDUhhiKQcccN1MkqKx
2Uc/sHKIc5Gp4fxo0zmsA0ACH4ReuVYHENE9EfpH7V6/ktq62K4O8SOxAo/lTYHeT0+K+G3h+fwj
3XnRmR3BS4CAN3KnJbDzqbhBrp/zXJWc4NQ/WqZL3TY4oT0UqJmYuHUiHUw/tJ6BanvQQfEHgD9o
H1RrZkLlOHahP2UOzc9U5Sx9I/lPbhgjknB4/5+ng50smaAKaTTckyVDiRNpgvsOysKxl/qdYWwW
5weuZwc83lpw9LHUcKtKOz0C4Fls7t5z2JwaoMFMeWcPc/eM9twDEbb8xglpqPgZIDeu2lFoygOE
Q/7VBL58g5H37fTbO2wc4OoFl1VlJWRILQCgbBozXEbKzBksy2N2lWDc4dhy4tzAM6rwUTWUcraU
Elf6QHhY9sVLiwKczSTGAyRmWtWSiTp13N23stNtHRJdfgE+oQHO1QCczQ64TgtCNWLg4JXiTQdK
t0h6lqauub3wNUYKYEFVe/gcZaVuyyBnv7tIhxfAOXmq+lobgCgPxsxMJPhMtJr7onDrPW2R1RLy
xnmHdV+El021l4dGg32kr1tkHsW6GYhZQ1ZKL8kgXgYWl8kTzX/jlTYMQPh46kcDpTSGKmsNc2SM
g2xOCNrGho2ball4T0klxGGnQtlfA1dCb12xIYdTzcvp3uuMppem+PX6cCnDw+XoEdg4YzyPGklL
pkRyukajf/5hH9nyixdkPARiqawG6AMzlwN4RsHIldGXw6BDVzCGjuDEA57fKY6VHd0t63ObGLwj
WpMUqOZD4L6+XMArH5fDAf7/QcE5SdSl8kmIsRjM8Aq3gQwKVnZJaNVieayy9GSu40R5gWFGWTIx
JfMpKTvFJ8TmZ0XxnrjhOSIqJbwQB4jH9aQcmu7em7S7qkJpEiI3xjoDZiFlHopJeG8WM07BSAOu
Mojyc4hCgZHdPHVWo9DPPZG7kcu/On6S6HsO2gZ9fIiCeJc1xjwwHFYfbhRLz1s09Nl+U5NYkiuJ
uRO8L+fKGi+PcueP8qmTmN0PolxMVfMlT6rjb36rdrQtgkEaWjojjKOvrnt33HXbEykredkoaJ+s
NKqG0QfuArgOniww28wR6yYpvECXBV5WbNj4u7KJapHHCzDK1W09oxzHnBQxJnH5Y+OTJe6xhsAN
qSdE5yX/CZ8NodyLhZmDtftwyehEir9Kph5yOlJ41TRdkC477dKrhT49l2XApJKgiWQ6uAsI7o6B
1IKx7kE7zhZ/wOTbmhMevDWGy0wShuI8lHf/JeduGdcgcln0uknwvE0xCYIETNeZ6RTDpxduiAeT
Yp8VYTKzACjcjhFEnTIATIrtupzsY50kBRqaTU2anenSe6QZ+M78T388vIEiX4bOpJ7T4NWOck+y
PlhUndnGyxOd84RoGeA+/bWUEEzaY9804JA6telIUJhqROIruumZuWMM0zP3Xg/t6ohqjHUmARD4
DQFNjVvgKH2SDCxyBoQLge0kuI+ISOOqS5UKE16yHKa5Tsth8p6LcxEP28bDnR0S+VeBff/mjf1l
BVjGxU9tVMgFL3hqiToYiLgYu70ZIMGlXfuDxXZO7WaypY1XmPhgimtN4dgah5qeWBt6HlVzg+Hi
dvxGBi5+0GQxLql2eQtpTP9+QojElxlBZEqgQbA2sPdaLGvoY5OOWWZ/FcdxW3BeWDgvzAFqeClX
N9TMsomVfY1L8ONL/NlDHfCzIpl4G7p0RRPPFcHXHZOTtIewR3mQPLYEtJ++Z2QAhx4FkFoujlKp
Tm08BD9hcA5gJ9mw8BA55OYY/oXYpUWBps+ZM3QS1uYRTYKb+eDKbeWYUOHElUs5VOdeSqwgCR9z
/ppDkncf2ja4NcMNKt70fNvlNPYnBbVggIyGeCkFfZFtn/h4bxo/Q3QRwJUe3cAPU0miDeyH+SIF
YJbw0W15ynF09ojDovcWj8Y+SZOJNYOc/2pGO0do0HsrOONEF5FmVpfWW7Eq5WWcHQg35uskw8cX
f1hpUSVUmHkHee6Nk7nq/ME+azPRo+jysRvQkFdaL3pKUoc/TWg3Pj4R2bh/57+Lb78DS5TCV3Jn
o6ByiDQk2xWJnvIlEHC7AVsS4vOAGipZ2xX6RAbo++Mf1k3RBKFPLlUBhcFgJulUHULGvBA5XnhW
uk4IIkBTYK9qxkKnVmDIICisfNQrZDlzX/jAaE1aQmuVcf+vKX37DfLUSNuXkvvSMk2CBTbOYjmR
SzJAC9N+knr82/eXXlipqfAp7Ryo0GUSEyqJUen2Xs7b/euEKPwuKd6Vq9LggkcVMHtRQ/WLZxxx
w5IfICabqF2qCBU6tCpTmdFpEevSiTRrDkRk+fYHWShfrB4RtbdU19L9SzoaK6nFOVD6sJoq5uD1
2NlAOTatl29zxy2/pucwWOokASK2JMpUPvwJJEXFQ+pdeNOk42X+lxJnyfN1pp12uGkjwDlbOriX
x1Oy3AlPRzPCkN2vDXntA70n8Ept1pF5VU2n1kxBNN4bxy6vcaw/lL0DabbopCoZIJP7/OkblrWB
cBaqdoAwQ2K4pIx5P9vhzF3O2eW091yvXE2DL5bE1GQEC4f0eiyqM7s0sYAOaA9Y/lA55/9dg92b
4oYHy0f0ACJ0ETNdPRR8Y7JznriJAU8sy4iCeXF+46TLoAk7RQeTo4sMz/Oo6FmG9OkracjoXhOs
UZj73602EowqxD9oTxlLHdaxe2UkB2sZ3Gf/wAns3+/XFzddVAka+VdZrJkNtJjHL+buvtZJGAD+
QmKuu7fqRShgCtXpRQkfMbW7w46rL8cIhHp40gbwHCCZl/xZLCIRltKzHmpiVh66wpHptp0+AkTm
9ntxJdfgve66MCYwQixGZ9xIwoZZ8OxQfUBabeVFfqngiUN3T9fTD1zMV0PjxNWvrl5mtWLwPvem
yGYQg2+LJ8FF90zf+WnlH2si/rX/66VyBinbVVdoEaDy3I5K+RR2NNjhRnFnzCh0k9w9juvxykKc
8w5qTPJ6n3mTBdbUrGasmU/C6XTukZyNGFD5yfldnsY//eTT9N2sQvw8Oi4GD7Mq/4atYz1amtyV
5SPpV1m5eM7GyXKh7uIoi9E5XsqQH0C3gerlfWLaXE+Op193/PIOBpSVcE2ooFRoSnnj57prSEOf
UM+TZYVKiGqtUlHr1r8Gx5hrui8QJekFRLv2MiZ414IahfBxOwt3G034ExV0AJ8App+onQY4JwPu
ffTR35vbzTMNQcoGFiTsh2Do2aOTmGm8EwAb30UaeOjJ4C8RtEeZ9A2nVoinqvUaMqvMs0bsm7Nl
Luz+YIQ7f5uje+26isjdQIPqV+SgZzfTpCqLhfLMK5JVmG9069S6cJ+NP9KGOPv3OsSV0xiT7rQn
GH8dvDvoeS6q6M8P+VI8nTHjJxhcupKL/tsrBAWtK6+Ahjrdwza69v3D6smqAPEYYrtHxgTA5h6p
XLpfNq/XvE6fFel8O6w/hPIpwNxIdUyAqanDH8dkpPxcfqOB5D6dhDAoQCCGtQiK0ietRkfRHzJZ
X+4tLcIzFSXTpsdnfbf4V/1SqfqAIqnAwDwpxov9wzt9Ry4t9hfzhAmz1YdhnZPc/b6XRiL1KlhT
PF4PwbqFmrekcFeeURJUHz8fQRtHvvqH8NG/gZ9z+fvcQK3dT/ImPnH9aMgss23TTOSwhWUhpLUA
O57a2nXFjYsMbChGSihxGi/xHBAUNJXk8rzqg99xD+4C7dmd/X6LAl7GbCG3A579nUnpZxbyGxq6
OyxdkVX33CcczRtTrtwBiwzibLbYaZzAcQr2viJeP37M4t8leyY96c2N4HIJI8znJ8MyLCW05ave
obEAG72YFUtNuPrNXWNxVAvRqbm657jx3lI7dyrrAKI+Ig+QdVQPazR1zy+M2wrJCCUpVMR3zqpX
Mpg/QU+VZJuuxkXgdrBTfTHiML1DoZHIXXrdRZm/e5oAzfeonxqIsgJOezIVx1H01YOBLTK3qVbg
fwRdSjjIalFhP5Y4wouHAMVLEBRD2gRtIIh26Bmr4PmOAwpRIcmVaEqOuDK3GYvb04G1xEWB+I4F
zUwDfJcF08hDN+r4nMYfju8XGML+goicCHjgc+zkaPfjwB6lfCRYGAyXX45/KRDln7cPwtUmKxrC
LI6O/+/OycaZAEHpAGILNbtSJdpDsXid1+8cRLkRKmwunvW6d+/D++aMbSHSxgQD8KzAJz9Pk1KB
lywJSU1913ZuSFIyFfjhPnJoOyX2dJuAGi8DgHdsR/RoVkrzKeu4mY7Yc7N0hll2y76MKiEPqeHP
DFjV5TGGQOcZTUMPBvlLybg6qnsGmL5HxSNJe6IkggzguyFMdxjLGRAM7n8Je93N+CJawaltT8qT
qdVfI0g2qHnilp6+gRJWJ4DjwHC16RXyTQ+ReimhyDVp6MN7OL6q5+Noppz1cghUUCUiMqGZojYA
N0TBdcHYxjAmWPn+iIyxljEOjXDx+cK+P7SAJl4T4zGUUEmyd7RXs6qO8K4eheePnej3Mu2f7t5l
argE7b2bW1yB5+IdlaNrmdHHesoWNYICvNBZUM8mcccEsS8jzSQbZpk12+VcGxk9Kwm7hHZvJYxY
DSWuDqrDT5tvjBdiTgU2ctkDYY6Y1VBB4UnWrswDZCefiytTN0kHXOabNik8cNrplY5KNQ4r/4sI
iIfU2117VTv16DRDDhdfj4tQUKu/72/Ei/gcOv3R6IoAMjzIZHOrOc4iY/a3ZNYPqPjTRozr4uxa
dLBE0TOD2UsvQZJZ9vSaZ/omLWWV7WQpCyXdkT9pIXC+Y81mlgx4OzoO411tmkvcUUxzKzBKwmuC
yyB+OcztfBQqWfGm1HJrMsfw9muOUGuWdRg9JJqf1Wmu89g0W/T8bO86Jx7sN9DVykJ05d5BCtms
0HFWCDWfprnSvad3WkoRhgbiqIB5PLlNcNI+nJ1wLWncF0v1VX9AM6u1ZdosJbP9Y7U2W0FDZne6
MPp5Vo/bC6d+RZIszgdE2D6xxjNURwgItxxqAecVmcKxGTyjP88pMLdhkHxCY4wCNrgVQ16nR5++
CG+bODRNPRet3HTsjX/4VvaLGcIJFIuh6EGLdooiqxlT7dNdMAttSuNFRHQUffcIlmV337OSFzPL
HPzTw7vNj0wKnN+UvN39G0+/5aL6ez7Risype2Yna+moUvD7eM+ovf9FMTC1JNFsCkzdZycjPnqM
0Xl6svXDp8uWb5vvOCH8jTVEASl4JhwVaqHMnJHOEatIWoQymOX4OArU2VruBtH5PIGpNHsNLqBA
OpxKOpfe+kK54t5nEobxBbXbL5xPZXTtLZQbkNCFM1hOQkivHYuLEnccjhg/MmowW4j/HFipCJYy
rUCMUTJmwoue58PL+zN3Qj0Qb9ZVoStPK/7y7+OV+4oyS8Xtd+ubwidIusYJNYvJD4gbQEmiI1f8
DZqS3FsAQXc4spsbK/c4R1AQNqXOBSEBSkiw3evAQBMqeOmwkXPU+IZ5QJ7rBb3uroItwZivhq3B
omhVRe8KIMvjS0gC+u53cJxxq4Os8j7aDjU9ZndNleW1OJQXTbrC0J5nbEACToiaF3MWi8k3V7fF
DpjWl7OF8N/mp4SRJoDGM3owvD0KupurrUIBM1p+Oj7tqAJGsGGSSWSFSKgalyVbSLNbfsstwHWI
8SZ9zF2mM5R1w475eWiJ2/+lKeSiACzmoe2XvpS9ZW2Eqznl7uA7ZbAk8g8xKMfXu2H86ZZzRnx0
VbnZK2Xj7tpvsxCW3HmtFwUxg7WcaQiy011b7pIiZmm9gmtSDQIT1MLROe/u0sWJW+/HnWRa50Sh
5BqB5EcLfmCfVgZkbygjJ23FmRfTJ/rARHi58Mz9p2mWVmjjxBRy35K+l/ORAjRY7z/Q6TMvSP6S
q/rrWlRSf3QQuCo+hoO7FkNI3FzIUe/dPz9xeEgvk6Fz2W20MexLHcGs5NDU8y9KVy4sUA1+Vu7g
2af7OA6Zjs5jyARtHjtDN+VSNgI2JZtAg9Qffb4h+BHOGW73NY05ejexz4lBlV6nwdHImVml0f5L
4xMRDHn0+FIyPguepUKDo/XW4ycUW9Zrk23m5ZuFQICKcZ/r5EGlppxYGTIFURoq5I+w9LdhKJC3
PjXmHM+b9oAq9hUzGMYhLLbT/6EGBjfdV6h48y8smpR3u0CJVnngZzN6jJCwbMqT44enszbwjbTg
GX2yb6bbfHhQAkCqjErggh17+06J5ppHzNuO2TLYSOcFxdQ1T8ggRCwrr/GyfTdiR0CAdKodD9YY
cFxhY/CUfxNn97Khh0Sj9FOlRhsL8Uq3jMeAR8GtELt3SW09VwlXa9NwK+JAV1p7LFNDa0egCJbW
s6Yo1/EeLEDkNUj1D40djV+WR8SwCsdyoANh5KqeXwgdZ7qQ+okdhOglXfQB9vUsnau0VnwMlFU/
JMnT2t3CCuXeHY0n2o8XtMWhl7bpd6kYAdtFRjV3ak2aRdoo6JLdcih8yx3Q0GsHwkUVep3u/g8O
/9oGey685Igw3Cntw76s8ss/HU6vb7YtIN0keGWEDMw2yrHB1vIjyVuroBd2zwJswRTwy4re7zB8
SewiIOo0krN4gAT9ksA6LzngqbYabH3Ax1zhua5FhQ6ck4NJ7SW3ruQpy2GPkIiNJhLrAbLUZe7u
5e+bSfh+w7aQMQpt1Ld6IqBHxrQapugfrh5jcjCwvY3B5rB24jmq8jiAjVRdDJYzCrtZAzsULj5/
bUekVSWQ+SP76coz2b3zaehFc+Yj9tXHnocyPbwhnC3THvqx270T92dCNqfaerJ67z8/Om8mnUjQ
uu9tXd6GXMTbktRxZuqYe3aHYmA3tRxl1AdeVn/TJXX6HXamVl1ZRau6KuDoiAVQByNFVm8+ob8m
BYzsNW6vaCoiodbTOPOl2M2ScqKKprcrJ4wWO/OpbfYh4ifyhb30XnI6PY26AOkfaVN4uLzvVy1/
LoCjiDclFTs6UdE0dpMmiyeEsK2fkYcA+RpS5pwPayAUO+a17cIXp0dsXaT1LJ0fx5RxDIsRJyQG
hLmYtiXHaevZYx8yRF/SEjss9vbgAVvqFMcQgl+9UoGT0UL2Od75atbBUPctX0ymytez6AB096uh
+ob/nP5RHZCKlFTJNAwic4YpkuC+o0sPayNspw1Q/+Dr8w8rkwfisC+r8dPl+vJhZrnI5Z42ZQHE
ra1Ukh1OLD/TsFWJZMeCqO6S/q4w6NWn+8vdvsonMsVVrmgTHT6DVa4k5fg8rO7OAbIAHIyBOhKC
Nad2J+k6N0bvF6fj+fcCdicwdlqd3xS9wQ8BBbA3CZViJIAtq0Y3XfkPRGE0eIVUMDhZWs+/hnD6
4hkamVVyA4Sp+uKZefNGv/PhNKRRgMwaUZ22y+sHPVSXdEZmCuZWOutYRgb+nAZkfbDd1EzzRLoo
8HcNdp6YxrNZMR05DQroHgeRBh4OoCnUw/ck1xQQNyRKZV2AshCm3a7Qtezth+Cm9w8myxP3muOi
anr21Txlfh1uXzxH/TMrS1cdwXKvacWzD+G3rpyTqIFeILj9bC9zmBG7b3U6iMCAw/MapDzU9KZ7
9XjEyEWbKouavpQ320Qee3MepR2wNw+2Zdts99uezdjKX1MXdiLbvSU4uxeTCDwQrh4eklYGzT5z
6mhS1PT9lIZfgw30pK8QxGwZUT4nGh0YhlZUr63sumzdiw9JDk7M16OiyGOSBahnE2/8FUmvzGMQ
Y5ipUbFMTn01ujdcYtKuhCV7YuoZ2GZQZ+nb6Q2xbqEuhTUMy+dFo6LSHHxGdq4KD7k673IXJPKd
ZrOi506a1GwCEHlo4dvw9D71sDiZaszIYXc8FQpCOETkqsius+DumXCAx+tCFk87TOVkiUy9QMZy
RgmeFDdiXA+PWobGwXwC58t5bDl+TMtc6HF4POaTNzlyOc005R3KZaUF1MHIyaq8VqL8Vi7sD1sL
9d8bRbFDUL1bG1+csvRQbxFewQ43W1Zg1nlIeybN8ADFOANCs+95ogNpyilmIn6BPnDDXkHFQkf6
pSdIyP1c7WFjqf48Nov6sV9678XHJLybPW37NsuQ+Cq4auJEV3kQbWByd8KX5s1XuSe/yhaYF4YN
5AtDJWWtZNqrWALAutirk3adgZUXf+SZYvnsKZe3D/iMA4y1BlLMgykgISjqlOekCYfkn6timH+P
92KH5ux7mVnBFbTImWjIAGjmcJpySqh8oVwVnOw4ld4otte1gLzJcmrsQbaFvu1FxinN4G5ptgt1
IW9y5Mu3J06kQzHkBvRrWiTMBVQZGqaEEjSYGeyZwqFjqyyU+gcJRgBjvMJeh72pNCs3nfj4g0aB
yVW/EheZ9EBJ/Vhn2nRp20bAYfdjM9KJIvjO4eMirJCGC0SL2H62XU3/5Zigq2pH8XYvtPhABF5c
MRr7OKMQ08nTc5OwlsiDVru90lLLvYEvbvmYtG3/QPMQbb3UvWMf8vJZm53+UzoiwWZ4r9frAJSU
a6355aSa4h1pRJSKIfQ+z/5Nf4Ra+d+ugVkHvpOEHI37MJJ85tyuOOPu2uGjLp2Xhb4HnZbycw2m
16bAQf402qEXquTUi9RAiqcBAVininJdFitSuVnPxVRRjNT4bwAnzkrAZvz3RZlkl22OIIkScVHK
0v0znjm7Vf4A/nDYaHuXuO9yCXF7jNDMaTuUCdkqYaZWEVex8yWRrqYC/e8DdmJZ/S40ExZTiI9v
aPsow/m7Nn14Tk1B/3ZXGnjp6wFTmlJ6owXMHlx3ZdVXu62IpuZw20trW9lD1kgCnLAFzLmbVDWp
8pjEp3VFGSwcvNmVdsEcIBJfCbl1tsYOQuahRRy3sUIyvKtSOJW/zrCStCD9ouruj2jOcxcXyIAP
BpiuwLs8+CV2HdCOVB1hQCptG/a5vszReCBfFtZuuJ2DJJmVXM5+NTfk18kln7p8A5zDwN+1OKR/
r2i4s/yRk51MOHaDM53nFBvKjSNFtd9QqhOrxkI8j5qiWkqkSZWf8vdcwbFyIfvOtQ3+In7ZqP3M
TZDN5kzIZtsWc478+8c+M4CSC+VbGohchwyZGLJxVsDziCscKYCyMT2jfk1lLMO2jPRvrhwpTyyt
cq3ae7s5FIQn0Z5v/P9pEDRYFVsiYog2DV64Klt7bsghx6sVti2Aq+an0IUGNUKoxHobmFC2m47J
UK/FS/TYpHLts0YgM7sX9H7dHkigHP4IXk5FqdF66dhfE7+qBYP5AV3ZLaNmnDmEAeH9D1mOJAdT
DzfDdm3lKwIULc9O7s/GBx0DxLj4FtXctJ6LPhkFcDv/NhnObyzR3BHHEeTT3rqrkwC4AmFzrAj6
8EjvdbsoqspPH08sMUwJu+YAq6AutecAc3ykGZ3CbmwJ2U51eLAFsdSLhg/BWzAtNfRalKn6N+ET
M5Ama474ZDKxngbKXvMDuk3o6hCPV57tCH/7REn9JEnXwzffxDSYJpy5JBw81egMQKVGesxkqYFk
+nB4Z7uIM4bw3OlEfVio/EM0O0Cw0YqA6MNpET424s7C40pKP0frrznViw1UEPl09RtoG2LQyqe5
YoW91Eq2OMygN1kMXawiFLTm8OB9LTFRRlIES1vwqbQlTjHpk1Uf/pw3dtqOh02H3XkEMXiveRjP
MFXj4dnimtkvPveZvIxt06IlHZBAhDrZIK6+iwKS+4qpsCeYl0VjwLqZk/VtBVyJyVmjJww5UOG6
em63fmn6Pm5FwpxE9ei8KWM7QAgXJDdgpLD1NoEBZbB7K4Uuzbft9YxYwETJr08xoFB/ixkbe20/
iF2LITvPKqC4i+bC8gqwo5dCs9evFgdr/yZW3VyhwKnnSQehrtdZdpKvxOQIgVUNb2AQLhadMFyD
Gdh2dt0QUWOcd3QjNkRS/bht8/keD6MVPIqbg649UmLsKSdeWhnt2KorNJurzMSSrB9CRlgzmwMt
COexVnn/mg8jbgDym4ARtaDYexN7yyiJc9rhzSZ6fG/zv9Ms51K5OmYmuvWm5OTuLcGyiMpihZpB
Of9RZojGmi3xdjkwvlxVcEobP5h0+K9YS0VXnfJN1cYFadXZV4cshBpZz2+lqCl1o7pFGiQElJNz
pYOyT5Ic1Lm1hMBuT/vawYe8CSvQwM6NvyJPYo/Le1q0Y1GdWBNOo4MnobinXfPyU281xylYTZle
gV78WmFOGxMitvKMhlYyMOcILjhSmBnVejiTJlkddvBUeStSuHvQ+Gb6Zz/KilH9EpzyvXviEvEp
F7aVRurjaT1rC0bqm6G92FDRBl1OGXTy0Tfo2TTzt9ych3Ia9MQPIOPmeObwpTybFPqNy2jk2RyX
3ljMpSOAg/Id7ngbAuOpFA68PfICKYug7G6zGyOoCoRga9WZR2NyWiDlJuJhOfau/lcuyqGURzT8
oJVZQQq0k+001JfpTYadgmbzqyO0W8nchjeYtl6mjdO6RmCjmu0wJswyAZqDATCYAycSQsWl6PY5
sdxSLSfOED7eEXvASArBhWAjunYd8ZTMHYC6Pt0GRkjT4fjnhC7UxaSSBNWjmGVYcGRiWCPCBn4Z
Aa3aMHBD/+G0pckv5J81mQLgdlaWsO4c16fgNSYy5oaSJH0YGX6Kk4kyPx0k+3X+EchLF38zbPbA
qC0bQESyZ9/v6FY1SioP5YcAyUfBQPCAqoEzRuKQfyK8x1lMtTASQHe0yAqxfAJ/OfWrZIuOERF7
v+V2Hgnbp5QDlMrFD0YW2BgPSmU5Rwv0N/+no1hlmLFH+anlm9K9H7FYMd7aktzrFtxGnZ4u11zt
dOki3gAhNJNdTt3OTrbYC+93Js7sRUMfBZrlQ6/q7BUQI+iK2YLdUFYuYiJMX90Xd5nijzU2T3Su
FnWJKrRLEJ//ydJOAJlm1KfF/G3nNWX3tg7LKVw+M3qxCv3pg3iqpHTHKOfYSj1uC3Zt/I60wZuC
K1o2KwtwlLe4KSjQAaX2hGFIhQBE1boqzKYjR+FDqKQEzyZ90qifo1RyUJC1MZ/1DaWEVQf+w0Dy
yh6sK5b2nzbvMsiWsa6+OpZmIftIku3qgk7bt5q3xf92mSpVD3UUkMZn2cp56sfp17wHdNChkzIa
TtdB/ntnVlKg2/TNKK6mWF9JI9AO4vhPJlH5mf3RPxnA+BXL68fjPmFFy774INXkmJkWvUIAsvk3
Maaplfz9n+8JiFu7xIver02ru+lt2xtfvyHdhP/lcAZCcmj9hbWpGtkkuN6n0Nn7AJQ9Y4Xpgc6x
NW3/mekH8gnqetnRUf9defF9TweBmsVww0J02VEwyCXjLfUnRN8aAc2H3UaFf70o3vdQcMh4kbOJ
J+Vle8MWn/3H5UveKasyo6gdzGnqeXCXA5ssdE5sH6fl0Alk5CUhc0jZGUSh/tEJjGWW+F0E9quu
HdptQ52kAzICBlw64FutRwPqowangBQv9ukb2bzN17tPIylXJnMHjaz4Mx6yypfo+dQ3tW60hNca
YFbIc4M49DQLj1UZyGAW/y/0n6w3rUJ33BcfLQAQKrj3P6zFagUOp8xB98AYYa0JFlwcUuy6838t
uvdWhyv8osVPYQl1T7PVhnKkEoROlVEVNtPahULdHJ6MI887NTYqysleGJhPdHz5IMiKoBGt2CsQ
oii8uG0rN4aeD+gu9likOnHhQ/Tk3R1KNduS1k5paJe0meaHcDvawYCNkAsX7g+r8G4Lp4IlCr8r
CK+9RMDew3x4gZKJGz53+teY0MDNw0/hy/Q9HAfjmKYVZaqTAtXrHSEjQC5kaHUB7jCivGzzEG4A
BByMzJjDyvmPc1yyQQ0pF+QxLJuJW4jXQuvfOpBmOWrwKxCTYq7CVOte0wyhdVbWaPC+tOQ8fL7W
/iJfsca/+SxGNWgxDI2LYcw3vA9dzxsFE03Z7hTEI6yYv0wASHcsS7AZ6PxnomacsKFYCGuPeKq/
1ttBLGNyH7hJC78tt0ubVy+wLasiPg2QmDNiHhbkJsJfqSLm2atYkkaKjjctQPapmiZy1zJhqGau
Y/H552aVJ4dxZVl4M18ruLRbkWfBn+YLhdVOJwk6ctzDihvajvEr7hy5/TP/3uPJNOrRqyX/u/t1
OHCJTxW009kVVMZQdO+9M/2P+x4H0YQ3CgxDDIs6lEN5dCCHlfeKyIkuc6zf+d9t5f5UKPqR/hcn
yElXk7n5cADLkr4jBS4KESV3ixxYcfnMSvDbe1HWkBgjlSaPCVDSBi9N+xanvbpBiwL5u2X1P1v8
r9HVipY3wHJju8DdDLqisNqGcH4Pe9cuKVx+21k+TKVRuCqASlD+ks9CfiQMUvkhcoWDEFfJIYeT
YKi6yk6NVjRYZ9vOSAeMTdcGdTIjqHhlXTlQioxLxL9R0L860Md2EWaurWAzc+qQnDXr2SwVYPiO
jf/5xRLTCBprZEOmSYZt1nMIAQ61N/KGBkaCVhpIDevUk82qi6K7IK/SWZ8/WT++PgvpzHjMW1JX
oftY6Bide3mfUijTBCK0svK7sUr+57yYglFFZ0oiEu6wK8xkdpjBuqIJOhh9RUZ9JbZZVwhHwpDk
FqY5I95PR0CA3TmRkf/VSP/m1wuT5Nb9Uj1yGibAxSZarrH2HxIkUKy5Onu55VRYbEQqqbccQLS5
5gFZ0oDvchwkJfZa5PXI/E+r5aT6oKKKKEIDBg1/AwZWi2VImW3S9miKUTGqW32n8OsYidZmNM6c
aqE/DhRZ5doSVYEoXHicAK5sN1NHJ0nzXrGzhTIlAPPrsYznpAjqhZhCvkLrRZkypy5WbwIHcvuP
ibk6GWKdSUnUz5vhluBIliPCRRLtVzCX68bCrqEGTYebXftJs9uu9AmDXal3uAsLvZZEC6YDcLOT
CDKBiqyerQPT2P6s1o/PRwketpKjHuspxdX8BYLLXWDXsRP39q+Q3deLuAdlGo28qSss/VpWgnv7
0do/6W3IJeNffah0UXaTOVhGlNYQSm7WsDULNG3KZetWgJzBi+nbFaKtB2vTuvlygIPH/VK8FAge
VyJkPuwWIHf+MilpA3CHPoVspOb1Tk68NmW0wmB2t8AdUQ7XdCzERVQgfQvg9FHbRtPvlGLQWUES
eUGYkom92fg8eJKY/Ynwce0eEKNPNs2bzOTbzcudI1fmXE6rLdVAMOyj5unpQ63OukOfkBARSmPi
nqLAt/JDnYq/B6FY7IzIOLp9FRGMVdUZsTYh7dxnyt18PyNNTGeUOH0CC6EWSWy4tFZhCpNeX+y8
MQXFugOZR85Tk6I2jd2r+cOHrbdmYbBvyjcphvNoCu9VtM/VCwxDCRxAWZqe24Q9xNdeK5Hslwbe
Q+Y+zpaUGBW5nrP81bGQVfO+Pfc65rU9ALJ1y4O3/QQkHZtO7jkvrZFSdON/HTLs/bTvBUFg99ga
4nvXcAXCuCA6+XdlpsqURna3W46FDX2/2lCxfvGMjhJnfC/y46O5aFlWNxA1ZRSsp9ReKhn67sfE
DWHoejs2xgnVh9m9d0a+625l66tbAFD5dQi16zbHcZXmpaT/TnNnRhNY6Yi0c9CqTQ+/4EEQ0mT1
XiTIqM+GRUxg6t4MANodLu6BA9JkA2535bgAuDO9wf5UV2ahGEe2pzTn5GXa/TbBd0n8cgH2NBdq
3TXE0x93MLjZ3v+gvT3mUfF3IXhnJCi5+LaP6PN9MU0sAhGPViHrFRYg9XLK/DYcnv0+5YJBIF4u
ofsu44l7P/8YmtBVBhCJgJQAOWdwOJqGvZKBl+kva+D62FYa+Fnz1z2cSm0xwTC75mBCF1nDbsW4
pM8BmsQPdYPHLi+5+Ud5lqkwZHIPziIkyVi3mrlpBTKdapRzfNzV77pTWl7NOszA5oKeZ6J75U6U
ox/BvdQK5qJpHhHrDxx3mXCCI3mRyTIlPbeLtcsgOwa01flBvXV9d9OxctbuVXou0+v+IFcGyyS4
W0D5T/GHLjNS/Xjtffvi2bV+7QOK1RyrwYJphy5cyBQbejtW0RVk0VYv9RNh6S31cn61xjGPeRbU
RYaqbCVjCw+f714rHDmfKvjGDYOpSiWlGxzi2KIEKmnyxXHB2vY8dddE8uCljGxY3xGu4nzeumps
sohaylVZguAb1zMO3VYtnFu4ax2C0iO7KE2KzeNLCFI7u4K252xZo1ktbpYQ3YAC2HmN9VdDVPkO
aJU4CDfOv4afo563U+8ue4yBjnjMVdT5RBmFPMhnmhG2ddbijQaVPcQfLgGsPFSLqTeD8m3JE7Mq
2+aUHJXixB3FY3SNJ4u753ti6XE/SGCtdfZczpKEkfMOPgKEEqsO+VELIwdB3/fDCp5zrgqvZlG1
E2EzgOmccwKe5d19BVF7mR6n4THl5VrbTVUzs5DYyI5xaMRoP7acZqh112GNE8IhWp4neJk57chn
s8BSAVxSE9Fvs60O4uYxpVH+p24aSCiN+9FXqdHme0GdVBHmlUwAo5DQnCrATjDFtfj8sBtnHRIO
APoVgGUmRE7IfwQUSt0VF7eAV8Bs+DHX9f8alAsH2JPQJyTa91AHUzcXUjX7DgL3cR9ExKnUoRjN
nKig+aW668xb3iLubU5lHOBFfCORhYSnyHBPjcODejzjiSDzev30Q9bYT9+YBZXUxbX9rfeihHZn
wp6c1bcw2+c++hGKkj/NU3KXnj0FcWNeS+CwywLRntnPy1ze5u65sCwUERa3pl/Qa8LZm3/UCUto
aSrRTBfIgU119fxlkN8dPxIbNrzEj+C+Ka/kCGhkM17SwzCJ6MDfwzfWz4uEjglPInAYkrs8o8BB
tbd0A8+63+v+D4vmuNgUn/cjpBFfI/fuZEfDZ2075gLf4HLY0vJ9+hFspq5hFGg1h3elJRQTEETq
ITskgQyQ899Gb7v6STKswxnjQq9CNWz+bewH8Tn7jH+tZvJ7C7u675tcsK4qG2Fch+5587bZr/JP
wFWXXtbEZrpMxfoG/OM9SpyM62QYnOFCWDTmo+ybT4FAMop1sWECRNmOJioKxqgMhRJzHWpg8ZBw
dpmg7Kyab/BEI4ImutTNtUydii2YqlYOv7sZvR9FCVK0In3Ym/Xva6bIQX8Ce8ofoT60+ieOnSwG
FoHyriFKsTQ3BfjHyYqvEPyuyKSQg/z1pvchiq8tHb9BlzFRrLuybdnLSr+FIKv5KeO74+16nKMH
N77u0T8FmHwhMoyyxS53gp22PXADSOs8UT2e7pqVV5D0ZowjQ0BGZ6TPhRNVGI9PskxGigouSs5u
VYtQ/gpXE17y2pSEtPlNMlhmFXx2/n812nLmDkLlBC5a+KEi1j6FTykCuQBmRltHWUW8aTibsy8v
PFo9iyG20i5W+8LNZKhesuOS9ymq1CwdNiE68Qwm3bqQvPzetnFHVz/1ZvRQwx3QMIlUDPA+i7ON
mW0Dz2oNOutxGR1Ku//9KLOLs+1PQNcT3CX8zqQ0rNN631B6VAePK7pOKCvxe+bBB7ujIwrIJ9KD
VfLEaHILrkMD+q4ICh9hOKKBPfAUY+NQlCY1sjBL5AHO2eSjwtZ+QhSIv88t3eJTUlHV+jfjhJJ9
QOPqx4lybRS7V0yRy9tKowict7caIT9uIyzcE9ve74zNQInAuJGb06KtRYflq9Ui9sDXqsHP89ah
hZGvxwPPkja+qgot61vLUWVk6/JUoADgx8YrgvVScgq9jCTIatahsih2QZdxqU1zhbSwCM8D1GrK
IAuBqQAWzUsAPy8nPusAkN85WUnHiENRm+LIGZ37qxkERbBGMuWpxssz5nf+qMXlfnd8kdswxsA1
uOKT3Y+lVSiJIIplmhocbmDJffInDNKRmhrTN0lEwMgimQpv5SD+FF4nbOoQSUMCEGhd8HzVvKKv
aMSgDNb6n+loGHbvijxmUZYtUzkztuFT4eavG43kiFgUwzcE6xpzaCVjAZVFi/MwA/C90IcHN3P8
LtrjOUpCjZnPQVkJywJe9mFM+Cl145tF81F7cK9TN7Q/Yfe8FOzTOjuddM8TMazFW91V2HYlBgrq
bxKF9CYl29AlIu97W0rtJZRYUSAivheVYuAUKDjRq3WJU3mukWnteuv3hipaeMQL/RCNSjbHGK5k
kfJWSuyFFXDhlJ6DmLtDsY8XiyDbsbXaHwFM2I2+ByT1HFt+G5MDR/sMQXZB+kjM2odJIXXUCdXk
9sxSkO5IHZvGKdNlID04FIBiu7bOAFXZu3PGNGBk+oJtB+zriRJwkEgnwWYXxzgfnVp9Nv8Mt8wz
d19dAk1GEnIxj6KIUZnDpWPXiEcMadVH3abmal8lLD1I+9u48HLxPvbP6vrd9j7ODyMA7oCdn/NE
RWLuB9EGKkV2cRmgG+tHpMmIfvbr2Jh+EBt+t1jOYXV7VuDskAtzbv+AThkb3Lq6F3MoZDc/fHtP
C1SK5BIDGXZuAE1kKn7DYLbCvef6K4/v9hmUwVeElIV7ycpCj8AWWXq5fiEPi6zmc4lXV7c7ztWb
8qSk5FzsrFr8t84d0bgChErirEzoMQ9deYkpPXurJ6AEiFDrS1wL0Y7eZcMWhwnxcF+lNfI2XR0s
NgBa1HQcsWierIwqUP6UsSQXbxswQ+n2vi5VjJjK4Om61JhivVQ3cQCkL1eM2HqNmZH3OISGwLDI
xi3cTHlw7A7AgO3wsKnbW9bpY+5FaIOKKsJSDH5ejjryfY4GHdWyiyXOWYL2bHj+uzzyOlu1pLzs
mFzfe/6e+FxtcU87SeLh7BSvJ/BXew36su6wZOhW4U2vxX4jB9NpYLM5vjXMDAM/bMjGd8veXfcR
vqzm25zjgp6dnsc+hDcIZslNgYJQ+uJpJj52T1hLWQ8ZkVth8V12gMRwbUdCK0fIFisWyDlxAAn8
RqAd2ksJL2LUFT0ka+WZuyLEpHNI64mpKcpzcuIwJG4zjXgmi8jnaB/Gw8J96aET148yU71W6wcn
1U3wx6CwUkpzLEyNuZ+KO7nVivcqGySEsx8iyUCbDWRPQ/HCWpfU9a3zqU8/POqoONIvFVeSLNOx
eK/gjISwxZLF7O6ZYFbKgSHs24//l1Vo0ZXQUMTxQTic+Sm1X+ToRm07wElnWF2xXok4dfhrUiuZ
YcF9CSQ61y1MUgX6BLk7jP30EObZOVpzagflbx1YW4/d+gZyVIx6/z4J+/IFtgYD8Oktg7Dcy5j4
LQT0JVR3sQIL4B6yhlrVhf8SnNrt70+qtbriLYd3c3xQWhu9jW9LF8CtNymDCCchj898F2z/+Nkf
6U1vGCGAyZauLln3kpiFE9582u9QDkMtCzd4g0inIxz808UUaKPjHDopYKdmUZ0KK4pWm/UjNori
/7nv3ZQk4+tN+jCypANSZwDfOeyjOuo6A5XSOUboS707WXeoqSxWI0JRkscXa7pTspIBEFLVqpNJ
cf28QmdnG6DBMvnZMKpUz7oubtNDxTxkF+L6RYI2+e7jm5ntdWo/u4gPiMjA2Y8LBHSXTNWmaUHD
KZrHlNTaLZex8+RnxYXD9GVi1dPKdllc54V4gd8thjErr1kYsgDlleNQSzf/ynDlbEV+1AYRy/eq
SYhgN9UX4Gk5yBI7NsQpptWjJHSF/m13krI1cZuAIPh+NkiMnfGQUb2UCmbPzb6o/1qb1o22tV3G
EZSuBXLh9Qvy6B33s0rQLmk+9MSHh2qV/A2apT7fL0dI91p6Q/84kcTcpaadSAkdVjX22aUyC3B8
IP+5LNQu/RscdHtKUVBx9JYfxjB5OcL1pvN7kg9DLNFMxR0bzJKrKNTJjof/hmTEGhUc9SBxtrhj
SMJKo1pvfq4aCpeI4Ciu6qVQkKy6ru9zQn0RAwXrXFrmcQgc7lHeIZ/zdWXNXuvlzqgGFGq1bE3Q
zvDRG3q7IZfZorsT+xT3Thv50knZUgY+bw7aEJ+rqWCGPDO9BsgmBa68WeIDPL/0RXKVgW9ofsZ1
ltspNDUuZ/Zi2f5ViFtJIg+RuXFQ3ZpSWbF0LpBzs8mpj7VZLfe2UAP+A1MGP+MS21Fq6YBvgZH5
Gepq/T35Jy0hEByPvQUR19QV6gV1mqjd2w/Zz3MopuKGD7tYW25WfBpT7/DmK/dFcg647iFvQrRm
pYNFKKAudHWpsscSZPImUaqW6it4HO6yam1pZtiioNO0KaZ0ZWqXPY39dbF7pzU9uzNrfWpK8rrf
iPny8LRSAWzUAfjtuTpsDldjEcITLwYUDfXWtRgsyUan59ziyTnsf1/GOYnaSO3VsSBOfB8lSTfX
8SCgCnho+JRcPG/ojUOm1KRnmsLwCzo3p5Q9QLpSzMADMAngVlDvNMr/HJsE7QvOKKGyD18moxaX
cC0NGLooVWo763P1x6SFxoyDJgi8/OTBkPOxqk+ssODv9s+CxfCwvPW6zJeHYaZ6uOulSnj7ym44
z7CSeG0SZQgM2fZrENe2+MkE9bpcxpnIdX7qFYcvqXrwsuLZqbXof3ASC4UyoasNXx59t7C1hP4C
oahMPcGky9yS69q0XSeyjd3D2I1G1racrY0owP4JdWkZGbFXC6yaXpTy4EowJ3KTW/31apHkvdCE
OHijYmVtH4rPBYw/v9hghnOGdjipvgf5Vvz5CkwBn2/DFJgnk1hWyIphzIv0hCg+4wWBpDBz4mQU
5y1ZK2LWS8542ohVtdNejXbfHhDNEW6rn3zsPj3zoGsI1Xabu/21B3E0mUUTfDUV3BGtk1k0QSPB
zjKr0ZuSObCMrkGvecByCG0DjnSyGIpX2tM9suWX+8UIj2rLBi8WcprslXWtYD4Rm4KUUJJLMCc5
Cuz8+oWmBNZbJb6WJljl2Cnh64gtJurFX2r8DJn4HUsMfW7ratAYasb22RnSEsWAtwK3SvarEcSL
xWar1iMzQyUzw3tB/E4JGcs1hWVnEY/LgiuaQLgiiRS/Lh+qb5r89ivhnby62MlhA5nhBtgm0K8x
SkdyiUuwn2YNTtlrMVOrbIKSYSEjLyFAQ2jW14BpG/S1m0qLrsM97zem7UJCkde2JYhhRLPRTSAj
3AXl+2hrlioCpoKzwqR+AhqAE74FVk0b3Ri5NnBxxOpetgELqR4npdFR989LUd7qeGuRsS/5mn7q
vhHwigNosX+MM/Dx+EL8F2GShjEwhMHHX5CZ5kH+PIKtZXb4ERW1zYqd+4iSIcq8VIZ4WNvOdYFm
wh3bdBvKgzt0AG8UGYBGY6MRsKN2S+gqZFZgvWUwMZ2HSaAiEL73zbtzdzQZAhKYH9Lxnl+QUTJ8
VbB4YPApnBKbzcOmxK/Id+baTg5L9uNyJ9hTqZm9/8YE5FcniNiPoCMNyGDGO7OMtYN3wNHxV/IW
+AD7QNtppFoDRQkZetxMdF9Pxw1WIwHc5pOABcCASEwiDdlV298KqVDnek+mahIwsK2rgEgdlH7B
sTzW163oSrx0M5JroTv4SjDmxDs+rPqwT3FKScC3+U2awGBals78OW1nnBO0kbvIOlTum2544tOW
N4TWioc4IVSkFBzz1U6yqulXA3exfW3W3qQgSlCGIaH6MdzHfK56PboOwVCqXJajwmR5mEwCqEU8
bKUGtI4/JBjdCY8PVwFAdldi3YFmnDUELE3MkOBGFfnU+RICJh+WiOo4hHqjMBtjCdy5mN9ifTco
8a+GKAIIrI4yMDesbaddB7u0VGAxRXGj4E3e2Y/9QRqPZIHdlAHVCIq6eqPW1qjQwC00TOZhFkDQ
gq8YqEjlS3a6nklubz8yQG2TmCFkN7g7gcLxMb7s9h6pc0366GJmMjP4vDdDxxLajUON26kGFHZg
YfpsECgqbsqFCuzVgTB2xRiHKvOpitmFo3ODC/RYQa5O/NKi6iQRuDWznoJoh/jTG2v5MvbCMi5I
EvD7ZBh1Pelw4qeL1ZuzhdsTmSOBJKkG55N0DedjOLNeDNRCg7/IdpkC7+1pgMa2WxBv/J2hbmxY
X7w8QTdP8XKKGtFEHFj2azboFHZsDvozo/tz/PxKGxNhNVDvw8T4oVvS3LXLVvsHOzPeJBpuByyJ
hgJbTbbNswFZoA9WPhWvY5kKGYmLaD9Xv7+AOTwJ9tn/7k4F1CYvJpZC4q4LG7yqFRNzj8YS/Beq
S8H+Xb0Ea7T4AYYP6S/vYBGmVtbL2mgMtl0hJiKLNh/UPMNBJoFBhMRAP7Mwo1o1zUXF6yMdKaLu
N0GtVSaEhGUGln+3P7680Jxsl41lqO2mcN3XY1m7aRBBKlFO6HMNcvEmqOaw6dOx+SA2XSMfP4G9
Z046UKSHrV70B6KPEBqXz1dJi2l4Nq86Go52kKY+28sqCN6ezywTiumctqz6qOmeRngW0yPfMatG
v/eVPUnxLnP7McI/1zG6YJjuojb5MM6C9GQ23AmWSMPluqezFak9vXNdjNo10E5D0l8w//n64OTD
2NysoQw93IU+wwnJhr6TcH/0dk8NwKIuYkjnHA5Jkdi/fQmhev8h92fjhVUyBGckv/xIys9kOkta
TfRd9sHp1J/LUfbmSATp/TW682rGXuG5rNzxb765QhWXZusIvL4sxw7PLr+e1W6UqDleJtiPR0JL
7H/2jprO7+u0HANFn6+4GZr/O6z4HgGBc+1DfATRk1zDJh1eFrmWnV83S420xaCotAMOHDTk+1Qe
Fnydhs6pp1T4lpbquQ0Lphd90fUFu15NyrkKetyYPGLoFUU2O+1/4BRwWV0BX4ARuXqTbkWSAShN
gTjL6QxWzY/dGcQZrECti/8ogM1VMIfAnBNCl4Jp3ttApAHlhivOAs0EQFCs+oEdEKDPeLuiaOL5
9ydQDqiGy3gBhjSg6XiQyhSwEodNcuNRnGvQrI4gSCl/47fmU9aC4jSxJ34jQV1edlDhJdAiOrjB
K5eqKH22qi3YfIuqAznom+RRdgDf9j3hbaWjSm3Kd1TcYrivwHq9adNDtbFkrj0VARcWyEtdB6sO
pf8LH02Dv/rl7NN3h56ROkKi802rufVjINvCMA8fGI4x0vfY6IOnah9xeSoL7+2FSTzJbmyA96HN
IQ6zdKZYNJ+UY5PM/3FAQMiiAbpWq44azitSHZwCfRMSB2DeXJF5js7avTGhtDwKTjv84lxuMXBm
sYlrXkVtshHxVkPBXakR6q22bmi29WZliOHg0sGv9NoUpJ5U1k0wM4X1rJdYrTvi5MHZFAbdWiDS
Itj8hCWtK5eFhwdLQ7YHv/N4+ACE5LFD+kT3VrbBh/K5Ikq63tlywBz22jd+TuABsT1oyzsoZcob
ObDJ42vhwdbVPSVYpPJ6+JiVV4iQSQ2+8+Yeh8n573syJS83Hcool2nVeSThhvLSMT+dYs3tNYbj
NIytsHq93ct6UlKxtmysC+E1OM541/b4wTwl61UK8DJAYEvUVGgFzNqTQwczZ9zf8hCFRg4FE8Nn
3bTd3l2vyW5Tq25YSiaRaTtxNotw82AcKB2iWD0O0MV2pHN5sn5TS7ayXdEvCpAAklvJgJr06rUm
ytucOq/rTV9nfDe6lujGPNn7E1/r95BtFW7zGC+4kqaAaaLGBLs/Wu66YbnhvVS7QCj6hT//3pkR
CzC9Y7ILs323yiHDjSnAD8w48xA7sANgCWOYzu5pb7x0fkLULF6BMVpVL/EJlWbqrEYkMOvm3q8D
ub8VvWSZovwPZuSOyzSMveuG3iWm539bnsg/Oyn/W67o7WorQsMtvFRA0HYWAwenHKaVkiE/aJUP
GBN/TRsVtAol6TyLC+AyQfgysXQfSuFyIccJwxSI8gT9oE7D95hEdgg9HfQL6t2iKVJpWNtd8bNt
PQ/iYIr2+j6rZOZl8L12ukTtpQXJ+jVyqsHpprFRjUoqPjCe5hGw3NfTYBnwTHmYzadcY+9mmO0l
YKfC7nqgocvnl0zn189bqhIoErQqq7WMUA7LZiXBPlawpYW/WrUt1d5CAaksuYdLZ17rYR/5Dgk1
onGVkb/qwW4HMohi2z/Y69646RPTOUebRUF6XF3WpwV+x9XkVfskfvjFJJ/3WvY5wvBekvVyZFTZ
tSdooA7riWMA8QCJBAmm7awtkKldladyQNsZATTCw4K1PQqMLaqyeNGJ98RuXdPSFd4S8HFziNXm
jgWA9jcuDcPA5OlbtVLrry4eA7os2KvZJLB/fpNHr7l322hWmiej72yU1xU6bdE35dJdUrkqOnKr
8XhXbx9/lDjv4FIaWxClyLnvkmXUfhCyGc6lPhrQc0atVqK4i84jDdaAB/Vcqk5rcGnjDj9bT73E
j5uVFJC3WET1+o5y9n8NrGyEXeyuB4qQ4lxcT734cXohJRpf4xZpVNeXFm2CoJfUAXeRHusNdnhb
Tfc2Tj3JpGosJFL4ieAuGcQXlqThtWT/hl1HgBC5+ig5HcEYQKehPxtmqDMOzNhAL59BeOFQas/o
Y2SfnGUggOsf3VPkzeuPa2fB8dj/fULahEMnXuJu5FsooBtWPR7z7farcUiKcSEYYO38svnwOFfq
rOuMpjA4aUcQbrbUCjg0bO9UpbRmCI3kJz6x9eIe96jry6RvmgPGrR0jDHg/t+sqTfF3YLYIdiVI
ZlAtPBotw91VA7nnWyu985n0Uga+8ctUNEr644o5EC++aXb9Neo0fyDfcJGs9o2TiZivGBGqJpIY
FW2GOBi206yZ7fNLE/+2zoeiPUpG31xJ8cEl5gSQwAlSPPHgJIRGtAUjyrlt9BYQuIb9vl6sTMyu
ucefp/3oepAfizJXTk71YcLvsH06xrJ3sh6/f1L5j1AJQXgFZZfXI7dfTEu8Gu04HxFdwb/slGLS
mwNShn3w16o4lm+OC9zlfoIzR/Zjod12UbHyjhku25vF69BiIgbezkRwVqs0leo2en0DzxGZ+/4u
lDBJVYj5XManb4Uv59jhTS9+NMgazi5ScNjYhh+dgQP4Rl19VzoH+xhgQ7R1ikm/GoymYKE/P8a+
tivIQJo5pT+Rd8t2avyJg0w/mOJoK3jA/d1a9vgnP7zMS47CJddkdgH6gPBNRf4VnKJ7mjKHswV7
M8pjv5QEb5xM930iq6BFUjYJsiSUSpIMWsRf2KAEAyiwt4OppIYNUC4txp+XUOqYVLKrYXuuQwez
NpgSmN81LFRDeN2iX8LsloQzSfsnXyV2BzjKhHXwPnGFIBeyQqkOpcpvYT6La4gZpCNESOwI6s0C
hmMeXW484mPw+TTfndAkoYUB/0xMQhbjt33dibH2VK9ojRPxOFJnZGrMyuNyFf4MjJoNLPvOwZ1q
0lhZ1RIalHbH25alzJmo7Kdfl2D13Bfrqi7AOfeW2ovKmIB2T16YMpJiSzU7Xnk6qd4imst+tmnO
QuGhgHifxwdY5xetk7Ua3T+Trw81p0APVogd+jGHUneetM63CaYiEYAVahgOwQZwqv0+Ou5wB1+3
i+vjOO/JS7k4dfPTWVsPzQSk22poy6itm5fgvX86QfSYbADWcHans8AC1FEnXyYX/zUyl68cZYp2
FnBe8ACUXZ+uTbtkzpdyTuXBIaOEJDFwbeqCfm0dwgMrR0qyzQFC5PjAjPIQVzlQoaQosCiOr4Z2
9ziTAuUXz1PSUgBubf0Olhm18Zsh+8ym4wB1gRvLQQ5oiVbaCJOzDSYU8D3UC2YGef3Lc9JXGP+V
FHMocQAPm8fexKoS157Opu90erNprfT7HuoOIA+eNNqL76DMDgix6adxMDLQeLdsMXpr5+hNY3nT
gge+ba68gDor6H5+bananOfro3W1eNQnhhD482hQjDWPZNEgLmfux/LECLUFpgBlogrYAxWgvWpA
gLkpMfXCrcJOqnEMAxHO6W6/UE49t5MiZlYJtCkdR9Ht8roj6qTeDqYq9j9bu2HMMVA3vR77bJHJ
oJ3Ylb5SkGK1VeU9krjq85bwao0k4N0n/zd0iRMkwHWn1adtM2dSsKAOxE5KiybgSIZe/thdrlcl
sz0J8nkQ5ZvuL4gQL/zOKMVj46IEMvDOCwFzNZ7HhX3TaCOlopWCpyokECu7skki9OkufRWq/7uM
bAVMFgg1qnjxCmGJtMDPXmpSBWWoJzzve4V31LPhhu32b21SlhiawLRnpzgRxvxiSr8yavn17s8Z
RQ5IzElNx96JCL7fRVjSl51Kxghm/spewMCISuc7aOu+ZDjkrpGCfmbM77rkK1NzleGG9Kj4dKz4
L0K71GJHAPBuOAn5W2hhGKUeXTKcObF8Lh80jSgixnsHBl5259e+Nk1n+GQsmJPdJ9EtMqjicCaQ
9LhvgaTVwuHyq137OPAiUAMEZUYr5pUKNLgvtfdF4GoS5JAoPGxHC9jUT8Zj9SZKNJtAl/vrd1RI
Ifo+JBFvLfq3T9EDTPA4xB9YPtA01TYmk9Fwt0Mch+7oW53+CEb8g8OxT83Znrqft7+WCrujZqbD
zTGcP/5XVn8b5cOuuB2A01er81DrOPlNR1OD96lecm1sSDx49wKQgMIjz3OpK1ZU8q+RewOFj7dU
v4TxqYCfX3SLwcE1NzCy+48JgcGnEPDXZwKmupuZswwT+JmS7ZjQzqsdSX6FL5z6jRMTQ01O7gij
rXosNHgegpHt28j10oKRUzp3r19zQMzg2y+tsvwu6/Ey5AkSA9rOInd4kQRCJKynUQVTYxsJkNHn
QsHCk9DwxYrhpfO+P/tqBSFH2sBqUsaxGBdIqwbBApZuTQU7xlyueZDn2jNPWm1+604zvwtNeStf
albjhErpe8njFwON0/3Xd45RS8/JKJVSVVdMjuE8jdrr2Hm7YvS8U7f8DM7nXg+FT0EWI4I4U4bk
T2Yiy4oIOEA+an9x4JeSYCrmPbdwt0CSOOtETnvXwgEmz6gkt/yB28lSrL8o/TlF6NHuCV74ucKy
/htnWFrFO/LSOk1irYxcnmylIppwfE/b5xRuGAiWph2eLkBZEMEdEWGTgFwZUqTrdpFWV7GMCzk5
T/Lr16x8jTj6NZGilPJMDtlpmHzZjIa9bl4BmqMyAHOBrbYvGHT9OPcpwXTqmmUbSwzqoXtk2FSD
SHGDZ3CAdwzCuTH0uqbAxWIqte6GCT6w8WnPRuNZln1QfnMDum4y5H0eC5u3DXYFrgT2Qg8F7RJg
7odyhT3IkIxQLBF0hMi35lsJNEGDxFDYWkC//76oDGMn2Ygq8bk8qlQM0GMC8+utMbTkdSjB2s51
LK+yuDvVBC7/rZTED0PIli+xbJzxZHAHJZ9AFRYBW5aSpjk03Y+TxzXXbQHnRw0DSJDmkoE57yXq
ACWuuRyNECFbbHUisi4wj7JviRetxSVlNTTLUuQgQzrsZ/9UduIAGW4V8R2XlIFnoaho/mb/7d1C
VU291jZg00TcofOYewGdxJ58zXUeI4b5EzM02jzdntifnpwbeH7xP/W+MXNHnL3gQr0iQwmohCwS
SfxMKD9fiCSuRqGkDz19/yPySrFdvDp2GVA+P8PMmV0mb7STaT5PJtB8qntp0/zA2MxRMdin21DF
FA2hz/bFreeflOosS9jbeQeMA+cgMJSodcC1qwR46XSxv1KBpcjpk6TVgIUosXZokvfjMdZAarQ+
CcUNuOCiy0mOyfcG6Yn1zED1IkdwWswVvJEKADsGugvXYvzDa9vYaKTawbH1ek5K1/LsZpqem2Kn
PiI3IDNsNQYOH+MIdZd0HoAT3PIGkkrnBlDtwJFEEenoaFXZCDWbg5IzEqYNVYQsaapNy09sDl0a
lX22vu3YZ86yp4T719CY+PkGkNSIE+c+FEu02TBwBaqN6MtJW+MCXXO0YeSwEHkybwepmb5IH7OR
aa7HvzYqRfNl7ZjowUkt2/phlibRM2+NlMeNhSgVkbH94tDxyrzIKrN1zK81HbzK24xcbVVHBV40
TvIYZAsTt1dqJWwMHZKxR+sG+WjGx+tQfG4+PeXrAwL2/gOeSJxqL0s+3pLC7cJLdfcCdetPf572
ZPoeDnO9wlwdrEEQftnwSXezt07FqAKWM+z+ry2nZMZ0bg5KhpM9E2nfZ6SjQiu0rDMhtE9r7M1o
EWYqUnQyBsHW42R3Q+XkQ2969D339JIbQL8mnqq65KIaoKHhU3s6wnsMlv1iHcacBD4Lcl2lS7am
9M02ijMJcL5txn1OQHhe8bb6jSO5JumLNYfKFSd0YLfcDeMwKJNspC3DD3V6no/nxVHPIbLUw+3b
rvkHf/Tg9LkdSy9TmSwSKK6a9DB8zNRFh8fkpyi+rJLhcfrNKNCMhiTxTlH8+TJUuK779boUmSOf
4zuiyCD4Zepo25N3K6aTzoU/IBvrp+i+FQ4Q1fO7euE1g3bcTBkBjrKlOJhfA3Gzpoc+LFJYKliA
7rkb/BbFWrB4SgUSv9YZ8Qyqj2SfMxsbhc/krSVbn0WHfBRd2bwLb4DnojnUN/2vEEH2vzuufOxf
cIlp8KnMt5aqmSS2mgrmIALTwNG45/ttdw9iYLnLP71lv+YQHc2B+80x5W+/1EK+MU8GrD3zDaE+
5NlHM/WLU0vRBVTT4ZtZ9effCj0xoEYGS9P8tetv1uYJyGvJAXBnGo3EnDtbuo5VYiRpvqTqfjHo
bN8twUWY35erIWUNxG4AEK49oQPGOpbx2WYu8rl4zli5aqfROGueO5wXshbLCKfvtc0xOf7sUhlZ
Y8DNoqmDlYSGttoaTOHRNMc79Q43yeXgc9JptT7XW4qvZxNAPcOFvo2/glrClcbQHFe5U+guElD7
RKeglkCnM+SPh6y0WDKJYl56G73Yc1d4YtjBIrIpQCNVXXAs4pS89EzviWPEcZTlYi+2car3V4n+
oAgdg3i89W9vbIE0VkXSSpeS3Aqtai/EzJUUG0Y5Fs1n1EryZaavLha2F9NRz2ONfoUcx2bnOvxR
tBOeS0g6QemmQZbIkTt5M5WyWg5VFcCp5tO1iBdtJxCrszdmH/4JW78YyuknOP97iFsvac+q/X63
gaj8EJZz4RY10H0GRfJdX/zXesZej9wK81DThhhjGkpT3MmLToBv9Ib2ZDnIWtUoSqmg6qzYf4B1
ZirMdQLfEfvmVoeizdO9TFiJUExIxvwH4ZH1l64a60cLM2qFWbipbviyZbzgg7YZYwETBxool6tp
vStuWZkx4HxSM2IP8ic9vjH20bSMJm3Tw08NFVB85Wsjxz7s41Dcz2mduHDm48E1h5cP2kc0YBQf
zoOYmQW+5sVMbGQCuZpq6GG7u7qz99JeFWAkUpNv3m3pMvVmRC1bIq2iu8M/2wVW3/ded0jHdt0o
RHixGMo2R9FiLCXOQPZ4BU3wi01gAi+VFXInqr696dLEAK+FfJ4rw8hKR9QPZGamytJJ9AfD1vFc
YP/Rr0VPS5NP+zYRtAeMpidZmNFtrAghCcTcUGdXDsVUg8iSfBl9/vHhKwCPaNeuwjBwIoM45Xbh
fuGalp88zotaLYDVBs1FaNO4XBRm1x+RQJb2kti/1rvyMKrPwT5WmUiX+ne6QmvSGiIrgkw/rMx8
HgoImXYIpEHmgbt57jO1+0oFHudatOA9sIWUCFyjKb6XcYmOnYKhbrBsCZz0mPOrqcThNeJBllXZ
JaYgmyEbiULp9D+yQle+ai0abVcg4JM9jSvJPdJZhbrE1LbCgNd36SWDYuZImvlP3t8Haolqx9Oz
hW1D0q5dTr/LmFi2l4z9AlPMGkZBQl189V/f9gmHkobB0qOIJGCdPzRidZnfkqWYsNvGgFmE1gV6
kLadD0WN6M3Lz/4Kq9+WcMYg9ot7pWXBigBtmh7RTgb1wzLHOG4BL5jXHhmaDSDd/+WSLsKm2oC2
eygV0DJASQb0SaDgkHCjScA64x5nsuAvntcY00oO7/6vq9ZKNcLDHU+4yXriIaAZEiPXbOeuxaJ7
gT5y4WdcAsuTOxZURA9RBhu+22MVvjNhlKyQcWJYWSrICsT6WBDnhQxCq11jsEVnwFpt9TOV6zVU
h4p6vBtvMIFFoKZjoKFNGvWJjQ2RUahKUzRR83jkYRUJKddK4exFX+FhEasjuBHD5XzwjhsKmT6B
VbRZWDundzNKyR/68P4wJLdQCKOja4KsXyM9APmucY4YTsD6e/QdIO5mL1pQTwy+5REV90wB5pbk
1uPh87hHEDptwEtovbT1d3zJYcUR2AevM+Q0zgvWql1DWPNgIc+tC/RCrEGr4qYqH0K/gUo8a4oy
ZbQVFWg3XGtRaphiwLociDxTzFqiofbPW3eOpOxsA5LtIoysTDP8A7Ln6MgOKuLZ6BoLzVcuUnlJ
68U0OZRZmqmepGzX0TKeNBcXh7PWiiumm1j0b4bYyk/TsziKvrWWLDQl/QCZhMTAgp8ZIrHywb03
tHSlKtmaUvH48vfWTB2Ls8mGpKmdm7hMauTuDym21FVYjNzUqGQYbEY8n6BYRcSAl6LsWjYNSJEQ
J10O8Bsp76yJLciH/A50EdHx/cugi/KqvbWXeD1JijOdG2/n4SMcKOGSLcQqnRfeRpCOlkiZutw1
ueH50Dp5vvmdQFlwKIrB5A09ANWqJNshMWP1UhzbyCotFRFm83RvgZeb1y+W4SgJJhJEfOJUeHhW
WS8XgGiUZfMheZcKPYNjPqlaQr1uRq7arfypk3LoDM8E9xn+I/ysg7ihbwyHEFmR9Mu6Nky86VKQ
edSfJ7YmSdWsW/pApPHUGaExGrJSx4KEPcqU+vg2fywCxI5BFnazOS7pFBss3Bip7ltdZzQsmWYf
ZEi4gAY6PWi0U1OQzbxkgcvVMqTopwKCvfafnWzDwQRqHJz8D6gh1O2Go4BHY0wzzD8ZEBpY0DSq
UZ5u63Z2tyLP5hqsYExUsGSyYyv9KGIwa3ENlo1rdQsJtmb6Nt8r+h4ELYSzVeVAXI2GUusC8lLw
R3ThAQZWIy39HZQYZk6DN11EGm23j19J0k+HnBKE5rtEv+qUSsBUUfGI+krw4bUiNjjTI2D/xdgF
nfsYSVvadVIJJCjBeiqVQxtwUVePiNQSr32YHJJyFeLutcju74j9SkUD/otGP0TdZ5NY3EhdWZZI
9mFGVpr7yCO3l4VPBsq5bZg84Yh8CaseOqA22I8aeiqKNKjMQZ31KBKD3LC2pAq7Nwf9HxaDRcNP
53Gx8UzBiTrbE8HegdhJ6fN4yWU0vfmk9W73HEgJo4XyFLMCZ0ywI+C2iSRvgVlv3excaD6KjPeg
f5z5gogqWjPXDFnIEUq7SJnC/UXLz1bfV6v8H2SjPQMuIe04EhKNFFGYSqwkLAtvW4cUtsfdEzpm
lVHA5i466GMird/8wZXqzUdLfa2hdCXU/jafvwCZyEevRZ48xwLQF5PSQXLfwYJzl738Gam4dNEb
C8M0E6wrjPJ+bg9I55cRE03bEQfxrSx0Q/tL34BG8xgGDlQeD+yx0PrdEEoFg1J4hLaslS3NVvsC
2lVW3rxCgZF+0l+cFttyOc0snNk0+U3OzGaBqcGx88fMZuCr7eJydt4G4YUd3YNx4RmMWdRlf5rv
uapmxTvKDqCe2VshlAWT97LIIGk3zueREFOIxVc+82jSj+j3QDiq08rYQtn64DzMeOYFMpEmBKBe
qe/Nw8Zh3aoWaLe8KjKBejslrBSYpGmOEDJyEgSHE3OZ8d93mtCv4kFDOpL5lJAFv4eW5EFv7RIi
3x7OrHjLCpcTnXOpMreyHGfHbrNc4WVF1gUOh1oRZc58qh0d6oLjy0kr6iFHQa6Zog5crQZGPs2O
Vyc0WUHBhjoQUaRnlCORNBo5zsA/i8gEp4OseR5yF7N5kKPNrNnYoO+oplrc/0MUTaiV2Guz+kz9
GBH0qJjWO0AplEFIdxnnSdA6K7tJFsQJgaR6saxU6ha1ZO3NuQiDcRvDq2Bw7z+HfU8vu/5K+Y+K
w5MJXBP18WMYtnxkMpXWAKVz6dK3TKXJh4qH47vB3zNr4ImGiKZd7mph0JUMUXzEn9wcwAdN2kek
c3CjbCgR0zjymWnf6UBODbcbcGAcUjCr8L7kONihQZ0iHiSSdLvmjPcoXS60XrrDcwCIlIVZf89e
zQ6IX9G/0re6U1a2XyIUw9TvfU/fdp8yAIoD1h74BYE65baPQBHSeYrxHQlXdSLfaMfjJ8fQCcVG
WuSuDY7zMZVctut2NLO8uOZyvgIZ8XW1O/3TYpsNmC9MsZcIZJu9wtNcEV+MQtHqW96GfJwwi4Z5
Bo3oAltpXrvq0U8ttzITJ3tIdI+hzpZcahLZmOQJs8v5g0nNvWMQGh5dMD20d5F8Lils1emRvFW0
9BOOHU17x8opCRcEYuO1Dy7fuCPcqyzljYSikBEfIMNIOHv9NjRDhbW2qjoFXnwDwDNjVdvvd2fm
RFCgMLP0fY4G+K2VxSiqRRXl6vN3zKHlNf4G2K4ISYoseEkR7Eyduj9R0pee6cd+8en5Pf7Wa/3y
P0acO8Wo5wrUfHkuguRszUTFfLILPqpMC0yzAi9moAsPBuLj6ZrURd/RlgIivm5wbDiVMjZ7sv/F
r7KfNAkLPvIBGLuhonNXrox0c1HqdR4fn6PGZ2jEI4ODD+qqkW/FNzlxdGR570EkUlLwZG5cp+y0
7CNcvCM6D4j8REMPML+uMSZimcoInb7SnIpaWvI/GrT1SmPxzcklK5vXyqUMjs+Jb33O/+cviDY6
S+cGzEvtnW+fPhQnE9X6n5iXADz1fgC1/t44ja6aZq/+0IrMlIZdquv9oSFrzkPKP7Ul40gjlSJm
vDWdy7PoDtA8a/0TB8arosbN2G2EVtDZPlUx7LoSImmF5EB9wFGt8B1k+m2y1oXvRwUYIe69Q1h8
u24OD5/zBq23ff77tfkft9lN2wpc1Fp/ujuXbrrD7Ww6etftfifoYnGJP83c3RYjIAHXBQp/CSMM
QFkDnRYSO28Kjnsd+dYestO4rTt6G0Wsww4JFZNtVTUw7nbHoapZeGAOYyvtsc7UwplLyPzFIvJI
v6zlTgRXuCrOBINAkOzfYP0NT8TGNZLbedcc8Y7v6zhX5KTK0HlJruO/IxIf4ou5xNtwJNesdWF5
KnPuc1bf6K5XkL+5M9TYlY05QxVSd9NRaXW0VI1WtXjoqXZdqL/XXaPW/+eb7t952L6WXOTQgrMT
0n9dwCD77GwhEDkVytivCCLQXuqzWWxq5NhJQAbmHk7wfgHHbfa9429d2mrwmDeAY4xWKy+7tGj7
EFhYtI+Kegpv11TA79qVQQoOhTpfvmg/rLTiARebSXl9isXTwfovpcAoIS2py/ZsthzvvUf64oQw
UxtlZpza2hJ6jt7xArOCfeSaDUUqVxqKZTBJo6/6jUl4wIyGqKh7/ohazfm80opuqVFLptVoAj/4
oV+HiRAg8K4ylHwIQmlsFdb4I216PKf5wEUuPpP8Cs6Lt5ShVlHZ2vxH9+yYHbymKXYF2yE0SN16
LEJRaCQbCt/kr78M1pelYB/AXZFPGs+CzwINtbmTy0Roowff0n6ZXIaKC949nHdbLsMCPm5Q3Ilv
wwLDYsVCW07x6qzAlANriN9D3MwrovK2rxZ+bGyGH2bMPQCm6cn1Q6qdmsy6XKW61v/YxjRUixNY
fyoqVVadkWYiF4i8E8kIV+JKnsWrxVxB35ympMPrvhhRI/O0FnRzXqJ6Fadu21mLK1UFc95Ivnht
iUTFD3IzFtkXs2l8cC0sZPMz4x8rCvmFUkJA14XKzSdsBqXslbeCPMmTMh7VYI39UB8tlTzFU1gX
LEmh1aznZrsRsfJvflBq4mE94w5UIc/XGDqkrHuU5uSeWOVhuxI383BRSAP+ms+tIIOhP2hxMld6
h9lcIDChkgptJRUC1ZJtA6EzgyoVQUlJdPl8UTNjO7Ls7xZNw3ctNdmu2ykKaBsbBCI4XNm7SAhh
StRPO8OR8WPScfAoDPswfg0FUB3s+DYzavHKeI2c+o99PW2IeRapYdetQJinQeogpwld672RaEVP
qmNfoX+f+yBFMvFzdJOxkumFraAOCbBKEw19zbPwjTEiTHEbW8WToy/01OlNst3F5AmaVa3UqcNx
ttNBfxEmkrBJNEdJonxlhfQpY3qPNkjLx2YOTg8vKbnYocssUtqBf57mwfFA374Rnwn8bwQ12tGD
KxktvUS1vHB3Jz/Dvm1bBqbXj/mnFGDsVGv7bLVEXG9VXw3aTRywse1uqb+UISPmA8kWNM2ShPxW
RPwS6xo1PQzr6sesrOFVlmwCUcJSXbpDtUpUwOW1Yx9LIS1FV0rXIujsBAevk1lInuOknzWNGzRR
1J//g8oiXxTrxj+BspdSvTIcMmIEmv4US2UhvQJ1gD59x8TUCk+0iWoA2I1ArglPJBk9J1K4IFIj
a6Et6wIPPKU2uAqrVZDUTH+ewN+Qa6g7Jn4+BT9931evhvlJx2hDWzxtRTkabmASx5UpJKDEyguT
OXcBjeLwIRxcffIBU33we58ezyqig7ah1t8tNXJgSyhTgEq+qPgLHeoXEamgg+NIrwTRAm6Kr9Zv
7Hn2oHEQNDw2vr75zl9pK5XSJ+1Z3zlzlwxDvdsN07I5HlkSgyv5NXCVCoEIrjT7j7X13SpYgqG5
JHcimj6Rdp/5Bh9GXqnf+K7EYE2SPFXkUAYoX9a4fg4htJkGan0qyCXbGLHigwiBSl6Cxag9CeoY
xGZ5D1WQCpT1dQlZdc4WnLVFiPenw3TO9DnnGEl9SVt2zFF0mUPOlns1EMm8BrceKitlBW9m9PeO
sqWbmzOczbOgbu60GyrQhWp8a4zdcvvD7HVoHNM1haP9+CPM8jnNDO8NszNXR3VfhL9IZVBtZa0A
/sM164FBSDRjd01I86/2E2X762Uy08aH2m8pErOQpPu9iSGzfaIktqpEnB/e9rUYkbHfGsRzkWBx
3UFO8L6QOn635xIkJntw3zzKF0NGeE897W8qWUwXb/89XYgWZKzKgQEvq3pzIaTVXYf20najWzTS
8Y1S4GHmEad4Y9HYAt7n9ChCxB/EKCmG0X1gRyu0H3rya8LoYd+DlYoVMHjypHfj0l9a98ABL5tN
ngzUMpDhzmw9gz8eoY46+ZX9mrRtNvbZTUhAshH1ce0IPoExq6MK9S5vRp5Xypz8bnmzy3mDMQtm
HhUeHnSbMG401C6bWe78XHzY3VUV7/rse+Oln8NW4fSIyUE/Pvxw+3KB+F9nCW8Lb8cdt+ID6LaR
Fo4dOoq0mXGuubj/hb4rnvd7mmT+14gN7GygBFmW+HhE4T69V6tsb4S1JpxR9PBp/n6dGeB121v3
bqkMmUy+yZuuzgPXHn4whpiJlKzx4XMjz1GRo6ihMKnXSeempIEfXT1m1z6aj9iXv6hQITXDqp4F
OBDa1HlKmyK1+6HigQG/pnRkXNTsXEuV9+wVGQhKpbBCXPcBVtnHOpOn8S07Le+XcdhSUldQdG19
60c8B4qnlHFoIEDVJhH95mgOrS7jcaRv8RrNEuIrpHGzgt2h4TybAo2oOz5FfkEBT5S3D+Q+titz
TQDf5YdaExk+SGlTsNdSpjsJNFVWBjlU8C7kfR8S4eQimNG3bVXPoYvTlesP9nwEpS2mKr1pO8kf
AlfhQEUjyJymVef8JbPBNCCjq6OinqkboMDvcQADdyKATF0rM+3PyvEOmdF6MpR8cSYGWH9e8jUe
Pi/krTjuVGEDVwywkSDdXPELGx0lHt5nRsHxnHyPoK2NYZBnHP8C5n3+vcN7CQc7Hh9mCoRW//Uw
+hUmePwczJr+MO9V8nuD0ETVIw+gtFLh9kHRJ+jc8Il3D5CXOqI2UUYU7WRy7UGS68CEDpTppuTD
f2vhZCbgSmSmqtGpr52z1Eo1j2vl+Ablru8i8TEhAS6Nbon8w9lX8dJ5agG8gHF8JVHYcMkc5d4C
bKR6aR3fJyi4sKyxoD5RliJNiFH3A2WVe81a/P32tYZyJnfs351HXfyqlc2RIIrs6SCKX7F/m6Nu
ytcRgsVcYqlY6l7XHGRel5VqsSoH5xQgO7MJs65TQvAsR0kHFBQpopxyxOpq8s+H+DegKEUGOpFl
XmOaAMXAIidKTB1xp81n7mliWMDULEtfY2QlGh+p8VxxCRoA8dtmnDQ3MPK6OsSLRzjMh/iF1N2R
DqFL6DCQpHOBHqHNgvExofXPxGDrDYtsXODWX9vQNihIEcJUp9AONR1/jk/uAEPUc+TK9QMvVRGr
NNewmYL5FJDKbDP5cV5y6iV2bIbBaa1lCC+/4ej9BZmdmmO22C+uDQhpUaSIRQ1G2/WF0H/VP3Po
5Yg25Cfn9cKoCelmnU6TGeSWCMT5sTR/dhxqYEJfFzxA3D+XauayqMkGpAtj7cMNjHOHPb7rOyW4
1IAqC3o5660NaFfnzo8fGk7K8bOzCNQ17v9twNf0QbMnAw/+7whWN2MAiHWEJ4nCUF+uf+EIWA+q
HgiuT6WIf5BNTQ6BFWXg3tpvWNhp40qxd/55kMjYYUx+RPQAFYkIR4Jc9wVjYzN0pyIDtplgNrIY
BNheI3mUjgkAYwgJkDoM6Am8luRaSlCaLLovMM8J9XFrRAlPwN2QerfYApwpZ/snDSCrM1IF/PTK
XJC6RTxrJuzphZ2SOsCQiIEuZPcwZAzCS0/LJQkiOhg7E9pbfKbTp2J+iZulDI+rqUcwW7AZJ/g4
i7DiMvMA8AxebMcOVC4nXLQ9p9hgJYsJ5PWr/sgOft4VryxVYyvfm1drox4nRudHeGcJZKVjdBU5
HZMAkay74jcE6qnUgprKdfyUomDcNKxJU1wqvyI1zwSjGsYzd+OZhTflyyIdQoPmmt8Ede7YaX5N
l0oZr+IABxucS+jwCGv2/fw39eUJkAZYOpBgiw0bihflIDxwx9f4yZ1KQ6KZXDjjyYeG5BFt2UrA
HZzMCaCosCa/Vbk5IQi+xBiNy0YrjggIkf4q0tatw0Ew/wMYGCBFt06ytVbgTrZKw+zL2XOYi+El
IsKXeb/4MN8SjFduleZCv3kQRR8CjZnHf/8YhqHz0fd0dGaMX57yJnqTvTPz3eCmgkn7Bh2b/9Ap
Z+6HBlPsSoAE8Y8800U9gfFf/gstfz495yvc9s9F4XU/VEtdW2+FqhjoxwQv/XoGk79v2YBjqVEW
IJZ7Ofd8WTYuY50YZxDm0KAXieMWM6UmaMu9xmWPX+w5Al0BCaRx7eOc8HmZrPQa1SWl93CWhU4C
L8LFetIndjDE2itDeEBNM47LEW9DxgD803wPOuYcHDYokd/BwqGZtTGyrB/kpga0/KZXW9U0tMQh
aXj80kGwclbjdqYFA+iX5Wviz8CEBIz6EYxQLBI5eUq1/6AthVqVNaPGmnkcpeEoNchP2yEcH0ND
21fpEfSnjR/Hha0+I48eivPqPWj79wNy3nPyfv8ZU9+MAI/AhtU51vTeWLWSYdXjPEVQrRw6BV1f
klhAiVm8E0OB+vUsxcFo9KUc1Z11XhI82MotZfVSLnDjxrY25tcKjox1MsIHkiWlfVC4i9zGsfPB
ykwiMwSE08Je2X7DGzdtu3VLhFTZm/kA/aTTRSE4F4WaCTGgj+bCHqHJNTnloI8ZXkwDR96G6GtO
5sXA5c5o1wJgPqs4jqOFBeOjIYO5J5PfJ20R1lsdqTp89K1r8mj1WSRTaVvCRNMsLg63r3r5eaUs
v3vpLDNyJK3V5gBgNPI+t9oMyakLK4e9r5Gh/bVRCxBqESdepUY83YSEI0r9BmyfTdPBTJNStv35
MTSsYbmCrM8lvYSR9j/uGuZi1j/tkuN2HAT13lOe2mauplZb7LF3LlW66CRtojUv0AHKKDeMLgOd
3wIthkKI2Er63bA7wVrFzt15ZQ1J3QjWtM6G622de3dhS7DZJ9lHPx7O45NIK0eBw3V0Tlre1mlj
eqGaSPvMzfuVvbUH49eTXfQapIvkeu3ft/aMOLO8CUUWLqAgxC/K0sCOZFSi8tT5V8L8hfxY6JQh
rpjVfs2priVlWz4PPwithl/8XRZFvyZHbGFmrs0L93bVKKpim/+F7oV/LZ2U0c6Lw//EUYAIGVjc
UL4HWFjQgY3efLryOGgY1FkHRx3zipYz74SE8x2xXTVdl2fO+a+dVnnVCauagz3HzkQMGFLSseVH
ZlGAoGMrFtPJqIOTPeaR4xBmykrjenvJd3GTtMiBVDqD+w75OKGAOaAwVJrskNNMwEL8s+RJNjTL
juG6xXqOc6Zsy67iO4sxnRJx9KoRnOLr9ePXDfp32iYupj1JyxOZ73A5UKfkNeS/DoyqX1H2z1yz
6ws07Qct9BSJK89Pw7tBVo0NZHxhSbVvUYxWG5eCp7e2To8d4JdYA8f+AintbDQ8HwGQ4I3GHPym
xkf+sj+IdJqNrnNSCvn0vQRfnDr/1dphBh7WjB/5vTaueXbBVP3RGTIfqndjvamcrR+amfXjognk
Y+uNWRNk2Bh5WkOV582bsfqjpdMxZ86+3fnkr9t5gxAWzxh8/GfFqK2iIIHB5tqUbRkT+SM9b4AN
3CIYML8aMTt8vmLRFAgHVwxBLT6lLhK7ATiLZ8LWRCboqc11omIPaYDiHP7Z3diRpUEPLwHjpkgL
LFDrwtm+58VBAgLeFjM62GiqNFFfnUUxCkiD7MtdwJ6itz9YldPb94RYPK54ViI2FBhdfbTALVDZ
68GV/Nx4mMg3ivCbzq6HYng/xZMd9CzYWXjeU1yRKOFo1CnyB+Kj9X1XfmCv2CrOixG8S6gsAJ8X
8EEzS6nQHg8aBhKprXi5Gy2LnOfCVgcdAHm1Gn7DO1Ao0CrH3UXOjffSa+OLrAeV7rnQEXmegFYX
6WahclwYecEHFXBRJ4KPGqQDduR5Lzueb2SfW2ZPEzjN+lKVZL2dqigDD/scWNgEPZ5rZYW/IrXv
22dP8wFSjeTm2K0+SgBc18K+K/Z4EYpik/GZP5GiBTRW+JId35L8KvqFQurC4uxpWBbp5D0KuR7c
RBlIhaXwatH/XiLegebItreZlTO4uc0ZdXDXm5YxiefBnd+DYpDxMaf4uCCDeX/QcV58/WRpqkMh
dE+DNoz6f9Yw/ANZ06+gxwMGhtxTanoa4HW8MfxovmW/wHz2t5npYCHThXXR8f89y6AxyrPYTHwZ
D5FucfRiwgtniKytphnGp1XNgll8BsA84ChNNcAc+xW54qvMw7SxcvhJfVZ9z4wY558UX17wb+Xz
7piR9LJM1sLJZYudsDWVtts5x7q2kSljFDSiwZuCGBYtGaK+UUZN5kdE+BMsZNpnormYZQiH98zx
5Og++dh3ezeHz9GWpvbj2fr+8mCIyaV26gh4bTtbKtWEgDytfGw122sEhZXjOWBzHqBewO5SWId4
xuJ3ovdqelr7p2LrlsDCTbgONdDnigdoQO4cJCxRVxBoQ1nQr2wBELg5p8204J/14QhGuzmUFKq6
10kFijdX9KX4v5MaL1tucQwOqTzjddp9xijzsCl3FYLl6hGedR27V3jps7hK3k1y6ZqXU4BcIcVb
IRU/ZU79DnteUVjRFnekYL115rN2+NSbNHPLYsK9En7AlDAkmcpQclHS1ogbjICd4PqePGdERVBD
xpEqgxsfO+Fnp3jytxwxTwY0lCAWe1EZykpdUw9JYtVQbgAwCmQA+OIcrz0QssLpvIkT51n8BC8N
NHP6LkCByBwXOK5of2fDKXawWmBRJn0k0DC4XT57GUYgQSgHT3kgIqEgGyt3UFdrQ20Gr3g+iuCt
vGU+ZH9pBSGyWvpaAr5JhLR+734G5ORMn3zqWU9K2F/LhX5lLvS3F37NSUPkRbwLKdww5GNEMPdK
aBxgwiZDOwzdR4sKGyzpGq5WyIxvJX/9M63k7oWzg8mczKV32LVjoHLmUcVIFt4rqt5PQ9pSDbyT
jr4aL6rLy4ipvjtqhsnz7nhLFvyyYZPcAJiaC1HM6LffW0QUvGo9IUHWhKsbLPBQE8db76rsIkII
oTXOIXNVm7x3CR0/3Ze1O0JOo+3wLOkgn832cKf8wMasaKAVD9mQxlbMQiULzuW2GGqGNy2b5jmH
PD7x1mTN1YyflMELghxI/p/qXzsi4Yhies3b9e1XhVFfe7f+l9lgC6uXbYqU4PG4J+8sI0topuCD
V1R+t1KbCq014BFz6kuhfU3w1GMcVkD8tinb8fCA/PxLD4O8cwEbu/3/OIEb61w8DbvHLESwLWf9
QuJGTp7WH95BceFsfcQD4kdWutb51HtNsh3+oS/kiNwa1reNyhhVZ/bObgqSeGPvNiBb9ytNoxPc
bryb6ZQCuxHvRsYMoZY4w9mc7nFVaTRS1sQvRQCCHjiXaORVBUHmMreFERj2cuvV2rknIJr/vnwN
aCOIlg6m5Mb+rMg6LX9OsVS48bRip/r03o66+zLzc8L0HKsC1Cb1VUz6txPVzl+aD7ts5PyCPXAj
nVVeiYlc3mp35ne5EQf5OENz7X7ZfouRy6E6lPXzy5sfijDXc5NFC04fu6nFgfRnQa88hRj5xJKP
8vRPmIRX9Cgk3jvkKyPYio2ytvwzS10nl+aJl0bMtp6Kk5IWB8tFm6jruB42HuYpIvyLCPB/tof3
rHM5i9RfabsR8tg/baES9GLo5A5Xeq0MIIQH5HoiZf4mZKddSqjlghtPJFc5TerRAOj9fVk17axJ
HyqirvJheFADD2Hu1amE5bpELWFbE9JzLg2z2fvXh4+/2Wk94ZkePRHE1dnpFYsWIGGgildarBA1
odOSLvUlIZ3WyKCelpGHMlOGrKdfyI3cZpUUkfeZptkseG86q/qDmDI4ahClQ+bpMb6VD7JBd6mX
5aIVpTBl5H6KQXPsKSldtf7EbFBO/sbQHALu37l6nhtk9OvfFED5y8Q0qexgpLvSX0U/Zlbl7e90
uF4N4uwXHmAkAhMW/m7bH11TmXImpfhn0dd77Cgp2Dr44rIhPmzfVH8XH+e2gN3/j1k3sH0QCDNT
MAtknnRVa0ZWU4mC8w8M55M3UTxqzhZrleE4AcFGrOxv05G8Xg6ZqsciknET8+As+vzKEH20qi6R
yPspNhNCRek4W2yQYOE8Xe3m7ft4vC/92zORgei/CcheGfs7HF5ot0PVZKOj1HqR++aLhjIwf83/
YMoW4GOnuQACHUSemLjsYJABdY3Wea6/oa61g1wLc6uqIV51U1GQSXSvhtXn4lF3Z3WjugInlXgg
glXk2QxXg/E8y2ru8pmTTh0TGsSqfc3kWV1WYq/dNsHjkmoot8Dii3x00OhEQ3hwI9L0b8fnWNwf
P22y/hA0Ruc4YdyKP1vZryUSlIW0KMF7f9c7lcqxZyxwIeiYkKTLwNTfsORy4gANlr5tbbSc4Di1
T0BxGS4yj52qzJ6LPOk/xdl9I658IPtH+CaB2Nsx0KiHpXllyQOJsQ5sgj79imyUjtYBWUyf8ohj
9fekx4F3LqNrv/XwDuZMMhhgQ6UFNYtNOk8rZpA5mbeTH0yeRoeSZIaDShBStqvajIEkBJR9+YPn
mm+Di0DP8rzWyKoEpmLO6/aLf2klYTQjNDhrDbmJQH+pDxibs98aNeC/bI5Os8D2nBLYWV/2s6LC
nuivS4emxqzXnx2F+j7XDEbx0tvuhEO3tuzRBlaM6IHCP//CDR8pdeR6RuBmYEgAv4GWTm5wahB1
eBsketCKHreVhifedMilg9yW/cXTceS1cP8msFP9VufxRNpNWeXWaoJ+bz/OgIyhUHLosCoFlhbx
BiWIsx0BROjjq0jKxvzNMdFwL/fYeIw2PVG4i4+rjlKRQvMV2sicfSUC7uzaWXyhii/oJRLXFrc3
DX+HsHEYsMFZMONlRSNzI4tZzbidrVZ+52fNBI8W1BLLaE9TNznD71iZQu+EGJQ1VlvN2lltsDk+
wBfmlpDkUdBlsWIr/y3yRuUC7nGe6w1aXKW5A2yxYm+blCmgoJoTyimWh4A8Lrxh0HPgGXjINHvX
byPNPPoI4VU3/uf4+6hPssgiJVPa+TAhoHDmGUzV3rGYNempis0KwoI3//8QtcvQjtzG7PN2dXMQ
1Na4/yQYtWM9JdwwqbaZg0WLVfdehf1iTWFytdz3LbwGLZ6eJDuX/M1WBFf+0I+9iu5jX4nl9Fai
Y0Gh57f3AvsuqH8RIo+INp9sTudYfuhQhZwQZNCD/e6z3LH9fFoSjOktV1DS66P0WOa+lFUQvFtu
sJmw6AjWUtfbYNM/jgbS/46VsPtVG8qBDe5RsOTsvbS4D4aiJKyRWBYBdgQx/IYcbuwhWgDKLuyq
atpohbcuStGw+Ppm11I2KhWTpGV4veRJolyW3QcLdAWKqzEYQbseVfRP4NOsXb+lld+0dYPau5t7
joae1ndn5tdaVrz70WV6E4tTM1EN2ie76HdUXzp2ihNQRhSs5JrnyT/eBKsTrUQLOtuRw5b+jUJo
MOWdtmKDDOu6DS6dmLUePG5K+8XiCyFFrlR9pkdPUfeZ1uMwBmu/mbcyZQwZNyLxH9wbfdcOz6Pp
N2DZOedzdVk9po2z1n/jBG9R9lN7dIH4xlrHfjuDdX57LflzNuA39IPvwK6Xq28tqe6i/EEzNraN
nIyKVMRLJsD7IvfgHTWi/FxWxRwswJHw3GUrRCEBb8t3V3sTxkwMkVlImyfxWd8pJm87DZonNUWo
Z/9sWAvqq0ViLe4Q8w6o7vWAo7Cbj/c4pwQf0tzOXTLTBSB9gXIJIkKgTf1jQ3W+ZdrtI4Fa4j1g
mh0yUl2fk9ROnJtoy8IjSpzCOw8Frysha32p1HILzgKBawBgf8CTUvTrCaHgU26h9lcT+ea8ufof
sVIYhTGtk928P6Wc7gbVxNOaetfhTH36igmFCTUB3Ae/c3JuVCwh9ZUlkIUAWY2xJagNN2zcG0XC
FT0epkYJAqiqL453QN0WN80IFTQZGdJ+qJOn8YwaS6rXnwDJ0T0/FJSdMlCnyjN9sZoAETNqi/vt
sha7vReDPgr/kabxHUgcXToialE0mzxDMzg6DmVmvlGccem1YghuYV1POVEqkC8PBfNx6LnWd2Ew
CcUKdX5Y6GPO+PGJC/x+KfKu/bniR9/WfDWmi6B+T76sekd0o1Ux+q+73GvrU+/JvPZD9Gu+xWKo
wA/VIky1DYWpq9CVgF0ay4JJuwqQYcxpSZbp4HXb+rEukCmewBJbwf5Q7MRklpq2hbGf12371skA
PIlUyZBjFrksTxpLBFhIPUEi5EBttEE2Ha5/8+DjvxEOYrjwsUcBWgkM9RETHLjGuuwlGf52tvGa
a08OlkEcgEYEYTRp+DNHo1ap4a1KmgynDKdswX/q8DJAx2gSjnt/i4+pYjrcT17mpYm5nPYcKDVj
S3PHs8LHh+V1OM3438CSnWg9RVD9kNG4Rwufjt0t0isX6BxNNCN0z62EVGIcY9xLtsYOapP/fpdr
IS/yjdbcp7psxCxi8+sQNRPVvYNbB2VqqhozfW1pQ6rJL2Vup4GFQtrGJ80kPg85mEFq9qzSiy8H
HcReEuW6pQrqasX6KqOh/L3uXqicfN2mYWPejA1x7cmdKDkc0J5tYnx0mjgAf5jDZHsWjR0e5TAY
N6PwgyT/1FLKjeRYKHFwXh7DF448y9tzxs22LWY90JxqaUISV5gazUY9YmPFQJrrWsyKk9pLXMjI
jsKt5TaZwXpn7KU0FXOCU28kikFSp4xhj9UZ+WqiJj9aG+bkC9cvsysMhs7d4Qx5fZSi+xDv+yNF
EtxDrIz4XZhsGHxZMqmUa9wt80yJROmJaJTWWyzx91bSt5BEqdm5/DqAV9DuC97vhYkm97Mq2HSQ
0UcFpldfpvZr/mIirDBOJHCilpeOHYe4fsAtgE7xE5YItHO6itUbb+8o0b5LdESdKpajlkeQ5zW5
ZRsRPgn03EvvuGVWJv0+KHtEg0JarYY8LG390xZhLUqDPu2bE51kpnWu5qhMD2ID8QzunD/JLFaP
ayk4XeTYkj7CVvFrIKcX9AgbvvI5pf7NCVs/nZg2FCegE6pqPS4uAdoJWZaG8FYjAxvcBGgknlQt
B8PQ1HLIOVdcnu3bWMPbP47+pvXyOn7iubVVc3XqTUs5UltMX0fG7nOvnarmCh2JChCz5uHmnTiH
w/Vf/8ge9r1BODk4xJaFVsh114yUbdoqUHZi4YPHK/c06klgb52OxIRcNRZx9N7fbLHOWORtnVN1
X8sVomibKp3B2L2BKpoxdBFm4Ly5sAvmwb+H6D/DR5QsljUxp31p1wXNw322wP0hzLKEdMApMtry
xo6C9wQwJY50buQQ0o2fYlAtgplrcRuk/7j902e2ZxkHuyWmd3Pg4wWVl+60vJOEcjY7/vpyakUs
BY8uj6mJo0u4pOJIZH3TsTsEtcx/9LZa0bI2FEI8MU7fjLA00JV9BZPcrNeUm9TbIXHrLKA7n4SZ
kZy8ZRTh2b10s8g5BAjWYzJxDaLso/aizFYqSLl6/jfni6KRfZCkukedhnW6uvHwS7weeosN+G0S
XkaaMyYMZGVb6hkguxKuzbhl9cEU1/kyxnkvU3FiLYM5a4R2wyPAlSFJiUmcgzt+JPydC9wdMfuj
jHCpMDP2JfEe+2SmxRYO0SphxS8eZJZoxF/mp0ktpQ2BamaV7Oi1OiBxMuiBgmf/Nz29+BMpOVjX
GVbR+bGDqpLGO3EIyan3b/Uglg/kVRkxxCTt/PIdGfS82CbIrxVAe177iZAIuCieI1pwAalBLjBl
hqRB+uzC6FAR/fQ=
`pragma protect end_protected
