`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FQYqpdKSALcRH6m+4qu1C7nBDJVaAkf74yB+aakpL0L1uoyBihbjurePOc7uG3Bj
zdNRXtCP6q3mEDYexEN+Ee0WWvWYp4gbSokveXdWe9va3SKsG9u6L/xQgSAI8Day
3CbxswyB45+YoS2M09JyYfARiZ4dzf0mU9fJPfNTHGk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17648)
5rv+aJgugLfNh97gMk3zUTwvMEk5knHmLB0SHWJM9u5uMzTYspg1YdJS+yK3d8cA
4aaKfniElkJ9cnaZU0aiDvqMfb/4QPXHXaXn2s5BIzhI8PdoghhRAhoxekkka3z8
D971dtdsoGey2zTK5R4OZ8TrxFYwGR0wFgNdm+ecM+CHwjO13oE9vSCs3t0mYo66
u5T8RolJcB6g2XHPLplRrzszZWagdDk8P16tkNVeZ68llY0W/Smj7/qvi9ohq9Pj
5FHf8Vk8pM7TiFmlZoImeAdvfdv6Rfkt8kpHgEfFFX3gUa+zdAdul5OZSz9Ugf8l
d5B/Y1bd2cdOQRouQ1az4AwRpBvc1lv87mUbp5NXsws6+3ERMvZympZH5l+LdfM3
LnGFpPepVBOlFHb3VE1MdHTDiKEyBfm+DhpYCghkm+ISTbB6XvEURGdDDMCCZBmR
na9aM/m0/jPGasH7nptRf/9ueWxxXehgi2BxM0c8X/3JIyoZEohtK3asb0CdLFqd
I6cON0vJqN6VlOoRp0kuW6I4al6QziNIOPfFYP4wglwg7k1wQ05Pmvc4L0+vBpRG
AFDnH+F/2roYY8uq0BKlFzEp13DlLgbS48F8fNFvtv3BtZz6TlcDhKvQqtOd8Pdr
G4qJrRCuYygM3yR69J//GLidWEjlAE62lhyD8z+deZ3zB5PvmqIgcfFS69oiUVpr
Fpt9Rkms0xkcXk54rZwtISMtoU11Bea8X9XK62mwMkXFR6A1gSoLGnAzXdF4s3qc
UlW0NeoXfDQ4MiNP9pXdRM+fZsVmsJT8etaYspxc8nEjMHsydlhKf3G5AK4NOqpe
9VNhSbbjH1xrmAYw3pTEN0pHQCJTJZf7mdosqeEp7FTeqoGMdJGSLK59WteQAsWi
/eeNyUB6vLVkxwwXJtROyYmgskxZvU7MxUWCNHNVpWm2450OjsTHXGhb9Ar8brJ2
PuVrXblB2kwnXL8bEkOsQNBdMrqUhghCoIYjp7MuzlqGecxG/XugUJzAcFszxu2A
DxNnjJU9j3inFBpY20mDe23IWRqHOYUpanGqz//D6R3NuH2GZ2/v6yu63kY1hAFN
mzkUbx/Sg5OHaLtoyPP5h6fBnff2JsCTlLlsozaEFW1afhS0mofj2k45COKzKyAE
gsIUKai3yN50N2szMrPqlQdDRxCev59KEGu+hrzq1nHmx+F+9BN1R/wYzFt1QngS
Iem46itlp4w4rHgez2mrI2mfAVxewMweOD/L9sNzdReTnh2lYr2nP5COXSChg5hw
0CQ4esLg0FN2546wS8tu4N2YiangB1L1CW/D/hMSi3eaQbJCTbV39HNCWrSGFRPm
B2NmZZfvHtK+FUQs0Z6gtLCsvKHACE6zRUwzRgt3LadwTYLLb35Knj1oahhuUxA9
gbNfIPzu20T5Gp3I/odMVsC842myNwaQi6bqCil44mWF2taTqBDoVg+JYMfqlsSg
F7siKgSrdUEvyDkEmWJz8DZ2jxXZqjubRhlCj6tsB/KolLBx0kANSGAQDzSoB59T
LubAE3yK/3gm4uPR3Kuuu909oewfoDD2r0yKXgeyhEIggp2Mv8hNYJyWzMVyFC+o
qVr/v+Thj6x8a9y9Yn4BnBkSVhwCqnvBBRdiigRub084Yfu+haNgtJhDuVe1a0wy
xTbyaaS6sZLKJrOIWtl9Y3c+JVszRYdI44ro/O0QfkQk9MWpF31Fyf5lqP6dQV1E
nO+0+XzyxuingaSM5BLnDvsyuLITygvXwOtaL9Ro6RfvFYY/Nt5kjOPDL4e9O7jF
1w1jBT2YhR1s7eVq7Skd+DdaB8XmPeQhdkQL4yOyj8pVIYJgpPOd/ng6MnklVMH+
GRNAUAlJIvHPoy3KXJEKqHdlrKs3lSMjL+wm4cCIMF+VI0duA0QywAVoWdMSUfiO
zJTXBbDUeJKUoYxe0weGS71pxH9YiwtywjZHaPNwbEx8mbMZ6vdrKTjydVKU28iC
TxmvRRxTI8QVscH9GEungj60fXo4zbny7YtwMHHhKj+XZv/4bQNxWEYY0Y1gDtco
eBCvsYZ4GTClBMMZoB1UGvZD2s/EfZS+TZqt4q7wANH8vZZuevZBxS0UUFYz4IsU
A1aFPefylZLHrU/a2TLTmjof00YEOoKXtdtcrirApWx5e/9SxOdKFaVxLgH++b8U
pxX6s/2CNqyXJyyEiFb4z3OJzqKFp82lWoR8JQwmm0NcltFiUoHcZFY5W/b6Wxa2
CqD9Kv3vugNpAKTPnAAhgh6Y6vVBA331SjPu3khMK6XgTiyXL62NdsP/wo8fDAhQ
4R6U0EulEQ1DCgzz1lWzCN31jz8GE+PipLg3lpyabd+P02g/77O0T47guKk7HkI1
bECd3dfZ5Ye59kp6xzzYI2NN54MsL02gK5qlY7sYS5GgUXkqkexQYffAJpmcXKMQ
WnUBvM51UBcxITbxdhjUjfQzkM+h6e/zDeMDCKaDvFWMIy+0V7fHdVtgT7XXUZaA
3ALf2b/y0Q7K3Kmdi4+kWM5NEnqA6UdIl0KeUFAXsjikgxYLrBMhs7P9UHB8JiWZ
isaxjlLGGMWw+lyy+n4EukMjP12B2hnI0xYPMZ8eTT8Hywby/8tad0UB69SPsKBw
3gMb1nSxvaYQeth4xHspb3O99TvDh4cuiIYfdRrncWCtaRlyjwQwArt/Sl89dRNa
LJ+tfG0BU17GA0rk7jUS2CRw7/lZX/SBRazrYu8NFuORnh4zeLMEy5DqSfdSI70c
nuYgXr+nS6DRXGDVMWeW/LO9tq6B1qzS7xRkn4obusrkS/K3hfqEHZ8yUwhwEC5h
d76FRTMKO71dLYWOBraKZ4CsHKohW6WjqYaZMXBn8TGZt7Aet5TxvWALK0Acw1lu
SXBrt8tKcA5z81d9w7HLTkvMpnfC6bF5QiKikVp9Fp/tP1dbGXTsRZr7oJhH4/Lb
p2deJx7E5aiU3MklFLlfVUWCL8F7KUZurjD47GSKOh7QpYKVjGE3IN7i8YEynfy0
bh4OMjyI+Jju8FAO2ur314z9roOnJ2hr+1nbQoG5VpPczES4/QUq++cuC14rj/ah
othhm+85ChEDchf+9IDsxtqWre+F9iLzxFK6ZGGgNsvf9smVX/YRmvO/TFjsYgRO
GZfayROLf4zTDm3ic8aqh5YtJjmfCzsKPaAuq2yt203KTlWfSiTJMxzoxHCuwSEz
IP9bGJGOcB+6LDXFdiMDeqG/+RRp0kFyRX/0HorANtlEUWREOZ70u/VklOFpe1PD
6EcBY6sDrpEboBRTIVNI07cSSY7UQcWf0lEQiNkhDgvy6BZ52BarLEBuf3kY931i
P4N+So2RJ+6Ve5i/HQA9FnJem84TifYQl6nVu6JIapBvgH9Az+RiONp45YzW5m0M
Mo27yHY+YEZog5zI8zlk7I0TisMrzw2Tx47qQRTKbs8G6i3GJ3EYoV5MRmsqlOeN
x2/p3xlXx85GxnMOqvS5nx2bQNa5x261xANNu8RLDjmM19Wb/TO1rAlvGhkJlxEq
/Q6zxthbLyKvnqpHYSkoSWm9MXzC8lWjVgyAwLMcHb6iJm8U2aduMzmKHs4WlEZY
neQYejhk0w0yIFI+xo521HaaLQ0Iph6qDPHcLkvFqF6E84qgNNzPGt1ezWgnX8ym
mT0E1NXLbMMv5nGUEx13L6ylgAQNfXs5Us2f9dbIVN6dMvRwkcOZwSosAK1Wyexj
aOP67m9LhOddYa9dW6UpGLq8PY3PEjHLz3w4xmLBL8jdhInYY3KF5ZDnsonwEarX
25fTeDMP/W+3NMttj0w1pCYBOK9Isbs+9AiTh7wst1zEF6UJOvA5UjLuPrFoJxKV
3op1d19uqi5D5mI1tleEj0pF1gMYAJBINNZznxv2Fi0GpvubuMmXnVWCvtWOJrTk
NrCYn/LGhGMob1nJ7yXClic+Zx+mC2l95bV8VhJwIENz/66fxFieD6ibl9xz22uQ
NbPxS2V6v9LDTn2CrLuSOttrKfaeLo6jxFePTP935OQVrgmspfHDsZsVKatQtgty
HDn/7I8QWr5XqkPhj0QhCeL5OZlP6fYdn0Fgr1GYxBGjiHZP5V6bR5muyHxPAi8Z
jIlzcz2wuiYu/SeM4FBoMb92I8lQYcLCIVgdA8pKL+M5GjGzoJdaZ9fgTsBGK2Bh
IKvFdr4mLQPeDpROhNHGUd+zcjXuZxbN61JOjuQpkfUl6CFO0Kg7al4Pd+/i8wgH
kNawkN+D3yuE+sCxVWA3ZUlkpgOf3DLt3cXTkheJsp8usHz/oMokdpaCTNzdT+i8
p0IJJrCyeqrAsC8sxwAbCcVesFVS9FjlyzvrAqSKpQCWOAIPtHPBGJi4PNOhnyIg
d5jg9oOJDit26ZryAeY6/YxIOyk6UB/49N6y7vIzJ0tq7e/NRLD7E916tBkUaKwG
qW4yYUqFQ3JaVOWK55ZMd1EKvNYEjyksPc9qTEtG49SvGz8RnEIQe6BNpReIW4As
HnI8/7GUoHQfzHan7pipi4gCKxqHfzlWC2SchS+w44rd0BEFxs9kosD3dt+YsC9L
UJ+SDLnAr/gtDPq8Gynud9Z95f3WapclhYDAxmUBlKqSDaDAzhLxvLNX/gnRldW+
65GKpnoV2zpv6R/9WL6csNcw3dMFsfVRL8pj+eLmMvCe221vC1yh7Cfq8Zf28TbI
Sye31EQevNJfdTUuVA9mwRX2DeCMBjjRjGMolgb0l8ifdSXqlpaUxmSc4R0k4kAS
npZHrQ+teXBPy8E/6k62AX4N2C9h4qUl8hgfZ421DbHLIjqgx33dXcjOaLIb40NE
xyCpt9px/W+JsPiQmeFtpEirFm+qcN2jX+gN9FYgcf0TV8L7805sxhb4TeMVRjwt
oUf3/bo9phGX7glNGkuyjvSE9ic+mMaf1rZfdA9dGmC+tnre6fqjHkI0A4z+AdDL
QPr4oqLa4w+mpVjqHoEihW84ErXcDassDQjBot7qy6+IW2Zwg31lFG+j0OQgI4nP
yq7mrXfxQh+7XNJQlQxoKc6z8VGyw7M4bX5lLO74Iy2/Icd68o4zigkYPjVzu8lb
hLRo3PuVayhJ9tHeeeRCK0nnbNVF0JWrPPCFBQ3x97NMx3v4kkbt3aH7OOC2Xiu2
jsN9saFEOydRqTcQN4fmOi7lFNfIfPUi3DLK5ZE/lAfYAKzAD4wKCYh4X953Cm9J
eoMR4TV7OO3PRvZdwPXBM+HfvKakyt3lYYU316/llIGSSr+ni8K9CDGqw9x07qp+
AD4ffF6KoSLVud1mrThm/M7SkPJXkyMfToJ3inSnaJM2bbuSkRTqw4ESQG7ntTdB
ZhjLAWqUI+Z921urvsYyqZEMz9iR85yYc25ca5KncgJ+lKpoP0CdfWXEvw870ZgM
/2dofW3gFJgkCfsZK+YXIy0EE/NoeaNfxY8V+rnEU3V+0cReDEILm2xqHhVYBbgS
J+E3khozjRPelp8nFDBtEgjexjQLwlrPI9Eq+ggu9vK8M4yp967xe3XVFlcK+JxL
K59MDyK5ZpnKXPTtulsTQ4KnzWSgAFe5zOB391WU6dStq46KCLcz7RGuqbDE4V29
quM944BAK27nJQtjTEIP1KPwGIHbCjFA7dlZO8pz1n7ahler6mXri9qHoH5y6KxQ
0lkvvw8wdMFOJq193VB6uIlLFFS8rDLundj0elgSwD+OLNQN6MZ/7GMy5/QgUjB0
1RjXotgrWO13cjMES+nE3R9PwUM40hHY1uuJpmPWCsVaR8jpSqZLk8TXtp06RKm/
F6HD5U3PaUz4hg4UwdTntawXJCz/pgpnxZiAdoGufKLizJOs43l1mpEdU4DlL9B8
KaBRU4RWbhsOAwpGMYLglgysUyU+YNdKi7tcxMQD7QbWckhYrTczxBAp8DnRS9xO
p4SOZePXilYOuEm0DxIv8JlCwmar0H7DjvABpFrsDm67n90JrFFXhfjbZ1CfEUJf
rcEYT2jxw9/xhMWw55lDfGOiFwbGS+6Q7TPXfNs1fr3KnKGTPb/9xeWHcfsrwXi4
8fmNk9rfQv5ld/Qx0HG+RxEDLpbP/aF5/iqqBGRk8G1sKkrdqEvEhORVNh2BWbe7
vFCWVUWDm70YSeWl5a6bgsxw6yF2ime++8aww3xB0WoMV3E9v7ccu4kY7PwiNLwO
8ZmnzZ/PFpt6NqzZgyZ4tZUIZseWHdHIusuNfvf34F0+db+PE8x9VyDaGeyz7om1
xv04uuWfMszMQxZDywBZzoVoYVMLPLdayYyKG51eo7PU8XFKx5NdDu5Izkcq5Cm4
sEEQcbHHBM+gY1dr8xfgyH+HEJ3gCezA/uNhCrdWonxXCR7Ukrzq44V6oQeVYs7d
ptpJttO0EEwzzHeLpiLy4WEmz86m5ZmaSb5XdcIvUvlUIPzFa5aKZMWX1KcQe0zE
cvRs+X+vLTcPgvwEMmpHIuTc+0FSS8MGnz8YLZeK7bYcyjIL9nTvvmfjrVConN6g
ANRF4jeRjR9udAL98NCBL75oVQtSE2bWjZaAjNKYnUoz2ObLyOIqRu74Ya+is4Ap
Dmd/Jo1PFpOT3foUJOiY0NNIquxyQLVTXkioGByv763ioUnnzLeI+CUk6q/wpjny
cx0xfezT/BQNL5uRw3G0oH627eRfcdeaxWPsCGpMduPrCw50j1J7PRoZQ0IJ6dsR
rsjZZmt277fz9GLWw8ciLevMu4+sY6q6OC2VPmU8pq9AKPOLjfr4Gw1uhLsmgkdQ
VvFkR6XqXoS0N/VSNfjOBriQorSaKBwJHmTMIJjB0qH2ubmKE9YR45HlIhtksPS1
JmBaC1NaemZtQ/jFRV6vmW21t+LShenA4JY8/aRZJK+vPjxW/RAGaNFPhXKh/mij
289ez/6qXqsAm8TPXvHiSuKBpnVdLsRmzCKfKUMe86CN5CiHtX541W9T4P7G+c+W
TtSO/jFnjJ6M+e3/m2ToY7bb3FhlNbl3FerzuweDbDhLs6yOYKVQHHXUF0LseNUU
t1bYxVIMKRnmkQm+QXXx7M2IQCKesLXX+MoaliMFluupny8qNC1XpXrzUYFR8XVK
3h2GW0crP+e1QtnUYs/8FvWW6eDPxXS/j2Z0Y9TeKfnLVUrq5uz84URvC6xqSz3e
TTMy3pO4KoJbnHUjCQo0Nohpf141WaEDDDr2gy7V6cYe+1YvgFjdql+5FQ4fe2w/
+FH7iHoMtFHQ1WWPB4la1pRaKvq60qS8+WF0Qy+ZF/MNIBwNuzeZIDDo0ZJBv/AR
XFBNL0ZAEeuFG/c1ab69osnP+yAWLisukYmngGm/OYWKKVEvTKOFYPhZp5yQJdVm
oQb7/vCjCb1r2M1fjFmmBNZ3z8oYWGKk/I30Qq/C4gQEKcPHJhUOD5oO8MhkVhRA
ChwRibaM749dNeLjcHe72/GCyyAMaLBf/jnbllvBWnVZTXmthowd6bbuUV9TL46R
Oqdh+VVylPqUpuxnnPkfBjy/7eFsPaKqA7JNx2bnBwv7et3Mzk52Lfe4+JjHzXLX
vPx6QITvQ+30WTsmlAlYwZdAMrSLg8JtLLMjmIaBJZIPb8nmkWAJo4SxQMaiB7Pr
A7wLzfNF1vE6/N+PMH2PX5KggVoyq7awVwjIjURNJEBB4VA78/KwMvG1y+DxVl2/
q2jXJsnhYWydoqSsFdfHYgb6IZ3hdPgl49SdIrVTBXMjnAwt32Iv6RO9jPXQep9T
3D9vifFd4/z8q/n3OiMFezJJ5vOK0rBzpbBRYtE3wFQZmab8dSGjFLMBC6jy+xbB
AIQqPu+AmiO7Lxs24CPiRVhUZWSttAumSil0mAGTl62GLUhwuZFT0gYwTY7zEFs7
cANTHpOwEeHj7UsRQFyPoZt7i1sE/G3qyrjvtuf8X17ExHO5hGz7lmQYzok4SoV5
LHpczXuKc2gJKoxjoAevrjQsHw9T69kOyiOP1ygULXMQ9+ra49bD+5FFgeaG5xb2
UX8b0tLqUp4Jtu1ZxDqKD5CJOKXvSQ1HV60Hbyc0TzZVA5fD5L8uZHT1PZ/C5Tsl
UJJD2Kf4phjCL+nzvAvStlYzWc/NkCYVQT+veYT0Mq8wK+l0vYZlV+V6yLKdfGkD
+zX5LDxD7fIAlpcnXNyRX9AjucIV3LPVhQ1w/gcJnRydUiH078TZ16/HxvLxkvm2
VRhhQ96qiaOZ7sTC+11LE4jgjcPGiCtRjDoQNeSVTYSTQpJChjazi6909ffsIq9M
0nd0PF23LhiR12ZoRM6FH3mSBnyl+a8lceaV9Dsu+HIO1jkw/IW30YhiqXMm4iK6
U/ZIkVpSIhPsoFYnYeyshTu8TXn5zPe+vnFVIqd9CPZjfS0mmsx9n7GLZg7ngOXj
0LVrhuVACkeXk8kXxVCYm70GASOEHAElnS5v192cEI/sN9vZTk4MVLuPuS7hcb55
G7AEEstofN3+ubi02ggRjUKUl7wOb0i3g/pk3Kaf9OP4dfjOke7zpaF6ITGn8j32
IZ75nc8fiwiVufVBfZVw6d8X7dGLjuXCsVh0USNtzS/cWIaz6+gBE+6dXgrvq3w8
VMvStFgM1B7GiBjfD0wMtg/NIybwH3dPgL1bGaaIo24ZXPVzRsp19BUBbYDaps3g
1uckesKIpTblCd53iW4ORK+JQLKM9dojvmXwC9eEOk1Ag72e5i10+JYJs189L3W9
v2LyxbhZYciJ2iOJcjK8uyoS79U45yJqe4qlZ0GdLg1DiSQaoyghIFgTAvkAxpZN
z82ku9a6Yc/6iN3qLIKAIwGit45UGv6GmGDt0b2MaFnmPPt6xKMEd6ClJ/zRCS8d
E3tGEzgmTSD8SyZ66gLMukBWRSHLiCK3zuk8AuezuMDQAO2Jo4Vd4QTFOb6Tk3T8
SV3ts+MZyqm1MQ/+Rsi9Li3oud8lfjJ2v6dVMJ8hyu11Owq9KeS2HPq36pYM/QyS
Ee8Gi2CKU67rRYWSKaleFbDAIQjQarmWI5NrwtLm0Gb/4+tPCyhSWKouEzfo7ppP
6p385niyQ4qUzsaHbRZu8Si5ZSDsXFH/OeCx3rK+ic+VFrl9ppy5YvmPQBN9fbSs
LXak0FtgbKFlcurZso4ozUCUCHRT4MT5Ncn2VCVKCRwCUAXBBy4DomeFP07c9SW9
eMRDAfRp396QoIpCXgZiPhx3o6+CBwRU8y+2RQTFbubZC9iLFK6g01XcAjt38SwN
LcltqjqK/hCfEU5ko5i6DSru8Fc81XP3f5zEsuyww+1bdRwGBaYJ5YQx+HWEVIyQ
7GZBpqDWJXewCxWR6eJXiX4NoZ4Ky+ObyMncGRMr6+z2iw1+M+Q8wA57To6s4WWZ
S0lwV4x72/crNfjTemBQYbDrOM6ppDctxYqlk/QoVlB4JdDn4ZAn3nFHVCq8HcJL
u7+nIJvSVIMZR5+pzGJVlLqYz4pwW31aPBlEvqM8o5dknF1+X+QZw8P9cmJpwKoW
nWd0R1ycwVqeNmz84eUGsB/VX3mL/UdsQ0G/abs+0U+LPfehvRPSx890aDiA9PFf
kF0h1NJqxh6/6z1bINSgjquFUOqjGFURTGKtlJJwN+TA8W5cURWqcgVZoAUjsaJ8
wKO5AycCZ6pOcAF0jNe3YRIziYmH0RNVrwpm6orV/8HpuNY6yZEJfZjeSDMRV7zu
+nZXyFERPhT8QlO7e88Re0yLkIYl3L7txtrVAEEV/p23MEw86NMsue6ZA8Sh6iQ7
daDMQZ67zDRsRuvIKr59OGWOE2xuu6PlIlxSxvJvjIpIU2RyCfKQB7xRt4NIT/W7
5VDBOH3liQChH53Kj7LMzli0ltnLHnvaj2txWrms+Rkoi7habWDf/g9cwKfZ+9ip
uchO0ySVdZX4QNCMNZdIXVjgPfyqwpl1UWMWkYWS4KsSGMKN1k4QgWedf1evaMje
HkQt0QMAQdadVAdOo5TDc+/0ZBaylH+hMMKQZ//EnKexINxjvk3QPkMPWohyX9Lj
Jbiie8+AJCF0kOBx46KIWOCkSPzVafzAV8z+AdWE4QxwDGJs9KUcmidog9x8SdLW
cwx/isaZ1B6iCC6nPsorZFNeYqZ7zKgur1rf9okpRkQLQo43CQ/l1Ey1oq3hENuv
L7dOOkXexui9heGqChBclpyr+oCacKZ5bdd3R7TvxYOpBcXnjN/IOUi0SgO9ToYc
GfGecaILqO9JAcVpguVIUGPhhj/2JFlq6pacShlMqZNW7DbG+Lmlfe3GiDJW93Yf
+t9HSkl/g+XcYpkUhDbfsywLNTaDaLV9rqhGQZiFN6A8/B2Xdx9+KI3Pi615xMFY
tbssGk5PB4I3bUNFqdFOu9l5vhXZOLbX/epOSxoOwDvAyls723BdCBqiVLOp1Mh8
N0j7+Z/4I8HVWiSepwcrVxQHtBEQNfivKQVhkPFNUVMiLjvNr506Ps+wHvSNm+H5
51apCF2z5cxoOuU1s3Rb3zyEspMLDst0tXK3rl/DgMz5ZN632OBqNa8QBVnn7PmT
/S54ok3+qxDKaXSyyvJX3U6pmCP/UirAfikyT+NZAocsVXRF5rPeGoVjBF/PtSOd
FRGTG/8is1yayy7zjOmz6aSbAvv+mb0N+xn+ov7vauSPTkkzHYPquXNlEUZJ5W3X
/ce4FMwRmYH3EpMmvujxHZr6z4LZUBgFpPbtSRKZlrUndO6U6Ot+Kk3OsZrujLxE
nUdYNpadioEhzSDhRSa5msKBLFpz7LvAa0siUGw5dfYOUbj66Thl1dQo0PY5dExR
V6USnoJKpG5s8nzSRM3xpP8abyJJn8U8xLP5HEktbMC0j+ct0dfPnzf/Iq3N/MqN
B3UcwV5uVVIElc4+dgi1tykJ9lmZ/C2lANgPPV5iQR23lfGLZh7mHN0CsNsqd1g4
iknpV004tyOWob+OqumenPtov/zmAZcoNFcT6gRGlvdeoA6bPPuU+hHeoizgE8Cx
ATbqZmdygnz6htnMY0Kc3x7he+Y7rUo/M0PcV+Fp1yCuK2OEG8h2RSCYc6SQXnPM
4ezb8pAi7I6vQjxQyePhtwzbAl1DvLgQI4gvmn7hDieQlB/DMW9YUPQfd254yKfJ
ms3q6jptVWhawGwqL+nhzJRKTrW4fW5VT6+9BtR9yAMqLDBO5o3jXZ3b/K2VTcb8
OsbpKXX+JhjDyrE7JxHeHWKWtKRyERViwFxneIyaQv6VPUCzkOLEK922uzB3QNwP
0J9Ckz1Rup1+CvssO7a+nra4BdbOhGgpmLJJsrFPFfsRO6kYFR/BM2l0duWzkBpr
wdHRR6Qqy77ALVNlVGcq3NfBJd1BsLT8xyTbyAwW768G6w5h7UP0IwvtzdSVDRMs
nCa4jXBy2SwkVDHu6Kza1GTLrEMp/GjfrFVc6KezC85ojWvnkm5hoX0gfu/VaYQJ
SeA4df09wboWvj0n1Mgyxr12c3F5L4jCHvvXQKLWaHgpPIaT3pNs+7c5IPTGSzbc
NuLV9b9Y7SyQEwnPzInqeEdh910/ERLvK4UF5Csnwqi0jduuYNPisKvo7NZvMSBy
cGvPBYMXHMurmg++KbPHSS6y6GPMjmeag5DAqtZKYEzvEI8BR+tOC+Tu9FZeLlo2
KONsC1/RY8K4K511Ysz4yMyIz7U8NWb/9I6I6Uq4QEFuyNtGwQXbBzMqgn6i3R+x
tDcXxl5ddvMYl2Yr/vDWdcrmJ6ZhDYrQBEezXVQRl9lR2LJZXxUm4HRxJ6Ec6Scd
Ilr6kaag3NUOtdpWii90YMBSQOBOxkLVb9XTD8nMXGee4aAJZT/CoSMckCki1KF9
22ElsoohcN3n/D6zRlXIO5m5aliFZPMb6+hsBXYIRnpL45Eeh2iIa/SWlduBlrI0
fy3vhGKHy14kkGltCEXn+XCOTTW8214qSx4OUSgRvkyNn8pX/lAJz8vw+sdrRmJZ
WyY2chg4QV3yxxtbZpiHp6AtRVvghqsifKFq0f17lA7+E4aabYJUC+bx8j6pLs4D
2ffSnIg4DsEDqznjapw5gKnlFvif28HCsG2ZSASZvu2m7A7j2Q/HIFdMCEkOEm+z
1WmCxYv96UdxqUcdj++OjyrLy0W5Ftx6C0hTBV73BTjmI1B0koTj6jHVZ+pBQmZY
0l2Q2kmZV/HOmDnN/5kuJSmVRe8QpH7WAaxT9d9fOM0V2tSr9PyehHpTjJXrX7oH
YzALOTkjOGtJ0oU2DQn1d24ji2BtQU0Y/ttGab6FxslVF+/thlWlPMSVIBIw5wBN
KjqBmt8zX/9SboPT94Tjgw1jqwYfmP5vjwdBzdSIybWkmdKqrqNQzg1tXVBDsrQp
718qIfIRZPKHVS+l1l8cWoHOqv+XR7/puXyn6TFZCK+MIj2/wpxBvWJqZ3YyRZYx
QtJUgAmXlNknjCoe+E1GK8GfaVxdrPK5hJ017K1gShRHYCvobcFR4QOq3b4W15l+
7a/RElTdx3n922L0rAuiECTI1C30PHj9qf3XV3uVR5UTIDAYUEwjYeQoNa2Ps6UJ
lsYMpaBReGgugixXoep634kMH1GlXt8LTPycTnOjqQqGs1qpV3Qk8h6IERbTlevg
ZEYLuAHN1HEebdAizZUIaL61GLCApEDLm5yPX7KXaPYbRz0qea5FaRy7Aoje14+H
4K5eyTgVHe+7eMWbyrGQb6T7Hlw4aAmt3T8IfBr3Z0x0i/nMxG7u760uxc/uvxtS
mSCddyuRKfiNlijse6GS/jo/t/lqGFuO7ZjmF78fg92UJVNu2YbzJwUV51n9qRx/
5iZX/oQZ4pED6bEzX4CQj9RuVf7hbpzHNC1DhKK9aFYaMd3tTjTy8lzl4WtmGeaF
RCoy1sqaFEcUEuAOOV2CRcgBaP7e0gvojirdQsPlXSNOxLgcC+keXM6XUjzcFw+D
mgUi7z9dK84KfrzC3CA/M/K+uQwL+8KyMbzzvSq2iYVb+oGLFRUZs6m609oayrkW
DHXXwvzZqBZnPogu96ZuRYrPCNjoGlkPyuzdDAVuiJhKukyTDvlfZFLzH60iC0AB
C3VEvEQuLp7/+ueMZr0v7rs31Lq+PYTkLx5GDrnP9+J1sGeu0nP2wDTyh78zF7ic
SIGQEAW8CIUBI4XDRDXPVSrbnES5f+Rtj8JutIE35lpPNxB2oU6WA4G6Onbzk+cY
erojO7xIrqs+ofczQxOaJqiqnN+bniMcGHg94p3FxRwtpd9qMBVvMYI5raC0Bp0/
zFitgrmixKQl5qsOssLC4JNJZ0S+W3NXqTZ9GxmvCZe+yGLtXrPKvgzBLo2mNV9T
jf6DMAZdjhQ31E5y8X9dqL19QioLDxB//RX2Avu/EajY3GvsESGXcnZ+0AFfuNaW
BB36K/ucnEwojkfIFcaRDwGbLEqlsSFKxkDleEo4MXDknnR7Il9vwwNlyRESLy4u
DQ3232MvpDf2TnTOuMitSIAoc4E7ZvoLn9Xvb3MwS5YM9JWnRUgnCdcl72K1zuzB
WHZHNmhT15iydrioIQrtTS3wqS/IACq88rP1w5AsNfBEX33HWggICTDgY3CyKJWL
Pd2iawNcyQk3VDawhMgQJVdT8gky08p0WR3DbycWyFPbwxF9dMSlVdDUoMSl1Su+
P15VGq1yIBNy/bmmrYKnWK65uakS7U64Nrxtk7gZBqaaICZzOav4+O4oJG8r8PMT
7SsDWz3Y4Iy2NN/jKfmTc0Di0dcXHXUajAHZqImYaOXq4uGCkTKPDVeKmKByaHMf
1TXWITEwJk0mvsrpLXqqh/IuGCSQbgfuarURegK47ogRkj5zNoI6Uj4v6xjX0HBg
ZHey2oxpc14XSiQSrsHZ4tDcKlKcPm5U1AHt+077pNEZsc+R2Aeo06vL1cekDskh
xhuXh1g6/SJRbP+zQAKr9DbH9DZPwhTItwxlaF7vQ9DKBn+u0cFqRLKKtLlJYz9n
qQcbPEeCa5P9Pm0jowqXLUWmrdZy5tsiLFnE5+TmASw2BmaxZO3bigcaX+JkiUwO
wKIb84oXLij+fGXR1mwUnuowPxVcFNYoYwr9/UFCgc2nXOrTLFr0XVYk0/xad/DX
iTt+I9IVN0MFQ9cQGTKwRKRodKXitjkmA0uY+PRbos4i93pK0MbP9O8uRzulv9V5
f4/Stbox7usPNhREaTgFFaAltVtgzaqwsQU4wTzp26O6xpbfmVPDG2pTRNRIjeUu
f9HxLN4glqY9IwEwNTkEMosb7W9uSI309EhtnRQOq0Srq3olUabGOgzsi8rS+EK7
87JoyjJKTcAb33mEhnolkPVrshSw0/+hM+Vt8JCzh1AGYbtt0/BgWY8CNE3l8mHJ
SBYEjyknLcdlPNdAgrewfziEKdBiJwsQWlUzfs9vzH80ebWc2msJwrBw0nqB2/oT
g1beGvaR3EtFTkLLxJix1SFafAYfKlmL7VEVG1FKYllaiXy7e/0bbvwnjj168Eo2
iOyiyzby0jT9T6um1qkRH+FmbSOdLhUmQWWXAqtHsz7/IrOhKVSn/o9QGilJpaj9
Nr2NmWkK0AwXfs4JhTcZWrQAF866wEQoGsA1NhOQTC46GTxQ13nc5txICZ7xZN/c
yW7jn2cXRshSOIAkF2tOhV3hLkGmlu1rYyyadzAI6pLhqfYv/y7fRvd5PSX9dpv+
J/EbepUbOwkOD+iN54eFn3nKduZHaPFXDKKEEMxogpLjfunpB7yeDA7pgAS7zPvx
KAFlpwTUxtw1jMe9jnRs4iHXmhQsVm0eV+gO3XEfcxTBGO+w++m/ZFkNLQ2qWC9P
/OQP1dN4fEKcSNSSFBFlNdrnE9mkn3udGMKR3aO/GH1esZQs9yX0zoCkM2KxCjzK
8xaSQ6yG63qhwDGUPK/4ggahB27eLJwo2a0ANZqtCkOGUZySX8HuqcM99/kIZdT/
n6qlJ+HB4nVIO96A531s/rEjIOezDwN7t5N+TqYl51ErEjrYnkS4PkQOMct4L9YX
A9Rgt71ud3v0+4Qhkg8OvLXBtfIxgy6PX8U7LduU66n1P23itiFZYLi/CNkedgsb
nofJg0ZYgjbr/KoPLqSNcgH3edaz2YhGssVhwrQ/SDSk1hze64eKQX4yVMTfL8D8
Pu0aX7n9+EtLCgretwdHw7rihZZXXgyTbexQl4ulZJfBofhTYEZnPZxt3oCytIx2
QtBO7w4kVCHnIIT2sTzKNr80zDbwzRoOHCasQZ+XzdOwoBjgkplQiUC9l3STMsgr
IZ+YW1NVrPMQ/I2RyzZ1xpyDFkcPxK0maelyGFhJaY6gmRf2YzEUXxuhATcVX00O
6+Lj3Y3b/ItyKTlVrsboXUD8KlesO5w6DLxoiB/gk1Di4qAMGvAWsN3tvqimnnpN
eiZNzkgCCcW+kl1a4pc8cyPJuFFyTC4DooZI6FSuZs83CKQdCz53U7ACFDuF0NyK
+BH2lL8+IXwNeUaGj5WlbhN6jgwBfJ+6cAs0JFNODOAyz9SGjyo3FQpNUzvwKREb
oS++5zT0PTrlEdTi4KVFHEWO9eA7/KFjbz9IXc778g9rcLU06LIPIWU6vEZf62II
9RvDmGkE6fufznTrRUO0qA6+7+lx5LJAGJyZgpTQe3tdaXBHLANPFeWBBNjJZdyz
3cPgqIRReAthuI+1X5jlm/zBExh6oLPh3VZuAE8PHvWHjmTaCFqOtX/BNI9d0kzV
o7shvE7WQo1KM6AFn4PlfHM2yTx5DUrby2oq/OUSRt/3P+s5d/7vv4zYtxdOh7cr
Mr9ZTZJm9d9xILSLH1lDsTs6p2VjAdDtU0Qcfa4Qs1Li6X92592ar6YgIGWMZu22
10UywkKzpbLQDgiP5qgwYz+zwQ36EsQGobfG6OPP4MswxG2ZCNJuHM0b4vG8KRrV
YnJY5vmk7EtDq6ZlCMBiW9POjmlJBJYxZu6FeAN82GHC7s6NoU38+gknxASLQUrU
bHhKBBdDbDsRGEOmag6JAqIDBRE9SELJv6HmWT20EXkx4VZlG5jI5++Ip5NIr5qi
j9x7FV5M38il90utPA4O1BaEXc5w73lCR0h5LP9rv4+gsetsNEzTiBeEI1peu9Ln
JJjf3SkYY5R2xZm6aie5T0Aep2uXMmWrcdYWpv5UOUwwlzGPZzPuDVwWaZlauHAl
a7pjfaFSEiusu4G12eqO08dq4El+HZ9S/AJKjVZxDFiB2fGF+53bH3m0y96cY8xX
bgaTfCbdsUx7JjP6La8kA/dfRBGoN+v5UZgA+39x/4H+k9GBbrTu1Bw4kwf2JAzM
QLw48mtGbs86bMm/egm0pOJ+aUqyxF/D5XG2raYy91yVgMzE4e+3SPkL5+cYPB15
wcU+9WKcVfZ4QpkcOdoX1os+i3aGcJSG1QM/P4xlP8a8t/JnXGlDxIGLbt7/oud8
AB61nD0DqWBqpBEKtgKnZkHqupK4qwfJPW1/uaGbu3+N+aW6E3fQMzuGz4km8RgX
2tDEfafqez0oUFgWPztiB54fFk1S3bHnVAzeSgSESaEdz0sSA78ZJEU7tuGzYuLk
N/YCNQF90oJoRZKcFkzMp7zvhNQxCuXvRHB0docbsUviixC6YYmvO0uzoUNeRMOS
gdT+h7OgC0jhwEjyK28AopGTmQu8wtIe/7VQGkk0dfKXReMIqUydOey9DnllKJDB
JS010ndZ0dTP396ITEzNTeL5H3zfFRVApHGYg3b2ufFLst+NtJ3JpRL4lVbuxzI4
0OKM0Wbdz4vFP/Q2777a7OGOF3V+cVDK7L8/ztz4+Jgzu6yghxWo8HQi9r97Zln/
ayL/syC51DRDDoCkHltZAfHY+a1PYfUFH6VgWZIV+oqKsmY5hoBp3JDVjNsi1MW8
KaeL8rdwXnw83PlUQJWtek6fhxKitaKNKik9QQF7vw/S9f5EG1ltecX6gAr8Lqvq
W+9VtWnoGNLC3x4P/dLU77INdq2yf1Es+QDwxrM0gq0Xl0IPwjXN3N59Aba8KMi8
1mz/qgERDeGBd6fjIDqiPe4P4KpOmd1eiKROmUpu9ZAPG16UH/hiKIJsFkuGZMin
EU5f4KrCQfV1/R2yqLs8nR9ZJGBcshpkxAaPO3EIDDKzrLHCNqt7hhfbKhyuFCoE
IvUUo0T2IX8uJcw9j2ch2tum+Dx4P/iZQ3GYNBQHyOOZiy9Dcg0xvxB7TgNIBgy7
dqSKUBtvsTnHcpYX5JFPI4QbgOc7j4HZgaNpcVZnS8NcLsIyQdHvBBehypfaEU92
0vYyQYZ7MzFe1fUgve3/1cQmjG4N3227WzgknNGD8xb5yEFJEBcUYd0H6S/wT0G5
irarDlmSU6Kj9gz2eQreIbgeY1iAOM5HnBLZZ8p7gzqwvl0yQQbc68aXZ4kwyFVe
jWG+MoEKHK48gqnzdwC7cICYvml0ZQtvEb+KWotlnB6Dm9PrDcZ5UUtaFl5MThHn
y/avtmHNPWN8oTPc9VvqlM02iR9E10d3z+fEQ1DYwAC41m7VAfRDcZSx3jMDkKnE
Yzawj0bjpXorO7+rxQu4zWJFlWRku2l6pr9iDjCv/r+Fxg9WrJ5pmQuMIf046UNL
rJkagBt/yMoBu+zcr01s43bNQTmAWUxZrvlqfv9mcaqrl9bwCOylWLUuiS0QefOh
7Nej1oL4AeChtW9p+F4p7o/Gewcm01D7F2Sc8e9BPGFG6KWulXFdORNXM3qywsjg
1lEB4GpgduH6a4yJpXkfSS67i+UgkNB/mpDOVRSk70vCTCNu0bIrN5KAtnU7bn2/
dAdO/tW1mu5/SafdsK3zECfkLKZyfm4UTREpjgL8qt/AGf1vJ/px5wCwsyun9cBi
u0Vm4LDOJSiAm8P/mnrPhfAjSfLP8sd+t38P6q3F8dO5xSPC1N9douV9hltjrEGs
b1yNKyLmWwZzYuo4tUIVS85q5s2iUk6Pm02CPQolJ6zbIH/VuoUmRBCYygRdpOg6
BvNNTlR+r6X16KA6lxO/2yXBdGShPs7HpjqXjiGQMAecDzbLV8n6VCuMEDDhzDk5
IPU0vHPBGjIz//Gusl4W2aDdqVday5NS7lz6ovBO6vVIfYT7GS9lLzK8O6FIaNG8
hcO691HJAufNw6F66N/XBPYCeA8t8HellD27cckX9GM5RS7YTyKRYrBOe1HnY0iq
oQ62tJQxmQ1zoico2KfJy6QvMuNCC5j3lIU0pz+WY2ZmnMMG/NemGm2aLFbZ+OF0
yCkgmHYT4406S6vM+hvGpDQV3vt9GqR8h4hfizfuLoerGUAzU+jmzaE6q+IzWqmO
0f8QLSjCg+0leN8ou1RFAXrkhF5zkOOK1RXdmSpYKCoDtXgUCLW13eDP1b8lvuZ+
1GLd5tTIVJq9qZMxIrtV01+qEwlAidJK3Q1TCNmRLYYHllapo2uBJNmGyVuiMVXY
24sN5WZrqOPUfNdxCC10DOgLYOp/+edo9YGusCOkT947f1w5Mz0PqjRsDEFeZYP/
EKiKMZsBUMbgN68+xdssQmCd2LIev6EvO2reRegJqhUqNe7EF42ABIoTeXtkXZ9U
EKs/2yxihkZieLaHQrnsB86PQ9OO64TUXtu9MQReP9t1HmO2v6H/94pdYlcfYCkM
r994LdXVZEfgP53FlVKwc/oMo120hDkHK4z0HG66qEcNWyUus/o1b5garUMiQZEt
dZA3vUuTCzul0yeH3Zuz3IN9YldG4tf4k55uMhx+y3R+etrhLY2amYgjIEt12vQj
OXyqLvICMHVmv7YdiQDCjEFNJnmPcuAb+TgNP2ZlwdiiknuQ21UbYzJvikX+/bLe
l/kGK5L0T4uJfDPZ/zqjeS1GYMxBI+l1yYv4VlewjN5Vg7wrYWh4o31n1LFenvKF
rzbA9UkmPQPKIwypq6Yl6jJRsngy4STAD4wyuL1A89HpFaGMu2g8JgQBfydx7OXu
iIBm6fQGqIDbJ2Ftl93IvlOqNJZxIToy+7XTqA8kMwUGyFAkjonByKE25h7xJPyz
ed5spRppB1FIj7m64MUzKe4dhGPsy+fJzQm4sBMuopSMe0tA8T/FXQuM6WjZ+NRc
obTjemxuFA0WqYqBIWLqCbfauHUQwBuZRhX6bZ6gQJYrwkgZ7dljLt/aq4DQNaAb
JnurhHsFH+C4pjUXy2hZ3seAweTyJ3nOQguiLELhnPtvHaWZDtLw8PjxcW1KlSFN
LnVC/4ILfVG6D2Gw03NiWGuFKbNdZ+yLeYIz1YYqRAVeYPPRUER+zj3WGuhWdVWq
K4Mv8rWjXv/Whd/p0Jt01RUcsaF9uwRZpQijlUKf1IO1A8kcJOPK1LtATS6lbThV
KyWxVH1V95CKkZMHhCg2R5/XPcaHTBM8AmM+QlrTer868oalGTbFMWFN8mIXjGHs
0s4OwileajRZ68wNPLnnJtIiuqdiO5PeH5vRKOG4HT6Y7QuuSCBTYZrI+Djk7Wo9
D8IFDoJNCsRdXQNwlAM/wPuLJRA7Rn6KMZ5LzJ3Xk8rcDjkWstqi4zfb2KCFW07O
9mjjR2DlzWM8Bo5l3+CjfqfL5p+mHmlv3Ra9h/Fi26+yFPzziIZLAAk0xdbZUZL/
/l1z69gzP+3BNLAzDnM0EJPhBYOEA+TSdrKs+7CkhsIbC8IiB7Ki3TK1B03Rbqcv
PGNGHDlneWlqeVS/ziJ4Qjs5sr9+loMkEgKpY43OG7GOHoREBQrUhJDLpH+i9cF1
AvQ6u9iFZ756CPzqhuSrGNpFjPUkRgTQhbfijCwDXthLwo8Kgonr9HITsIB9TxrA
gth8RUzfGt+4JNNBIBUOQz+oKi0W+BR311n1OKu5Q3S8K/j6h9WCiMCpqH26nxHQ
+FT6xJq62+X61RpIeI4L5GtbapFcuKADKSU+O/9fIYVQyFgiQEjFMer2f1ZzitF+
KZk5ry9Zw0EeuIdbJtfe7EWRRzzg5enxELOhtIEnjPCq+xB3GEB0TR/X/WO5DSqt
W8Yq822RxsYtaaXfHHF6yTgW92yRHfievcTujFeUhx+Z0FD3f0j8VKWWpeQxIxeL
q1rWO8Lxcf6MsR/Qj941AGczvyJl6/Ndw+PeC8tWP061S4VeFwG648epLQlc2zNK
AKy2TyFgOiJKv0P4qjlRcd6+ir30emV/pNOY7SLD8LSVG4wlUmHJg7rsgUbLp7rf
+gNC0PLtHC1CA/v1PgxLRzj72MVYRHEgewEMcUsswzkIV14+Dsv/8Ajzd36i5jBB
7V7bkx4dNVsi0ZPltNgbAgEj8g9/TjokSHsDhxH5yjuVNjhg3kO/hs2eZbWcZJr8
KPAtBwP/1p5IRIzFbWIIkrMsCoFQUTykTvHLX5njqKEEHjZfFxf3YYUr2DY0OcmK
lCmTbEpEW+uI299ZNdag+oibHjeHktSCZie57llYMXGOC889rYdmSm0bkLXXCbt8
dIEHBPamSTZBepeo0xiBrjofjfUMEKNCRF5ZRDXjLcNvfLl9Is7wdgvXkKbup6CE
eJhPolvl2y9Bv+oiTavy2bc5aWLi+AZlLcYA8aaRXYbDSNhw77swv9CQrboerq31
YiFlvGlppUlbvpcrAPUF2LmyvtUbAbLBHOFCU2pa9pppJX/p6SUbI9zdP0jgI2Rd
vstqXzJuEFPFnCkjoc/d5uss503w7v8KvKtIfjJAaJBvg3trv0YZo1VGYL0GBaCz
9GwyCFU055dwsca/QU+yelWoTUSGbkZ5d6miv6Q9/mLhoOR5iJ5VdHQYPudVE1v/
jfqvfSW+sta3Iyiub3OI8eXs4AQAEgkdMP9KTquCn6QAjzL4v00oa3EqiLizZ5f9
fbIqXxT8KGbxDEosm1Bf6hG06jbGaVSxbkPCvrMpnTYa9D/S0gt/KjmiPN0tcjLE
YBYH3t5wNswYJgMeOjCX6USPvmwFGiFmzpKZph3L9hteimn1vdXjKrlmhgNWtuu7
w6KfCA0xGcqtclfiZTXjqLEn663KaTktzsNRKjoPLdGdMNHotJXWpMwGq8M++n4b
QeiFdDpznUoP4Tv5c0bWshaxFhzoVcvQ+9/ZQdOlvSunI41328PqkwwzWocaMmf0
cjZ34BepDlYFtGhzStJ+XTs009FpNp5tqyzEKpVHNghjrDak4C26XPMNIcR38TDL
5TqOyWWHleGpcV6vloXo37LqqqlzeO+/NeF/3VwruWbX0b7lvcUCDgHbX5onpbH5
Ub/ZwHOAdeCSMSTJsHFtkN4Tm++flF0hSExF0hweDbdhiE4oZdLsm9Vyna/62m+N
/UV+1BIyn+g4uis6Aern/GwAkFwaFbsIZVryNBfF+ScE7F7IkRN/0rrHKCvfDooZ
bwaqaOuUE8V3JiTUK67Q+dbLUhL4m1xLm92KbXv1cPGk7wpstbAz/fMP/JXamHUu
eD81ZFvNVwj8zkU8cG6D33mrycivhy8osrJUhi57J8WjmEgqhQwcwu0WiX0PuW5F
CgptU7SG85zTFQ7eJzq+3TWS0l7UjLP58hGkTRc/2y4IcInZq1NeJAKUcob/Y1C8
Vxrtle6B6/9wZwZWfOKzWFlLz5k4EQjKj1NTaIbh63/Hy/q4zRTMUvpjPHCiGucV
bzv5M85WwlynnuVbkBtL0MNBWGsbUJg4XkLa1Ju3zylRj4N7SSg2PAuGVs5cKemy
I93LB4Eq5sNiIPf1RQ6bloqRoZkMV+0ATE8nFl2fVx/Xrwpg1BSq4ZQyKQ7u/ANp
YnD1Xg41+WWnr93PlqHsvv/mGcHt4vLHdciLnqDAtgaSqBBWfIvewScf4BWFBU+w
wCDz922R4pgvdXSJ6B4A6oaxugE11gsVp6ZtzotyGWHfZ5TnPrAsPc8r7YAkCnWs
8GPjwyCYidFNEGaWCCj4YJ8HgVvUqmMzL4efZS9GWGGA7uEuB5BB5XKtU0nskwGa
TkBOmDLVrTx/0SQU0Y+L4kCgoEXxex9WvXftgSL9flWOBZc6Nsb6ZPmM/BOm2o0i
QnOpbpt8JKSLTMBhdQhPtBLA1j0dBBp2ibLy7RrWWNcuVdLjgjI5HztrZpV6e+v1
cKid9FCklxDNQDGiM917TV0wTU7yRF8/NflUYZikZ0LA5s2oHPGc8NpIXs2KfQB6
8W2f5rAIKdLINZpxqL8hr95VUOAZVwb8qJGhBGJAk8UYwoQ6xm3QadMrub8iYh3T
j9BvPTtB56hSLk5+pPTwN7LRoFQQHMBCSVqKM1pSSM1mro/Hw7nuDyYzaFagaA4W
OivrSb2PsA7wtIJ1QQfV9qHcTiGqO2Y/bJCuNEJJjt6wglgnhWrtmapCSXGDonL/
pxCup/d7XCxo8eHmnu8S9/o7BAtTaZmbO60xnXvjUG4RTIm1BkptzPbO9BvqwEkY
frTLwtONXaTDU88ev9HzucObiqTCsN+jNyTUGVwhMTqxAqYstRe5EItA69kHJTV2
iUtjsxlpX8gS4eCbokH7wOSyZqAEDIZNmNYzUj9m4jITmOsihw0Bh935ssH4r8jJ
D8ICtXtoZaOu3drZid0BROV9Chx5qTHGLVhVfK33ucuB9D8nhKbX5Gjhnj4hTqH7
QbxsUJuhe9HRAdqGYtceKi3SmZw9xBzTMkxPO7bkTaTnZYoU38AcEScGFge1PFxt
M4lotnvKQCU2HmMOPVhKDvBAJDbe5wkyWyC0ZbbKGombaDbmliWIqh5gE+XmGYRh
Diz5iq81/kd9vQDegvLy06XF0/rdqUnFXlFJEUYjOH1VaEkET4bTFUO8dmYx0byP
v1vVHAgpu7rn9YPliXFHDn+dxITVBUkAGsjPKOsO39xw85qVpKy6lP1sWumjukyk
oVYHOoBDJ/hN+p6KC8gdg3a4wgf5jnDewGYppb6M+k37lraEqiH8N6Gb7TP+qO4E
+spnVVSFKwCdpA6vVKS4iHr2cTmNHms948ArGkQbrh7vkpe8bTQzJ1aXRHMg8qO0
0I9h5DO8QQC0e7c8XBIN5sNoOzk7avwqqvidgr8xMvDaoK7ipmpKErE5RTXMFq+7
ziR446VIWC3U5dkWJLRr+LAQEU1M1G2eSdtj5K7Mf8iYky7TAd0oLnYcWNmF+JX9
SLaJpDhQCzbG6Uk06pI8zn+n8vztfP1wBHLyPULePX2fwi6NODdmBq7e6I0qlbsS
tupe7hVbUUL8zEaOxf6P6Y7WKxp4qgkZNgRaGDTbiqvI+1UVEqaFDC7KcbABXPJp
qM6vxYIF3vxFSF1YCm29TPtkqQA22oCIUlwGEGmNzEnPzEmq/eShzXDr8qGeZ2Q1
Bdqfmb0A1m3MRUVr0AL1I5oP7ox23FiiUKdTyG/fs3BXUngmOseABf2N220MmVvE
r1vIvXNw3kG7DKGF7rWbqVRL3Nu5Z6l4NU2Da8JQxLJA3HGekxI3VwxoaH1yXnO0
RCTuznhaq2Vt8wwsSdiDJ6eQVpwZfHblgLCVYosgtUTZ9cImlk/S++PhSOiLYfDh
CLbw8zK4+svXNGu2go81u9kSqvHdYTdf6l19tnuFF/uyKC91sGqmPIv+dV/DuMyI
xbI/pDBphwvLwP8TYEEO95nSGRo6BW3LjEaCdy5YOTeim6mR+m//KJbWsagrGIkd
XdptPMJ2QPcE6e/lJ2PJjAP4Dyto1qvwhmYZl3vgZdCY5odkHLNxCH61QoY5h1TG
vj98exY/BrX2Dz1+asQsef7Qiy3l0ohG86NAkLauXagdJSpqRv6XZZxaEOh475oT
UBNt1nPnr/ofVBBO0tMO/31qpPTAq9hxypgWG4V7+u0=
`pragma protect end_protected
