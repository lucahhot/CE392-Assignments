��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�:����R���9��Hu�0�/N�^L�$a�Z�p�P���'��x�ώ�~���o)�ۏFp����E��]gwį��j���T4)z�!G�L��/R�@�9[
��)�� �~	��U��e�]�����ug��Y'5�O��u�e��V�&�h�f=��$��z���@]�{�������)����RN���0}��ik��.hx�m� ��b"��>�����
�#u�s.wd�g��kf�pyo�9S*"&�X��
�=��k�&�ZqȧB�T�̩�춞 ���{?��!�$S��ߦ-���F���+Qֺi�\�v}tV����jnL{�s���7P���
DJ����-����&O
�i"}�/�/§���-Z3N/:�)B�1��0)E�P�O8�3�Rpwu��Tm } �E9t���q"y�'�rO��?�4����)T� ���i{ �I�������r$�;W�C�l	SY��;�����ʉνq]Qt�&�@A�Žvd�q�¦��j/��5ł��@ʷ�3#�3�c� �'�X-N4�ɝ���w�X{���"�G��<,����{L��h��Yx4^�[�R���G�AiX�gy�ź�������Rh�6���A
�__���
ǅ� *h�[�Ï�O��Pd�!�������,J0
������S� ��[�2��+��$�!�W0�r^�LZ#Af(���;-��:�& ;l�����)ڻ���ئ���ؔn�u�%NP�k?z�%�[] 8����G�D.v:�a(��L(b�@��,շ)�Q�0˶ �^rNbL�c7�[M�t��/韭��A�O�E�ւ����Bo���4m�e-���7b�:g�t3:i����?��4�R
����3\�`�tn�:�L�ɾ�c�$�m�S�t�B�e�i�k�i�Ci�%�. ���Y�C?�T�º�y�uo�Mׄ��~��q��B|�z¡���	�U/x����ff!��$��"n��鱗��m=������2o����D@Eqf ����T�]��&$,������m���m,?�5�'���E"�n�3F��� T(���jIS{v��S�f��y�ex�T*x�ڰ�Ă�|�vZ�W���!��,0R�Gr.��)z��0��E��e��I�˚N+cIhk9@!4�g�U����;�i�]=�Lm�]UH|��y�"�M��.�XktK���]�0��t��y]R�J_q�ߥ\��̧��k�a���ҁ�蝮��5hi�j�V�m0A�2��؉�� T���Z�@3�(&�������C���Pp�VT�; s�	u�^ֱ}*�_�N��\I6����;�W{�߼ط7��N�JS�<�����a��t����~�!���+8Mj#�Ξ��LmISh��<Թ��B���x���I��ػ�k��QƱ��ӡ�.�2�bvaXU�
�~Gl��Í�u�J;�˓��%�\��A1�U���[����
<>g�Qv�(�j|��9^�V��5�O���<��xg8]2)[���H�D�^�<ا��k0�{��&te��I0vVB: �oM�Rt��:��2>z/(����ƞ�`ͥeǉ���$f�w�+9SO)�(�ޏfcy�,�h�_y�M'�=29͚좞��8f *\"'/���:��������)}ܟA��ɖ���U��0�sa_�q��#>�|>���C��αTdr[��?>�|��tKE�̜7�>��s��g}7��F �_�F���'�)��`�.�q3�E���oH	�z 6�t
K%oG�H(y|ٞ��L��Thދ:_ph���_hZlZ-,.&�����89R������Y�8����M�A�,Fm�-�M8"����%H7����MS�cq�q��d6
��L@�#me�}/���Nw��+�DR��$)W���!���)�i
s�\��E�E4��	�rSѼE���\(<��Ȧ/*d��|�s9[�\���n.��i�>*0���~k�/6���򛸏E7����I�
p��Ui�[	�c�&|��1�	>:���b�;N�nۙ3������hc�-��M u�}[���c��@u�K�a��`f���D���3T�	��c9�:��YWd'�r�n	ǥ��!$E��)Ҹ����q�<�8��p����X���_~?�[?H6P��<9}��!@�O�S�
�,�T*i.`�H�O���*:z3^���!�O�p,����N ��}.Hę�Vy[�nvNh5���Peg���WltH�.?�f�X�ն���,�����O\/ �
\J00?�^�3�΃�H[(�}�\D�3������r�a�S������o��͵�/�|k�Ȅ�u��Ŏ�.-�$��6�:�d�=N`���aF��J����IN�L`s�$�����vsլf=�I5KK��>2M����5))xk��jvx[�nO�R�����W��l�G������C������3}S��9v(���$Bw��\!����X]�FN�y���b���냠�s�涗���A�Gf՚�?l��L1��h$��b��=ʘ����~�PH[�)Z}��|_�Qn��;��flʎ����:�9��(l�@���S�$�a�
w{ϱ�+H�|�ӌV�H�jg?��t�9!����y%��WHԜ
��k��=���K�8/�j�[vw�/[]_��p�`GrQĮ+��?�8�E'�������K\��N�+.^����}���|6��~�M۹��Ff������<D�yP����v��=��7����%&��5J���)���
KxJ�vQVXAK��*GLWkxI�`���o�p!q=*�Q��z�B��U�d5�C.�ruG��M��(4=0g���V�`F����O����)K���N|,�⡃�?wdck^����&��H��~àbW���5�Iz@P�����6��ѭ5�Zr�dŁ���n�\��F"�S� =�ؾ�Eb�EU��C��� ���&rC._8��klvy��E��0��_m���F�� ��ް�����_R༮�������5��rP;��x��5������y�B7��M���.T�F��跜Y��G��AA�eD�����獘�4F ����M�4�e�\��ui��+��t޳��5�/���8
^;I�F2����|�@T�`��I��M���F�z�"r>�������9���8��a��r��pr�A�����6���A����J����U`�lEH��'U(�oHA��>&��i�.=n�>�:}�g�(�nS�j�j{�ج�U��W[�B<N�pw�������0��T�dO�MV�)�rl6�O~�{J�xU�m0�#rҝ�p<%j� 0@݌��������9?E1��dm���C�<�EjULz�g��S�}�_���/ 8�[.�觾
a�m]dY.��U;W0~����:����ш�,4�@HIH�Z��U��d��c��H���?{�h_��A�(�ݺ��L�j�����®N��ȳ�U�D)�F�q���be�@������h6��>T��F�?�X,ib;��?`���LVC����x�J�u��&�Q<G�锜���Z��8�/ɜ�U��OIv�:~��ș2��TU���Ò��}��}��r��Jc������51�Р�2x�J�a ]�S�ecW�@d�U��%I���*������E���>w�ǣ��#�71�f>t�͛E���=)��=��f02Ɩ#�N�%��j��ˤn�1�$��P~;�-�n�)3��_r]�G5ZW���]�+y>`�~�ZՆ�5��'��/A������6#��Ax��qI���@-���K���G���
L����J�F�mQ���4���v����crT�4�3Z[���g�r�J2 ��ԅ�I�[��&9׉�
����S%ǁ`]�"�(oFܡ��K�gw
����W�=��e���g]§$�'���^��Do#�!�^1xi��1�N���%iGt����N+�с�<L����D�Hmq�?�L
�5`xS�gM�ad�o<]���F����F�
C/��͕L�xh����<q$y����1>TG���L��9s!�_t���.9����i*�@��NA� ���*�� F�M,�**�����G��m;Y��<����^H~�
�����KS�./E��.�?�G�~�9%��p��f�P#�j@ǒ�D��^�^��x�zN�ݮ�V����%G���
S��VO��R9]C��P5l����t`��m[�IP�v<>�ii�&M�d��.޶��>�V�۬*�s�oz3R��o뜩�ҍԁ8v��V��*�g��êZ���9tENB��h3D�A�T�xX]j0���)�F�e��-!�3�Pd'j`>�~�De�����lq@?c�9��gO����n�������X���?��!�)O�)Y��6b��s�1Μ��΁��
,�ѵZ��u ���&���W7���rƎx�ƥ�_$+%�h��t��c{�{G��r׻�E��+lu'�D�i��W�t�ç���5��?'��pГq�'��\�y���#샞���W�y� x���~��ͩ�l�>�D�+����XRħ��YD��& �`��ȗ�w����ro"cTGd��W�}�Q��d��5W�Lr�72\\�6���V�Է�W�ȡ��^c!��3���̧͟� �.�r�Ei�%���J��
���\�Kt�R\�7nC��C��^����K�y[��v���I�Z�{W�b���]t`ے��d�e�πf	��#�~r,����} �B;6��L�ᬳn`��r�;��:i3������3��k�وz�}���E�������t��+:��տ�?�4�t�ݛ,�c��VW���p����H����
\g�lrxV�̌wkz�v�lrQ��ri�L7�ʮ�M�^	��~!F�$5�!���v-g�,��"p��J��cK�ɛ�#���ҰH0�j�� %�[b�.��N���5�C���d�KS��e���8�u�>��*lO��%}kҺ*/�	�r�B�+�z�/�lVJj�V��2Fq�.~S_������8w|kHA������kiR���u(�~�,g��ō1}�`����x:����@j[>q_:���l��C��X��"�O�Z�Pg����\E����6|Mؐ�ī!Ip�a~!�%e|�M�U[�>P��w��u-��ֈ��/��Q��`�X��j�\9��Z�2���@���m�S ��z��ȇ6���ѡ��ѯ�'�+S�a�k=�Y��B���ӿJ_Q�K�n�Ҹ�n%��`V��9
�`|��j@�G��'�[�	c@��ۓ�dNB)N'n!l�G��Ѡ��$v7���O�_
��{�Z	=��JR4e6�ͧ Q�V�SZRa�L!�`�KnW~�A�c[i�4���-��̧A�Bj�#�?YxJba���&���3Z��B���dj9�'-(���>�/j[�&�;�y�E<~l��a������~+t������ex�.�� ���X!�Qi�
r������@ti_`x�<�n.��Hر�}�����	a�*��DƲ"���}�we� �垑�w�gM��o���Ț={���ݲ섭�$�/Ҕ"x��U%[���^��{��=�z���/��o"���6Km& ua	w�uQ ��=����A@�����v��;sѼ�`r�~3)ĬɅ:�s�ݩ�����Ngks=��ն��9e=d��F�����\�p��������螿N��5T[6��"�b)� �JY�AM��������z�|��37\N�{Ág��4��fq&%?%;b&��J�陣!h�F�����\���nW��l���5^B��9W��N��l�ځ����޷��I:�.��M���Ns1$�2u#@���d�1�-�6��¯��� \q/1*����'�w�H���s5:҃�N��]��E-��+,D����
m�Qg��È�sQ1�W	��3c;��V�0��&ٽF�����a@s��O6�f8S��F)U�����j���Fq�X\�L���R����YD��8���K��I�~�@�;��hs����P� M�l~C-Ή&7#�.��zO��٪������*07��},["0��Bso�1>��GLd�I�R����aѸ��_X�m�7��Рi�t��a&��v|�$���$�w���*�QKב����WOk�/؛��TC:S�$��C#c]��Y�,Oܠzf�������E�"f0�Y�� �Ż~ ��XE^�-%K�@��eם�IDZ� �՜�9��} ��RUZזړT�m4���~��RYAү5�D���'=���⸹!j�W�)�¥k�f�4R��9�Ļ�w�:|�V.(��#(:�a�]�iu�5��#5�oĪ�D����sq�t	���1��i��Һ�?�a�_�	�T8H�nW�G8��>��4$��!��Zb��\����H����|�K�>{���ʾ����_xKs]L���~��1&&O r��U8H t����Z��7�3cb
x�%��+�f�jnqqo g	վ���`�u�E����HR�=�4P)?��Ǯt�P^
h�e773��]�oT]����|�϶0<���6�WAe֋�p�'�V������b% [h��qÆ��餾\(|m��i
B�~u�$�1\�%t�Q�|�z���K���4)�Z���	(X������L���v��{�6[��32'~�m1r������(h�����տ]%a2%CD�)˹��VDO)���Q�g��ȉ��h��� �� 
đPjz{�r��-��G(Y�N��S^|�}«���P�ul�]���OCk^&,�_��,>x��	�B��nP(��m�z�R�������S/����4D݅/�o#^,sn/��u[�@��"��1Qod��8D�Ǭ�0i���O��V�ȋ��֊K*+`5z�)��z��=�È�W.ce\)��v��U����!Pr�b�k�Yw�-��R.JY��g��������+�w�����,����\a�Y�5Z��E��P��Ra��<�R�V�$C$D��?��}���F�#��Ց;{�X���9�T!=��D��籊E��o�V�_7�_J�#�y(��p2�@�S{P[�`݇�� z%7�K���~�4X� בx9:m3�h�Pw(��~�`kq@�al;.�&��-<��R�'�rz�3S|:Gd�bò�(���N���dC.# ���Я�L����fE�N�z���~{c���/≯�}��v5.G��1Ɵ��-s0[����(���ʬ`o�����V�c�	+c���o��o؅�H��[�	T��%6s Ҍ6���fEǑ�)�E˿=�T������J0f-��q���&2�ϊh���9%$p�[y/��>�5Sg;�^��	�����~R�m�-i
M���Y��c����[Ҧ6��{�ʭ�;��w�r���F�u���v>����%�h�J�6���"ha���	��n�"�v�d>qV%;����V�F��|@�q��1���A���ſ*9rT�#Z-��%�k���L?�*�/����K��H���i�ҽEv�T�8�MqC�T1G�ed��&���Qy�p�E湨D�[$Fk�C�a�lMCZ�7VT��~�|�Q;z�4��@ԣ���C�	�i��lG{C>d+_5�\ `�Ʌo|�9�Q��ˈ�v�p�z�N��ڝ;\���5ŀ'�^�5��*��>�>b%r��R�ei�a��3ȡ@�5G�-FV�
�)dα]7���"���J�BS����Q��T��JM��4�O�f\�4AhF+��m��EI�AE
��h�o��3~�?8��'.e���֟���J�w�|C�*���Z ΂'�������cȿ�����e1�����E���v��tю�^0�m+�f(�գ��� �cK�������[Ӥ� %  � D��m���Zh�D��fC�W&q�p��p��:�qӋ'9��b0�I��ڥ��4�ΜX��B��-7n��=/�m�< ���e� V����'M�����@�G�����)�!Ӷ޽�Ў8�Z�H� #�|)n�ԫ���UI��N��n�	�Ơ�0܏\%{Mxx���%IE�(y�}ә6vD�Mx����Ơ�"�Ϛ�4P���<�9E}�͜��I�7;��������Ƃ���o�'P͗��ڮ���S!o�����E;k̼t�������Ϊo`!��~q;;�J�'����DM��S.t�ȷS]dKb�֨S#zIS6)X5�d�p�b��c���H�n�KA\/3�,>2v�]a��}�|����"j�����%/a����f��U��=>�|<S�E��y��c��+~�J�"g3S��'���%~�e�W��,G�)����Iz%g'O�MbBC��%�Wa���ȫ�
|єT�ky���\�1#C1Wf�� -�kV,r�\��i�b�c��������'���w�C���ϧ���V �K���.9�w� *߁ >�+C%;�xM?Ii8V�ħ��F[���h��y�zI� OBQ�N����+�G����
:Z���}B�嶢3T-Zw
Q3�����t.j����T�:��OأE�M�nc<.s�F����>�@n��:rY�#{�G��;H��5�Jr�2k��z@���r1����i�
����� %�>)��0'�iS�~?���c.��q��W�{_���0�
��fE/ nb�%��,1P���5D��5�;Am�=pdli���btCa��>i:0Pݯ��#h��x��D�S�Ջ�\�a-e�K���T	J��L��;T�>|���Z���i v:�w�#�X��s�e���O�峗mD������d���b>�?��&��G&BNŸ�|�3��)&����m�朗�m��c��VQ���pD��o%�Z�V+;)P�"��� �p����g�4U�/ �Y��E)�R�24Hw��9X�#����_����},]�[n;��u�T#�$���(h<y�5��ƶ7���9���9����$Q��ܧ����"q��ج�XcL>?�L�m@y=�"[At=�c2x��(ӫ�o*������R�祓�>���l�&L��|���Ԟ}�!*L�2<�m)�N�W���u�?AHp���*[3�72��
񩦯/�!����B�F�A_��=	�l�-���_1@������3S�y�����@���V�d-�K���(΋.���-]�b>��7�j��Hki���A�ɭ�TK�]K��#�YB��"-�\��O��e�d�W���x�0�u$�����o�{����yW�n��ĝA��D[�������i��G%����0_�Rl>J�k�4������~�"�N�9w;�u���HU���Gp_>7�_�Z�*8'�)Lt��K9�os���d��sh�..�T�ު`�a���L����K;Eaڭ���@^��6� s*�T8�v�����tHV�\�{$=�������ˌ��Boe_*~}p��X��$]g���.f��d	��|M�5D����Q�(b��V"��1h���'���~K���i G/�����@��A��":u}q�p��D�<A��|�[/�S	Sl#��}�vʹV+�������?jS0�{�;�
�K���
D�M��y��xt�(x�C���_�w��_�nJ���c[�]��M ���;P���l�3Թ9s�c�R��{C����#��"b�Ekx�W��g=��fL��~�/Fq����4�K��;U���c�C�W�Q���"���.����B�S����5$޲������ӉG��;����o�Ά�]�>�%8�gpHw�4��`d��7XT2���\������'��-$��&���ՔT�4�� j�\�k�)y�����?�$x��7*h䠊dTQ�;=?� 9b�}����Y-x�����
�S|�W6��Tz�x�̮Ho��xK)5�k���b����9���!4Q��I���q^�N�FE�w�(���Bת�ڕ�D8����X�˓{�m:���%���<�����L� �K�G���J:�����ʳ;h��}GA��o(�Y|r�p;P���uP
�6���� ��ɷGK;�Ȏ��7��n�����$s
Щ{7<�[b��c����)"�$����v���Bw�G9����	Z���P,t�>��dƇ��BY,ctSC���y6[�m�T)@F���L��1�&
��ǩ�U����0�<W����u��I?�J�"��yΏ�2�a�~m�䂴��zX8�ܦF���D\cj��w$chHȒ��G8���x��_r����5׭ڂ�f1�ߞ��^��a���I轟d���K��L/�=z^�DJ�K^ܞmΛM�~�?'�v��鮖\Ϝ��䅇}���{�b�]�oH�2�Ҥ,W�h�v����-�&2ꑞXL8�qȆ�#���N1��̐lp9dT�@B�
�D��-[�R���N�&��,f�-D�vO������j�S~X�o4�1�pR�ޮ�����K\av_�iU�׭|~���zVtn�Pjk�Z\�,����I�\>�t.iK���y���*��}�B���*���������,�U�炙�|N��$�m����R���fi� ����3'տ��qu��Q!!���,۹2� �)�ܤ+>�� 8�!o��L6��4��Š�����M~��Ǆ���-���-p��v��9���J���8��w��1 ����M��f��ݮ���_tg��e���]�0�#�hGj�K�@S�⁢�&/Td����C�ES����w(��F��Ԅ�8�{��%- P�[��7����lL��Z�o���Le�Bh,P��֜]d����gu"�2Nq�_s&E�?}�w3�\S�b���B���|`��֬�p�(F���D���_�=zx:�4(26�s�� ~���A�=D2���� ����"B]���T����>���#�Z�v}���/���ګэ ���G�1�R���g���I-�\�:Q��/�@�ᘆ��;jG��w�E�F;�{eu��'�CZ���P����m��,�$��}���G1'��	�v���ƭ����7?��g4�u>�|޳�K�������τ���V�A�6�h�P{l���:�d�2;&&�ce7�aBD-�;��Z��$��O,!W)���V�I-��8N�~�5�lh�w�eF�k�S�Ty6+yl�t�Vz6sB�oQ�2T]$jAfD�F]�w�øk���qs9},m�;�U����Հb�EЪ�d��U猭�in�g���@��%v������Յ����>�	<�,dT�Qˋ:�>O�y��_C���IRq#�������A �<�G���g������%օ�ڸ��Q�n�&Y]�1X��XuKM���}�q�$��h1mP$����~C\�Ve�e0y%)�+�1KQخ�L�?Knz�M^K?���gFr*o�>���E�>Z����Yi������YD�5�;���ݯ�R��R�y!?
���m�V>@>OG|MWpf���|p��48��������bx6ew%����>�+�h}R'o��-n�|{�8>/vrA��{1�h�iK�C#w�V�a\41HcP���`.f�uc�6D���9ojv {���!�騖`���Q�ޣq��nޘ8/���~��U����eq2��C���REw�2�F��Jd���Ko{#��u���K��HHȵA;�3������ia��o��!9�z��ꦚ�T��'��,����H`hrpr�,�[yn$���2�f�E�m��-�O~�L4�o����\�o���@��;����������m<�}#�GnewEm��9w) ?V��K���m�Luq�T����;4~j�n��9�[t��+턅���XO�ę��K������0O���N�{�O	&��L�R9q�nCP��[ ���ܫ�/�o�Q"��͚��>��XL��g��&Ş��@�h��H%.)��j�,�I˴��˹x��(8�F(�}�i<O=p�P<�;����'��3ί��G5J���G��z'���<O���guq7�{ �8��(�CD�2U�\�!�7֯���:XnF��3�.)Lj��
��:�6��
8��~�%%���G�⼚�����+��4�<~��n�ӿ
	|��7�p\+vMjʽ��z~��rv+�sT�3ۙi� ��S�����LU����^m���|/�?.�'��h����i�1l��x�H�-�Wg��)J F��c�xP�h��������b��ʭ�1`�u�RY�k
ƅ����T������R ��^d�|�~���� � }S��
�@>B��6��C�:�f2��r���W	R��DkzG�f�y���ĬK�:H�&���{:�y���3�i�Iw�����.�8N�S�-7Aa�q��	m!Y�sLI��9k�u��ف;*�D�������#fʚ��4��@�}�r�9T���u���ϯC1�Ђz�����A�F�`ު���ٺ_��D�m��vh^8cC��2[�!@�t�.��ڝ��J��=R�}�Mc��-m6N�����$i{mm��<��v���k7s#�֟L�fJ����J|�փ]��]**�/5o��g�v�hK_�%Ғ�E˫�9,�S�]�*�2�\v�OB`�(=��]�vo�˹�>݁�㢘�8�5��*F(�~SY���^��BM�L�P�O��ƍ ~s�E�'C�+�n�kw8�	�q~�X��?�%J����\�����c?+C�Ӂ����(�y�OE�p����ꆠ��}K��Й:���Y�`���������b�N3��g��JŶ hP?�p�M��(@�O�>�
Mey>w���/91��3��kGz��I[���|��BG�cf�"R(�M�m�ٲ��m`�	S�	|B�dl��}a�u��rM��*t]��Vh�����-��U���V�v�?�X�n��*��pm�t�I��F�c�N��w�,�e�<��k9�5��SLo��� /�z�6��;��y��j�k{���'��$6����1���� �*N�<~�,+&�yv�4����'W�d_�����枠�Q�����K�f^�]Goږ8���v��Z�x8���)����u�c���kO-�hHQ.�蚼It��0FWbso����R.�ܬ�Nm��O_�ā'�Hi�ݳs�����h�D���^��J5\����r=�ý�~��9&�3 ���A��1�����d��`��X�<�b��EP�S��[G0��ʥrαm��Z�F@�������}���z�yٵ\��cD`:W��O��j��w?�V�M����69f���P����U�v�㌇��H���1�%��R�ɹ���ǃ�_ZHp�W���U���n��
�m_'�A���,߈*X�+�k�%�>'y-E�Rt��FҦGI5��b�Ɛ�I�ð;��m��ޚ�F����W}�RE�3�@���0��~�W�Y������B8��H0|�%�]��x��N�JH��g�m�����F��H�g -��.�����a���DZ�n�,��<y��u�}etpT��#�H���1�����4��p�G^!�9H���
�\��rz�/�;ͩ�����ڏw�����n,���������֨T�6�	`�t�m�W�A8P0�m�(R�R�d_����<�ĚKGun��;�9m�H�����#�Q�`Y�Q�4X$F��%��75�JS58#����ɴA;��C���^�ʄy��C�n�wjuK!V�	 �N�(*�|�i�oz#!Fإ޼=GF<Y�-f��Q�af�Z��� ��՜4\]K�m#�]Dt����><��O�cA8��Df�#�im4����X#8��K~oi�RE��{^��kUO�C톺�ޘ`�$K�;��}>�I49�I�{���:d���"x�m��|�+��k����	�~ʞ ΞW"aܑs�=Պ�J'Y/�''w'��]�/���NSv^'�{�P�H�\�Ն��B���3�h,@K��p�D�b����ƻ��< �OnnBE_����>"�=k�y�u�?~�=]��� �4�0��2�:�	�O'��m��LHjrmO�}��)���d��>w8�8���hC�Z��J%K&��J�B�f��-�[�ч��/��f��d���j�+XĨ��E��0�Aq�7��"Z^s�k���6͍�� �z�5F�'6r'鰰}����a�3>�	�de��l�D�<�tAY���\v]�	��i����~i`�ʝ�0 ����'D��(Fmwt�9�1{-����\��)�6�y����88���~���a1�5��H�%�ڻ.$�|��9�P]���a�gc��l��O�� ��GK쇴/�������P|�c�#�Q�%��*�Low����$���ۤń��0_�+}]R1G�v�ibm��y�w|�}V��B��"ʑ�)�eґ��cӈ;����(wIPt�r!���J�ڥ7�����;�pl^D���PYV�����g4��k��>�|�Fq@�� Ѣ�-b����ݺf�Pl1q�NxB�_�ѵ%'xa#!�3ȟ�g��Ֆ���
D �cJ>tA1zH#�Ⱥs�!cF�AQ��H�VY�z-t���h��=�Ơx9rc@��̨�3��ONCF,�1����= [9���ђP�E�_������i��qL�	�,2
yly-�\=�ֈ:� J%3��1��/��0C6K�l>�F_��Iٝ:�bbw�"B@;FXs�� x�Sfas�oo/Sh��h�W��L�^PZ�e���!fF{�m��?A}!ȉ+�*��[sz��r7r�N�̔���[�4~w�MVj�C�2t7�w�O
x����u��N@��o��u4�R�'� ��<e��n�!���V���]zJ���Ms����M��d�c]��]z�'9�d~'���w�ʠ��Pyĥ�8������Bz�!�y#7�S?hF�S}Z��V�qn��cw>��q��u���q,:��>�Y^�K�d4�5N��,��2��aa.8Z��}���a����x:Z�i����	�Br+�nv�T]M�2�4���mp����َз�t_���(�K
�Ud��lP����*1yٳ5��2�cE���NJ�ki��kd�.���K���`MY)��v�(TA��Z�[�$(�5Q�w�m0��o���2S9�/q����a�&>Ei��8Y�*('� ��!��n���-3��İ\!E-�Η�C��Z�dҲ��ڊ�0�WPI�x����������O����e�X6=�o�y<�#�/=��3�$�Lkʈ�ύ�(���?!����z4��IQbvZ�G���)�������0�r���jt�Y�'�}��e�JvD���`/<*& ��1�˂A�槌�R�a)sL�VZ!�n�O�V($���@�̃p6�eʎ�0ܶqEOl���r�I�z�x޶��G���1�|^�^y ~ݹ#Iv_����Isrk�BL���V���tņ�Ay���}�; G#fy�����"0rf��kX%<��P�C2���d4U����*�N�I�:���}2~��1�tc�,�Ԉ�c5}#&�t5��贽��v��+��kWiYF1��M�����z��1n��j-�gS4�;�$Y1�"��)���3.l)̈́��_�1�s�G�\n�R��1n��gŞƦD �2{g�ugU����sZcF��|��,��Ci� �.�.{Y�R���d�K߅L�z�uc��0t�	ǋ�v)�2�·�C�B*,�
���Vޞ�x�eE�x,W �{Gt��qb{;�=&�m����l��w��mU��Nrzpěmί��`�|�3�"⁫��?'��M�KZ�3`������.5i�W��U��Z;��P�MˊaJ,�.��ǑI�/Z6Ԅ�k�B���$�v pe�x78�Q���GD����:=cU��L�k��a��\�t�D�#��c/�`��JI��Q[m���ؗ��0f�^_�)p|������y�N�f�u�<*T��]�B�p��q�N�5H7"I�o��B8M�r����A��~�-%anO���Ϧ�B�+����I8�K�@"$3Y/],
'|�<��kL�� �\�]
�i1r�hϴ��f�S���ߡhxü.���!�,��ʾ3W����=w [���?=�O��_`�j5�-,_|ּ�Drс2�ۋJ����.&�Ur"`s.F~����H�z����b|	�k4�q<W��D�OBF�ż9�����`�K��;ӳ�Ib)�ݔ�U�O�?b��[$�K�P+�k�G��U�o+��Nh0��Y��<M(ա��&mO�l/��P�Nrr�IRv}�׊4sq���R�� ��yL�����i}i�X������0�؎F���f�W#���^��V/�܌��L��菮�Z�n2X6���P�7��X�_�*�����:�i<��j^)�9B�;i�'px�# f��M��N�ءށe�p9	X�)2�v���w|A��x�Z�atǝb�@��]�=�.ű��ݕ������`�i�,��i>��p7�;NAH�Q�=Xjj�.��~�e��D�n��H�^tQǊA�H�$#�p9�<��o@��4 ^	ԡE��3$!��r��1�I�r�O㨯�z�f�H;EÜrU�"pj���/�t�����k�-�9ȔlK5_�&>����o�>7���0kRT��V���8����s������@ϡ}R�Y��r���HQ|�-�Z��s=��c�6P�!}1��"��n��љ�F�IGݓ�|��;�ϋCɣ�q5��Y�=��^�u>S[|�K��䛑#������m�N�@�,vO��6i�q��P�踾���t;7����W��fࢵӖzNQ�{�qKyx�9����:�bݺ��P�zu��TCq�ӝ6�g(�%� ��*e�9/� 7x��	��/Xb�|�X=���'jT�����@g�����d���yZ.U/Ŷ(-v�ð���q��Ϫ乾�Y�A��6���=Q@�֩U%��yc0jw����^!�ų�C�ȒV�#�#�s �V�TR�^�$[������(�G�_�<��
M̤�h!Qv��������K{n��?%3�`��Yd�������X��k3,ų�\����i���
�G9��*��C�gˢ:N#�=~쎍<!Eq��ZߋI9AɌ��9m�d�S.��?��w�GH5O-͋�!<�B:��5���{	�M�qQ��l���ot�ޭ����Mc�}:4�@D�6X]$����۩8��,^AR[�c�� �{a���NB����*�>�17h��Z�m7�I��F�������2��GA�@��C��o̔�P��a���[�f��ױ�����gK�����V��GB3$D_��!��'�e��q��{6�m�^��m͐�`��M=ȥ
�s��{wV�v��O�>][������Ǔ�`���&k���-V;�#�þ�c Ȥ�+U���˫w�C�*m�*q9?r��F�ђ,3
���,P��emV��&���X�F{���-�|�Hi{K���5l�P�P׋�(�*���\�b:�4[��{g�x��B�Z�s� 3|<�<q�G�������1�k��w�V+K�uVA0����,�%(�T�^��ڕ�'[�Xz9G�v{2�y���E�gz�3t��(��]��Kq�E.�uW�<Ei	Z�
1S��aصx[�<�׾�{BR�3���}�@d�����G�R����@�| ����G����#Р-ˎf�*&�ު���i��ü�	B�}����Y�AB�wF�ޚ2Y��|�X%GG��ݖ�� �U�ܛ����\��� >���2��W��nɬ��e"`LR:��H���Ls�B�5����de�B:�&$�'~�o4��U{N9
km�w!8U�Tg3��o�`��r�+�������8?��c~bn�K1�veI�~"I ��G�����D-�l|SΎ�B��D�(X�V
� �f8�BrD�%� �7Њ���IZ�m:�:]bת�%[EM���(�E�[s����V�џi����!��f1�����d�����>B���5�>L"�ԧ��pc�Q,-?�5x�\Q��܊D4�mTo �*���J�R�\MQ�W;�NWPZyq�}I|H�]��Q|������Q��e�ǈ-Ek����~���R���9���K��Č�V�ID��.��N��+h>�	�f�DIi�
�����;�^��#!�v�Xo0���Mn�\H¼���<#j��	c䡆� �5s�^�ƈ���Z9[�-NA�Z���G�
����1���C�s�������:@ڝeכ>Ҍ�8��#�f-�ē�p�-X^�B�8f6s� �El�XIϔ�������,�b�-&q{`�lDwq�߄mrp�0�NMV
-kf��w�/�M<Z����f�5�5p����*� 5�䭬фj}�V�׍(ֿFc�[�)np^�<P��& K�a�uC�L���:��f���Y���c�(�7<Mt	�O^�)[)�ZtRD@5&>>LT��ꩴ��r2�4�����+�w+��v����1xd�n��y�+�_"��A���ݎ���X>ĉ=G�r���U�	Y�0���A��ձ��i�r�z����a7�{�`�T�����ա? 1�O`�lW��㯭��cqT�o6���'`��	`���L	N��ʹ6�g�I�ˣ�f�5����1e�oDh4s]XD�l.A��=�)7^e���;�,�0� +�����_�4h��phQ%E��c��*��q0�F<#E��<�����1�E��%���(���4A"ʔ���|WH� �/r�HYj���Y���Aa�8E@�oS�66����މЗ��i<�����Vi�rX�u��>�ry=�F�ӏ���Ue?�3ſ��gQĶ��[�Q5ER�=Z0���s.�Z���>2�29��X��ݯbLi _\Q�Ը0h��)�
�e��{l�QǰS�:dd&^/i��w�P���~ɍ�L�ur�/����V����_�xf���;u���\���4R�D�"�>凥�y�`�Pފ
�q7�
��}�g��s�~�����ލ�/6�?^Ȱ��kڊ��pC�}�}%rf��3!wP��7$ڙ�Ģ�C�T�D~�MA�����K�}�݌�
p�'u�kӱQ���d!�6��������+�յa=��>�I)��m��4i��y�'����� ^G���!�*ʏ;�!!tJ�$𼜘;���E�X�k{*�	����AYާ-x�NV��w��X����Y�q2��T��NA�pP�����:�=�ԪN���I�c6!�6���ԙ�.�(Ozw�?(5�j��iX$Vۃ�]�^�����t�'T��}V�y��s�ai�~��N��-=����jX��U�K���`v2���D1�F:{Rj�k����T D}l�\i_uy�{L�d�S��3m�d�{��W�s5�̴<��.Y����y�􅌋�zpB�8���3_��r�G1��bp�#�wy;}v�'$7�π>��`���q'��/��`?++�|NwF�s�y�Q�pH[��^���IܗՑ�҉�8q��P0�%4�D�x;���QQ���kM���o�v>�G��Pϼ�ZY��'W�+юNٜ/���Z�~�kO~nO?'3^�ꛔ��g�:�[//�qm�{?D���~?`J�0�#_<Ũ7y��K���}C�}�'#0N�j
�B���\�(~ɞ��/��ъr�{9��j�["t�y�+�;��	���p���/e���<^��S`MR<ڽ�F{�^=���.��4N�˅RЏ�wގ�3k��[��z�D�jrH�o�ȕkm;��f����8��-��~���͕�ѣZ����}�����~�@���Ǯ�n2�۰�lhK<ຶ���[�b�����R&�dx�v�y��'[����mC���vM��y�a�����_�O3i+�z�����i�3��8W�&3/ۛ_\X�	z��K�&�MS�+�5!bN�K���P�������i�!�!3k+C�

@\3����D=�R#� �f8�!2�{��x�2٧;D���En��2�c���9^H�བྷ����\ ]c��S�&�3���Qwyb��J|��ḡҖb�Gή�v�	��!��� �{��J�����h赛��`��y��d�������:�?g�|"��(=&.F���$�NX2%�S��P�3�*����pL�Q��9 �	_����KA�� ���@��c�=B�U���M��3�K�f>V������͐hGem�r;=<�s	�1]�ާ�ig1i�b���O�z;���5[B |��O��Y��א�u"60�E���Gna.���K�?ŢZD�[�=�F�_�Z����z�
��Z���H�lY�c� ŊM��.�k:4{� �P���}#����Ӄ�bW��oG��ʽmB�����*Z�u��TNQ:b#t �g����ר_-�]�d��Uy]�!EV$�9�G���0qy �;��e��P0\X���D��&�/�#� ��Y+��3bxa����S�U�A!��;��q�^�;��@NzX�P����?����<�?�C)/j��pBH�?�������:ц>kv�ZrzZ�܀hb�Q�L�֨T}D�o���WI��n���d1�ԕL�!^�6i#�{`0�߂�T�}���3m*��1n*@�kʘq��}/3����6�UI���މu5�gA(��p�@X
�Cw��w�+�"T8�l�<ץP�AF1PF3��tD`�����[�l�o��`Oq�b%�_��-��1cl~�_Y�8�̓�&s��"�@���{��v�c��ŗ���	���Ks�>\�=�73L �����KJ�VR?�x
<��6X�I'n-�!>��S�<�$e�q����ս�L}��MM���|��l�Y�٦C4����<�M����ѝ|f˝鐉�, +B�Qy���S�����1_�u��l��o�-���SLL�h�xŖZ��;U	�J(�8`}��̆0c�x��l9D�Ao_�O�4����������C9��5��q�(��AKQ�X�C[�}�w���q�_xIY\ ���B۩M��J��5�p����0*�}nά�?�� ���tFKn�ܧ:|��+��.ں���0o\�<�G�_%�WjJ [�.����Gts�DN�<�r{ꂁ�X���]�F.�/6�9y]�p̸�.��e�S;eGU+9�㞚�VP�N��Dtm��|q�NG��=-�,�#w��RYZ�Ͳ���0V;��g]��S5�� �����~'[�Oo!���e���P�Vf��<�$��V#U�ڸb���;�`j��W )��w>��&��6���OS�r|����7ݑ�q��˨���)��l5j��w4-Ǌ;���r�q��;�)�P���R�ɉ=������K��8!D\��Kk:�`\+�ED�������O�<(ɲؑ��7��8${�j�>��6�(�l�,e���Q��h� ����0L��W�\�K�s�xU^΃��`I��U��X�-��]�����U"=��H�4��v,T��C��Xd����(K�;Ĺ���V���Z�X��EU)��\d�g�:��Ac��rXH�҄�N ��y�����'���Z��l����/����{tI�I&��4��3��g�ڞ���#�L����X���~�3?7�B Xf�H�F%^a�q�u�xr�Ǽzz
�\�Ű�]2��D��6DT3U%�p�E?~��F�� Qռ穖d�"]�K�|M�︹j@ٕ�>:��D��>���8`���p�n��'4]�,�1�v=
�\<u��S�ƈ(���۶�D�� ky����m�ӵ+��T�$�d�м\6;Q�d�����Je�7�(�5'�׏����O�_�ǡ��B�o�Q[<��������UKΓ��P�V��c'�%tmJ����;�A��Jw��+0��g0�������8E�� RU�K8������tZ#lp�X����g��mA�1g6oO�2�}���ұ��hۚy�\B�N�0�Z�>.�آ��A̐���:q~c��0ծ����u�[�^� �U�v0�Q��-�M ��9�{  L�Owr5aK֣��@#Б��E�z�c�%x���i.-A[�Ǯn�ݎ���L�+G퇸�Ѳ9�Q�mVƁ��h�ӭ�im�����f�W�|V����S����
������kS0*BC���PB�"��u".�N6��&�,o�FQ���hFS�m׭���R "���Uz�C�Lc�-�f��}�8�:�V��ںZ����,EV�E�Pe!�

Xn$˷<�C�7����Jܹ��:.(ByC1�cO��Sz ��IW�B}�An�1����I����X91�����W�FT��6�a�F���w ��1��������ȴpt@9'�e�iXVL��琠@��4�;�8��yb(��@%(� ~�P��s�
�@U�C������gƍ�@�%^3đ�'���c[5gB�d�0�W��u��|��)�]�yD��J���{˶��֗���#T�ݘ�dn�;a��Vg�q�B%�h��_�L��a����//L�Qy�g+�#+��Goq@�W�m�����Ƅ�M_��>rve}��@�sy��Nn]��[S�P/�v;>8O{�6	1/(�np�#LQ-]=q����~>m
L���[!�^sg(��P$����#Z���kR�%#�p���>�E3�_B�Mten�h�����gE{1��㞅Xs���I}Pޫ���L�V�ރl�X�T�?����ߨ�3.�/'=�_Z�O�,�ݐX4���dp�da�{頒�}����4[1��e����>�Q́XDD����}�T�n��E��kK����F��ς�T�q[�潷K�}��$��_�m�K;�j[	��/��堂�{�hoT�����]$rءl������_��PҞ��