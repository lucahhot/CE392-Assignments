��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�A 晶���eŔ�4����A�PQ��T�����cSZ�Ed�\ϓ��ۍ����Sp����C�6.���.���A���Jľ�wB���6����5�?���^�ɟ>Q1ǔ�B�������ɢydټ���\�g%��9  �r���cGw�Z����ۇC��Ȇf �%�۵��I�i+ihvg��eU�&����^d@������ҍ��$Ym���@��`I;<q5ЬM%���Ԧ�sʌ�wSB� _!�GJ���-pR�wo}x~7,�T9��
��I��Μ踜�BصŪ���e���l�i�T�I?�"��[�165���=L��܇�=��v9@�=���N(��J��v�yE�����Y���2R8
���V&��`�#X�׳��1���ye���Ӂ/VG��_���ɑ�%��C����ie	ɭ.+�O��a��P�~��$�I�yYl�E�J?_��]UL���	�Dd���8�c�B#�מk���°�m�؄:�ʛ�ob^��0l7R��J$h�Fj����(���q0R��Ե��r[�B�К�oa�� ���r�@>�qY�9;2Y)��MTz|)�3�p53��v�R�Ggt�8�A��%���k\��(�R]��\���tj�^1g�X��~>�O�C;<�A�0�[�J^� �������\Ѫ����v/?�+4n�/*�8������0�-Zb=���j�aMz2���4�����o�:�~�h�:�n#�T�O9�F�x�a3���u��@���³;9��"|����:�fg��l��PǤ ���+�M���50&���Y������t$�8��PK�Llσ1��V��{\�C�9ѭ����Dp�cԃO��9 �,�V�DQ��<o�[�z,[�S���j���70�7����"־k�"�ż�d�.��ѧ4L���d�XG�q<�B�W9�!!�S��GC�u���J8 �#�!�}V��un�Ы+CI3�F��JP6��E��I���:)���\/��_A��3Ⱥ`�dY���F�G�����G9��q�s[4�O2����	������B�ܮy��?z,C�'Zy����M7?9�'#˂�c"�����eG��q��?O�kF�ǠE����>D{�װ��������H���T��İ�?�j��(k�C\���_%��ƅ���f�ԅ�T@�{ �����J�����w��j�r0_��A�G�5Ͻik}�o%R�S*��6�^[}g���Iv���Q����1��q��{�u@q,JSN�N�o-$?|[B���r��|(m�S�D�:��_b�i��Β�����R���a�g����2,��Г�!<N����oc@T����08��� �R��k�霳t�����P��wʘ�B'��8C�5f�k<�<�$cmj�����������Cڃ�b.�A }v�/�CԐ�!�V��ɳP��I��!��G��r!��1'����xϪ2Љ�v0\�Z�~�������gP�����4W:{���tf,�6-l�m�3xYHv݇"J*�%�PG��C��i�ym� 9u*��C�i�A��8P*$������"qЁ9q�F314��z���$u��9�fqRrF�<���:=�YC7��<�UȰ���_��)����s���̻�J4�X�� �t��l'�%+��N�a�3N�}	�H�/�q0J�+@P����������vr�9���E�2�����j~���/0���r�~��[�W>V�W��W]�z�ݪ�]����v�b���u��VضN���sS�}S(o�7)�t�W0��`���a��@$�J�օ���4����p�u�n2�%A�/x��L,�L�Ruw�X� ��ꎚ���Â1ؔ����skuq���y4��~|b��{LRΠB��Lt����J��ĭE��uQ�N4���N^='TR���7�w*��sZ-�U=���J�H '|��f���G��UM�	�:Q�:����|�EB�_*:Rf1|�h+��*�lI"�J�C߄�=��b\<��1����0"j1�m>FSp�\�X�ث"���հ}��ީ��֏�v�����|ĴA��(� B�io�S�ԇϥћ�ʰް���UX��M+����i#�V�r2��W�C����~yù��*c��3Z��a� �w�Q����w����!M���]�!3���!���i���3%e�����}�Xgg����$&�>z���#�1�4m��G������x0���2@��W�M$颋�8��JP_��\�0��u;� 1���%�.�(�'x&��Db�l��V�5&�{�l��ק 9/� a�������:��E;��`�ǖRj�B�U:t9�z���St�`������^�G�?X��
[k�z}���6�F5�d�n�����箆��(��yra���Ir��p���52pK�>3�tw�֝�#��"
g.y}���`5c�$�b��G�}w}�j��Mu��l >/~����,�r8�PXq��\TXx
=I��=�7��zMrM���h��LZĿ^p��T'"��Jy��'���ɓ|�����V�Uq?��a�%�t���O�`P7φe�<D����: �Z[E�ڍI��2���F�5l��O�9$i4�^tc��m'��Ђ�J%�v����(�[J�l���Y�RV�����׍3.��7k�`z�ױo�������l�B���/񙇃���9��SljP���� ��ґ#Yn�N����H��}5�K2��_S�X��,]#�������Vg���~'sy
�/�ꛏ�{���uq�kq&��ƥW;j�� Ig���jQ>��鹵V�����/��'�ז����\lA�ڀ٪f��[�OتU��*-&�a��U@R/�2�����i||U�*D��W����c����؋F�ׇ3'����z@l�u�6H�q��+J9{2=�(���G�%����E&�>N�V�>Z�����ym,K���-��nr��?�m\s�O0��VǮk�!��j�+t�"քm��Ʈ��?��'�i�۔$���eD�����w�-]׃ֹ�_G�4�{,�l�U��꧿�	sU��g�O�,#�SSi7فa���*I��ee8^Mk�����)2t����h����6{�y���-c�ܖ�>Z\�8��Zhtj��\���_&8�lƸ4~¬&�*����qu�7iY^h�gȪ:�vG�v�'�:lđa�ő����S�Z5�KrA�C�$~)\�����oW�zr�+}h�Rj`��3J�S(��\�`�T���P�*���Gq04��2,
H�r�)=*����]�B��˚�v�}@q����K�נ$-�b��䉏ZS��N�0����_�N?(��,�C��cܳq��ea�-�}+�Q��G�Y&������[^���$�*�ra�1��fJU�`Ą����g�6��.�YT�^3�-#�]��?�2ݺq[�W�y�+��_ޟ���Ĵ 9?h�起�������؀x�.c�]�Z��Hc�+���4��5{f�01�@��zĤ�*|���rǴ�K�	wk��
�x�&�:�Su�_�H#���SJ)bxdˎ��a��������L�D�A�G��.��,�����Q��9�ْ�޿}o=��@v�(S?L�p���4%E`!���c��Ek��΢�z������a��-K½�7�Ș�:񎶯���4�7��7�r�n�8r��U5,]���rg]ڳ�#o�I�Ac=�'���59�M��HqRIG-�Ҵ8����3O�TqP-ZO���6��`I�SM��Rh7�9�҄������.Y�)
a�_c`0��Lb#��S�P�aA>fq��-G���U���5�?2-2xR�Sbm_:�.�]��J�go.~��!TN���"���@��2iz�h.�Co ���~M{h�ѐpE~�EG��-��sf��t�n���Wӛ�	����?@L.�޲͚pP��D�;{�uB��/��G�8���������RWd_*��:Ճ�Hٯ|ݧ(��oǤ���l�/�(~rm�T�ށ�WRo=A���|��&��l���׳��W�����a84���4��]n��d�Iׄ"�;��3��#�۾U_�N�#L��=TVk,+����|�1��B;���K���.�^���2|AI2��t����i��t�>����Qd�௶�&�G<)��!�1���e�8��T ����Ԙ��.�*��[{��`���1������C)2�C�e�2PQs�f"n�ȵC
���G�z؜�����^���<!eڱ[�����[đ�5pc����0�����4�$R�JtI��  �y�d �����.�y�|�/p� D4\���1���T)o�T��J����}.l�����d�����h��8����/%��܀�AYi�{j�7��������(��5c�:8c��ìy�=�>����f�l�N��<D7����
ʙ���[�z/tŻQ�� 쨓M��k�֖}����6��P�E��.�x.�ɪ�&c�h���!9��BZ�� `��t�w0�&�`���r:���̲�^�F���*�A��2 ��}���h���Y`yA|��H�� <P9ۢ� ��8���ʳ�a�+��j�ʄ�zi�TuZ�><*�"��"8�:d/!��[��S�ۥ��b*O���{QR��{Vi��riVX3jUf��d�b�T��)�gk��j�ʁv�o* r���#ƨ�y�O����V��G��lǽN�` (��yK�^�6RJ�k���D*�e���>�6;�2=Io��zP@4��j��2rβ�_�o��=�D�2��\��/&��L�U��]E�JCa����'5��WE��i*#�t��A|�J \'4���3� !G�D9���pS�Մ�!q3h4����-{�/V�cP���t]��u��͐��%��3�V�A^�jI����2�7�Z^��w�f�v��r)�</c�ؐ}#�av�!؟B;G(�������Tw��?2��h��,�/��+��C$���v�&�O�!F"UG�!��p�L������~�Q	��,v�B�Mc���d�Q��$F��k�d�4��>&F&��;���b�QC;v4�7g�&f�B�˚����U�q�0>h-ۧo�?j.?�)n�S`�w�F#
�E%
[�t1��ć������;���ڟ^�H����р9��w�|��w�����@�|�2��h�f,�9t�LUuN�i$�XB�Q$�-{.��젓�5�:P�ѥho@����&��6يY'R�*��.���Z�ϱ�3^5��ž�h=K s_���	�EE�f�ؾHxp\s�|z�z�ڄ��d��@'D�,na��$�O�7x��!kB�N\[���`G���愮��dҺ��%)&S���"E���h���3�B����(���WIq� �&�%5��n��gw"�1�Kp���9��]ՇͣpI\x��cv��,��M�`ef��U��R�x?ת�C��.�p���޽��*)5�PA�B������O�G�|@�L�qc�$�ʨC�6X��*Rn!������m�Xj��0����01	�^��ξ�u(0Q�SJ�I�U�dy6��x�UU��c���~/�3L�i�ny�C�m�V����{���؋���ZԠSv����c��7K]`�U����!�1j�I�3u[¢��VY �街��W}��K��vlel�Y8��Fq�kɀ����.���9�ȋ��佮�4߰�K9�ջF��uU��Y�Pg�4_�4� ۱o���͛�G5�������ÉaG��Ì��&S���m5�_�D�������sb�r�C�y���Mg��V���߬\i���k����CdJ�گNk�١jʠF��޺X��FSJU�Ӌ��w��<$K�1��$����S��D��߀�I{yU~GK��׬�
5���I���#~%H���s8����B��>+��e��U2^��b�l������չ�6�I0^���=I dk�N�k�|�(m0o֤��=�i\P�=L�z���e�%Is�c�u�Du	��.�g�c1}�)��nB��ߺzŜK ��|5�<:���h���w8�ʓ*�H�~ᷟ�����	rxoS��;��-�OI)��
9i�il(�-}lG�c�SB���k�~kV�����-�S|,��=�:tur��1��2�t����v��yتS�NL���QVx�ۘ��ד��E�W�u�J���ɠA��n<�B�F8�5n_�T��1�����_��At@��G�w]}���ƛ�'����ؽMds��)��/${�&�g-�'&�M~��O�z*]g;�j��Y����D*\ϳ~��}���o�a#�3�1jb��*ZfD�C�[YC��	�{�%�z��W���dU��G�;m\�b�*�#\��$O%�S�M�L�����-; �)�S�ߋ㻸��>nw��[�c�?��LR��Y���݊m�ź�ɠp�,�I{,�W-�<�Db[�ڧ�V\
c���WI������|I8D �U�Gs��*��Kxc�,�TʒC�Ѐ�ư�YkF��^��y����`OA}۲�9��Y!Ʃ���T��A�Roajsf�'n�^&n��َ�pW)��Ib���:�HY

�-��$Zy�Z�ς��'TŠް�&sZ銩D��{��]��c�+����������S�6ω�E�ܵLǴ�hT�#Αu;����߇�x}N����DX�pmW�m��OT��h7F%x�n�M#y�vv�R�>��Z�K�
gy�~����ҍ����_��o��&Q��Isc��h�N�ݜ�q��c3���#��<	$�:��/q��|�̉,T;�U�6%��3�W�V��
���Ҷ|bE����.����� F�m?eE"�:�]LUY�1;	�'��}�*q�o�[��;L.٢����d�,û�n�M�����r�H��K�5֍�n0[;�F'	[�5$>���#�1;2�Y���p߶!��B���D =��]&q��ߒ���)*���K��8�njh�ߕ�q[��+�Po��ܪ�?Y��y;,ˏpϦ��@�l�<%��g��%��Њ�oO���2������^�&�|�3������̜�L�(x��"�Ty`$�V��ɋ���q�ma��Ȳ~��H�'��v�C79�[Ҕ�}�1`�X7j�থ�QS�kjġD� ��4)�E~�wF���YZ�%>�T/��ij<���w�0X�/zT��uo+`���c��R���A{���OU���! [\�+)���hJ�]��+ދ��>�r��hb�AM��,��;Ye�4�^6��Z	����i���>�[�̛�ޮԂz�@��;�Tr�6gq�L'�9� I,ׄ�9���<��gF1��g��8ވ~:�f^T�M-����[dܺ�V���5�tfT׹�[���������Zּh�E�:6Pz�}JG�:��Ґ�XGN|&��<v���!+hy�nS��H����z?%M.������Q#�C�w�lb�� oJ�w��%�{)XxT�����q
���}ؑ��)�$mTՆ��x;H�${D�[��=z\w���\Ά7tи�D��	+��=t⍃�(�"�������V�[��D.�E��@�֗�l$�6����3��6ʾx 1��������e��mo����C�|�۫��s,b�Y�E�9F���,�`��
�%\�	[�5�?��l�������7r���U��v5�����N�yBg�)�V��x�H�����W���KB��32����cp T�^�w+�]�J{�:=J�d)*
%M�P��H4Ɣ�-26����qS�X��0i6ja�֚\w�a���{�`�ɛ�þU�J��a����TgRY�[��X���P�N���T7���4��Vw��,�`Mɟe����@ �or��&���5F>'txyX�Gx��6�����ŇZH�Z[��K��"LƦ�sIʤ,���`�y��_mR�ײ;��S�M��ݜ�*g���u0�ˣ���M�4*q��}�F��k}l(�����c��j���\�Y-�f4�h2�0%P�B3�v�^$���^/�9����ܱ������v�OΘ�X�b��j�w�Q♅E���F�Ȉ榈N��)�db��g�#a��_�էM�짧���}��3Тsq����ov/k�p���k�6]��h7݄Jk�;�M���헍��;���dC@�L���u&>�%1^��=��qF�/2���o�ƿ�X��fpaCi�����ߐ���WL�^�� ]����}�!�@��TI�I�_I4sr�� �΍ۍQ6��ݓ�E�K�(e������৾�Ǻ�՚��4͇�OV|�9�ڡ3*��Oΐ���9T�*��2��n;=�@n������`w�2i��$R�TC���MBڠ��ƊK�t��?�h���(�
-'���@��T�Njr��H;+��b�-8l�/T��Q��Z?��t�^�;6(3z�G۪�>���O��/5��#Ī���N�p5��kaa���׺�W�.WTI����ĝ���X����p���z��j���]W*+�@-X�`jם��_���9�ق)�#<��Ƌi�	
ᭌl���\�����E�u�VBVתƑ��;I$!Ģ��n$Ms^|��є�������t���uI������"��u6���ǿ^�������)���A��$p��b���3���/�%���l���i���qf&�����5�^y�W��v0���~fN��bH v'��j�6��*s��yc��&Գ/����_�Q�2�k�(��,ᙊ���c�x4��P��>����ХS��t�v�;9�u�����L<N�|!O+���\��#� ���������ىZ��T#Z��U���^�/�+ʲ��PK�<qV��W�CW	-���]�/�#7J�L*���S��9&�����юYq��'�e"J������@f}%w��J�B��=���RϾZN7�{J�F����?�W��U��'s؎-$F-�y�m�e���ؾv+Lx�������=m�8��⏎�a����$k�`�&iw*��%�VG�vI��x�Ƥ$6��_ј)��YD�(C��9s���z�BZCe���rY�1K�W����a8y:v۷��f��¹���M@D�X���lZ��o�Ul/���\p�S���A���-�B{�xˋ{B-����~��'�C��Y�ܻ����]NK�D,����e\>r�1��� 9�<��(A�����n���T���A�grۘd��9���$-���dy��a�
�@��w�+����8x>�`�8��0:����O7Kh%�^k���E͠�t�Z �����=B���W��V�>'5���;�p>:ȼ�̝��o���.�����8d��$1-.ϒ&r���]A���t�x�+6���Hگ�s����Fb�I��Lrn������+e�~��/�M� I>2��N!�H�� ?rU5��F ����yȸe-_�����Q�����M�t�HV�����Ä%���5iZ���io��f�U>�`V�f�	F�۰K�Tpw>�5ٗFI��&8��׎oJ,�!�F�\wb��\�8��*�G��*����5��!l6��h�#�G��,�y�������-�l�
Bz���������p��8Aq
Y��@�ڃ��ӻ�k�=Z�)-\�A�*Y�|ʊ�+YXh��h6�G��H�o��.kGO����}SX�P�'"���p��`�O`;!�p�:���җ[��&���6=�1�j5�^�����d-@ ��xq�:�Х�=�lw�
�FB{��t�>�iP� ��y�Σ��$J�Փ?#��՞�3�RYp2|Ǉ529�(�w�BJњ2���~���Ɯ0�/�^@�_��'v��j��Е��U��|��װtZ�DP�L��>*Z�ep
��e�0DpY<q����򇳛�<W�m�nY4)�h��� ������sMy����I�fn��U�?���N��dX��T��)߁�9�u#)���PV%�,<���a0>D}�&�Fe�ޔE1�<����R�?[+� [b������N6��0���[�rW�A��x{+cA���}����0c$z�g���*aմ�^P+���I%��͌�j��}�4��<�4ރ޶^u5���[�ŧ�+��+�L3���jh��p�q���q<r!$�\H		���ũ���5�s�-u�+؃Xpi" �,��F°��X��k�*8­�q�WZĦ��;E�.�*���'n{��:�V��";�|O�%�5u��^�|��ɨ�)�	�/ll��9�+��T��~������'���wA�f�/Gjnf��ù�G�ϸ0�f�Ur��d��׹	ę�%\�N��i$�($aX�:��ͨ�.Å�
���k���{����	�e9�k]r^:�T�6j�\t�f,��3��P/�j��(4j�~��Ф/�W��T�����C��������b$u�OuyH2��8r2�p����A!�0��G�;Jު?g����~hiV�r��#����ܫ����t�\6A�A�T ½g9�V�'�!�_k�f�5,WA¡,�&�,��K�?n�Y��j�����*!MgJ����8E��A����h���>I����G{�w���T����sJc`׋]�S3Moɽ=�V�J�?�7o�!@�	�s��B�3SDp��0$(�60�fqok����$�N���lS]�*��$�����9������]������e��Me�Or�]���!u	��|l���m�u��h�MQ}��2.�R|=Ш!���9%�#�I��@�����L��k��;O�;1V�Ś8UK�+�i��Mi'���W�N�����Ep�Fu�Ї��: aqp�f1K���\��v�2a�;���`�	�}X-4��A0m�smSɕ;-^��+��Y�72��u�OMhkK۫VY���5<R�J[(&����� ߖ�q�Mu)2���������J��4�+I�@��7;AS���^ߜM?
<�ц���eZ��7��y�Q���������Q��
)C��Ck�RFY4p%�c�0�;ꥨ�(�hϑd�:��o'�XH�\1v�Q��`��=�9��n���?DKX�qX�!��sR�׀�`�T���h��y,az�^�o���Iߞ�1z=���4L�+�q�Y�xds/n���Z5�����2�Q(�-*>
��n���P��]3�F¥v�Ŭ�
B'�w�bw9��1}�ށ��S�1�D�_��H*&�L�1���WB����i����v�s�xC��q�6ݫ���`��/Kf���6��nga�C����6'���kU3݀h�t�r��-�گd3~4֠��6�V��<��)S���8�_ s�:yF� �h�����P\ő�^���伇i������p���h����9u0�E��z&���6C�/�۔�3�k���p�St6���ҕSEҝou�#��?�䴸�}Ѫ`�s�W��}����~�&<�"fX�ӂ��~�O�~4�G��0o)���3��N�O�d����b�d�v+)�%�PJE�9ѐ���Dެ�w�B��'~�q��|���2��B���&O�?�n�3�,�jOr�5��y]�6�mmJڮ���XOʲsb����i�& C'�s�9����F˩ފN}T�P�$TdҢ]p���
�^ &8��oY!�C��f�`҄"��ʱ �s�4��f�������z��u.(�h{O֨���u3��	����x:��Ή�j{���by¨>)f.]��t�(��ﺐ���Ι	��Qr�\՘�W)<�����C_�q���5sk���91e^=�[N;���
�U�䂴 �Or6��(�,�胣�tX���S:WG�s~�������~�"����}�ɻ����1F��K��7�5���S������*!�N�&�7[��޴0�����?D/Rޣ�:ɕŽ�>�Hg~c#�#
����-1IWwr���1�%:�bIл����R$�3�M�T�r�7�:��߮�;gt`�q��=K�JPf6_O\�d�W�730S���5`��y��U�F���<�1�%��^u$��~*k��q�Hp`��Ilf���c��`;њ����l�vtU�a<ZPh<;��CtC)��(	c���g�wt"~��+���PyZ�Lɬ;�Zݏ\9��H�`��{�^$����g0��~�-9��#��Jǉ�f�Y|�jM�q�{�!���DF#�_!]�M���(N�O.D��[	9-)�N!��f�ì*k�֚h8�EG._,�#��C���[�HE�X�-=���\�鷮���CU'bpKe+0����P��O���Jn�1T��n4��1;6�$)����Q�ń��p�J�Ƶ,�� >�?�q�'�ĚT�	V%��X�w��pڻ?�K�V��L���B2'Kv�y*r�5z^�h����e8��&�TM�����I9��~pܤ�h�+�ū�h��ec���=��T�拫W�a�U�����* �����U�EF�y}��cSDNփ1u2��%��B!�jQ����%zx�\�l�#�C��[>�PoOu����Xi�
a�b!�<y#��e��vu֐?=�� `�Ԏ�/�ս�Tw��Yu@�����(H���?�D^ŭrwz;�,mӒ*�y��T�)+ ^is����i��|Z������+r���q��4�����sFd"��u�|�kuth�h�6t	�!E�!� UчH0|��>�B�u ޓ߸�({?w�{��=��y��8zD\(t_�\φ*��EE��N�P�_~ӅK��%�"h�D]1fv��HN�W)�O�n!	4�(�����X@(�۱(nH8����
�f��vg���M�A�|`ϧ�մT<>�	�C����;�{@A�б��/�4��F�s���d�����3U�	�۶{(K�C9ܵuN�=Ԡ�U�Z�#�&�6ިX(d
Pg]�h��n�:����F�5��]@�v�g�UI��0���H�Z�u�2���h�sC��� :#ӿ�\ߤ�?/;v�'%M{�v�G��<����"7g��;'��M�����������x�`Ђ�7H�*Й+y��_$���]��ՠc�/ns�η�Rz<�]2F���	'��oZ"{�z�MX\¹BS�K.��ӿ�n�M�2�!S5���q" ���x��,O,���&1Y`��CLe.�밪E��'$�{����S2.,�bǘ��͹��'8҄� Lh�������������B���w�g��N�n����!����C&Nq�s�� f�<vɀ(G9J��&%ؐbD4_�p��	t�}�3����)�$hܳ�x k������I�A$=�g�!��w{Uk��4�� {�룵��e��߄�[do+���(�m��o^�5�Z�+�w�U��;��� �8��a��nu������_�<7��`1;�kQ�;��y�/-]�ua�C�.|�3�����p�,X�+����P�!��v��]{Cc��v�e��j[@ى�ҵ�!&��5.��� jbZV� �u���r9|�YC�l?B΢��MY�o�)V���]�#(��Z�c]h��	v����H#D�,]��R�.G|^O�D���i~�����|n^����@y@�L����0��
�CɯlB�0�FXb����;[��r�Fw��P���񱇩4��#�{	�|�+�Ϧ&ҽ��j��aL�,S*{��4����;>�(>�_(N���L�9�#�s����!d�1�t���
�!dc��(w�6Αp����aEqʈ��L���iz[i�m��
ſ���OHe���g����{�u���؇�e���6��pT�|��
n���ϜӬ�������X��N���Z�S�:j���\� +����',Yܘ�n�x<��CD��A�Ypa�2(i"��9�x��o�/�;�0�y�) i��2Cd�B��X�R"e`� �D�*�x ��t�x�1g�L��GE[�b�����5韐.�2�����~|��5�������k���e[���P���P$r�@t��νA�{��fӡ?ĖW����C�+�L��X���ͳ���zY1p����W�K[��ǎT �N<*��7bȟ����tF�Cb�R�<��k��Z���S��ݐD+K�_��ޡ�����3��m�;h��xn�i�xo����ڔm�(g�m�Z�M�Sgo 	r�$ƻ��\n~Wx�9S�"��=�*t_���������h�xV���`qƨ0�b <�<�p9���d�+���u�K_�1�����j@�s%�:�W��ԡ���%��n�a�[  *�yVr|x�0pª�VL���u�*����D�x���V[U�\��P�GK��{,Of7Lc�>ZR�Y
c����ꈺ�`t�d{?��vY\�t���`e�}5�z�}߲�Gk#T�3��kk���W��-c�9w�Q"�j��%�f�WD��[��ݲΟ=���X�L�LD\.����#|L�c��M�M����Gߙ�-}���剭�)������םj�S�j��N^�x����`NʺO?�q^�
��$C�!���;S�auZP��I 0��ϑ�oɠ2Z[d�8`���vI������!�
�%^�M:HO�I˓9������H#l���A�W-IAY�mK��&3�is��m���ѥ]:< ��I
)�̽D��[J��ȷ���9Sa.�1���5؋�0K:��,|D;�=�N���5�׍�Y��sI(I��m�*��'���׆f[g��+0oe�=���@��,����W��@"��୑ȍ�e�-x���Z�P;Bz3��>�G3����iH[%y�:JU�K�E�v5��!�c�aݽ��Q~?�)������Ui����kQ��+��}�o`��O�$9���'ç��6�9�P�T�sڧb<�;{�ǯ?�K,	 �f��Rl���5�Nk�-
��A�f@Ѩ�
�]��}��� ����դ���J�Ϻ�f_sʭ�'KȆ.�!�o:�r���(�-������Or���#1?ub1Cn�T6�e"��K��$�Һ}Y�S�z���v�S9�CN�ܔ� �:[!K��v�ܦ�zo���z�Ж1�����*;�o%��6No�E:�"5�*�#���V�M��'�(�)���Z��L"n���Ż��1��d�\�ܣ��WW��*�¡H��S��m�J�����N�!?-��� V������<r9�jW]�A������]"��úc�>[`��mIo�lʹ�R��&��JF���1?�.�Rt��@��bʯ����:+p�		]zl"
���5����64���(�})���c����`�I��C�v�b��ȝ�V�028�l&`H]�7�6�R��vL ��<���b��S!���y2�jg�:�J�3����<���N"��ٻS������+ও%T���;~o��6�L����w�vt;�6����l�m(�t���<R+��*ER�P�|�$��op���t+j|Qq&�(��@��-�Ǖ����7F�c�����(������{�z����u0�A����ZO�LV.z5�'H�|��� |�"Z�2$;C���
�J��`�P�ձ��Wz�i�C���B����s�o'-���w'#�	X�5�j�$�E�N���uѭvos�ؐ�qtNa���G��b���M2C�������Y&&�Z����������X&u;��0&M:?V�O�O铮u'�=��k��3�cT�o`븅�`A�J��l�w���g�����8���)��,۪��~�����=�Q�{#�]f��ϱo�S������V�Yv,@�&��Z|�=��� ^���w�쁦�����}a-{�]�a�v��P�RO�.���n�y�m1H8V�7�%��$Y�cY�]�8�Em�Xvb�I���6x�}��9t��	���˼��4/��Y*3���
�����n�onܶrX��<w��h\��˾�Ҳ����Nڭ�P� ɀ3�%���{t�#�b��o�i�m��I��4�5��z�_����3�z!�����H ���h_vQ|F�_lD�F��8�n�e%���I�b͜�!+(/�)LsQB@z�Aƽ k́62g��E�E��mh�����I���0�6����'ͩ���=���Q��}2�����)�>jԈ=�h��ƫ��P��Tq艥�>:Bm&k	ۂ ��0��Q�q<��V�n�-|����6�lW�F�*`Ц�@�yq_����W(2ΐ❏�G�'9W.Z�`Q:VL��gK��	P�.��W����h��_���R�B�<\��9��>�5��2�!�uM��z*͖���!=����U8��z�<4�_SÔ[�y��H;4&9�a�(s�r�[!�w�Wn_loU�э̉X)g�tze(�M� ���@�&���>Y��MF�����:�e7�l�Cu�:Ggg���-8B~���+��y�տ�^NL.��`���(0Ѭ�n>G�Y��^,i�b��t-�������5�$ȁ��хFKr7� ʬ��'L��h�P�r�!��9a�1z�7�:#��,���F��5�co\��`	��Y�8�պ��'o#Q�TE���*̮���@��4���Qn/!6� `�_�	Ͳ����(��D�g-Lf�#����q�����;R�1j�A[B$����^xP����OA�u��NQ4�_:21hۙ8�/��[;bl��I\�/T�GϖP�6X��5�����=|�۪��e����"ބ��ab��Y�0��4��4w��NE����3�~5ͺ p������	��ԫr�p�9Q�Fµ�=?�է���2r��{B�)3�ɧL�I��'�>bj~����؃�t��	�!e�X��&��Z� �B�'�ZO���u�5`��^z���F�z��{7�����\�a[���c�`�R���I,!��wn�_�؃.����#�?&;񵮈&w��z?����@�g;�<Ƚ.g�O��y �V�_�աg*A`4���v'*��R��an���K��[i$ܮӢo����}��jc��4HV�q�k�m�DU���-7�l'kb?�N4�-/QV����6r=Z���3�] �y��C����:{�ŕ��^��RX#�#"��3
'�`�-�֙��j�����������K'׎����r���o��Zf-���|\���6�U$�$ն�����:���·w��B��1�b|�zM��O��#׮I'rR�<Y�y�'
,G���4<�mԗq*Xq!ࠏ���x���}�6�|�yݘ�Qv<���4۫AZ�w,y��Z����|(ӵ�y���۽�0	t�yW�3����FW	�-0]l�_:֐B����'hw��x&Z��&�Mn�9���zs0����ш��1�g�_d�"/m��ilWZU������d�)Ъ�#�9-�Lч��5�lY�8�r�L,����z;����{D��Q��� �]��׍f`>�[ ��Y*���q��\,�yr������p��m�%E���Q
P+�=�� e
����3�$v]�4��%�mG?W�t���	� tGTdp�̵���8��K΂�4���ߌ��z9Q�Pn��\���T�iǜ�(�nSb��{�fs�y���^�ѴUA7oeh�&ș��/�]<_ ]�z�?S��E�*�v����쳣�F��|��S���<�e/z$���q�|X�w�w�ᓓ&�_�U?t�Jۢ�&�Sمh��D(�\	���.�Kޑ��Y�j)ü���P}H��j!ď8~zY�i��;f�׸w:n�qG��7>����a$�<���v��㫵��Ts~�������o�"��-*N|'��46�C�B5�f��Oۯ��汐�my[�_c/�q��<���K#���T.O���?��	��$1��GZw2%�5ľX��\7`��x|�q����:^PRvec�TR'��ݹ}){���o�,�}��w)���u>�*��O�,��[�Hl��YxFE�5;�91�L
f���tA�E��9�ç2L�?��'Auv\=k���4E��!h�*ڸi�q��M/�Hq�<c7:cH�}�U�q���^(R�-��U�$��6F�0h�� �g��� 3�^A��{>,/�j���?(-�Y��wD�~2K���r}�9�å��P��C�b#��$SnRY08	jq�݀�q��j�wt�o��K��T�+�=��:���t�f��a�Ǿ����uջC+(�^�	ݓcQy(f?�����n!�kiD�t����?곲���𥮄1�M�Vʽ9���w,&)����2�:�:+@�V�柃
�&��S0v�������Okd����$���碧5���D~�:�0G~�<��V�BÎ��̖,C�Nat�9DZ�ZQ�H�*{�ҝ@lÂ �4G1~�N6|��i�%>JGb��?{4�YL������oE��/k���8þm�Bx1s��M��mej)��î�,j=��eV�)Y�>`�A�D*=�E����T�BWʞF�5���@ǉ�����~<�8���:0n�v�j��i�	�x�n����j˖�Q,��+@���t[���N`k�L��Ѫ�q���ҝoY���3!�u��ubq�=�l(Cbw�E��c�[ROLu��F�>ܦ�u?-����]�������tF{�"��hc���@&bHڎg1�á���O#d���n��ǡn8���Ƃ��:�:1�r����ӞO��{/W�~�|�w����ۅ��bh��͚��p� �a�-(��&�ꢒ�G�B��7eܖ��W��I >v�� �r\R��r���W����Jm�y�x�2�O�Jh���JdW���%|�����M����A0�k���(�zw��fx/����5��s���S1a�����Uٹ�g�[�Mx��$(26�]M���Ɔ K�\�ۮ�@fmO[%������}Fbj�B��Pd�X��i�Eck�:����)��c01��-�4��x5��T��f�����F�'�l(1�p�TR��W����U����:O��苈��f��oCe.�1n�#{��T����k6��~,t0ޙ~9��#"�F�%����K�,mLsщ��P��.�W2��D��jZ[����0��Oꄾ�/qg1�Hf���+��JU}��[&��G��������B����j�����Î�Ӄ�oat.0�펕p���T�]�m	��?b\��D��o�ZvRL�G�5��l#��9�uL΃r�J�tf'i߀��^���-0�,��3,�U捴ߞڋ&����~�eb`��R�q�,��TR$���5����0)2)�9��NS�u�VVJQ>Wj�dd�����HI��>���Zq�>��
�
���(ߋZp�-���`z�~�ٚ��+ɲ�iƽ��W�9�����F��fr:�j��i�#t��8E��$jh?K�U޷?� qm�ҖY�U�?Bo�C��<2��xh���	XYG��a�]�k�es���:n.�܈�t��,qN�Lۑ����f�3V>���ñ���6�.��-�4K�E/�?��3'�{{7�Ż���\�N?=x���
#*�<�<��驳���H�@�OY��/�����K��>��2��'���a�y6�@Wݻ���0{P>�
��COg�r�p������岈|/r �S�ن����ԑ4r#T*J�`�����;^�X�T�=�pOd���؃3@��̤�f����	�J��I%���dO��f�`ѻ��g��R~/&��8C�jX��M:�b�7ӟ��c�nܲ��arRGCJjJ��g�D�zϳ���D���X�q5��-֋_�2*�)���_�Yz7�v���8i�g�EF9+;���Ջ�q[�aB6ͥ�����P	�>^�\
�,��k��\\�����S�,	/����X[�0�O����"��e���`b��EE�����}U�|L�l}v��ڇ�<CN��y�iE��1���|��b�Eѣ�"�� .����/76��!G�)���dmx���к�Qz�s��Ɏ/���6��(�{��i��_���y�T�Gm-�������8f�z�_T̽ub9�+����4���7���5oƸmD�	�+�����Ag�W�f5���+ZXzg��=�!%i��h��L �_���g/M��pg�Z����6 ْ�G��CI���o�qo��?�1%H�$۸�z]V"��}z�l?i��.H7�.�Iu����
��H%���#������%\37�#,��
��7(u
]3A��O7���6% �rwN����Զj�z���%A)�f�a��<f_^@�I���f�b�y���r�Λ���@�(/Љwf����� }�b��~��a|t����s䤩��b}H@��zй��cK07�������z���;���Q~0)�4u������WD2*���N$^��I_���(�m�5 Ͱ�-z^VJ�P�djȿ���Q�q ���K8����U��AɩH�VI�������\O𞔒�i[��n��R�j��u�\V�p��,��G���~��3
ׇ�IM��yI7�kC�t|¤K�.�� �W����%�_i]u_��SE�X@��U�H��{�3�h/��Ҷ8/w�'��Y���$��]ϝ�dp�iTcqPS��T����
��_t�Ӝ�P$궗��͙ "�`ۛ���bBk�җ��w�I���;��0��z�?�m�(ԉ�<.�C���8�௪qz���Ԋ~��'����?j�0��.;�?���2���D���mYI's��g�� e[��d���Ԉ�R� yM�R7\'Ok�6���][###�ر�
>6Ѧ�TaX��#Os�v�f��3e���f8_y�P�1��HQX �KY��W�'������%�,���
�����u�bـ@ٽ����- F��2z����{ �.����rg�)�^(滭_Y,3vYGx-��|~f��ҳE7�R��q�݃���Hsz+d�������O��w}��yes����ق�����<�B���Ǟ�ƽ%�%Sӂ��V;���mX�ĕ�;��9�}���M�P��+C�m?<͘�6ˏ��ն��r�:	B���9�3Yg!��6�y_27@�is��F"�%ٰ@Jg_rh/�$菎!��H;�bHƲ�O1hߝ��|T��&P> {��o������/�h�}?��Ĥ���v��C5�)��vyE�A��BX�
��4��oW":m�u=xجu�hJһ���w2��x��9���|���9˚U2���F+�_�@�4�Z$�ܫ���ԏk��Y�>ݟ���p�7�a���y����g8���i-+UMc����R�Ζ�<��q��J��.<��3{��������#wB��Q3��3Kh$��V
"��q~�GUj[Q�+���+�t�l�@נ��;��H�P�Hn ���Inn�4R��L�i6�; 掯��wE��ʱ^��Q�	h�8��k�U�r����V$��ԅ�k
� ��C�kX�"��s����b��ry����ay[>sS5i�0#��+��e���1�Ʒ����p��)�}X���#�l<��"�?��[�h�;-;��hg����n�Y�1�.,��+u]GE��q"��O���$�xb�{${��#Ł�����$�IbO#����{1e����;�Jv-$���}��V��>:���Kq�^���[P��ؿuf��DsM�'�����7�76+��d��6ٷTi �l��2���3ݤ������+#��r����=�� >�S �%���?W�IOb$j��N}z��'�9�Pڍ����<�W��_v�<es��-�=���M#�5��AOϲ
)V�
C�}��F���*���_�k�f����&V��9���!�a���[!.]Ĥ�Gi9�V1%�>&`���YNV�!n�0�C���Ck�[������=�*���o+ď}���	�p����SH�ˢw�t��.�ֶ��H���>��񋭵\�,��O�b~�R��r;��sn��Є��&]�Gn���N:�6��c	�%xLڶ\L7����Q�w��\
2!����#�*4_�b����lGݐ�?����(��I<{g�h���#�[���i����"dL���r>�(�ʗ��͡�\m�O�-���e��H�Ax�:c�2���>�ai�/ˀ~�;���a��ݝ|�΅������;Ə��T���g�A�fd��օ	�U��.��U��G��_���S�|���]�`2�2��|�K6�@�'�G+N.o��(�?O
��P�z[0�c_Ni �fp!�pũ;v����z<���0�8�-Ul�>IR�.2�5�2���k�1�s �k���ڮ���� җ~���GN�ó"iU�\v),0��O��X�rS`�n�5��������j8���5� ���x�r�X̀ � )�@��H�9V������n�����dpŻB���<-�����񦉳J��
�&���'1���|>/)����By>d��cU��1^�>��iq�=|�� ���>��>�e����>(�\�Od��["�����M����W9 �����h�ay�|�m���n�\�J/0`!��*BB���5r2�bTC�TI�\dT�M>=��w5n����<�ѽ:ٝ�%���Y�(�^$R�����s!:�oi�L7���o[��shjsK-�ޓ|�2����cx���������R��28�k����W�J�ͣ��IS6���c��f ���gw�7��Y�����2zH����A�b��%C?K��X���]�]�k���с��Zz|��$�6�ל�j�ʏ�������#⼗`�_!aC��A����`��Zy���/����c���Dxx��֍��7m%��_ /�)wݑt���:�&�D�.=�z� �,m�3m�� �L���Y����(�V�uh$$FXS�����`͵�8�V`�� �Q�M�yùǞ �/�o�Q��_��g�y�R�
�»i�A����]�>c�����-D��``$���m�rAW�S_����D)��QA�9V��7�`�)��>�:	���KA��ÇO.'�v��nQ���0���� 1�Y�+�C�I�����φ���WZx0DJAk5����2��H���!
�!S��Hg�:~�[�
�3�N-��h�6��H���`��Q/�K�9�M�|݄�x��}��O������5���	�-P�S��y�͏"�.^]������V��
��m�ɊEa�� �ǵm�%[�Is�Kh~�LS�� ٗ�`�J���! ���0�x���5)/_���0J���7��ԑ�-�F�4�)����꺍����pq�U`�I-*�p�U�-�(84^q�ю���;�A��F�P�B���>w��cR��=����m��6A5Un�ʌ)rǶ�����6�f�*>��l|2(3bM`�*�p�&妟0�����S�."���T���WHe��5�;z��܁V��G��M��
.��$G�����en�Ÿ ��=��lKh�_ʊ��6*�E,�qQ���3��ǵ�m��'B������R�ъ<E3�s\NMipZhx��@�w���?��{��B�5�U��x�O��M��B!���r�)7}��ј��1N���O�	/��*�+6��6�(���]5�Px�vR
��*;�����D��]U�&e'�
�
ff2��×�!F^�����ꥌ���,4�%�����\ՍD)�������=��cnk��Ufjv�qLzƒ�Xb6�lY�����ɪy���$>h���w��O�9������P�9~axw��E�-O��V����W8=���~�'��9��Y������ʣW= wuO���'���'�-,�&o	��G"f��"�;2&����!i�؍�����1��0�+��_W��d8��I�Y	�z�>���)c8��Ss�ՁJ��t��u�0n����<xQ3c�����pU����`��6##��R��3�7Jr8��a��<]��������>~��|�U�sD��!{��W�8q�Q@���"�>ʵ�^X�,R�x�j�(/�fJ�1��E��J�W�;.\�;�/$7�o�xB=&��s�H��U�ʔ:�ęj{&�S8´|{��O��Xl>|2�8�ʙZw��B4�s�Ps��h�eՇ���"�&�F ����dj�@ޠ��B
:=��%�H�Ȟl��*��_�M��U������3��A9��~�/�q'��#�.�@�}�i�.�X*���d�R��������VO�4SL2ڛ��K�	9�3k�/
q
���<8��̊�2����S��
�e�㨛5.�YC�b5�+zr�6L�G�~��~dvr�����T��Mg��1Nf�B�<�^�Znh��-x~��4 ��7KO
��:T���T�4h(��Q�j"��J�.n=���P^_&Q��P���tl�:�1N��7���Ԟ���C���
�I��mv����#��C���:$"=V'Y3�Cw����(�>����8�B�G�h���e{�UL�1�`)M��35���AS���%��]���U5�ƺR�xd�s��n�N�������0���2��&�;Q��3I@��]I��	m�[)���݋�|kS��)��T�p"�F#�&��(�싗h#+�s�ƪT���*�ٞ���#��6��|'�sd�T�U�����6�H�t�y
���#�|Rj�T���&�{~���ξ ���Z&TՈw<��`ة���Ͽ{��2��u�\�q���Л��x�� .�������0w��|ľ,i����b��xAVL�k~d�;�R$�5�7~�E�=��,#DK�&h�H��i�4���B�Z��c�y,m��|��a���8Zs�Y:]#,�^o.A<��ȓ�< `�)j�q0���:�7wR��*�<*��$w�kcB����	5R���2T��_��!0c���� �C�v��J^<z���?�hr����_OU�\��@�\�����[��"A���B
b2^C�&z�Ҿ�H��%
ó����x�q�,gz�db���ಳ��R�<��]q0���C�S���L���:��#y�-7>�3 �:&�e7SS��%_"�;���IM9[aВ��Y�|$݄�Ԛ�N	��2�h3���BK�[�����Je��G��Z��f/�t����*�n�;3�L}F-��2��r��jJ$�o��顩vŤ��c`������W�s�"��n����4oǬx �B�����K>
��$�Qy9�D;"��`�	 �A�["1�q	�Պ\	d<5kʀbz�U�ƕ�D&���።�z��K��
�{>���{�$���(~�֥˳m������r��
X��l�d��v�h)���2ƃH�\!y,J��x�#�|>xXUÒ��v�2uK�4�CAI�r��]�����`d��7#  /�IFEc��EBw�QB�l��


�`Y�`g(�=ѯ`ay�H�k��p��/����o�hN�>�<.Ip���8�/��L��ž�~:ݞ�mvQ�G��v!�fv���3<_�\�hǮ8��;�<�����[c��O�wm8� �%��z�BN�:Ǘ��h���@��6���ހ�������!��Y�I2��h]�.Ki��?�{;:���,I7D�2	`����r���^'ר�^���H����Y�k�\/L�jG]�MN����)�E�i���os�Rն��z���׷t��oEc�(�m�.D�i���`���;��n�<����OZ[��cK�8�^�A]kҠ�Ŵ�q���I��;[�9�:ۆ�Hŵr��E[/@�z����4D΄��(D]���y=]^��4z�]��c8z�-�-hhaS�V75����5 Iq��#���$�]oX�:�A�#A��+	w�t/�t��K��疤6['��G�?q�@�c�B�r��,_���Z�����zl���+")gk7��[Q�|{f�%\���8�|��$��q�n��ʕ��W+�w�Du�E`j���g]%2�k��ӧR[פ�=]��1
���%���glͻ�j��Q�
���J��Z?�b+��Z�]��:�ďE��� ����V?�7L���z��w���H��,�kBm��LB�����.qh�-��@�6�������*dl�Y%M6���*�(��Z�752�Yk���?�8��趒7����b�4�_XJr����So��?��~WF8[5���aV�/_#V�B�yx/k���a\5�m�����W�R�gеTlv�|>{����>g56�Ys�f5f���
��;�O	c�*�pJ���b�k6��]��'�����'Gw�h?���kP�I����T�%�串���]�}����qἒ�'�C��X\|����	ɶ���D���"S���A������E�Y����p2��{ �+P!V�װ�F4�ܽ��t���q<��uB{���\L�(?N+K?"v=v)qF
C����$�����&$�����	j�lw�zax�O.��;�k���S�:(pr)t�N�`0�l�M��ZJ�h�m��b�ȯ��A��`�t%r�>hg|�X\���K5��]Zx�v|K�#���L[�*��M�r��~�/i|t;U8,��������SB�G�`�$���8&9c�����\ܨEkD~��	_m��i��A�8����27�__cJ��,�j�P
�FX3�{�E���;̥��ѩ�:@��i-r߳�b��lQ���=d��\�a�H�U2H��ʮh��lZ�I+^�����Wn�Y��&�����](=ֈ�������ԧo}�ю���� �����R�AGZa|]��s�,��~%S��
q�a\u�./�Y]m,�'^5f��5����A<���8�6�pT�[-�K��X<���J�D�Ca���bJE�p1�Ÿ{�4[�Ǜ��,�t������j�w�ק9t�¬��2DȲK���
2Sx!�9��ŝ]G�y����GmvF�9��LQ�(X��k�[\S`�Q�z�[�|�-i��_^��e�<kJ¼ܚm���&s
9��GU��|�r	4���$�Ń���_T$^� |�B'2�g������INiOZ������<Y�9�v��vDԘ
/��T�eC"��>c��u����	��'����w�����w��n��K����1��z�	e��N���}��7�$����g'3��x	_q�-��
�n� ��ZZ!M��������w�)����Ͳ=~9�y�N�.�/e��u��G+eܶ�����|z�%�yբ�z��c:<�B�6��tQQ�j�8��t��r�½����E ��9>(��E�i��ƴ4Y(6���ăRIB�i�`t"�0�\�=5ft�-�/[��S�R��{_q�&O���s�,0�ۛ(�F�X�&)���P�Y~�9`{Н'$ �!a�.Y�L�`�&3�$������jQ,��^�B"K�i�[��-:,�iݞR�V2lNt�|Շ0�#<�m+�d�}�u����ؽ�M ���g�`��g�ב���]�+U�[�!tIɰ�#�FP�MZGkN[4K��a��f!B��	��Q㑕Ma�wY����P������y��Lߛ�ﾛ����֊��p0�-��'�@-cY�;���67�U���kR���R����_J�՛�5H"_����d�}�U͢�f��UXkZ�����������#IRPu����o�8��G����2�T�����n;��{����|.LH�sh���<�ۮa�	v�, ��
P��p�/W�t����y/���~��`A���P����!�gp��e$2F�+9'�#ǅ��Flv�	~Л�V� LN�b+J~kg�i��u���3�ɑ����{����k����/Ѵi��+ �#��c]�5Zi�RiO�np���)}���^�0���8V�UVra��*q��I�� �qኳ�}P˱m����a����R�I���&� %U'��g~�C���	��N�vG�؄�\]i�Qy�u#a*�T������X�/��/k=
 
��c%�d��ֵ��ŋ5`S}U���J��؟_,�IR�/g�+��P��;��H�?�*3Ζ�3e��t�|�)DD֞�5G��8$P�麿b5"��}1J�}Dᝎ?�$"#��]rz�#l�g���dKc��R��R���0�i��>* Љ%3~�^3&�?���f�NH6t�D6z��1���Le�g�#J�����֙��7��ݱ�wbaY�C��Y�oM.��3:/U���e�`-^?`b:��������Ē0՝4O.ϪK��Bߡ���n�0t%B]-l�)�� R��];%r$Z���Z*������������"K{]���>��t���j��0 �<9q.l���(C��:���έ��u �|�� �>�X+ր�`��,bJe�N���q'Ă�q�!/|����m�`|�.�Məa�**m&H���{T����8|k���(n���u�����A��=�|A�c>I}�K1�8��Xݽ8����3p��0yv9s�UR�V$d�{���X�Y�;- ����hx�H)�X^4�� ������s���b�k��1���C�6${�>�+2�a>�?{<�Q����I%�/|h= +$
�O�Y���\{U^��֝�xgzU�D� 騴��$0�-�Y��!��«lÖ�F�S�U�Mth@���'A��أ�/��9)�4�z�t=�����Dy�������A�b��CL׼΃J�/��DC��hC���3#v),Ό��u�l:6��\�/����&ܽŮ0(�ڋ�Pͺ����FO^��z##~���'w=)�61yHB�˘/�K�c2�o�>��L�Ǵ�+�O\`я�r�A&�b$�t���B�p1-����dn�O��~�߭r��T�[3��*6:v"#ԭԲ�bmR�*?aϝ`e�oJA��(�n%����}�m/���"��UNz�@Z�
���j�22� ��3+p]B�������Z֏3u�5Ԗp�D�-��}�-Ӧ7�������{+W��Yۀ��t�?����TG=�
7�q��ܔ��n��$��s�+2�)�8E�w����Y2=�wC�3_�L�+� K#D�~��JP�ONf{�\=Ȉ7�K���VB�ٓ��"l�ŗ��P�D�+D"�ۋ��oa�1#xD|��\��Xԑf$���`2�h֓%^�l{&�jR
�i�ٲ$[6�s:齲�@��L�t<U������!"~Ӿ���1��yZ�MVSB�����m\ԁuz�8��r^f	m���9���I��A�-������=�7���IM-S�w�e�Ku�l��H��M�6=o����uG���%|�J��Ayvf���V�'}z�d$��m�Y�a溊��#�a>V��"&��񓍟*�����E�˳6	JFy>#�8d����T4�b���h-#��!�R����n,}Dr#"��n�̖�Ca>��lg���ȅ�U�`p� {l��(�ye�����CJ���d��%�oR�1s����r��o>,�����&�H^�!�q5�0�(�i�H�]a��X��2i��󫰴FE1�V�8��g�%�P�.#�����-�1spG��J4��h����XC���<���<n%��<->�K��JJ�xC�N�땗b�b�(s��8��Jl��8.�]jC�naP�
���F��6�����^X&�0J�c�??���!+��G��A�O�4�����V{<��&))�5��?�-狶<�~���^�����+H?~o�nh'\!5r�Fӥ�(�׈OQ,�^��+q8>����#��q[��k~��퇓�WP��-���k�f+E.�?�vq'�]�g�Bp=�+lm�����h����H񽤤��@�D�_%0�8G�C�{U� �GS�!��@�!A�u��K �p����yH�~^K�J�:e\�*�Q����8�������mŖ}̈ߒU����#Ё�x�~�m��^}�F
� �;�x���_��vC��29��������,(ǰ��L>,�#��]�sK��� ���h���h�ܠ�W���j�&�?b�Dȴ+=����N�W��!�B[�B��a��4NomC`W�|�p
X� �֝kb"�0�4݆'<RX�$��L˃��R���[.�E��+Co'��yN��a�)��.hD�~j�H�W
�8�~�(��܆0+�F/a �	#�[l�)�֋>E_�7�i��4�%HQ��Zը�?������Y�1O{e�����
�����HE�q4ǩ/�PSȂ:ǅN8����Rj��P�H��F�i����K׀dov{*���� P��w�o)+Ge�����cS�����>˸|N��WZd��
��"ZuD-t�{#�ː-�s�OfTi��ꙡx��2�|��/!�P�ޙ�1�Gd˟����z/�Yԋ�8͚vtTu`�i)�S��h� ���?HÂQ�N�Y��Ì^��K�>���{�t��-���Q��]7�<�P�@��*';���t��|B���9��*ϛ,9�3/)�HxL�:������DC�c��{}��]o����]'M i
�9Q�In��[Te���N��畹�xOb��Шщy1�����Ls��fQ�~��8/��P7O~Cs�aB��t����r��]�Pȭp�3�̾�p����4\�D��8���2U�r��@��4�����z/��>I���v���י+x�4�-$0���Ul�������¹�eXxe��25m����:f|�~U�K���;�d���V/�+hN9���$}a�xqz=dv@�$���z���U��Ķ�M���y��w�k���ԏ�˰��=��r��$Ԍ
*��q5y֚]oM��?�$d
@=
��6��h5�`�pb.��%�(�����	�6)[(�����Ӹ�۽�:�چ>4�;
5���>����~����@�a�,+�O����B��7������?�=^�܄�+Ϛ�a�~�4�ѧLC���(�^��ٿ7�oډ�cR���7��&o���el�3��QvL�F�o�e�
/�dI���P'�ˣ��d�	��s/�L�m��;��:VVs����(me�ލEG�W�1��KH�c�h�i�+ �"��4|��pi!��Pr��_caf�=�XO�3^����fg�{t
��F9�;�8�6��W������.�HNnr.r�� �.���9z�p9�c܎��`Y��	 px�q3�h`���L�Ѹ� �#	E?�'.�An0�:��y� �9�!K�4��Sn��H�|��I�uK�J���n����d�^Y�<�`D�i��'�!t�$�vn+�6��� �Pk�	Z�^n��:���A�x���ۀ��Ōl�_�H�=XOˈ�@��x�/�����U�ar��6�6a�,��|ouÞ�����W E A@"�����pl=�|V���Ex�O���2��|b��Z�R��f�fE��H��n g88�2T�T�Z�.(�ˁ�r/����L^{V4'^N���9וRl�y252�O�׳�IB
�_e��ȗ*�Ҡ@��	�)V�'�|�N֮����k��e==�SB$+X���đ�(�'QYN�Q�<�������;��d,���wsς����5])ǀ�3j��������Li߂��빪�s[��43��1ɤ��gㄼ!���"�Ί-L�x��
q���;!H
p:J�9#.̤:�L�[��A��8����fc�1H�6��m��\
},u��c-�'R�U8b��/�c�y¨?)vE��/ԩ�nF�gEi�⼖"O|�G�]l\Τ9I(V��y��.�+�ޙë�����!�5Q�eZ��Dp}���`�/~�*����������̍��g��QXx���O���o�K����_?��Rg{��XQy��T@@��!cߏ_�h;�G��u�b��!	�a����\<���$�'8�r�$#s��
%��OZӼpܭY�kg�:*�U�$ i�~%XSF"�2�C�@��Cd2��d�&��#W��o&�"�6l����m%���>Ď�{���b���T/��	�c��؜�Զ�������`~s�R\�h���� �s�t`�Bւ����e��ݚ��O�!%2'���8p/t*�&�p||X������t�٘;d�J��?31]����C�݅F�X�V�����C0���: �F ��V�(�x�� [쀣Y,�����;���3��F�W�� ve�5�a�_��uv��For�[�+�����Av��7�O8��I�A+[�J[�ZO	��� ��J�L ztP໐?i���m �o����wu�/ʁ���Y�W�cDr.�^�7hYVV����E��cc�ߩ�G�\�����F5�B�א��p9�j66��}�]TGH�%������~�_摸���#��ؤ��t���Iۤ�#6Z!Du����25|h��y�Qs�0��^:C�q��� ��`w6�h�؟Է�L�����@<��	}MҽR.�v�B5.���w��]��S�V�N��3ф�@����;Ӵ*�B�����Bk9Q��k�	��1��DV[C~�qN�:�ME��Z������U�e*����T7�Tal �>�Ed�\����.r4��Vu�e[�l�!���ն�1NBΎ��D�1�M�JS�?�����h�/v�T������ ���&T�v�#�y�W=��l^��bn��3����^��Ni��D* dÒbz�VQ}�Y���[�]�ORn�XV�t[�yi�ϊd��g� ���2�3��|z6dF��?Q99/��;���4��_�(p�����9Ce���gky��N5���ja �c�rre����~PR;�N�i�U��E3��1��N�"7��itU XQ�j�iS��iZg��v<��	��Ee˱L��/$��l�xd+A�:���m��x�;c���]uۘG]�H�;����Xv��5EAf��y�5��WM`��[w�GIAG���|d�*�y��mD�FAv��:��� C�@;[�[X��͓��m)�36`�v*�s�x?�]G�5y9�Q(�n � ��8v��t���>;��Bm[�j�ME��(7��ܬA�&`o7���qUyE� ��t$��_2���/��6�3�g�B�(v����#Loa,���>�K.�G ��酛Cw
L�xA���T�քn���-����q
m����ꙫD��|�W�˹2�
����*��M��j�g�eP�e�ٮ��)`i���̚Eߧ�m4+ýLB�36�����"���>w�V���=6���9�X��c�PhV���+��0�W�����oϲQ���Xf�����?4s����\5%;!�x��irwB�����:�m���v�«�r�!�G�.���7�ZA֝��%���x�(���[��P�'��������uH������ml���3NL���r�Nua����8&�NK�1�G���&�U ��KeaѸT	�|46{ӎ��P��@�$��8��^�'�����L����X��N��~�B�?�w�ëG�L�$Sb��%+�qJR�A�udP�Eh:���u���D�h ,"���I�'��^�R��6{�U.����D}����h"k�1�3�$c�D�;0?�,�|6.
&g�l�2���j�6�Eh���XG�t��R�M*X��tCȼB
�ҝNg���{8�p�	s�G+�@��G�\���ٗ/M*�����3�?����0������s����FdA�2�VH��9��ܓ̞ߙ�q#)�|R!mU��ܔ�V����>��/ E�A�<*�Y��#���Y�NqkfbW !�5�l����*�@b� ��;(�������ptyDV{�z/4�����9���iZ�ؾ8o���Ǭ�}��]���qA2�ya��C���"3����+��6�b@y0ҘT���<A0�@�Kp�V l�&ӳ4���Y�p)��yZ��V\�~� �V�F*ꁙ����'-At�[�:4�����s��j�N >�a��q��Z��mSP�v^���<���
�M��(L������~�F�?�m����2��MȤ[I	2\���	|��a��AlZ˟�\E�zF���hs5Ɵ#�?��,v�k\��\Tʤq��l��9��Q�Ư�I���a@��S-��`�g����i��9H���H�O�k�1^���C%m��SQ���0y j��Ym9���KD=ؠң,E7/fnH���{;q':�BfӀ�J���Uؒ�).�R_��LD�oKz���'�О%��lQ��X;��W��j����%l����.�݀��>&�%vwt��jH�^h2�jPL}U� T�9�ʢ��b[��mdGD@R�[�0 �Q��Nr�����1g�Rj�|�.ax�L��M֊n�P����1��׬ ����t��o9��Ï���A��0�{�G��25��hz�,T�[����<Ψ6j'y�>���n��[��I3��@�6�g� ���?�w����:�A7�����'VU�p�7M"�����"������B������r��v].���ߩ;sxy�� ��%=;HWV���y��Էn��^]�$VT�Y�w�pK̒�<��-�K0*�R�Z�r���HO�,Pfz��!��"9�Y���)Gc�v����<�-�_aX��ӫ��Y�v�y"���,{�c�O������X#�D��s9�Q$�[<j���� H�GhZ���U�U$��/�Dq.���1����2�d@�������LN���X�Jrns�'���l�;?����{�@쪝��-��bGŇ?e�VP�&�����s�h:�뙡��q^*��Jf�8u��/	�4q$����ΙD� 9#�x���D��D.�M�xȊ#�;
hX�h�P=3��R�M���N��I��4�>C̚�٩�d/�)� ����<u�1G��x��yM:��no�Z<�����X4����t
����J/츃�� _�J%%�l�6���M<�wSx�e�g�Ҩ�J^�%��XQ���ߊ&.�m�R�+��)�f��<'�н��~��M��r��1�_�s���fT�02<��X��i˱����`��8Uq����Nݫ�����4�zN��2iAٔB^Q���Y�a`\��e�W)�����/��@���RTm� ���<�X�r������:�	��f�T�+�ٜ	pޭ�:$��6��h$��
(� �w�|�Ҫ#��^��Z�@�b�|.92���Y$m�
A7����&��0BuH��FHl�� �����L�y֢�(�2�A6U|���P� 6���B���8��
�|��.�\��M+~�s@��^�bJП�#�Y��y"sC�C�^�(�PV��ə���O�~c�<����zi�fb��E�OϷ���f�!�cG�^6}/" qW�]w�J�"��oG��]>OM2:IT4n���9���I�)g�����(�"닮a%����i$�A�`~��}9���	�k1.s�=cv�u�bƮa;{<�� @̲*W�*�Rd�D�а����6[���Lo��p�6wcuq�VG�J]�_��hұ�a 7G�(��yx�f��>c�T�:���uh��w�����gn)g�����w�y}y'JBz��o�C����!��ׅ�=�7���T~5D(������n�<���fpv�v��؍��O����^ʅ2Ir���Tc�o:�9P�ֽ�c6�RY���z%I�I�F�?s|�>�c-V�E�O^�"ń֚N�c��]�J��ڒ>'ZbOc���p��+���,ƎS�h@5���c�������)0$�,�"�H�b^[�5��<�wQ��l���<4����[�o��xV�g��F�S�S����LOW�m"j��kOK�B��<^_���N���������>rjȝ��R{��[ƪ��P���/xc�t3������d�H���+`�x.x9�$��$ə��'���[�w�+Z����%l��yLw�h�.��(�-��3�a�)J�b�If�g����3/��s,p]A0bf=�����#P�*I��H��
E���e�B5�jx�n(%���Q�E@s�����F���vo���&�6�b��$�����Ih�.E8:�FS~%n;S�J�yTL�:���Y۞-�>+q9�-3Tp�o.�C�ѥ�s, cbPV(S?�Z�.lZ�^6~��F�Ci�}v��)Ʊ�1e�F�����ܱՄY���3[�[��ŵ9aB��@��Z��.|h�1H\��:�O:448��j�)f� Zs�{��M3�����~�S�oQ�C�jd�wqo\"��Lc�Ƣ1mac�~�$��u���wT���|��.Fe�R|]u
?Q�����,��U��Z��]�WU4W,ǵ}���}�/��hQ�^#�(���PM)%:�t�
�Lz��p�I�~j<�f��^�ITM ±��ZAlc�.�<z���}�>>ׂ"��V
�
6�ĬW(�ϓ��^q�hu`�L.WS��
-�S�]��^H~�p���h���4�c�Q�g�;G!� �l�����)R@�7Ԙ����x�����X��+|�C��p�=��J^��r4�7kFVB�J3��CO-��g�W��*x]z�����)?���@��^�a4FS�T�I4��}�z8,��q �xH�����W�5r#5�}U Ýd����Y��2ɪ}� ���(�Gh����{<[��F� u��@��[�x��U=B��w��[x�x){�����|�`���L���X���_������ʀ<�	�	kh��u���gW��u������Lx��@�}%�Q�������`��-��!�ݭ�Ji�^��l7� ��um+;�\4�;vK��'A�gs�+���٠�%mɏ��B�H�;h�=��Y���K4?/*W	�N����.�][h[䂲&�� ��цI���M`3������P�6�kZդ�\�C򖋸(\�(���FG�#$�s��ՙ����VL0]�;`�4����m����Z�I�^_8�CD���os�wߺ�B#���a��D_��L�����[�:���o]���eÆZ��SW�w�N����{B!x����9���r]ɻ��U�� BrJ�n���j�*ނ��(��)��@؂4b}�ĽZ������J�j�'�p�@����r\���i�"��Xjrda��6FO�~�LCR6���bޘ�s��ݢ!�ӯ�0�"���@ ��'Pc�U]	���G�Ȟ��-͇�S�O�)����mrWԽ�':�i��Bo����۹�9�ld؉oGs'G-=e������2���?������)�9pz-�#���=8Tq@BX֬��.dݽ\x��2~g�p�$:DU�[:"&�krV?M���c%cF=�ǝ���Ĕ��¾@��0uX_������O�k2��ՏP���o!�]X��j���#�.;�N���luŧ7����Ƿ��"���i!��
���F�H3>�X��h�9g����G[�	6�٪Y�)E�Rs�4b����XF�Pʾn�� �.�Y�^t6/�d�r��546�zs��XE�'�@�H�6��I�ը�h�>�}@`.,�{��<�:L�چ�6a�r@st�7Q�[X�t��QҰd�R©-T��K��[\�{֫+��^N�y  4��Du�[���dJ��' F��r&���0��\8z�aW�����G������s�		Y.S(���i�R�64����0bbKmO�[1�����Mm)L����4a3͊:��B�~�:þw59�,|Ɔ()����� �����)!<�zvn�/�:zך�D�u7�L�g�*�_Q����VkMɌU(��]�dUq�՜k��E����7��<�5,��%�~Ѕ5�B��ctn��]����N�!qt�6��)t�"�V�������n�+��<���Rr�E�f��n�n^�ңխV���i���0�Y�c�ʑt_p����d %���7��!ݞB����S�R�n%&x��᎖%���k ���:����X�x}D/D��-��E%^�$Y�$�s��;�@��t��T]�ĐYʯ�H����:��j��YG}.��1�][�0�G	��-#:-����[p�ʄ9)��U��y�y#`��~lI#& ��K���1����=Ȱ#�����4nh;�.mU�=),�=�&|���L��*�a���*�02jX���E����S�7I��m��tX�@l_�}�WL�-@���֮�����) R��Fd_ѯϩd�J��z �%;<�ᓰ��|b��NVmj%
���Kq�Ѣ�e�sNm�1�!z���,��?���v�{�7���5D��e�6���p�����wh|��z�y�.g^��"Z�>��<���|��v�n\������w>d���t��^�$@�K���Х%��Q]gR�N���I(������m
ʬ
̖�k��KD+U�4��A����Of�������]ʿ��Eo42Y���']���5�~�����h��E�&��^����\����Ȯ�ߖ&�@q6��7뒑�*��,���@x
,6z	w~�)�p��7]�5�9A��[}� ��j���r���H%J�
E�哛\��wt~@O=�J�hyʊ�i)��iZv���6ؚ�����$c%@�'�Вm�?ߣ`Ti��|�p�D�v�`ZkW�g��l�V�T��1�E �8I�#Ǫ��cg&��ǵF�Nǂ�|^��d�}?�7lȅl]c<�60����q{Atk�ی�ʩ��d-UQ�=NH���
��ZǓ�����d�G�ذ�6o����Ω/�+��ⳳ��d����/��{?�i.��^>�lL�cs�������֯�	.Ĵ�uŞl��10�r���z��w�{�̣dJxқgs4��a?\U��*�;�]�{��9 j��7�;]&�fbj�� ����\<Q�+�[��7j�%f��ƨRr23��^�"�z��&�B����ҭe9H�V�=�Y�:-@�攕�K�� �fr�S���*��lc5�e� ��Ni��jD���H���ke�Ж�[<7l/����(A��ܸro�Y��,�<9�[�2��˹�JS�b'��Ŝ�ĥ��t�W��XvV�B�x�1�̌Q�N��	ódY3�L��[�'W{<	�H��]uJy��_�˝ZlkǇ�Е�@͟:�`��]O��F7Xz�r�y��8�)F�QN�eܛ޶�[�g�H� )�Ԛ�衸���+�����u��$��/�L�y"������ޅ&�����}�����~��h׺�9��r�*�(x�#4R\f��n���c�r�qY�%C�������KTH�����,�Ɖ�_���Q�4'�g�0������}�P�����7�G�z����nbz�,ǛA\ ͚V^�G�����.�+"�x�o2� ��C�z@����B�q����Єͬ�e�,�Q�]�ڸ=�$p]�\�������1|�Wrr�:�`x"I���o���NPJ����F�q8:�A"�DWP�,O�g����pl�X�a�{L�<-�}G�i�7�:_�;�ވ��,U���C���~������w}�6H�V��(LV��&�~���d2H�����OQ�7�*�N�[l�=���H��.��pm�.�!��<@5P#��=��z���i��M��rF�v/d1��࿜���Vd4*�{{!#�{�30B�~���3�b��F`��4&{��w��*	���͎��1Jk@29Z�#X
Z�ڷ�����,�s
noI��MuT�J�%�
�`А���Ҡ�tVz��=�V�{�n�չ�WO2@��K8���c@������6�q�ŀ� �����N+GŤm�(
X&��#Pɿ��Q��ٻ�Dܓ�"�鶂��
ڦ�N�D��87y����P�v�w9C[��|�D�&-�O³P�ǜ��������
f�ZH�ԍ �=��u�u(���9i!�Q��AWo�R��_PRı �� ]�'ISBFM����pr�1l�(�s:�=I�Vu��&�UfS��q�%��>���P�O=��Oʜ�f$.7�Yf��Wݡ:J��R��]y��*������	QP��k_�� �>�X&���2�d���1�0O��hJQ4�lČL�rf�Rg�Z����Z��'��h��Dr��6P��.��u�x��"'%�K�����P����D Y�g%�N�[ �U@1'4�Oӭz���V�d�J>$V��"X���<��rd�꣋\6}��Le�B&h;�'�[:pa�F�����9�Ѡ�(�1�`w�wg�`������� �J�����d5]LP���nđ�j�� �{n��S������ǉ����C{n��\��w6�';��|Km�,��x&��ShD��qzsׂ%��_d1P͝�13�0��1#�c�	��� ���n�dS�W��1O]����۹�|��iu��^�0-��zt�k#��J��m����=0'�iy�Y����n��-�P's�-��R�T�%?�_�B�ggkm��^���~2&��X�W&tl��
1��Ҟ���@ ��~������-�y!43�|6YV�Nd�����6���Z�2���1[�âk �;�A��[�"�ī>	@Bl_��qÙ�C=J��B;jYLMJ^\����e�	'���)Y���	��x�P0/�G���$0t/Vru��6j�p��#����Q-`TrH�:0�x\�e�d}+�?�P55}��l��S�C[�v�ܿQ��y[f?(�����Ԑ���5gbeMěh�h�_[��|�d>�.���d{�gѲ��m;J�x1��}����4js�*w&�D����-*3�i�Dͪ���-��)K�r�_�u�;��WI���O�cG�V��Y �b�
��>��V�K���=�Z�{H[z8a�a�G�c8`"oY�쬪��ϟ�ő�\��F\��)���}} _�F�s�B^��/#�M;X}�`lu/�88�pG9x�$ds�߼����VJ;�
+\m�/�aM@���7'���0�)��@�():@ m>��gݖ4~�A��`��
��گL�v2JWP��8��;5���Fz*���gP���ӠrB{�����A�#�?;��KNAj��q�˽��$?�Y��2�ƚ�|<�_��`-��"b�n|R���l�>^�߮!{x˩�S����RX��^�f�=F�#�pƌncn��N�r�m�D�"r���fk�_����=9��E�ܹ�n&XN���غ�����2�#�4�f�"-R���c�v�j�z'!W�V(<�f��VY�{T��Ž��g-҄������\
0USp[�U8�]�#��t���'^<���[L|��ග�v"�Ӕ�~Y!` �7�z*q��r��j�vxw6�b�s����0�ZJ������W�`�3�ip��X8N��W:A��i]~:rc�r-��ݾ�n�&u��c����������	w�4��;@������@1��`I�z�r`y�R�Je,�QmmW�ތX"�
�T���#{���PMJ����Tch�O毋(���_4ķ��㎫���7�ȹ�(=_�||,e���b�s�E�6�eP�8���	�1-��(]�[�#�g���&I+��0��	���u��{|�4��2�:���QI�8��f��9<��w_�х>�!���B����mG���."���)�5�]�ծœm�Ϭ�b��ԓ敉� ������Y�	���<�e0�D��vL����ddC���Gd(\���j�R��B�N�uZ�~�b��*���c���og��)����Jb-o"���T�h	�xH����jHX�_1N����%�����Oŗ�+鬲>����R��A�z�Rƻ�	����XdƼ�3�i
��Қ5 P�L$V�3ԓ�?�q�k�W��G:]*֫���_�0�?�% �g���hԶ@�ps�4�0��!7��*�	�>�\�;�޲��h�\ւkTN�����ڂEm�k#YZx�ޔ�
�e�����PW�	�>�aF�ܴU�`�=�T���+/�>D=�4�4�5�+s=j��,�3=�8�Y���J`�۷ߟB�Z�xS��$�ΞN��J�A�K����*$(E0Q.	wQض�����*-
$e���n����������ؒQ}���l_4n]Y��$���m�2��ׅ-��&B��Џ�N8�����+16"�f���)�qeL�m���2Kݷ��7��-�b�~��t�(�nM#Ϟ���"��0]\��K�cdIx~��փ�gʓ)p%v�B��R�<�~�v!+؜N]Z��#9HN�؀��ՠ��I�	Er��T��z_`��7��?��O�ȝ���%ۖ���c���j<s5�� �qA?o���P�8m����Cj�a�iy<��bb�/0	�9��s	�F�����ɩZ�k����"�sF�\εռ�M����U]ſ1�Pr�a����}�V_&E�������������I����A��l4n����s|�seWF<n#��E�g#m٨ȞUT�!p��Զ�ݨux1��ܴ��@l��K��y�ܡ*:'wP>io�DirrU���3[{i����-n�5^�A����L�ufM�#��q�t�]4��5S���-�Ig�v��� S����G#��N��߱���NƸ��_KLDnCR>�����"�]��-J5<x} ���,0��,��ՐC��J�3���5�O�]1��&��w���-�9���b��N�t�����ےٳ,�L��䞔���[�m��e�n^�LU��\�:A��y�s��.�a��#��d��!G�.y��7@������OȈ�/r���R^���~�6��l@c(�/�[��W-S-���..�g��Pjq�hiB9"�~T��ý��ư���
PB�J�[!�h/p��s\K5�����`/�3?.U$%PN��7�P�m+g��)�N�'��ID�K%���w�~�:{�+ړ�:��C�8>��Feۊ&&2�瑂@`F5�������'�*�$Ӝ�
���G�N���;.Bi܉��!W����"�yVgD���������V���M�DU���������Ly�<�N�L/x~zc�'|��}E��UE�O�q�#�ɵ���\�]Ω��M'��w���g�XL0O"z�<��@q�,YJ�i�dCwVE��y�>��%���B:�e,��ZsRA�@Y\
�2�$N+��f�D,���}�*>��D��e����S���ϑ�t��'?�S�M�h�q7ɼʍ��7O����{�-�T͸�)і�y�+���vй,�@���?^�Ym�>�g��V�@���{�_�ߙP���uxnq�*O��gi#�E��b)���rn���U��]n���Q��7ZˍuF���՜�!���z^Ej>���[a'�B��ڧ��%H�y���N��8�V��c����?�^=�>��VX�A�R��Y��Aـ�~�w������	h	�3}����l����6W5� �=��?Qt妎�Q��*x�3��$��w��<���z��hvӮW�@Mc���"����ݗ���s�gۍ�
�Q�S�8CJK�]��BmS��~UR:�8L���Er��T)|΀�ɂӅ��m��<������S4�օx���~i��"��P���V������]��K@��^ <{&���zY�#H}r����-��� Db�V\��˨�������K�7����0$M�����S�Р�W׶��M�����>�WB�-J�T������R#1�&��Í�i`�<�l��V�w)��#����;�i���m��'Kl���iHx2�B[�Nћ�m�.`i�z~�|.k���#��w�,R*6T�&T��%��O�ݡu�O�1]��_)��[;��I�iϵ��3*�nyaZ6i��B��lc��!d��) �e��o<DXX���4d��rg��@n��W�|�H�lo��w@s���/u��~�F󏁴'�5�7��
D=3pDM%>��$݀���0��*�0.X4�!�x��ޕ�jq�e����z�fw�~��{���_ƛ���7��k�݆
��P�u~%_�����b�ֳ�ʄ��[��=:��-�m2P,�������"��A�A��e7�l��	�Lx���������yF�V2��=w�4N~w,�}��Ԯ�k�[��qGM�B�l4y+)���Z�����|o4*	�����HAk�gm�M��D`	����7E岒�-�ޕ4���P��w�|��>��2Q��ͨ�=���D�a��pl}\}�g}��I�E��;)�i��h���h=�%�R���ڶ�f�i��,x\ͷih�2�z�0ʠ� �LJh'�r�^�Z�e�K������%�m���5��ˑ�˹��'���4˭�N��q�N�@Ol8�n6<H��-05������!���%��z"Ds�¼EF�d' �p	v���g��i�����@g���b��]��>�KcM��);Ǽ��Yρ;~r�T�/� �8���x6:�H:�R�o38���������&�K���ŉT�`�&85��K��ϔm�iedhE�<B�p��f�p�	/f�ϴ�eAE{+2�_�/��ڠݓ_F��^�w��� (��5����q]���`tpՙ��;�Kq�|mv�d�������5���P����?�	.�?�aw@P��o�J��1��g�m�H���R�ߺ����(�d�.)+���~	���yW~[�s\�a��P3��4l�D ��@���NhM���tN��{�]�ǖ��9�u�B���q�6���j���v<�/�E������h�7~�4Y�~$�������"6�mP�9O���F1�q�N���Рf������T����b�Z����m�����6�� h��eXh�|�`�%��.ė"|�����;���S�0x 15�����{�x��������eh0ھ=�	�χG��I9�����O��H�j��I�����,��/N-���;
��$�f�N�bE�$���
F�� WG6�3�M�i���6B��Y*��fn��?7?��R�r\���@�±�v M�G\{B�$c�l]L�BsLj�$�;A���7l�|E\�V�j��:�!<z�W��ў�r)��.>�@�i�E���UY���Z�w����2^�k^���K��L��x�Z��A�HVKQ�[����?_��S�e�F�{���\/��Bo�⩁%b��F�/l5���u����*�si4�����9Ԅ���4BD��Yk�y9?q��D|7�P�_&�y���Y��I������M�������̄��N]����p>�v1M�T�.��󻦽	���A=£�U]��+
�Z�HAK���	7iӷU$_p�4��vT/�J��9��0��~�|��·fJֺ�r"%�R��"�Q.��l�F���6t�:��*;��6�;oYK�t�s(}d�z$��՗6�S8��r�V�@�ox��S4h�+���R��MbɲR�mNN�K���n���H�g��{yq�3�0�8�O7��䂿�zz/-z���m��}<-���7#�v����t�N\��)�ՏHx�Udo�ޏ�5�Z1bm-�ޗ�Oʠ9�VQ�'o����{7��Li.NV?�0}��0�bzwQؠ�d��X|�T��,%�>܉��hf׿�����F�=yu$�mL9�r�Ň��0Qʎߘ�re�.�PSC
�B��-�z���:a��Dtb#����@D�������6Rv`v� ���Y�$��n9l��sAMő���4���I*
��p��.w��!D��7�W����۲��2oG�K��[K�t��6�1�9N �㢚��ݪ�,�b=⿪Hj!��Q�t��s&-���q��Y4RGVى���[^��u�d�I��>C��O��<h߲��o��x��!n����뱓t�o�0�ȆJ)S]�$VW'r�P��uq�?K�u��>����m�]|ƹ	4=q���9��z�k(Y��8I'er��0�>�BoI�j���&���&,�5u�{u�?�	�}1}��A��A䙝Q}V��C`5��Q�?�c�f�#K�� r>�� o%?���oS��@z�OC"_�,���_G��\��`D��I��֏����KЂxg�m�������^���!�ӏX�.\�aY�,%�$�_<�k���@�jɲ�Z6R�Ļ}:�r��(����-���:k���T2�ș/�s����ÎJ|M�T;��Ԏ��������dS��h����~�uRc�6�(n82;WmK�Q4�ͨ3S$7��E�t�C�W�Y_/�k�UoR���0��'�+�����xd�*�X��Ρ�8'�J��E�\��r�J���2T͗'*��2��
e��̡Dk�K�S�`���3ˆ%)�_�#�&�EMW4"Ԭk�^YXE�>9�"�bz�	�� z����"d��!2�j�ۭ�[A�,������Y=�;{-���37|Țݥ���X<l�D{��t�pQ�z�2 �ƇʿX_#���������=�Ã}�t��}\�6Pº�?3�Tv�~��y&~�n��]A��ĕB�C(3@���n�{Wd�N����fW
�3[��3u��\����m�{��u�i��'�A��<;
�b�P��@HHG�A����Apy�..�K.Ck$����n�Q�"�����z�s^�G�+<�a.3+_Ҵ�1dy7���X��Cz�d���e+dq�!�i���Tj{0J 	��Ke#G��\�K��C*�C��'Mԉ/L'�4��D���^�pw1+U�ZL}%*��ad��E7��h$����?��HI�j�&ת	�P���R��~"~�|,�]�Yv�~|%`{��!x
yơK7Km��s�9��W����,Bc���r� �ӛ�����'-�V�#��H^��ez�nI�ΩN ��b�Us+U��Qig��wd���+�(��lZ=�8���V�G�b�����nOG饬OH BNӋ��-X�����8���-�Z�<��J��0�5��bڈ��5���e�i��)x�a��s�#����<G�E���e�1cD
dH����%8Np^!�b�#���!�5���)F���݆��<����)�H����0ȍ���t�/��K��T	���;�;xN�z���(/����Q1?�Љ���}����8��E�:O�Q�u�/M(����TG��_m\��ԜY�-+ǰ�&�����l���w�d	���ATӅ/F�ftܸ���S"p���z�KxDu�CA�v����s���B����������(-��R"�R� �[��3�e9�؀"����3c��4g)��?�!�c��N�i���[�G ��I���|�S�Xg;�(N(`p��5XX���/�g�g�	{�j�������B7�ן�@t�Q�%g9w�������h���j�W������}�'�:��\s\>(�H���%��y�����:MX��yь��啛}?:���q|��P|AY�>�0��D�Ne:juo&�|x� -1�pY�x�ל����V1?��o�A<k��c�x<S>-3�o�W�<�,�Z~��E���)ߘ��cz���v���?��l�jO�r�M���S�A���l*�mݞ�;��z��M�[�)RL�;p|�C��F>+�,y�b6|��tS�	G!��Xm���Ү|1�s\�����
��������ƒ<�sG��wO�!�~1�+{2*OC<n�ӥ�vdu���Y����+�X[���2V��Q$�o������ \���Y�W^�.A��_�:̗�$��4��,i.�p#)m��OJ9�ܴ@�>	�(E�ËH|�i���v^x��)��q4�Di�/g���޴�ZV4�nr��g��|8���jy�)|�f����]����(]	64y�sZ�U�f�a1n'Nb�7�@��I���B��_0D�Eѫ�e���7H�բ!*�]%.^Rn+��cSe�Z�{?@�A68��>i����δ�U��,����Ș�^R����0c$�c����$w��٘^���_J�0#��$sx����0w>���å�+1Swb6zC$�=�g�,�����tq��]�S�uY��<��8o�E8����["���o��d)ix�4����k�G�� ��66T�'�B����x�(����6�N@�wؗ@�{�{�kQ���lY��);\z�ȷ�⟣lJ���Tz+e#-���EA��f=`˧���ㆾ����vܲ��亥Q��9�2)H��-��<s��6�)�^�"xEOCa��J�&q*�^�����t�O2X@������_(�ǅ��I�m:i�%g �5IX��W�������̎���Z��Λ�a��1C�2֌�t3&��9r嬗{�}�ƕ��F���Rt������lL�\>�o��7�4<�5�����Z�";#>�ᥡ6﻿�ܕ�T���3��&��U�CM�xm���0�q.�'~-��nXR�9� f �́�BWB�<������6�f�np7	fÆF*��2�����pp9�0F�F�N��U��s@��Zf�c�+_7*V�������4�l���|6�I���ѧ�v�3yqvr �c�ɓW$=���2h�2�J��+�_B���?(�0�zT�Y!Rۀn�-S��-��w�����zB�����Z�6�� &�pŧ)5�Q�}�Ui+��V�/�(�p.ܒ��g�W��bR�*��N1v��^n����P}�M�����'��S�ďWG�k��s���E�u�_Ze/x7i>	���_gPN��\<&�!V��a��h�(�Z��e�aV#Sb�����o���;����"K55J���������kԓ���i�
Ш���Ow�&�Z�-�SqE��6{���|�*��I���0��F����g �с�;����ʸ�i�c����/��lK\�W�p��p�|LD?�dg�{�*���J��cg	��g��)M �М�@��>��C�s'?U��Eoft+��B��)��J
�.�c���c������F����ȱ�p$�+�|,��FC����Z��e�8��S]C{3J��M�C�k"u���s,����i9�˂.��<�����*�IB*�6����[D���~=�W��e��l���I�ܛ��Nb
��"���)������ʍ���F%K:����z��^��g���Փ߾������ǽY8��bz���NH���y�St�f�u�}b����O���h|��D&��|�-7VżR0��a�.�I�~�B>'�I�:g�k�-�F�_�&�|u�E�A�Ĉ_��0�my�[郊����Y.������zll��"r\�جfS�C<z��^uH�ľd*�8��`_H��Q
�Ƈ��%/N��]̴O�$<�H���4#=~<��j���׸�)��f;W��\ި���L�g�!�Pot�l��H���+���ا9ɝ�"�F#�l��P�d`P2��WS:��v9I�sj�?i�xgG��J��&��b�сc����i��1I�J�֊Mn�\�H�"md�FQ0�F^#�/�eb�����\���D*m9)8S�0r��|��q�������)�Q%���[X����ʛ����F�Y��L���@��Z�_9?v�,�����'cY��+���j�+���ܕ.0m��)o���ب����Av^r�tZs���d���>#'�E�5�gi��Ee]�Ԧ��$���b$���^��QɊ�V@Gx�6����Ӯ�(���;lpr��S������8��x�\	gqrnݼ,�56��I�:�����Ag�<+0��(�[��Z1�7��ۧp�~0O�B��U���¦�U˨e�i��'�͵i�_�\��U��XbE�gv=g��i+%E��.��R�y�KU��P�Q�B6~�#���r�~Y�63��afd�����{��h *��T�+�Ǩ$�9�u\z'?�������e,�2��GM"���t�&�A��28���U�=����t�:�ZFU����ј��ˬ�&�<Z�0��JF^��9�r�u���ҫ���H��:�e�2�m1k5��=żF���4���-���@�S�����Z��%��+p��uA!�D�T�>�qn����"J���q|ן� �L�CV<Dz��g�iH����j\����ǂ�y Yf0�V��!��+(�@.��b�ݳRS�޹�����ˣ�d�*�)�C�,����*��n~"0b	�"��dI��\�a��_:X���K�Bi��W��l�&X_J��CCe�[I�A2��ϝ�����-0V�#*����<>6/�~������9hyu$�+���,do��h�Q�n��9��Q��I��\�G�3q�R��"3#+�U:�`h����W0��h78?�>���NL��i%��䊾�1������IQ�;���\�})���d0d,��E^��{`��ϸJmuH�)�7�
R��
����zy�Ck�dn��
u"��]^��?�`uޙn�0�
(�iXrʼ��T15M��2�2ڈ"LC����gBb�.]@���C�S�
	����/dP]�}m�~��W��I�~�iO⏃���8W?+nb�y�qa�<���nSz������\B�dp1䏘��j�!�(M����x� l��
���1��6-p�F�N���r9�*�t��e��>�+�7��D \l������+ߜ?�:��"���CR��ZI�Ԩl�ێ#���ˣ*����m� �XV�`������ou�~�����q��L��zǼ!� ζ(�6lcޜ#ʏ�p�F)����Nҽ_tͣ�E���1�b^��3=.S~ۋ�߁�Y˿��� �f����F�?U�Љ�◜k~6BN!�a���o�k
�Z�n�o2)�xEe����A��9Kœ�n�FB��p1L�EpC0_����>�|QhS+���Ӌd:�?���q8���SKɄMy{BW��C�qaYQ�V�v�3N��%��pD��t�W,eP
��`�u<���Q�R{�y�1C��z���Π�ލ�GT%�i�2�GR*xj9�3��
U�ݤ,Y�'1��P�{��ꂁP��kހ������p�5�=����|M�)��o�%��ݤ�w��|����K,L$8���.�
ԉ������+U
f�(Ә�������&� Y�zx)0Xo�b�D'���N��c�T*�C�[&�t%����G������Elrf����ɟ���LՀ��Z��Y��ͣ	�L����7��k3NG����j�,=�:���ym��eoժW��_$'���J ���!1�1a��2Q���^BxZ}O���{���e9ao��St"z��������/E�0�b�/L���7��<I��}���-ƻ���	��K.����D���XX"��>~�`{�ߛs����=<�V�������&�5�w�~��n���<ȸ�^��B�@C� `�T,�r�]~Q��F��VED�U�e��b���wfN���l~(�"}H>�K�����<�\��Ʌ�Λ܆�|?lu�����2�o2Z�NR�3���Nت�	hjdٱdN �f����L$dT;��w g]:�߄���)r��5�S��~e;5�>�����D��n���a�������o�0��6Ff����D�Y��b�a"gvʗ�FO~���[w붣1m�K�*�x�(�*���+j����zޚ��}N.h_F���]�^��TkԂzvH�b�B�; �Lc8w���2;?ڐ�+l�J���;�#^���Y����I�L��}�'��]�P\�<�_�iO(5΀3��P>���O���з�u�4�2U7�P(c��~I8�y�٦� �"��ZP�x�Hw:O)��Q�Gy z�m�Z]�[�m���f�����&�i�%�ÑV�h0.�DpXs���zTH�4E��"^�F!Q_nh ����Us���k�vc���V��oQ}��^�ղZ1�1���ƴM�(U��i�^�f��ߑi��2b����a���������]7.�H)��u.��h{/b�d�iǔ4�Q���Qw�]C�[G.#w��ěp���"6�r���ː�����m�8c9Q_a;wMD���LSߍ �U��w�N�.p�Yi���p��fG����EH���&Yr��|y+�3Z��F	^�Θ�<p7{Nm�#X3��/,��y#sg|՝�=�qh�F��n(���n푠���c�ď�;�1��fF������ʅ����&�!�݅�
6q?ֈ�k���O�@��U%��T���E�]$�����e|>����X�ȍ'�,��]yh�v�5�5����ǈ�-~�[Cl"��\mXv8�uG�Y�#UYz.�M��UVܾeBy2��?&�S��Bdv�p�8�/14	hK�P`��FP	L��9Ta�[$T�^ ����EU��Y�$B �bi�ȠFvkB�M�8 ǎ]��嶧��=��&��^����YF}��Jź���*v���p�X��mXST�aǓ����W�Ġ�l�u��v��z�y�L)����n��*�Ár\�2�'�}65�6_}0o��Ƣ�B�^#Z�å��JؾuLsS5SR��+`" ��<��T �FJ�
?1�9,������R�`�=M��|�; 	O�R�s0)��w}'$x,�W,owB���.��������0z�&�<�1&�b�V�/"��	j���K�t��х�
����m]"�P����8���w�
��z�@�*�yצ���D��4{���#*r�͸�k�~�-�{r�����Sڭ4mi�n�JM��)b�"b�C����y��0����a�:dR?�G=�N�4g@h�wC+�a�8ili`H`�=�*ջ��y����X�e�t�e߁B����*���GN?�eD׷' �?��o����J�)cD�b����%絰@�1�F�^$|LR�L	�>.x[f'���Ģ�� ��݌8m4�d8"G��t{Ys.Uԧ�q-��qj��S ���}�Ğv�;�_��9��� v��V�������4)�F�X�!p0�K��<�uF���DP���|�1Tx��ؕ�x���V!�6Ҕ\Xe�|��� �*7�J&b��^a/o�� 	�=�b�&�L��#�������l ��'VM��f�gYJ���n��zt_!�T]r��d�)�q�)X�ݸȃa�m�C�/.��bJ(���kL�kˍb�&�ɤSt�q���Y�|i�A����E؎��I�CU�x���w��f��P(S0y`��8a ������\��@v���(G��|z:LE\\p7'e���
�Fv6o��֏Wxr��s��v����~���(�'�Ǧ�(���L�ֆK��7ƷѲ�����]�@l(\NfZ����H��(��?ɒ9��]<T����c;��I���g���/j���h����j[�<ZA�}1��|2n��h5��u]�[*��F�?�	F6x;��̈�*2��!h7��m�I�7�cU��C���Ѩ��#9�x���ko�c��	|�����=4b��5so{�]��w6S��v���fI���{�I<�b�w���{8Tq����ڀ�jLCu3^�^ء}c��y���jZ�m�'R����@2z-�U�t������é��g���v�;�����X����+�w�_�'0>�ײ쒷�0I�4�ԥ��故hNc89�������C���=��_��}3��"3�L=1�BZ��T�͜�Y*������=G)alS�ɦ����8\���,��Ge`@�hf���r�.k:�R�gn���,�-�^�r��.�)_�cL���8;�|�����&��C9s�:�Lu�*xm�:9owІzZ���n,�D���czݪ~l�ԝ'�R]%c���� ��M�k+u�@��CT�R�Op� ��C�u�@E� �#�og	Tx���W�,��2]��*j8�!ر��G ��������`&
�\"
�	�Jd>$�ޥ%�C�s�z������s�䌰�_�ut��g-�ٳ��r:1�nS7���k�©�o��xM�@;%. �a{���� <=y��B+Gv��Q�Q�0u�8i�X�a����~�N������$��x�L)d#�o�I�x/�j�n �˃=��hO�̯�T��z�Ja�_��������H��Mυ�5������h�roG˥UW�p�	�s�v�Ȟ��ع�0����ZSv��i�+d��ʵ~���b���������1��K�%T�
3��<R�Օ3.����M}wZ�q������'%4E�=:�e0d�j�Z0Yw셾�K��-��lz�'��N��x�� NC^	�g~���v�
eȶ�����0�U&��q���B%i�&�s�w���;53�n��}M9.�V����#>� )�Zժ�<$�i
+O�'�B���x��ۻ��&�20%�.V̱�B��C0j�X-�	��n�w��j����X_�<�|l%Ő��J�`�h���j+K��sy�g��v��I�h�3�$�i-���8�ێ�Qܡ��6��o����O�s�kF�:n/�n[�_VlI��}�@�N�N�-��ֺ�m��W5Z��FǱ�i�J��PW����<M��9�J��捛_�����Od����է�rjY`�FL���,�繝%�A"���_k�dR.M���_>P�ո�߬�|�23��ODT�rp�R�%߮H�v��zYp�H�=�M�\����6m���3F .�������J[���)]<YJ#Xch&�?<wh4.{Ch��olH�\�Qoh�p#�_�jf�Rd��;QƇד�k�@���cĖ��`�1d�v"P
���챨jkO� 9T��(1 xRw�Ӂ]ѣ����u�hy�̞�+y�/���$��,�~�������_?>��;)ԃ9�l�}�3�;��C���QIr��h�.�Z��2�X�$���<���2X�7Yؐ�'&��d�h%l ����λ�N����/a����_�!*x��a�b'@CLZ6��G���z���S|�e7N)�x��v�n�����U:]���U�5�9R�-��&+Z����N��K�ɳ����~�DȆ�k�+�n�m_���0�)$l��� �	��2*�+��R��R:\�ٵz�OAce�W�u'��z�!@H�+g!ٕ��wl�&S�P��~ ����Y�I�}�T	���d�����������3�d�+���Y(���L��Ȥ\zg/��u��t ��D�X���d�0p��2�eџѣ2����v��t#v(+t�x	������b5VX\f�ʴ}����-���ڡ q�y�?�<���:̹��-�M��}������&0�jM�Txٵ���Z�a̩���	������E��fO'��@w�|��_'Ш촠�!`�#f�<�U%�M#��V�h�{�Z�d��v�co$$��).x��1���Yנ~��8�b������`jङ���5ϥ�s��䂶�U!yw�w�q ���Iؕ�Y�ь7��PJ�(�"vee9D�64�p��̣ޛV�f��T����J�Q��ہO���ZCTY�$�
�m�:�4$�F�ᾍ9#�u��y���*i��7eG[�ل!�ȝj/1�A����ڞ���\L&,���g���R��������j73BC�\�����ag��E��]��CD�Vu�ҥ�3B����{�!AXE��3GT�1ċ���D��X��r}�U���9/���o8D���`�0B�"�;�5�mRl��VLH��e�/%�Әpv�I�K��b;��Lm˅k�Ŷ��c�aeY�!����'9�"�ZQ_/�i�G�b<tc�&�?�¬-�u�wy��,���x��HG����׀C
�A*�d�U��ׄ�ǻ!�~�uB�2�
K5��%\�L�"�L�2���K���#��ж{J�Q�t�� <
�������o,�X�lx9�M����A.��jJкw�k��c�de8[Q@X�sV��t�p����pe4x,;/L�C�y�*�E|���La������������->4��iՍ��]���3��4X7�޼;`�"��x��Z�E���q���F����_�У6Aa��2�d��.�q��Sw��5b�s�MX��d�&�Owwd�t3YՄ�w� �͝�؊g�k��/�!ʖwE�IΕ������r�0~q0��ϱ��w����X�t��x�i��U	M������ŀvB���|CE�!��ƭz�����-��dr���u��J��Im�ۊD�A	1��F#�:E��pPrL�Щt�tI�����&?<�}����N9
Z��[���F`p)?���Q�΁C;E�ڥ����z��7��}3��3��,�2�{������g�N��}�4�Ć�mI���FP�3�Gϧ���lI߸�R�����=�pM�.Ry�I��ZK<RM]�\�C= ����]~� -V�V��2g!e��~^:����p��z�Ռ��| ّƙA��D�fihߺ;i(��j�X8���~D���w0�4�������0Y�ُ�̩­ A� �g�!��(ǲ�|�x-ڣ1n;MU�2";�b�9���R�u���Z�0��?���ހ�R���e�:��E�<�b�ZE`��0���o<�u��]�Nm�5cV�#��9=�н�O�C��������R��4����	H�3�Ө�����S��5gǬu�G�r_<3�hK�
SD���FPD5��rd�UCK��L���<����s��L��C���>��ڢ74Ҙ����=bK-��d���Ce��$"R��/��e���Z�����-�{KK:�zԙ;����㯢��[O�F�U�V�
��ƍ͆��]�X�Ɓj���i��ߜ�!5
J�H��@KyJ4�EpT�}������a+S��H�g?�Q�?7�P���Q[�|����F�F�nj/:����Ft�w �i* �=��j��h;�UH�D�ƚ������H�_+a�� 'S�0�l��W5���]ZczSkʑ��_%β1ڽ�Vq#�K�<"w۝�ׅth���<t	�C�����&
*���p ay�;�!�!��3,O_/����<�4�_�0N<�4�*����N�kRl@�`�]���#��8G(�B(�=g�k��~���j��ls�b�Htv��4��)2By��ēB��ٿ�ڻ�YԓI�ʿ_RJ��2���}�y�K��r�����@�h�v	<������Eȼ:Ub.[���C�tj��=Kſ��rR���a��Ԩ�f ��FN;�	sL؅c�����z<�H����K���I,���y�U%a���[�^��/����j��N��' �*���z3y���0[}H�\�x��]�z��,�.��H��P;��CX���	�%=����h񇠲N���.E�y��3����b_Hs%wB�2Ͼ?H��+)X�#�;�G��+�m���3�G���[Y���.nr_���E�A�U�|y����9�O����*@�0���Zt/;��Cm������b�L�.�+<ؐ��V&��Hm�R-oϋΐ�J�aKb�H*.ٞ�(~�IP����P�f%�]sw#1H�3����Gi:�V4�7�K�Q`D9�6�}}Z�]L+���i#C�g�:�R��>�:6[z�ʰ�?��zQ@�k�6�oi�\��3	�����ē�F�#:���U��D�Ud�U����|��f	�ݗ�'��G���]�)�#=�ݶ�\X�&��Z���N�}&d���zi~i���֣��> ��G�*�d�+��7̯P��s�orN԰ޡЗg6�Zsa7�v�{%'����u�AfC6�4+��@��u�%=%E0ڠ�!��L��I�@U,�R�n�L�}>äM���-���,���Fя��Wz׽N2�M��%zL����r� Am����HL��HS�_Y�}Z�S�JL�J�[�;��5�]�e53ȘDz��u���	��M�9in�,�s��}Ʌ�¤��d�	���~�Ξ��t�v���. ���#D��TS���gK9e�?Ģk���{�����I�0�A/��6VX� 6�3��'Gs4"�	k���Fe�%���+���7D����C���ĳ%�Y�Va-�����O�<�* 	���O�-Ԍ˶Z=��RB�9 "&=�����A!_d~���s��o�L���o3�p���6̀i��FJ�2��jҐ
} V��?p��������Z�&��]x�j	r�o���z.���^�i����3&��cv��Ҷ��z��� Q�N��că�/h|�����+���)�LSd	�{O����K��yAf�M���}�?�����6jx�Bs[�vm��+)1�n��zX�Zڌ9�f<�к#=EQ�j�ֹ��!a6.�m��s�lY�V_��4�o-o�7d���2�A�E7j&tQ��/kR�Rpm�u�ݻ4�M�Z�9���A~(��7?�b�q��3��>���H���*���6��*��j y0�(Rrӕ����]$]��f�� V���?U�U��r5P�w	!���_�i�M�P�V5����'������yI��Z���~e�{��^G�"�{��RPl�WHp�8��֬��*��"�& ��X}�h*� M%�v8���r���xB�0cᏏ��'���k���M�T~bϚ�C��Վ :�������!jh��C
c*|7�OQEg�37��Mv���U�c���yW����#;ѝ��p�r5�h,���MLe�ry��؝���	��"��n|3G����s�DpT��Hq ]j�#]l0EɃЀ�u��ۓ+�SJ{�M+/���g!���3	}�\<'c������pd��ҋn�Lx��ARe�D�}Z���'�9����w����R�-���?%��T2u��c��D�>9�嗼�Ud���>>�t$�T�������$��U,K�%�{�4�/�{Q��$��-a>tn�]����6�{���梘��a7L��!G1<��.|�I�˷.�F�������B�-͎R#b�D�&�� ���cɗ7�\��ٷ/�H��n�ce�0h#Q�� �Y�]�
}���j��EB�zO�ȁ,��vT�-wR�
�kKe��)�Yz�"v�Xw�p��
���x �	�[�r��O!���eumr��I��r8�hL(��/�2�rWM%���D	9/mi������7��<���(��I��N����@�=,B�6�O�x�f���i�W���*L���
Z���[�[��7c��L^vU��0=a�$�������.?L/�`�H�Ǝ�m���Խ�y Gh�-��L��8w6��M@�nږ�d���fZ|c1�n�|������Ñ�#����� �z��a�fF	����3:u;��h��6�9&�|Dh-թ�]F�΀G��7��˭@+���MT�݀��?�����ݎ�����r�N�M�N��q�eYđo�<��=Q�>I�m��۳�$B�;����C�S@���ET�s��Yb`�x�V20I�<q�2�y���~��/0R�7�]W�+6�(��̘BUZ��GK��G��3ϻt��Ť��vƢ�k��ff?�g!D?P��G�7C;��:�?f���6�{�_W�G���b�F���!8�]xN3���@�nx�F�cw�.��m�w�	��o��V](����p�ƝZYz���e�����9g��uv��oy�~^�w�h�r$͡Ø 2m�
���t@��'uxO��J�p�v�����kc�x���'�e�a	��o�}[�;l-����������&T��T�Zpa|�x����oY�Y����y^K����P��7N~b��`��c�.4�2���Q>��b�1G6q��l��},5bOd!�0�C�D3��")-'�OjW� �C�s�x�m#�~�M*��y����:L_��&E
�&}��������G�@�����rL#�ti��`�R�u�D$~y�19�@hw��e�ݕ@xj���	 O�j�����b��4��[�kбf7���T���~��y���S��ٰ!ʣ��� �D�Wz:ۡ��Q�-D�d���u���3�k���ac���'?�T�Uc|&q<�B6k���ˇ��~0g�����0'�hA��5��{��vr-s��?�������)�W�w�(Q��(����[κ�$��:�*Ov��
*�I㒖6={f؃�6P�w;I��P�:��E��*}�F�y܋l��\:\ㄠ-��Ȃ��=l�VA�˹Zq1: x�'��*S��sq�.��[�)ĶT�3����:�7e�1/#b�v������WQ��IbϦ��<��jTÈ���'��cLn�w��dr�q�h�����>&�T��BaA�ꅀu4�A�<4�^���.����`���F��%9�TkS��M����U�f;t0~��t����_���E��N��fnt���轭�~�� l)�'�ܖ�r*;M1�[��h�-��NX��p�T�:���Yf�q(s���_��j�E�(2�F
�i�wC��_���W��D<��P�}uj�
ܿ�m ���;h�f��澹K}�'��	��@�>ˣ�X�d3烯������G���*��TU)^����gI�9�_|z�0��:?H֖�&���=����D^g�'��[B�}��
BU����e�bχœ<�P�5��]{}Z�@�g�ԡ�qb�����})o�Ͷ2���b�ٯ#az�����0H�Y)�8  ��L=��eᝳd_���7����ѥ�r�����>ƥ�5t�����?ҳ�<+�t%���|]v ]������V�Ń��]�Tfo����.�]�b*�DTN��𒶓��@9sY\Q�^�U6UQ�#�����>��&�sxl�Zv��ͅ5�\H��xA8�r�Z|l����jď�z�Ĩn�z0�D������X9Ĝ���U�S��� �6��xs�����=�&(�aR��3o�܅�*/��N��������w]K]5L�b�,��V;���[:��3���橉��@K\��T��Mۋk�l����C]�h�+"?߇���(7����V��߁�����	��鮢��'�+(���w�d��^>���(���}�U��-7�ML��(�� �.b�_��gv������7��ec	ultzȍy�zЗ�Ȱ�$��E����O<Ħ�s-��>�_�f�-��[8�t�4,(��� 0�+}�j��+�A9�A����w�~��x`���ij���6��7l������t#����������K�48x��A�ר�UNn��H�T��R;6'�\��zi���u$�t1'�fc�֏��3MT:�N��6�7;_tWd<!תI��,9�7͏��+�Un
4IX�!��1������e�|��#��F 
�0/A	w]�b)/6��g�a]n�
�5�'������4�"g�d�e���Pe7��@�����f/��� ظڪeǅa�1�S
<�3��z1��@�C�]1J�K�N�ml�]�xQ�߇
��
��1[DڦFw?
��9��z{��mf��)�՛����ݦ�C��5�ӎ*���8����5��x�<?X�6����s���-Ő�|XS��y��*��*S���w�ǉ\+�^Xo�-#��R�H�,���;�
P-/�U(��JƐ���}�j����7܄�)��'��s��FCͅM��\��(!��[YD�C����?�����T�KǍ�X���.DS"�J��ϙ}Ȓ�|�u,vQ��ͧA\rb0�����5
���2�u>���qz��eK���t�=�8 �,��V%f�JbA�կq�b�L��M퉿��g7����W�>X��hx`�H��N�&��r�Oy���.���I���e{���oӨ�N�0�Brf|�~w��ޏuJ���SAa��~�]����}�m=`;eu �1����n�c$�0�q��Ʃ�ʙF	1��
��V�B���5{)��$"�H���/���;W�����+�%��v㰘���4��l{F����i���j̛�}��!�@�q�.��':�d}�(*��2`��f�:"x��}����HN��cpu�+Pj~��a:�X�T���Ĵ2���'��k$;�,t�`A�iLBb�כ��iBVĭ5��R��υS��X� �>p�^˾;BhD�^��i��T+���:-��I�_7����fR�.1d��J��x�/`�7�V]��Қv�:׎�X�-̄i����Z�n�D�u)��jK@X���R��z�D�궊�T�ziR�Э�M  6e�0��G��M��p�z����Xɢ�nI,ߺ�i:w��;yw���ib�T��Ԋa����W:C�X����<SY��>�yz��I��!m����rJ�&݃aP[���l`����ހ��)A�̺�5��HqgErx�5/W����i �����D��um-];����o��h�l\�N��!�
�{��4�a�d�!�dE�_p8t>����r��)�X��H����M����Z_��9��7��Ă
��2	nrbpg,�]�OAc�����M�شp|��jki�b�rb�('��-�륮��R��ߋ�:CXO���L�h@�Q�,/�u{�)�8 �
\� ��d��?B~<���$�D�*nՌo�<��	���Y�	���C��rр�WÝ�����L���o��}:P�|V��@�rS��c��$��b���>�)�&c�G��P��b^�>��a���C%ljc�n0S^ȫO~���A6���*�nI��l�^�O*"s�G��ϰ��c���t[6@[�D��o�zz&_"�6��[���#�5O�Q���s��!t�U~�}�cK��\�'
Z�RWa0�fMn�)c��6�ϙ9����G��R֓�a|c�΁��G{\➫x-[���x� ��X����5�;���n^e$�$����W����h&f7���r�ŉR��Jic֜��Xs�vS��R���=��r�}���iW!��YU����s���CMAFU��8�W2����qc�!�Q<`�fq�nQ�pm�����ӿ��dc��P���9U>Ic��}�>o@=z����#D���RC�0���+��򲑯���=�0�d���d��BG�6�PU����J_N�]�Ś<��5�,�����a~��5(h���!q��0��%֎��ϰJ3I t��w3��w.���x$\�sU���#]�3~'ߢ���^0��I��Ǣ$��ϽJ7ܶ�H�{Bǋ�/�逻��������灳��CƸ�+�9����M���e}�nP$���Jp��1�M{o\[V�HՈ��Y�rԈ�na���
w܅+C����5(R�  p�D�Ǝ�)1m9�π��%����{z�gw���Z���V���=�3��7ʍ�7�@���~b.\&|W�[&/Z�G�;0b���=�1��+3�ߡ2[�����*��S�y(ʊ�+�� ]ūAR�,�ȶj��	�S���Ϋz�u�ޮ���*�%Q�Q��	6����D����Ϩh^x�kV#�>?�4S\���O��>[�D�{�46c#�Y7����Zr�=&;{����
���w�Ư�&��B��/+5>�F�f!��
O�B���1�q��/��HrXFh�M�:����(�^�v�ACŧQǃE;�X�\5ߺo� �<�E%��סb�G�a�VKÎ�b��l��Dc��;��r�'Ei���>1�cPi��w��ñ�)?�D|�F���S�R�+�p71�Y�	U}5^5U/ ~��X�wI���{�8�"�=�eN���F~�����d�2���d0��{.+�A��Ru�N������H�q��CM��� �j#,u,��=a���6��mMT뿉�8��������ߘ��nLY��n_�c���b�!��64l�K[˦�&��^F�Gy����R�B�K�<���(H�ĝ���9x�%��l�U�
F��N%LA��ޖ_^�&Go��}���2��OC���	wg�2*jw�7Nu��J��p��/�U���EaH��~n����T9�����J�8ۑ/��YW��mm��6l�4̞�%6;�8�gR�e~�j��x0}kӆK���ˡ��O���ҹLpb�T��yu��Lu'|{`Y���v�a��QA硾Z�R#�7:\��4{������<���)�G�|���s�5_
�f���-�/i,���p3#0�K�x��_r�[;1��=A��D.M�pǚ��酀/`�J����V�Z��5N~籏�Ǟ6�$ɫ�,���$S��e_����va{����(�7r0E�e���%��	R�}�5��A"y�c%ÍxWc ���X�X��w8bB��eQ�%��!wR{�!��Q/�QB�t0�%[D�1A�Qll@m1����i���`ѵn��H����>�7�ݷ&x|�S�y"��IV��V��W}�d��U�[�e<���)w'u�7�G��T���Jy���<dq�)⫉'I��,��G�_�I*�I�X�k!� <4��	�6�j��٢���6�-�Q�;��Ȃ�v5)-R1�:2���;�~�@�㟰@�ggX+	��k�oZ�������J]�o'i�Go���Y	��VYs8f��SlM��"Qr1�R��/�NcT�t\�*NZ!R]��1O���UK09t��HΕ4H:�&�1����+
F.-�h8C��~Q�ZMb�<o�EJ�~`��z��d�����؟ȵ�!�{|F.e�5���1�j�Ϥ{��MҰ�w�-u�"n�F�6�|�-�����Y}_�"�����9O�}�M��!U)u����,Q������^FX��e��e�x"�H��*ۓ�,���i�.��i�$�JK}J����H�#�,6-z����3NU��3*g� +$φ�x/�G�쁦�05�A��gx֯�O�k�\~�ũ�_?��x���b��$$�y$w� ���	o��_���Zo�=ѧ>��r��o"gI���
�w�<�j� ��<e����v�Q]����|qc}ğm�K��/�P�:�}q�ږd������mC�z�v��l�5
�&M0F�s�WE�z�;���hE>OM�z�f��2N�8q�q�9�����d�c���/�c�e�+��/��ݪ�;�"���ܖ��_J�.��)L�ĆA�/�8"��������~�m��\f@f�HP3�\�12��p#�G`�ٖh}# �[r�m�鄳R�T��So��e�Q��w��"0�ףP�[Q��`��M��7�N���r���1K�eqC��p�涣��\j�Y|oKx���7R����ll܀�=zH{i4�ȴ���ճ��	����X�p�{��#A�4(I�����ZZp�o�R�<�2 U���.v�c��لm���HE�5��\.)�`1�gv8�� ��O,�R��G�+10w�bI�����6t�P�_� r�L�B =7[+e��G���S����R��I�,*��r�> ��߽��L%8Z����{����@���1X0?�cP��2o��X���0�n��Th��P���6���v�.U���k�I~�kCIvI"Q8��xٺd��9�lRT� ,SF��f� ��3�r2����`t�� �zԠl6ߖ��B��C�Go�U��Y5ʟ'�O/;7�����J�,-*�4T$,��F&��?�:$�tB	���|�xqՓ�*g��I���!3��"a��./�:��09�c��z��у��-7>V�~�>���/�m�Q�s,��#�7�I�l�p�r�H�\�u�J��hN���[���^���M�E5۠������p\#�����}�,H��F�p;Ö�'݅T�����,��C&2Cr�F*���/��b�'��^��e� ���	���l�Y˨L�1/����S���4{�����7{�� y��[=eE+O8ӔkM�_HŒեB�3׵Q��@�2a���j��-D^:}~Pj�.⤨�M�0#U�c�Jv�a�B~_EEr�t&p�Ȭ.h�N�tL�ѥ<.VpK㺮X�88�.~�?�߬
��;3�w��k������s�l���lE��`� x@��5*P�	�dV�ͭ��4q���Z%1��$(�����)�$X�ls���u�U�ٮ_@<����U�p���r����w���y{j.?Vho�ee�S6�0K7j_�s!���C:��!~�_|��~�`�_��������;�	L}�n�_���P�.Z�5��n���ɉrT>,���)������1��L�깙�QH�g,��-䬕;�=��=R�|o���{8�wcI�vPF�I�����?w	�-�YlY;���.��<0�8,�=�Q869J�Xh� �8%�����^9���`��V��_��w��]�=+� B5�V�
W����b7reN�Sy|���p/�	�Oo�r�!9G���a?30�oBn&*؁)����I��L'��П)���fx�4���=��ߓ�"�ן���������o"~9E*����#�[ɑ���l 6��{%�/
ӦM��Q�?Ү&i�ʹ�CxQ��E^�kFR܈a���`����O+������ ���4L��Įtu6���#�����M'�J[I͛h��~T��]J����.�Ɠ"�w3Uӊ����IDߟ:�b8�g���9�˙�h�i��$>H��Y�T=�Pܐ���*�	��)����8���|��E�`A����x$M1��5��a�	�ØМJ���fB`C=zG5/�C��j,���Y{��]���<x��~^L|���?�g(e�4�R0�Rw^�M�ae6S2���ϥGӑ�t:������V��N���8_�%��,�'����a�Mb|�łl����~ӥ������X�MR�RR�P�j�L�ȥ?gsx�GG��r��$�ս<>V�0�5*Mo#{_~���<J��X�
�55�jỞA������?�|Q��O�	Մ��[�)�ګX�W@+��0��� &>[n��T�j��'B⻦�\00�qP\�D��"�i�a1�ܹ�^����N�Q-���H��+E{����LRQ��~��G݄�mP=�I���!dh�M�#����}eu��$8��F�,�I͆{��AR`$�����ө�Y=<�Cdc���J�2>�"�K$��V83eB�5&+W����� X��V���d~�����_�[m�>���A(�a�f�"5Wo�7�p� ��y��eKM����5����g7DB��17�3xO���*��Qԁ�j��=�&ܠO�G?eSP}q�o�X2+�Z���Y�3��U��3��\)�E��g��f�������(��L=-��~×J�nE�Ӓ���襡��&`��&�}U�&�w �ZWP�r�X���̙�ϲ۝�E�GJ����0	D�qA�.a<��Jy_/�^$�w�]�}1��5F�(k1�S�D�{��+�f�+��:/��h�x��(���9���R�r}���l
���,����32�M���[ՙKe-�[B8��%�ο����㶚M�r!LQͲ��E��l##$�R��{�
2P!�DR"�*A��������Ӿ���[�u�'ZY��K��Okv��9������Km�>ϔ�Bƚy�0o{�A�e��*�Ĉ"�$�KTK��^��[����EcxI�L_��ʖX�I��,8V��TȎ�臰@�r�s<���1�U D,�v����C3���q�X�"3v_@M�-X��V�{i�ƥ���x3x �6�g�*v�/2ʰ����@T"AY�~T���^	���>��C�Mб�p�w�?������]��E����w��-�����!�un����^�.6m�Ds�%^�G�l�H��{|U �Y��1i~>�iԻF�u�o���3�Tq�#T�� a�C ���L:>%p����F,��6�ڡ)yR��uJ��g��t`�6k�=� QH�_���lO0SP�ٺ��	��[4�FI#�K$X�eod�3�`*Q�n#`�,\��b��N¸�ዜ9��"�+��{���	��ϛH^@��:]��1X�	�N�n�W!�X3����N�e���6�C��A�,A[���_�L���@f�I��~��"B�2�y	뿙�d8�3�y��G��=eu\É{9���4e�}(�@�!�k��A��=?��\ڟw-���ds�4�ƧbY�e���ۥ���}�5����a�����RG�?�~ޏ��լQ_�6�D�3X�ݨ��o${���D@�ꛃ�-|�tF���YH��_���-���N����g����/�%��n��Yq��ږ��{l�~Ճ�dA��ϧ��!�,�V�a+���N^��B�	�Ȥ-��`��폎_� `��I��3��>��&�+ۥ�L>�B�" pЦtg���<���ևI߲}p��GTMx��n�qck�e��8Og�G��9G	sO�)k�g�K<����+���q߅����!0�
T�����v~ 0�ؐ{)��U,�)AA4�H#/\��6(W4��E�O�U�zh���R�x����,n��)�"zw 0?��z5�MbP�Ԛ@��f#��Z صT���� ��u��w�3k��PK�+H��|J��4/.{:�C��W$:'.�,��F\�92����Z�@���9��/|U�s�=[�Q�k�x(�;�1%rv����M�)�&�����i\Z�3���Y�Ɨ#W�ԬN{Q����u�K����m\��+[�5��	����Is��n�FR������Y��ZH���U�n��cT*�Q�T����"�C�;�K딂�L�Tz��w8�G��wL|�������CL�E�Mp8��B�+w���U�!��q��!�([2���О�eLD��4/u��s�|�{�v�FT�-,�'l\O��8��<gR� �@����y4�L��`�,� �MN��*V�����@K�GEu��:@w�{�(�<K��ǰy����7e�|o2�<�*^�ދ��Ry���+�;y]K��MOj��o2�>�ߦV�Rl>j��i��'�M��h� �	�[�]�0�f^�B�R�T�i=7�X�~ ��N��� U��RoX0��+����-`c��e���X�I�{��g��1���,����-�P�~�(�io�� I.v�ϺE|6���&T����`{��ң�ոL�����ٶ(H�&*�rM�8�׷<`�������m_xP:����ʆ��i�@0���zͶC��N`t��t_~�E}�AIouy���*��TS�>��?p��J��a{7퇜�j`����LX�}���M,}�	s�}owq�t���捥,��Q��飢����=u��g��ڤ,#*���ߋ-�a��<ֶ�$��^�9�.K9?�ŧA�1��~l��k����A
���=~Xၨݽ&�@w����*�r�K���XM��Cr�!6ʱ�5Ȉ~��P�26�l�����Ղ<<�RP6C��*��t��a����Zy�"ʍ�,E�����1-:�d1=�6��5[<{�Ơ��O�Y!Ds*�~����ބy#������x���r��� ����l��e�S��`��|�?�9�A3ާcuI ;�����o�G11_�]�%a<��&G	��UnJ�d�?��w��Yh�>�8�{|n�㗉>R	#<�	�l��Pل�O�� T��|��d��b����VZGN� �R��
Ӗ�="�V}S ���T!=����SY����AX�������:Ny������+-{H����1I92�I��X+I�M�N>,"�e�(��c�n�J����Y�[-C=r����r���)�E�u~�M(�X��C�tg,Q�_�zXf��6���Z$�A�XF��*t�)g5.�������;) �Q50��!̡LrT���Ș�a��0���N{.�yH�fʞuIӌS�{ڪ޾��t<�*�8a�y������K�TϥKL(�|�*�܎o��&�]�ک�S_���I+*9����L>ύo[��T��O1���-�^�ՙ zƞT�w�����2��"X�L�u�=n��L��I�h%�Dٞ����xuOn�zPY1�⭢4.�c������"QD��zd����!�������[�O�����~I�R�c_Q=��ɪ�'+���?�ˈ�M�0�V��l�FiL�`+��+B�*s��>	3�ۅ|��eNf�L�BD-�2t7�yT\��U@�QP1�>�K��~	���?m�s35v���B�LW{;@K<�4ـ����{5���!�Ā��3���<���U��=�G�?����w�Be����)�B$��E ��f���lA9x^��|_��5�m�M��I�z�����x��TV"�}M�N�]��	T�ڞ� ��R2ŊM�����KB��CG���WGV:�4)y*z3�G���n�^�����I'�[̺�: �܅��:����%�1��J$��)~W~cls�i�ױ��b	%Vr4� ��τ���j^&��\O ��fݕ� xX�f���T�2AWvA;�ԅ�sZ���&�d[���:f��>���{�P������M���_�,fQ�D�l��yĊ5�)�:5�k����%���iSsQZ�)B ?2R_Z�M��j�%T��ݫ��7��۸<z��Fѝ*� ����Jf�����R��v>����p��e)[�իw�O;��qI���
U��oPU�ؑ ��l��|���Xݷ��(i�MQ��mϯ.�ˎuu~��R�OƦ���Pm�8���Ѕ�IϤ:����W��3��[&� Ϲ��Qm���r����2,��]ĩm4D���U�x=<�����p��?���if��*��v�CA?8��Uo��sꂂ`;���֗7��zSc���=�����������\	�q�*��,�A~VkY-���mG>4`J��5�Gkk ��k�d��|�����6�56�'F}��E���RgY���?GOax1L�BLn͕ġ��Сo: �R?�R� ���ne/X�c7��S֭J@�N�W�L�י�Mf�X�Y�G�h�S��GJ�BR�%Z�s�%t��d�KV}���c����p�=.�P|ޜmxj2��C�����K8��a.n�y9[��7\+��M�,�@��#w�|����[e�PHK:�m�V�8�)\�{$$,=����(����Qz�N�_a�ݖ#(��/�Pl�0JS7Q��I��Z�)����]����`�E��L�������\�U��Ɉ�L�p[U���e-�G�I(O��H��?	��d�R��e�Vb���G>�Hq�:�*I&v�iSY�f�}�6���7�6�1��:�d��0M������>4�c��F�BZrn�|t�JSS�d��8;[g�{��L�44V�՟v�7�E����@���}y�:4f{��)�G������q�q�?o��IְGyǯ�A�BqޓߤA���uHN w��$�S�M,��E2w�!�Ű!!HcKS�7h�l»����	���9>�^l^AK�0���]��	wM_ !k$&:����fj�N���X��E1�Z��+&���r��P.�&���P%�I��E�z����Ak�V�@b#G~����"����+i�z`{Q�S����)���Ǝv|=��E�)@5��-�%B�������6�~l�^�Ow/��9b�޲�=�TC�u��/�@�z�h�7a��u����g���xr�|/��������h�����[t8����N���5R��b��;.=����o�����.`����/qqϹ�yˀ��ԫ>�6��
lB��g!(��`b�2>l;#3����w��(
���Yכ�#�ξ��u��P�S�W*#Qx��2/|2��a�c�T�m�FښZǂJ���~��D���9=�F�ףo 1�("�xı��H��	G�k`��?��,᎑��k=���j!_� Vg�cǆlT��0#�:�r �!�R�X�� = �8lS��9a���"���{�ۊ�o��Q%T��慜��)��G�XKG`C�Z3��R�B=�G�荃=;�6�
n[Z!&�kY)V"�d&���iSm���hm!{��̘i��+"g�M��"k$����?������>R�F��B����Y]�vlS�o��|4[��(�^']7+C��ʱ��&����s����gAx�{�Uu�DI]��j�Q��/sᅶ��T��1��[���T�e��f	f�m8��W#*��P�^f�-��K(2���e�ӝ;��nt�@�j�U'~	Q��
�����1��f�V�L��.�ț��/H=r�<�v:M�A���-��E-��<���Z��GW_���N>�p�n��g*�p�p`= $��/��'҆�w�ʓi��;h(ׂ���u����@�\d;n�Q�Vi%�q���"I��IB�	����B*��J�����t�*�J-X�-�&�!��O���aH#�I_��u�^	й]�w��Y2�Z��c(�!��1�$R2%!�^�1:[�#P�Ӡ��Q���Icr:q,� F��
g��s'W�_���u����]ʎ�S%$�H�.�)_|���s-�*��fH�/e�Q�cu��syNN6��A�<��#�ƈ7��{l��pU#m���n�K�����qf؀��#,�x:
4 V�ՇO�H~̒j��:��g��|�.K�e�Tވ<q�s����^��̦v�8�=[H�=% �C�VE�����m�s�vM=e���#��`�Xu���)�	�>������g�n�܁�Ce]��¤���<e��<6m��K��M��?�A����c� ��� v�&ǔ��p������[
1�Ot+��Dm#�>�@�4�XՀ��^juZD�K�t�����s�4�������e6�?���h�%�#Β3��"4xf�B[xgy0A��[`�G�ԭ�I�SL�� m7��I`u ����&YZ���6L���z��1��7�Sq[#ܸ0O���'%|�ҷ(���7Wai�2�-�~+�F��Vl���+��xv�v�	���a--@U���#C��dI�ۦD	��3�zn�E3���k���<I�@�
0�
��	;��ø�G9/�B4��Er��¹��lZԴI̩|E�-�<�#��)2�!O�YGa���_�[M��Ⱥ�
�4cx|V�,�
& /q_��%�!�rZ���ֵ󳾜7H�V���e�rsW�����d����N����վI1j�$��ؘ|=�v8њK+1�g|.��nfQSM��OJdC)���k����6p%�J�U0s��< �	�o6�I�~�3��$�F�-�&����*"nA���K���# Fё�ja.�VC���98��ܔUH��WO���Y��.墜=ү�Q2ˌx��s,������l�촎�Q�D�
��&�8[Ѡ��0g�,|{�qea�B����w�b�A0��'�ǿNn7iK݌#�C�l���a7�7r�ؐ�"�/��g�!��g�4�Y���S`E�ӹw,ݝ�p�B���oe�����BUj3�3`�E/��[�a)�s��^��N��\<����1U^�L]A�p[����jkF �bb�I�9���z�/�Өgq6n��j�v��Vݕ�e�!�{]v�8��$�?���>�<�8}����8��i�ƺ[;<�R�~�����n�m��� ������IQ�yy	�=�e8�?ɒF�o���Z�s#m#�gY0<�U�&�:��i>9<�R,�K��OF����V�Klu�%M��oRĩ(WQ؎�94���O|�D*��v���ldK��,��7k���yPSB��� �ow���.�s�����Ђ
|%�����-g(ȵ{H{L&����h
f�������B�ih���GOZ�g��2%2є~zr��[N<N��F\ ~p)��y�ͭ	j����"��x����"�*)�kgLqz;'%�k�?0�nIZ	g����y����4�7���Ts�:E�T"�g�j��:�	`�î�Θ	�xN:� 4��B[>���ߐ���������Ld���}\�mt�pK����m�CfT�����ZP���孏c		ց:?a���߃6�0����(Go���/��3���6����	ڳD�����@�$��tr,̛c��t����뺁P��X
�w��(L/|�:{NQ�$��I5`������(*�
� ��GI�Ɣ!�86�Y�L&�e*J��GHuO�w��pO2h-�`q�e������ �BT�ʰf��8��V���"U[�{�$���*{�R�1��ɍ'�eM=�s��"�;� �.�>P�Qޗ1~�'��ƘPa ='19�;�$�ʳ�gK#N�p��^�ĄT<
��2<���m���x4:K+K�B���bD���v�n7ۦr`�L6�����}f�+����j
��ܣ�1�����vm������io!�n*z��Y��fue^k��p]� ��Q�0�_�r�����wf4�����qU��D�ؿ�?> ���ڗ��+�X����z��We�&8�uvD�ֵa��ؿ�X�27�\���D#�����bP��VA�
Ƴ�?j0�����H��*`q��i��M"�vh�Y�r�S!cn��]�k�8Ɗ�Pk1���3��PD+��_H���7�������}�fn������I$�'�|&��u�{�m��j����Em�m

*�t ���~��v-o���E��pD�(eBa��O^��8W6�R`;�k!��f;D)�;{��ꁐ�3T��=`�0��U���_���b�:c��cx|���1�*����^��R���Cw��]���-�uD�t��$ �"G%���W��*)\�G�f| _�$�RAJX��K�I���1��tz$a3��Q�ii(`�kpkL��c��C1��K�/ʠߨW���6<8���HTV���*�
���#��DA?�ͫ~�h̿��#]�6�3K���W�wap��+��I2׎��&MX�]ɧu�ϴ�@\��PR�$��VQP#w'�
����q�:����en�_�Ikq�#r6�_z�����y�����$�I%�v��}����$z�v��NcØ��L*d
״�b�㦐x%2�C*��%Y�I���4n�O5���B�T8�͒5����z�'�|�!���߿�2�'�c�h�� �9����(���]��G�'E|nc����^6.��G�˂�d�:�J����63w
Ek�> s�Ɲ�x�~�p�SQ�]�,�|d�e�7G�9d���XrSN�#��������G	�-��Gv�������]ͬ�Om�BY)�5�p���n��4�D��(U���
s]�e�lc
��S����E{�	��J��6�R��:tэ���p2[�
��,a#��'}�F�M
����V�Dݥ���(�" �6Wr=�jp?���$���zsiZO�k�V`�
2�8���y���5�] �&=��t�}O�	5�>MTu8�-Y�h�����lEC���~z���(�f�sЉ�қ��롹��o�?{��U�eV�k�"6�/a~��7cڦ
�������>���v��A�������a�1�mc�"���2��Z
,�co6�.G҄��v�� �+�^H��:۳�$*muGy`�[T�q�*���ʾ%���x` X�p�߄kN�5�ì�;ҙ���D�Ti��}��N[�e �0�R��m�.�p���8<�y�/�XX���##i��[E%#�R���J��d\���:�4��j���[o�2i�`�ho�yK,&w4`r�Q�p�:
L ��ьo���|�]m$�6z���|h�Z�����G����t���%T큍��U'��QH�K	0m۪u�j��R[du�xy�+\��;��G$~�?�Q�S~
}@y������ۋϔ~KS(N2����}-9X��*{��YEɔ����:a����T�qca�����w��e��+T���S�����_�Q��!
�fE�Do�E�E��ɀ!HL�UXϬ�"b����Z7�v�,<�u��P�%,�)nM�ST�X�y?C;i���$�I-�t���Z8�Y����P0
����5H>���Xޣ[g��䫶�
����!��CnL�T���%��"N���z\=�e��$Pi�_�T.f!
ʝP+[�|d��>O��;��<$z8�� �晴V�H�FW~ͺ�Jd*�.�����<E"�@s�d�9Z� ~�]Կ�պ����ɂ��(�Eη�y��S��ˤï�\�����z��u=z^e�G�:�xT���d�ڀ��Q�m�L��qS��T)���2��49�~�ď��e�Z�W�n�c�3�畁�c)�?
[�\��� �0;�����'� ����VV7#���~��ǢU�cY͈A�k�u��t���U�n׾�hf�b��.�KX��M�1r!o��*�S8�Q�p�N�-��z ~\�ZS)�2�Zag���=-)�	K>����v�S��i'�mHAߛ`�i�F�.�V·j�G�*m2�uWi�N|�&cR�\����jtS'*�h.�o���}�\�v�Wv���vsѶu��H��䂡Us��B�����7ޥ�j����
�[��+��6���	d�����7���*�J/u���̥�
.�o<HT�Q�>y��\�"�����u���}�Ԕ�?��*_$o��<�AL��Ul�BҒ��&.~�H����ɸӟ:���`	[�"7ϝ�^_��N���a������[s�W���'�����\��!rSoڪ���Ț���3���7��ݼ�QSy�b>jZ��.Y
�0���b
�;E(t����R��i��Q���I��-�l?|��6�a؟#�
��x��O�L��K��O�c��6�fJG�ʚ\�B/�q�����&2
EJ9q)��m/�f)��]��]>�9Y�(�U���e��l�Jp@V,�(�}x�H�A��!z�G�qB�\^���,�z2���)#��(�\��c�%!��|���Ga$:�šM.\��o礑��������N��,�y�4#��6�	l��&d��!1p�㋔|�m�KζH�
�*o�&p���FY��6�#v���euѽ�ef/�|���\�iJ:ե�V{��\!ך�ѸD=/0�
>��]��}I�c�{�ÇO�j� i/�z���`O�@l�%D?���t6��; �⫄z�ck�c�Z���VJ�E&<Uuу�"^Fߑ�5oi5s�a{�bSM���� �mߘ�4XP�˗m"�|N��n��~�����>B5T=�t!��,;���~�����n���)�tg��z����l�6_�B6���7�l��.�<lI���R����U���`�~�7u����)E���X��� KbFd���!�ݟ4(�#�KJ<�E+�[�a��D�3S�ڽ�	�K`��i���m�p>��u�G���tT�dx���%:��-��%������3u����~q!���詧�?���`��#g/��lm-@��0 0M�Y�j�7m&�Oᨘ�o>�[#�D@P馉6�B�����@��=</�m�{��E��^n^ce@`��(\�q�] zͬ?�l�@@�B��7��	�F����$p�h;Ë�
�#�`G���f����Q�ss�{�������f���
��h%7�٘[!>��kZ.��6�7&��Ϻ5���K.F���<�v�ׁ��Z��S4[_"�n�l <C�.��u���CV#��"�׍�C U|����W��/��J@�d�����B�͓���H�E�����+g)���O�_8��|�&S4������g&Ep�M�+_��d��)'�2�i'j����^9
+pAk]������P��q�x#���_���&�&��wU���K^Q���L�RwH=~�dj(�p�z"Μ�ڻ�V\��-  �௜fCL������tClӾ2C����c�FP�ט�����a¤�+�14*���Ӑ�������Z�8�8N��ŀ��Բ��G�J|��R�:����Q�18���f_U�["�4�u
eFȚJ����>i,�5&@T����.����S u���.yY�J�挸�Q<��[�o����A�i]�SH�5}��~JWa�P��Ӟ�Ǥ,G�~_>u�� 6���LP�;�FJ�7jc�<�=�
M��߷.A>S�>�E̰H�\�;�6Nź⳺}�`�.8�u%^���R��3uT\jLT�`J`���q7�^�x��K4�k�f�v���U�5�<kK1���1یR�����tZ)�ԏZ��jk�\�<������\�$�e��O� 8#���*v]��)͝��C�)Aÿ�	Ȋ"�o�,�&:��O�2�0T<����c(��a��X/�T��;ڲ%&*t�U��� 1ui�^�$:X��	z�bS�,LV��a��n��#�_���T^Y���F<��t��{!C���hՎ�,u�w�AL�϶��Hr��ݟ�C�q��AYeW*�Q�Bh��Хz�H$G�Y���~_��F�zO[�E�/4�c0Q��~XHk)Q�-��ׇ��JHU���պz�OIt]�[��@�X�)�޵{�A�x�?>�;�(�!��vD�1x�Ro*�5���d��{	���8��~��V�is�d��ŠN��H�/��4�u�z���}S�Z�g�.��I�z��~V��>�4$7l����mӲÚ�YDmrԔ/q�����3�O%�/7QO��2�� �l��-�< *T(��^R���)�{��l�G[ ���$#U�z΃x�M!����~C�������(�	�4[g=���kC� mK���S��=%F���� �l�K��kj��%�=+��bwsCK���y�7
7�3�P��ϡ�ͣU��u�++K$9�$�Y�4�x<s�h 8"���zn<���~_v�(ڭ
��[��,Hk2@ō;T*
{Ճی���$a��UΑzW��D��G���px�y'Vۺs�a��SO�g���#N��w?w�5��
X67��hE4X�{%���>���0D��<��)��V� ��Ě.ӏu�h�$Kw]EЗҸR�	�m�6B��`c���XV��[����]:$AR@�pAL�"�k��
��則�\h'$C4$h��$,��L�N\��d�.-���VףG�'�i�u�@_X�H�T�`l����oz	ܫ�����B(1��IJn	�2���P��ڝa�Yi�>��[ƿ?_,r`�Ȥ����l��g�,�P/ -�Ij�A�0J�H��Mp���U}�#��w{Ɩ��T:���a�i�B�S�&?�[����leUp��7,�3Ģ���f��I�=���Pn_���.?ǻY�dBG��.v��^�b]���fY�aZ��������ZK��~�\Y�܃��s����A��7�����3��`��*FyT�klT*��H��3��~��xЂf
[��]я#�l��.rƳ�鹔Y��?d�k�%��n0�!�һ�aZ�}Er~)`v�S؄�mN�8Y��/a��H4������xUT:wUح�Z�`n�l+k(	����]3B�!�!��M�&�b������c���\h�;�K\�7ÖTY��~}Wq�v���tq�C3y�&}j�*{��K*VjȚ���`s{4lI�N�;��9K�uV����I�ס.~��Az�W������x��	��Y�����:���K!�):�9{������0AS<z��{8��JŊ:dEF@�7�{B!���6��0��h��ĉ�ZM��s]����B$��ªȬ�o"/�F-�:St54���#�b��1�~1�"V68�)^��S+���bA"P�-Bn�p���\[�-�rn�Yq��e��l6W�0�Hw����*F��ЬW��^���1�BAkl�6A/
:�0��\3EO~$�l�8y#���<�Y�{U�fR@h~M'(����v|@��T���k	�\�hA��M�߃�v�ָ�rׄ��u�e�kQqB� ��S#jy�	���cCZ��[0�������r
{�E�@
�q���8���'`�Y�o�3ک���B��A��(Q$:�l��6<7w
_H�&��#	婑�BSl�>-�n.]4��H�6ǋH�q\mM�k�R ��̮lgN��Ǽ��p�"�0:��p6� ���?9=���Y�k����
y�x==<�9�6sۋ\�� Q��.A&�gZ�2�_��hj;%GB�C��|�||]�N@rj�{�M(�Xw��0zӏ�����L���O���]X*s�q	)K��8�o����u�R�W�Mt\]���c�b���P�(=P�VL`D�pc�?���R�|W�m� ��Q�M��ു�L�3��>r.�7�&3G�/#�L������6N�;|��6~zb��W��m�w����ԠR�hG�Ŗ�h�ؗ4�$E�ѣ*wZp l>.����B�������?����?5(��}$s��"��}n1��z�bK��3:�R���\�߉�r$G��
��XB��L�ӫ��/cT)A�WbWmr���A��.��
���Z�Wb�mwls��
/kí��ӵ�u�4]T>��R!�D�)��������$�
LO/���6���R�
˿<��cT�f���^uXY�@a�?��b��yC����O��8�����Ѥ=儶�]��?���?��<�*���q��%(��@��1�~,����
�Sdy8�#-��O���t�Z��cY������j�C9G��$բ�y8E����������!�-����&�X轞� ���0���>�J{��
��r�j ��;&2��_��o�	�"�$�!��[|���O�Y�˭7:���/�tQ͢���1�h��O�-y^���e��XWWf^��GjU���1���j>m/:�Bm��7�{/)W�Љ���C&N���J����\�$!��[f�o���w��Cd����8V8��{\�ل��� e*T����&ʣ��H��M�'��D�Z�=��c�<����c�-�3�EP�19#�@a���$���{�N�,��g���~I�ӡt]@H�s5.��xxa0�x]�ٞ�d�Z��D
ӥ���oD+�����К�c�`#-M���@���%"Y�aug�S��X���ZTH4 W��������c�2*Wg��ڳ�]��T���8\��B�����ߥ���b�&#��*�sk>�b�xC+i�9~�'���P�<ު7u�C���� �AΩ�s���1��T����^u���x�`0��������'�R念�UN�\Ra\���2�����s~�l�er�	�ULW��f����tؐ����}�0e��%4ݚ�|��ν��lN�Ah����W�-�o#��ը(�Y�A��]�7�:λ��D�ڏ����d��/������n���\�奝�f80ң/5KZg�-y��w��A������
�C ����]Lx�	tK&�b��α��f-TgΎ.��Q'3Nw���,C�$��g�ю��ȚW��1�[�Yʛf���w: ���s�3��`�d�Q���J�.�D���ѵ<�����,V	O�{�h���j��&LwCsTq}ZJt5�䊨�ߎ�jG�8�:%qp_��id:u(_����J��6]Y�>Sc#��%XO��k���!翂�i;ek�J%�b x��3��,�`�
�4�N��|�?C��F38�V�Ĝisյ
wEql5<(���x�H6~� pZ�%yf��5��ņS|4(Ѫ�b�?_ތi�֊P�e�%p�CHm������2=W/��@��~ƤFql�p�V�`�P� ��?���]�ot�X�%�>k�w��MBݎ)N���?�p˳�N�Uy��d���/��T�e)�����E����|�	T�@QbM��Xut�sxݎ����˰<������[Wv
�ZY�v]���D#=+w�=�rf�=8���&b���su8�!h�Ɨ���l��4m�@,�Bwu���* �]O���=��D&��m���t��͢ �l)�F�X#F��E���C���"~�J;7��u��v]��l�?�?@w�17wm��$�i1���Đ�OY���q*�G��!�b3���B!���p�%Z�NeD@��������+��H�݌���-�l���W��kZ��F]f2���2����xj�Ib�I �S���=xَ偣pW�9�n?	�6�q���>�X��TlG�w(7;o\��� F��)�ߴ�HU��?|R���f]��%H�����9��q�"v����xU��^���)D�QH�5�{t�4��Ptv��p�C�G�Z|a��4M�M8b̿��}3��ɵ���#ģo��B��@K:��܅K�/C�Z
�5��`99����X<V��?� T��\J�������6��q�-�]�*�2���c���z%e/���#�����"^s-�*"�vXa��+�6m��=�}�O^Nt �Z��X_�P�K���^�B��`�&B:��h~s�p�b���}"�lC3sz�?���b�ŌBa�F�K
h&O��B,$�y7��9ch����)�{b��؟|��	�t3��)M8�eZ�+Oa���aj��.�:QFf�,:�����M��C��,���m����[��U·Y'�2�X<�	��(6��u���1Mn�-����`��7�D��jh��f��)����_�r��}�T@�Iv5�̛�b�}�q�Cz�x ������%�"ׅv�u1[Hlc��5�*����8��6p�ٗ�mb�H)���z� �h:zL4q��Wu=�~Q��ۊ���MQ�DH��r���Z~~����rϵ�����P��B@��L�>��7u" �r\Hvc̓��m&Rh�8�T	�DLo�����I/u�M}$����"N6ge�J؅`� ۪�(�4��T�~�R��H��p��i.#�C|?f�DORe�"u����$"6 ��@�%�|I)V�i�̝{��T�&C��v�@jM	����z�����8敳1ۦp�g3�nX���=���t=_7�]7r,c��_zk`\f��5�1��3�s��j"m[����cp7TQD����5��F+��F4ED�#Q.����!Kn�����9��R�@�_�d�e�����l�7�΄�&<��r�G'��������B6��0Ƚ��@�Cj�����:�!�[��>�.7}�5"[��mt�ٗ���B��V�U�pO�-�ӕ�[��>�s��|�S3�C8Q^��L��d�Ԯ�=�UՏ��>��
k�Z�����w�IG[x����F0�,��Jg�>^C¡LbCQىE��w��H9�xM�M�M�y�*���6��������% ����(C$n��A��DuY�^��y0�� x-���L��#F�s���n��@�p�Z\M$���LN[��s�����}�f�g���$q�a�3l�C�~sh/�V���7��B�e����R��"gL �,���p�	�Kp�?��y~���oQ0v|D�("�uDhl3]���~n�%�}j�m�ќL�����IG�d�����3o ���4G�c�wݿs��K��/�0�5��E�?K�`��`�p�N3��4��U{e����w����J�����Z���e����
��
�����>���:�o�2�x�2��=R�:e�*M����~'n����DJ-1���ʡuc���a=��53G�f}��A�����sA����uΘ$���uf�DL��|���ڊS�-��iI�&׍��S�Og�����_n��]Iʃa��Ǻ�>TTߌ�Lp�+$�lG�<`���@=h�ܛ�%�Ěגc�����>a:o�!��P5s���hv����Iry����?�-i����PH�G��6�����Y*�(Q��O�lfuPѻ��rE��P��%p�=X�Z��&]c�y�rɊ~�/҄�O����H�I:�CU��S���	�Ԋ�T%��Y�C&��T�w��ם S�/�Zs^Ѕ���Vd���������"�U��v@���a�e��5+����9T��%���bbP����0&R��tp��ww �^���u�]�����	7�4+
g����m�P�Gn�V���5F�~�0r�`\pE�N�V�����:hס�|��0��`���I=Vr���=Q"��Mym[��|����f@�-�4q#��Y����B�>��G[���Bq8�Q�\ö���>�v t��^���<�%-ꋓ��@1���k�)&�_.������)�i�?��*I�䩹�ͫuB٤���!}�ŸO���_� ��>׺�SY+x�	+u\�]`�`̮��1���}:�@N��zk�<���w1�(��5�N�>��&���~1�Ѩ�ܲ���:F����Ǥ:̏-m��, ���sdL>����g$��)���pTM�
ƅu�?�sp<�p�J��p��V�+-�JǕ5.��*�;x�V%��}v��MB~�2��R6�ހ�^����N��C:��J#���l4�Y�����l�����Y��΂��d
�K�`�~��
��^Ps�������N�4T3�m��c�����:��R��h(Ҭ?7��%�������j���Ƞ�[��\uBZ�ٞ�����Q�\nu��6BR��֝��&�kX02�NT�y���+yb����=?�F���Tt�}\�����X���	�Yq�R~C�v�{`~��-	�c:��z����w�s�b�en��*
QaU��u��=��6Ϝ֣u�
a,��gjU���;C\9f��)1�Y&	�E�g.7��?h@^5	}��..<�N�P�r}ƒ'�I�d"��ۆv��kTl��s�bGga�1�������l�1W��2��<����鷨O9n^x#��{��J �<�`8G�1rG�Ђ���aE��O��V�)t��e�����{�(����u��t��zB��JQB,�#T3�'��M�vr"����`ɋ��!AR n�O�^Չ��f�J�b7M��j?����T/��������5į$ƿӾ�z���W\T�Kג�����qW�P�h�/�`��^�A�a��0���AGF�I�6ɼ� �I#�\�˰Z�6\��6��:�n�,L)�H�b3�$(D6�����Gh��P�t�X���F^
+�Y%r���W�L}CF�z�ef��G!܇/��P�W�x_垻����o�rՊ5s6B�\1�Ov5U�B&B⟨�R#�GWc�z���{s���Fq�����b&���	�3�����h6jɷe~D�7\�B}$�6��Z��ꉾä�S�漣j��U3#r�X:���+h���>6�`襤H:�9iІl�Wh̜��"��҂]�u����h`ЬD�\M����2��[�4̊�[�}e �Ί(2H�+��-��|��+,��3�diش�.Ϳ��y��S���U5��&�y� b��k@�(��|a�<m��S>I�R˧�>"6G
�(9��t��$G�	r��3��T�8_�����H)�ۄߺ�İ�Q���
M�@%j�>/������#u� �O���u�}YT�~��x���P�\h,�>:2,�(g�EvMЅӆ^���� (k�^�#A��m�G��3�����?x�b�?R�8�Q�c�]��gL��E�#,��a�ש��bȃx�؟�'���� �UyW'A*ި�+o��FR\Y9Au3���2,$��v˦����kp����N��g�@��ݍ�A�Q@�q�;��&LAis:������k������c���4�f���@d8�E?dwlɴ���o [���"�t�#��}�1~(76�s4�	�(��`�^^ C�)B�͋��l���{�{�9��:N�x���q`�����?�u����'�� i�L������/P��7�`9�.k�G��-zt�C��:��=��[_�Q��)���w��.��2���H���ED������\�>���g0�S��>����$�4ʢn_�ߪl��Ps����;�{�,�"3�
遫)��\H�+h,��<��#t3�����:x��o�Ho��8���V�}���	����*��r9��Bߺ���f?�D7 ��Y'��4�O.]ϰ��<�Ȫ���R�oc�R;<���W
k����7|A@0N���o[�X��W�g7�
�x�������珌|�a:{�D��L�k��+�hgc�-���D#v�����iӈ�7¢���U[�d+*�Q'�Ph��p�m,��ӝ���i��d�~`Ge�:@��+=��9��(؅�'���Ye<Ž\tX6GR��X>��K ?t�}�vR4FN�U(��@S���蕁�	�ά�.�E$s�c�۽��7)�&ɸN���Хg�A�R:n�S���EJ�����j�HNؔ�%HXob���G��;
-����ґ�uc�L�z ukYL;j\oՀ@S���� �	�� ,�c`D����Zt((4vB�����˻�B�ů�b=m�j�6��(͜r(?BT�(�9/�+d�G}/���8n��B<V�wh�G�V���/�;����j���].K��ِs���v�æ�R�@Z"�:��Lװ�1�/��� ��=/}�5hD��JI
6�����)�ӷO��}J���R��/L�D7o%���MOOuo���1R���O[&}Z�X�>�oX[	?w.�E�)Q���l~�4��b܉��f��U"{'�`Ӱ1	�=�Y_~$v�f�gƑ��J�����(�d��b`��^<P$1e�w�t3��N���v+��`+����59ν���E��*W�]�����,W���b�m�cCbɛ���	mU6�"��|�����&�E��:������p���j*((�<�;��3����s�ϙ��l�XW5���d���Db��F�0い����$&�J��?�=Z��c�;���O�s����r�y)������\�����P0؊�k�z���Eݕ����!��UP���4�l��43D�6���7ؕ-·h]�y�0,`Ӥv�x�6���"|^=�iQ��[1^�/�mP{V7u<�z�`b�~��̸Jt���K�5�羇���N!���d��D�	_�5A�g�ijPt��x�^����2����لToa��T�s�,A#QI�s�8nu�4���/\Hg��]HC��u�S;������#G�b�^�e* �!�k��tm���tl���(:��6f�5��w<��"�^������.+'C��������+f1?����H�	]���T9�9�f+��h؋��3�/�m$�A0Uߏh��<b��m���8GY|W���y�)�5�~���k�~������]M;�] <G��_������3��gwK��Zm��u���.߂d`��!�O�)^�!�_��R� ���P���q$��u��g&��Rg� ;�ZF�!���D�����W���x����
c7z����_A�i@P�6�&��D�zE}��#�-��z%2[�TyHT�%�%�k�xn���;!�0�`p��	H�! ��+ag.'��TC����� ���O0�r����/q[9��Z]�����i��eږ���鉆� w��gQ�j���:}&�r�̩X[�y�[o�\��H���
e�:>��җI�+������_�{�b�E�'L��*f�z�8��H�O��,�������-bH\�n�HJ�$N��&]�O��vҸ�@n��K/�;���wgb�����5{'cc�~�ɟ��?DE��"�ĝ>��ѡC;��t��Y�6�1g+�$?��ږ�o�˧��� ެ+5N�U�S�8G�Ϟ�	ŗŏ��$����Z�&/H�a����U����xU��8�@�e(��$��kx��q��DO�0x�J��%P���}jùL�F�U!e�Ge���T2�o�|�u����C�!�k�T`������I��Y7F���G��ZjwE����{8����;�X�w�]�U�,�q�/hT���1��U2�V���a�5G]	^����༞��6Y�HĢ��׫���"��,�| 	e���ꨃ���gxL���G�i��� ��d�<���g�MӴ��M�{Q� 
"A;X�N�T�
?~G�s-W�v*��{%9 �T��%�j��_l���?�x�`��1�`w�&
�qN��5xΪ[�����/�	�,�8/��6�-3�2�⒍`�o�x�&���o|��ȃ,A�����`�����o��iܗ�
���UL�b�7	�3#b!a<�C	�0��anpN�����
�HL�
n�O��_�
p`��O׭2n�,j����%H�Or��%`/.g�Kg�G�P�8{o�z9���y8n�w���Z-(B��]���J���`M��=%�~5�@�q���3��}�4�G!���n�oM��SY�?v�(?�����@tj��i, NqnQ�6z+������Rݻ����+�Q'��4��!v֏�,<5$2`�;;�E#���!B=V?�h��P�P���J��|�]u����-{�zH�X)��m���o��%-���hG�����c�WY`�l@�\���u��g��NV���m��.|#���GC�8��A�J�S��+1���Yf@����DN�ǿJ��������q�J�I���A?r(%������ 1ɐӻwK!�р�=3c4;���)նKT�k��|hR�{3�~�6�V�c9Š��������#.eH·V;�&e��@=퀾w�%�O�Tx���*���@O�ú����1և&m�y�{L�`;:����U�bF7�����c��G,�!Li#�� ��>xO�=�pK��
�{K�UUm��}��s��B��(��'�4.۹_,x�S���[��!+Q���k*�WضPV�F�<����lN��t�����t��!f�1E }����)�=3�)���A���h}��&AC%�u�hM��l�����cJ�=ͣ#ºo���<��@Q�#x��ӷAd��{RmT��@?��Ź`
���΢�#~1f�t�mx�ޤ�Y�zu�
p�_@+�7q9�J�����*�/�.����#���t���*0V��>j����a�������ֿE8F�Cf���0 ���H�M�k^��}>������4���_�@zx�'�_"�c�i�Q�Ð��6�G՞kDT��{#9�����9�G�$�l�Ymk	^`O�����m��sT��Yߗ�E���f��V��� )k�2���U�H�.��m��I5�1���Ѓo���-[Odt}K*����)�Xcp������
�Zc%�1%��RV[Hٸ�:��65�xbM�ɳQ� $0g�?ռJ3)���%���q^��8��{-@Djge�wE�bPi��uN���"[ǢP��qON[x'Ph�%0AR�v ���䝍���>�ӯ3���2]*G�yX��ao��#��'}�� ��p�U�����ݪn=lB�S#����1R���f�������Pr�ɳ�*S� �:AӤ>JYg��J�� =��ђW\Ȼ�Ђ�4:���➕
��|��&(D�<<T�~MΔW9���#�8�d��ZTj��×�Q��=GI�>�`�i}�/�/�A�Ra)q��W>�b{`�� һ#I���a�6J�=!��Մ�>����;K���&��b�3�A��2b�nϦ�+j���+h���O,R��. ���J������ _�=L6;<}��x�yBko6�E�<3Q�+\��HL�?"}p��~S*����LI�(�^�NI"-�\��#�~m�כC4i��k�`���Q7~� �����Spn�UI��=�"��dj��YM�ꢪL��9wΛK�.����4��D�!�v-G�L�:e�6�о-������}�@�@Y�Ov/Ag���ƴ����?Nsk�bĉ�OD�vҚ\�rA��d4�	$��5<���ٿn��;��}p�]�`N�uU<��ڷ�C�
U����� M�36%(8'�\Uj�b���:�_ў�YmF�Q���j�X �$��Q�>���v>�]�	O���R�'!x��զAX��q�ظ�V���-U�K[��ь
�c"��%�$L�*Zrʤ��;���$��2Z19h�Q��q�/�A���A�Z��3�� v�.+�M�߁ק<G�֊��QoJ��[��I�Y��X�g7�t�O%���	Ca��Q�m��g�D�*���x���r���,�&V�5�+�w*+�\�m�מ�e�0�c��^>9k?�W�^>!�I�߭u$vk�n�ylܜ��tK)�<@�>h�l9'���0)��Mr$��nֲ�q�}n8�kt�g$MX��F���\"ۦ�']�O̕�7�O�qV��n�{�Y�.|*��hX��4	����eٻ����ʠ������ꥹ�8ĸ�o��*!���%:�8 ��>5�r��$�a�3 *�娀?	��� ��:tc23I�b*j��õu��
T-Sq�&�ˆ(�&�Ì�0B�X����`��#�qym�y���gx��\���T� �� �	Ð�Ğ	�NE�.�����F�ǳ�%��ۊ� ��1M�ו��[�]8���3�[P�l�����c��e_5~�o���nT�� ���G"k5!�K&%�¡j�ډ���&`V���A ��!��\׈Ξ& �h�E6�E��5u<�*A�fOj���z1,���q˗�y�ݑ��}y*��b�
N�b#/̡�(����;g\e��Č���%���O:�;�s3��1�j��F�"o����ZYM�Za�{
ڢ�t^?�O�`aF�ѥ�x>!q�r�s�w�D�+�X�znuSmj:����7*Vpۅ��8�e�\�f0�S9�%�VnW
�3�'ԕ���j�k��������b����XXk�����^����i:�ڞٹ<��� <d�6_
����̒�k��8s�:L��Uf�][ܾ�Vs�������&3����|bS�m����Q/�����	����ݝ?g֍�7vm5�ڏ��s�t�qg�}4h�>����)�l`��O�gAx����@�m���7�y�O#aZ�W�[W���>7xiҝ,����4�Ԇ�r l�{�"����e[����8�I2%H��������a�z��8~M��c�3]]Qɂ����"���vm��b�k_66E*�6s0|��I�փ#��|P䀵is�`��@�����7E�݃���c����6l<�hK)�8��	&�kU:-�9,4$�)�Ox��X�d@�oW��N������h,�e>Q��%j��S��	�5`!�܍d� ���
'A� �2��q���q��.u������b���H�I�b�2)�X>�������_xB4s��H�N��t{հ$���b�t�/,M��h5Gi�_0 M���nA�<�5D:�� �MO�d8v��6����C`���
)
��Sj���֩'��-���`��N}����`���ȹ�`�7���w�q��?'�9ی��R�!��R�o D��f0Y�"r�1��-�o9����-�[k{�'_wC�����o��<����lLu��;浡�����p.�]���Y��̊�2�FS�`| �o*1�H�&e�E/45��ft��'�gg��z�:���o]��d�B�� k�k��#S����i��'�g��Ԟ5~���uѺw�����g�(�E6%�r +�+�8�K�]�j�O]^4���fv-f�#���=�o�h2n�<�A_`n��H����X�D�Swؓ:1H-��1�h�љ�Ɩi�-����J��� YC���dT���'�g's��G���@6�I�md�{WW$�jG��'_\RE�җ+�Խ�V�5�m������`j��:����-.�Ԑ*w��d�$0� �����b�������pL�Q�
�pBO�g�a+��G#U2�QL[%ܯX�cK��K>�}æg�Ķl��?|-P|�@R-��71j���A7}�w��qC��tv���܆ڒ���U��m����t�aꡘ��PJ��Z�U���e;��{��5H���I +�C��c��q����0I�q: B�N#�*������n�J>�# �#CY���T�7(�@����l@�9�r�gv!	K{��g�]��K��.!G-�D#Un�	��(/�I���=C�\����p����|��ߢ �]�Nہ6p�J�p����V�pZV9�62L�C
e/�[�����Š'�R�t�ރD(��ݐ�bpu����N��#38�����P�i��u��*��d�=���9u 4�&�nWq����[U�e�2z�-�[���/�c� ���_����IG�@�(:�+����^�C_$�,ޕs��y�og�t�~�]rZ� ��jjH'�Al[
B��zi��4��^8fD:D�|q-b�����׀�S�=�c��Y!�/s6)��k�XY5%������a�*T�x>��[V�����xx��x��^U��m�ZV�-a	��!�����o��:!U]��6�И�� ����t���@�&�QT��4�w���1�F�~W���|�*�h$0>jV�W�y琶/2�����ִp��r/�Y�Ǐ\����2h��K�[v|�;45E..y&��ԩ�^yz퍲��hnGX�B�޶Tܵf;�Rg�f���衤�]��f�+�Q����q�������+,|E{����׀�����cG\�~x\[X$"6�'���[�&-�N��R�FTirc�I7�[BT\��ߜZ2����9s�To�ay@<	�F?�9P-�HpV�!YM.��l�� �οq���<585N��y���N�܉�m�h�|!�����v��X��1s���'���WJE��ȹa�2��Fۮ&X���*�Kݽ��#{7VF�ƨ_1ϔ��.�����kX̷�_�m����
Ad��K�L�_13:dE��!l~6���b�DB����>j[H�h����}�E|���sf8���x��n!�غ�F}��mDw�soU���J;�n�����ص�i����!��� ��َ�*u�u��Ҽ��O�R��x��]|F^��%j��7:8��A�+q�w2��6�%���5/m:�Y�1A�<��13�=�i~B�׵/k�� �
�t��Rl�&0��f<Ìα��kMr�N�W��i5����j�ni����Y���i���(���+����Q�h�i��� /���Á4\&|G{fY�WTҋ�!0+,8!x�q�m��R1�ϻ����ӽ�|�b~�۱ۙGCWu�%��}�>
������Q����vJY	W���m�»�)�����ծ,�k�e����7]Hg�<($n ����Uڸ�����!%�"�F���я�Xx�{���F��6�R	F��E&A�����,f;��/7�/?��� �Բ�ٰ���/�)�~!��r8Ұ_ljc�-1�{$p�T��̸҆D߂��GQZ���_�WA�Qhh���U2��pS�=?d�Ѻ�<��<�5�
�F�߉�E[�o�Y�^YB|Zy�v�Pɚ��9�|�'�HXU�5	��'���.>0_œ��C��9(W���0�?�>����8�<.P1�e�)yѝ��s"?���`Z���ڠ;l��NU脶�?��c���𭣋븕��2y��)����E8"�X�{�|��#KJp���5�/$kf?Ηp'&��V:+\�]��������n��)�/�0G�g��N�4��Ϟ���W��*Y``(y򥳸J 6N�y��#k���V[,Q@����NJ0v:%�q�	�냅?0+�.�.6��}T'��Q���e.��K���q� �gg|��Ѹ�O��P=���q����E�*����qj̓%��H��9iU��#�D�]�gB8C�n9$�V!��C�:F�a=�Q~sGd,^��ħz��:�g"O�@�f�Y��Z;V�J�{��#�H��
�=�Jk&@��"i$�{Jź(>�M�K5.���Nk
w�Zt���������m�������^4���3��fȼ�K���PC��L��rH�ᙳ�d��G�q\�j̦�gE�oȨmQMF�%�m��V�J������XRn���K!����sx@.T	f/�a�� �W-mMO\��Y�O����6���2�^aV���Nu�%?K�M�;����#۞��������]� B�k���8�ƅT�K�Гv��.&�2[`U_=D�(H
�Mb�`p;�5�"���-�C(��辅{��Y�cɈ3b�A�V��p������ê
1eV'E�	�/�.��|s؈�`��~X֒�/$p�'T�ȫ�$��Q���el^no�
�Ow�Q���T,�O��S�(�`I4�w�0���*�=ֳ;�R����r<�P{����C�K�딕��>ɿr�����z���e����HF�q��R������y_�A8��?�p�󥮘C}��[IQ��Js�<'2݇�d��y����F9��ǈ�h��e4�h�>Eh���mkwvxz����� *cL֯�E��av��!��F #�V�'�=�5L�8�k����0�|,%F\�	O"��d��l��+���p��mאQ6�:7}�o��[*�P��qA ��k�|�̅{�^	��|�/�S���q���wo�m}OZl>�}Ȥ�zw^/�� m�t�j�ʔ
���,"���8���F)���QI�f� <X�%���>'��yT�p�OM���Y��f�Y۹��Z{�- b�F��Mɬ���},��K��$	���&F�h)=�ŀ��^���F���ѥs�˄�S$�_O�ϫ�Hq�)�ö�ߟ�����	��ۦW�����J���_]@\�/`U�;�����q�m߈�{ErD�9�|���ɘ�{Ֆ���+�۞���JP��[lL4�V�1P�pC���r�&���Đ�8���U�A?�}	 ��drgq➻*P�2l��(H�N�E�F�ġ�[ �R�~����{�}�&�C�8��`����Mt�M�
���+S�{/E��8fo��58f��S��3z�c1�"���<�o�0�9�:dN~�!�|/y�'�(CHq�
��N��\ؑ��J������b3��%�M'���,�gH�m� �@6�T�&�k0r`�Pg �x�[�s3����A�����k�;�`�+�2�!/UX3}ծ��8(u#��h�H��q� .{Uզr��=��G船.-D].��tk����@z�m�p����"4P9-��? 0�����>�*�[��q�M^��p'}
�v(|�yiz��M�@@��Fol`����<U(ria�=A
Cc_�K�g�`]���%������Y�V\:��M���ٜC��/�!���#�Q/�Ddn�3�v�qh��k�w6'�Sw:�&��*5{#jp�7�|�ߙ�<�����>�����{����_5��`���q��t(ی��T;`��,So1���G1�1��e���� M'Y�M���(I	�-vtz�JG�V_��qC���ؽ� ���~^���(W�Ý�`:E��o�yt'Z���;-�.X<cC5�H�Z� ��k�)%�F�,��^�B�/I�Y;�=�����#��"L<���ҀX@�b\F���{�����1FnA}s��XNf?�4���X�rXVg�R���V;E��>{1@8�� //�9�5�M�e!��D@�s�d���_�؎=�w���R�@ݯ�Q�8�B57W��&8���'c0E�6�b�OD��$�qĔ�R��ˣT ȹ2m:i1���}��.�x�$���Us�'��g�
�w=o��W�S�,r�� �x�]N⒩������	N?�W�F�5�X2��d�U 5���ny���-;�w���u�wvzv�R�(z`(�*�3�N9��H�4��/�����M��΃H:<��ZQ�Y��$hyjd�fJ�Q@m��[%�v���z���r�%�Gݎ�P �W^�a�9˃u�M�+��V>0'A��X�E�����yq)XB/�3�c�Z�:U5�3)p12�����8�mhv��ƖK-�(� �x�����@T�n8ɸ=Xy��[��0�Odc`�sod5z�w|/�VU����AV׷�]
�2}v'^�4 ����P[�	e���I2��6��/Yjϡc��X�`�઺���J�0,�,\Y<qpV���r�A���A��$�ȇֆ�x��S���mO�*j�9��sW������~֟��.�l��s%Px?S���}���F�V���p���Q�z'Q�x'��o��Y%|�Y�s��IPP%DnG�%o�]aZx��ǃ�w�'mb���,����"����h<!C���inKM���P�2s���0a�%�Li�p�8<6�</*_�i����F��l���K2q�h������ ������=Q�aIv.0`7���_�<�w���J��!-����������%�e�0�8FV�!X���ԽWI~&b������OaT1���)��j@�[�'DDt�5��|�w��䡀�0��{�g��G�{1{ �ˎ���>��mK򪶹G���FǱ��0��W��J��d��<�u,t����lfH�8�Cz�S�#�*mvڰ�'��B~��`�ԙ��~��b�v/��}�m�./���Nᣱ�tt5�H�O��csG�t�R�%��QQ�8T�ܫT� !���ޭ`=����ٓ@��z����ƫF�VX���ʆ�#_χ��QGXAk���r��c�-��o4V�k��cd��X�u��**w�jE�Q��W���������w+*
gM����� n���%�j���� ?�� �2ÄBA�
���j�.��?B(����^�6ڐ�����)yh$.tg�ӻө��٦�1��4�#nh�7�o-�C�_A�j|G�dU�Fa�}P[P!�$�����r�0r���T��N����a3��>�<�^�9z��Z)'D��r"
 Y�B�15,!T��'(��I��XJ'��ݡ�~�����BԎ�&���c�6�4nTp�V3�YPGى^��: ��N`q���Tv�ˀG��_�]�0�� ����j���M�ݿ��P,y��Ŀ���i
q4}�8xN�&���_��٢��y6�+�>���-Yԅܤ���O��j*B�n�p�+&Zז�X��op3*��E:�a\\�����b���.�X���L���yυ���_d�*0��p:�(�U�n�7v�]�Snc��T�����؁�@IyӺp�S ����ud���$��,ӦS�i.�S����^SM0����n�w��e�wes.�c	����r<�	�!)9�PVNx�,�[�e�������}�}�3mJ�n�ϯ)is�-��%���~W�| ��_-$dڻ�NlAʤ)�aw�N\hv�ͯ�ħ�ݫ )<��±�
�}ɤ�m�c}h*��>:�m��S�g�4�1���jHe�̟�MFnO��|T'ƾ�����K�6;=����0��n���&\�Q�����"��\�}���U��Z�>��5�0�����s"�rZ����ç���p#�,��̉�rS�x�S�q�Տwu�g�<�[������%3�Sa�i����=l�n��e���e��k(�?�ٓ��/<�Ym�5g"̐#-n8c`��R����V��T�o�F���7S U��9���C�>�oRP��΀{Ĳ���3�ߦJS��{�u��}v���h*]@���%�'-MU����$�^2��\���^^֥�b�8��7+^�͛*��*�2��h�B������D����Ч�Ā��/��4 Ǚ�;�N�A�U����IOb�9#C���dV�_�ft͂}Ŧ��DA7����t��/rl%X���`�Z<�ђ��#*ʊv��5�G�ހa�"�l?����vC��k�c����_]�b�)Jcel�ɑ�?(��#���gQ�`�J�����O�|B�3I��Gr�__�yq�!���.{C��,y��K��(|F�����!�>)�3*`ל!��*h�mh������p������ۇ�pRp�K�����L�5�V���E��C69w#�K�_i��|5�D��^K%�q@a꣙��.��-�_�R;6ތQ��md�F�^e��$�fw��D��93n�j���R8��ʌ������Z�bM�S��'��AS��|;ɴ��(╇M�kӹ�㩈�u���������0�/�nn3ر���/��lq�F���Up,!١�=�,�C��6���Á�K�5j�iXcP�_ o�zЯu�� '��Ϻe�<��;x�sҌ>O��D�_D�`�)q�&�Ն���q��}�,���
3���o�{�c� ���щ,���}I`�t�A\e���<yC��������¬8/ �p�*Y�}l-w�7��鸄#H�q\��V��~V�{�µ����]Uw�L�܎ (�5�]�F�ƥh~�
����4Ѐ霎
��(�-�2{��$��9��,�Im��bM���m��(��i��#�4�Fh�:\`��m#��������i>&�L���[�/��X�YSKP��p}C��j`��:�gD��k�"V83�ݰ�Z���.�5����RHv
?H}�y?�>�/�X{�zbQ}���xko����C�x_H�����@��i)�:8����Ɂ��g��}��/�T���!���=M��N�	+����+~�P5r-�n�Ժ�0��ۙ�L�J�f�(�%{{ ,��0��W�A�[=K�:���d`.]Nx�]�A��X)�˒d�'����}fP���Hߒ�M��>��W���b<��9��N)��V�0�LU^it����ş��3�.�t����(H�s��X?��R����8�:b�1�����q�	��H�?s�y�J�-�ޓ:ľs���#�J�ܹ�kF+W�m�e51�� ҋm�(@�!��
�a�~2�%�J/��7���+N7p�z�5|�)���졉�qE4�!շ�E殂�^gM狑)HB�DPDO��>�x��+�BU>7ڲ*|
L���ؖS��4B�a�So��c�֪�Ӻ��"����;��#}[Z�lD$�~!��%��r��=m�:]P|�S�#�[>,[�gMb3�ƚr�"(r��0�|��[>���Ql$��f��s����մ|.��Y6�
eޗ.�6�������
�'oG���W�#G}A����XRM�LW��R|�<���I~[9X"� h���$��l�DǢ�	B�*����[<%���܂�GNTH\��r�/�.ϟal����q�%a��!5���`V30Ol����e��Y���}�E�)�+p����:�SI��UwHB뺆@�
y�:1
�6����a@~o�̨|ĔЗb���^�Կ p�'%\�JBޤɒyi/Z�살&� ���Nd
J)
��[�8����%7���?�ɞP��_�C0��vR��E��d��$�q3*i�������ׂ?8���P	MQrj��Iwִ���F r����+Eڡ��!����1�r�`k��g.C��7�T�E$��M�_���A���7k�#4��䬔��7�3BE��_{�I��-����$�9۝�wvI�h�T����^v�I�����"�է�KR��p�6=�B9�37����#2��hӏ�^�H�~Ƅ �?�IYRpCS�:�XF"$ڤ�s#f3�!� ��N	̹1|W��~����<�_��fqYn�g�j���M\5ƫ��TЦ�L�W?=I��n�`��n�2�j���r�ǥ�t���X4�����c��TiCڽ	����	r���qT��@�'~4�����E �L#�� �	���,t"�e"�"�Ü9YgGsE� V�r��f�eD���~#.n��8Q=Y֙Xxu��c�,���Wd]�
n�^�y0AeO%"�Q�:��_�b�w�
�S��γ�*(fcP�)>�I_�dH1]I*[�P!6�<������oȪ����&NfZ%�Ӄ,��:S�O���5/o}�T(�ۧ�3IT�o��r�2B�x��H�����>3oVE��)�u ͓� [g�q�%O�iFT�Co.CF2�!�fGBm�4�p��?���n���i,'�:`~�K���?�J=~����	�`�K(ဃ`VaZ8&����R>�.9pLe�1$���P!���Z��a�,)^��)��B��bD�fS�"��ot&L}��z��5�pោ�&nSFv�E�Ǣ��`I�� ���Q��������Y��2��g"cq>�S���GV*�k�_����¿�.�㒰H�w���=
-BG+�1��Kfu!�Q�l���gT������t�q0ۍe��ȴ�]�>� ���2��pl�~�1N{AZu2�.H�:b�2Ӛ��v�գ�����˗	�2�Mm�7.�Y����l�l@���Gd�f�%�Hm>�|f0K�>�ㅷzt	��^9z����
2_�����I�ۢ�ة
��)Q��A���7�O;�l!K��'O~+ل	V��xmr�*�bİٙ\��~����V>���u�ڳL�	�7�W�H�o��-��`�5I"Ywܘ5�F�8��u�1^f=9�� eN,��	�R�+�U���R��N�sG�'�����,�ˋ{B�n�:L`����ec���'����K��ve�8%��q-bʟ�{.װ��]/�`��P�����T��I=H���\F��c�a��\ �rC��W,&3��l
`m�J�k��&�����[��N"�s^t�py�,���W(���s�g�Q��	r7�i�0SS��_dܯ}�W5��&)u|����ɴ-���j��������C�{��ω��,~ߛ�r�x�Z*�uR���U��i�1a��Z�G\K������i�̸�X���VJ����fN2�ta���2J�y2l���:,H�e?����m�s��=��<�*��0.[ƙ��Њe���x���_t	$��/���O�`�>� ���:{ � �#���O9�_6�Z�_�o��i�=&K6���[
�������S�Ѱ���N������TG���\���)�xݩ_ �2���BV�H0��s.Ra�g�v���M='�}��OֻX���@��Me�z�o�y�/�0�js��uE�������퇟P��_���h���C/�P#X�L���%j�q�M �$O�	.�:��!�W2k��*9���7~!x�?n�N-�|[�d���';hܜvx>5����s��a�#��-��{F�N��"�h�[]�!�ޥE��ذK��3��5���,/7R<lip��[pzg��'O�i+a����@�[&��bǽ��f$Gs��A�U�P��HD�=�O�5x��l�g���++�sVP>�4r4���/����]ꈭ���uþZ�����]Y�:�;�j��1[���۳E�i���f���;m��D��>�3g��诞���o��M'�ƍ�ͯ� ��ߌ�g���4Q9(<�na�aQK���[#��a�/"�����j;E����[�I���[`a��~�ӿ ����Oᨮ�5�yt�<ᷰcO�Q ��T�3��:��[8?_��8���$�va\j�{��0�@��%u_Y�
�4��\��T�����B�5�&ֹY �\�@���+'�Z�/bO�\JFt�2u:W���&��UjR�c.���X=7�8r���[�V�ӑ�*��ӞX�[�O�%̜x��;ke��
��:�ء-�W&��ZFT!���pSw�D�aݾ�R��'٫ ӑXzy^�H!2�▢���F�{�F����%��[\���&�����x���1�O3a�?�|�h&�\����ȡFN����|���|B���;y���ԩ%,����Xm�B+�m��8q^����e;�4��41$��/I~x~�K.B���D�N�Y�@S���UO�v٫����������B��w�p����S"Zo�+#j���^�4�VZ#X0uOak�#HNEǏ����� 8��XO;��x�(2>fΌ\�s�ٵ.ҁrB�CI/���|��E�ͣ��|F�O=f�VUc��M�^�w?���и	��]���.�?�������[�P�LǏ��+���:s¢/�x����9�t��.��%N(� �+ ������c��Fz���`U�z4QѰP�T�3h�N��*m��+L�*�bCۭ\�`�)��t����(~�Hmz=�{��+�߹�#����Ǻ�F�%�I��Be�	tK�O#âg�k{�Y�����ng� j�VM��U��"�)~��a��Aʏ4/Rf�>f�����
�Q �����f��pi�(����;Ѥ�Kl���n �������,D�~�H� `F̭�XxEN�Ւ� �%�1+���6���o�����S��ԑ����"^X���J攦����WAd՜R�?���5�T�氢2���fWgA��7E�xe^�6c/no3�L?i���K�27Q#�s��}�?��kǵ����Y�Nܝ�������9���FXMo]���ʌQca�0W�4��I�hʵ���T�>��Xd����b
T�|#�0���6�s
��g ��|�'���!�?���?��S�ˤ{mi�~�oƀ�J�]d��ǑS��c�*�1����>�@F�GQؔ�:�����Y���>��E4j�w2�3sD��@L��O�W��(Ƌ�I��;-
�+�NUO�t�X��'A�<F�����6��[�}@���X1��ѐ��m���V�-;c�����^d\�\b����������F݋3���i��Yhw�k{��� ����ʷ(�|%�D�jA���̛����O�?� 9��%����R�5�!�����#⥦�Fx���T�P�/�aJsL�s��m���/,u(~CF���Q�"/�ߊ�� ~�ݢd����g~�u���
�!�<����W|0jHS��^}����]���$;2=�Hش�4�%��T!���w�f.tSz�KQ�����F�k����2�B_��#�̬<�Y:�'�ZK��+�W.(̈́� � =
#�p����[&<VQ�x6�hVP��\L�.����@n���+D�?pnc��+KK���I�H�w8��-*��f�z/X������x�%���|� ��QDc��]�Be4W�f��V��ퟞ��[���{�\��wyAb�����5���`�v�\���L��i=Z/��]����NB�Q| �uͩO�S�W������y���q���t�����k1u��f�W!{�.��L8�'a�S�ax!���i|;��a}Ũk��P���u~зE��Zc�1rv>�Rz�_lJQvƮ;��Pkͤ��/�|��G�}=�گT�W�_���F�L�R�{�|$�8`S����������3W�oI6˖ U-�����@lqwz��R�HwF���K%^ Q���R�mJϤ��2��Ras2�P�e�m�E\�Ȩl�c����[rz<H4��%)$��N	.O�(aV5TWL��+�� ��,>0LӘ��u�7�Q�!.@S��MD��їxܪO�u�K⨎K�Y�-xy^�$mX'��U�bߎZ.��l9d�䞼��ݦ��-{)�]͋$et8(�f�*�B7���=�d�r�F�
d�h�4���ࢗ]}�����ӭͯ��K�\��1<%]��T�Wv�	���A:|�d�#�hJƦ�kw�xy���6���ϯ�H{�)�������M"'�X@�"F�%��K_u���
"wX���8]�!
Wq�굱������^�ONbv�ZMzm�����|����J9!?����	[$-V쏄S�;��G0f4J�u*��x�of� ��Yf�@g��r�?
�X/>�����#���m-�}�w�����K]�>cܾ��l-��$t�mځ	�dT"R���J�}{�3�T{l�,�_����U	���6F/���C6�?�AM�oN�s��@�B52�ew�m��$B�?�ʩVR�b\�K�!L�&p��g�K� �&{:��Gc`wQ���(W���x��SW�JK_���$��O�ۛr��i)S��RO��7�:z��^���ہ:��~�9B�8%r�Z&�,�6�+�QŔj7��iC�sF�ˑ0�(�9-]�4/�Ìo��I�t�G�qS"��=�d]&4��0u���xÐ��H7�>Ap��������&#a�VխN��|�8�,����;��Ƀ�����
�:Y:z�۬�Im?p�G?.~����}\o������٢f�Lkx d�Pa�_!���d[��[CZ����l�����B�=W�q�%���h�`8.S"x}�?����x�;����b������:�,U=֒�
��tK�������M�+��j�Hj�n �H6+�+����t���L:���c�ef�z=L�\ȨK1ֆ�E�X���*��T�/��B�7��uR`%pƑ����cq�\v]��,x���+�d���0``	
�'��J���FoE���@�� �e-�@�+"�xL }`��-@�jj��P ��n�Q�d�4bIW���)J��֕���.e���b=OK��A������T1\�eK�0:�M�Y]�^/��YCB8�f���_(�2ݎ�sP6	���)� ���
��=�^��Ţ(�٫}VI	��Ԫq���R?�Xh�tt��G��8�^�j�C�tz"'�eO�Wt��n=��6��ʻ���t�H����%��K�d_U���y����:�I���/��wA��ќ�o�#ܶ�½`��h�
_�|�C^>���(̀����5���'K	�� ���5r�SNc�Z������8�˜�#(�V�]���7�(���9��?���yo�-�������@�gt}Ĭ����k�I=#��f�V�+!R�e$/�=�>@>E�z"��R���z&MM��A��@#$�Y��@K���}�QO�g`OH}��=�^�U&RJ}+H0���=�g��[���e�I�ᅆ�=�禞��=!@��\��i�g�;ѡ,7_���Z�s��}��Z���O�s���'���G�6q������Â"��<�9�s>�	���p���u�O�'Ai�3AsvyҸ�ʐ|��M��Σ���q:���.�������I�4�(�h8�	�$�	�=����| �j�|\��LW�ңN�En7&b�D�%�rI#�C�����5��5�R�)��mK�O��7ϳnד��^D5��X�fgGQ2k�^V��ea�k��M�+$����Vu�z2�����BcS��~BM��v/��L�\*A�)R��i[BHѝݐ�_9���xP1�x����;�0�����k�Ưw\��@H�fEqь�/%�8�g���~+[��������mkoRޠ=B��7�LVDd�^/p�q�|�����Q)C3xh,ɹ��m��^�P�_ᵽ���~��mT���(lWA~0l8Ϭ�)ə�E
E�8�[Ąbdߖ��"����v���Q��{��E�`>��ι\�[0��i�,E({��م%�8V��-��?"����a�6u�HJ+�DD"��<�Q����OH6�H�"���HH�c�uV��ǛF%��s��i�a���A�8TT32�X����J_�i��&��6��:H�B_-YA��Ri~�� ��?KrD�8\)��
`d&U��k�t�J�|hυo�{��0��?;�ޣPÏ>�����q��T#� ���	�
S�9B��d�D�/U�"��zÑgv�YֿŉD��P%��d��Jó�C� A�i=��G�m�N,���i�{$d����oEՆL#d�qx$�-���h��7~�9>tR�̈́����_"�7�"Zx��X��8YmO���*��Ŗ��I��n�$=���Qh%|df����#UA��Ett��3$xu-�����.k�\q	��xW,�P��&�S���d�S4����RuO�bu`��s)�4\Z�@�q���6(�8{HA�Ni�W��S�㉌ �E��C�8n�'8DtW%7�qoȩ󋨒u�Z�D�E4_�s�;b`W|`���5�I�>��I���0��Pvl����CW%��lMa��&�3S���>����Ol�3�> �}3z
^��i@��U�J�=Pگ�u�H/�oe�c�?�H�\D���l�%���D�m�z�8 ����7Sr���n�9�S��3E������Njw�*�zP	��/Q %
N�%��vnߟDk�,��f�U�|��weV]�4�	��oz���W��@-���@���U���T!�oY,�˨:����oE�nES�U������.$���۾n� XU`����.4&�tC�4�<��s��'��Av=R�S�{�/3���zxڧ,������d�]C�;z͏� KJ�=��F��-_�ԊJa���7_ �4�y�%`��O;���}
�O�C*VJHF�sb��\��F���R 	E�-��y<���T�?y焯��5Z�FSU	���/��l����#,�����W��Q���w�d.����G�����J5�&��A�*ȑ��{�����;|ʘlByo�'�r@�"����03� B�SW�;>�T��_����0��߾L%�潩 ��c�@��6ૉ����A��׊^�4��K�&�������oa���;�����PY��r��5���~�س�<�!Q��]����)��@~�Zǫ��8������a`wzvr��3�~0��y'^IxV����.���K�=��vx���Ƿ���f��+�Ó��=I䧯Pn����ޣjId��)��)�C�;B��åFIP&D@��w�c�̺vi�r��~���:�"݅������l����h�4����,=.kO)VTS�Y����E��F�������A%'�������`~�Ez���m�İs�'�sn�d��Z�(-x�k��ײP.ru		�0���j��4��[A�aga�RZB�#�h`3|�ω
�L?�ׁ��D�!�������ϙ�Y�f�k�� �����U��4K�eq���d��;wN�fXJ�)���Y	$}'3��h]�
�ڠk��Z! �Ub=��]ezL��y��L�}��v�C�m��&`��K��(-W�p+��A=�=�>�?'9�����I~#L�V��g\(�M�+,*��[E���@(���j]�j����qz���u��m��(PR�fNL�"�d�
@���.�~1��8m��y�-G�G�-�a�f"�;�����R�2B|޲?oL��&��8�#��Q��N���8O3�`�� �5���^1�duXUl��8r4�Q^��u�[*l����q���˛�:�xպ�`)
��?Z����{�U>-�4�0Y�����1�r��]CN.p�-���-O{�E�^�G-;ٱ�����U�!�%���&��D�
�Z�y�A�)�Bm��H��G
w��s�-�K9Y�6C�ާ�u04\���''1z8����3O��|H�:��%;�MA��^�9j ׸^D
_�<�)���*��%�+�-}���uҎ5¹n�@�s�� #6a\3z&+�fٰ@�DX���8�,�l8�i�Du�8�a�Np�&� �'���A�ҫڤ�B����[���0�E0����Z3��3j@��|�C �Ll���٤pXK^�Ծ!��ㅕa*����/+>Q6�%륙'���N���@��moIo%�h��>L�d0ǜ�	q��`:k;afh����!O����#�OE|��\��>�ց��7�ms�倂�:�k�2��
�3���-�24�B��
h���\M
"��;�>C����1!`w������e�Y�7��^��*�I �svBQ���xH/�~pv�EM(A��`[�F�"MI�J���Lݫ��kF�UԲ O��XW�ͼ�fcN!�J�y �r�����r�_r���x�~;y�ЯL��z�������ċ7��~9�C��u'�׾�2�W���")����^�N	�l�X��4g˲ >����r@���u*��t��K5���{H
�K��4�z���A�����1�2R�s��ZA?����!�-!�n����18�F1)ؼ��6( t۵��n�)��3	���;}�~���o�Y5nt��`��z.�;q��Ș�=^�p�ޞ-��Qb��3���*]-��:�.��x��[?����/���^�\H��Av:M<0BЕ��XL�1^z�Ϯ��o�NY�$����&i�D]��+��N{D>A<
�[�$��mFMn�wt89�B�Q���Za�c�y���g��*�`���Z��`���%N��Vx!U�$�5�,�5�Dɵdg���+�A�}�*��]5�Ϝt��f"4����o����|G�H��g�UƏ�nEӄ���${�<��"n�w�bx�G�_0��#p�gӣpS��]����_hA2r)�_+O�^w(��{���#J�?&lpQF�r��R��͉�FV��3�]�6�$�f
�g� ��`��S�(P�a���O.]Br�ꐤ&
���YN�li�g�$��G���_99�=�Ĉ@�եɛ�d\v�:���^^���(�Of��?h�0 :,��!�Q <�f����]�S�	�-�/E|��+�3cdj)������oJ��.�ykLx��Z$�(��#'�d�,@B2��_}d�?K�x}ܸ��brf"�����>�U�N<������ԀD��E����@)v� �V-kE@KD|���u�Az�R���;d��(��$T��@u�X�u�1��g���l�k�B�pR$��-��5 �x��
����sz�U�Zҩx^mF�w(�i�pּ������SI�;{l��H�BTtד ���~���K <�O��`VŻ��z�Q2�i�Kg��4z����8��b��I˔�>PUbE�
�H�[W:�ar�ߍ��:>�G!ﬅu���4K���g�p��fh��M��2A�*X���O�	��Ф���MF��~�j�8��Qx	�c�F_戵�9��ӈ[��K'�X��_���b�-[�F
ҰgV��l:V`��h�oK�ú'�>����H4��E��#Q�[�̙{��H�e�8 ɶCAWH%{:E4�a-�M�T��T��p]����m�{�Bbn��G���@�T�9*c��Z�G�u���~�
��ϥ��-���LCv���SZ.l�~�(����!�4���)��7�L��ء�%f��/�}B�{�бd��H�>�^X�5���jh�� 
y�o�U�\���ŊV˄��5[�� �����[���s71��VȝFA��k�ȶT���=̋�yHR�5�������<�HK��;F�J!^#�``��L��LA����!vU���H�R�pbU�R�]��>��nc7��S�	��\K����	8��`�L�'Rf���(�P*|��홋:["b���t�{�:O��Q�e@���zsMl��P]q�Ł�X \�a�����ǎ��׈�4�Q����R�+=Ҹ�e�1OY2�A~�����L@C��Uh��8<�����n|dM]C��pb�['�{����Z���cH�g7�c?r��̓Ri�Urަ���h�:x@�1���ڃ/�Z������2�&̬�Y����W�f*��u�p[���:I���'2�C�c71���D�;�!�YUU�zE^<U�2IP'���i�7t�����$
���u�2�?�����Q�WƹSj#g)�v������w�{��k3�Bǿv�n�߄����H���GŠ�����B#����q�o,$-L�:��Xc��ٮ�2BK�nj�ڂ,���
����Az�m\s�)B�`o��9L]8[µ�y2sR_�Kw����!SJ��&yf{kH�>��� �']��d����á�Z�i���<����ONq�Ƚ����h�=J6_�w�"�'��5me҅z�?��d�vYN:r	��k�e˳����[,v��o��}mT��5��A(x��O�►Y��/�P���,<n���6�8���*�s��!3)��죶��*|	Q�x\��Z��G5K�w�qf���xv��Z�<b��2O}���H�^��9��=����qmG��Hu���b�)�9�=6���t� /W�5ܙXѐH���/M���zD��}�����5��#� �Zp[�y�����ov�_%�SËB�4���~Mu5��<έ��+�鼹��G��t-̯�x�8a�}���������2cwlB��6�W�GI�0�����YX��� o��,��|;�;t���`r'�P���k�v��;�
[, �|tsQ
�z��t�7�3��n��ȅF���m'"����X�&M��v��BϧK������"MϸI���p=:ȾÙL�'��
!�?N�n�9�g���zn�ϲ�j�G����o�����͵�Hp�����Ӭ�H�_.U��j�D�N�#'��Q��7���De¥8ηOq����'��!�Nf$0J����L����7LN�iЕb���

�����ݎ��6�[�De�;'����{�p��n[���%� �<�M6uY=#�{|H�x�f}&"�(��Z� �l;P��0���~[ڗq����2І�/-�f�'ƚ�K���8�G@f���'��2
^�f��(�����{�����.�D�x��������#I��<��5�f�ǖ� 	},�x5�F"���KIN �tgD�� wʧ�{�cx�`O�m��q���僶#�y`���E�D�o�-#���4�x���,�c+�!��"�?�Ud�i��,+��W�&}���<�A�s����I���cޕ� M��ҽS!	Jd�A�1� ��9�=�E;�7s�|����E���R�� 	��������-�IA�'V��+h�� ���\dZ˧ޥ�E��S+���JtJ�J>��Y����nT��s���t�,!�M�?JHe��ݧ��#T�� C�y��or/����,t�.�Ƙ�7�nIOQ�F�ձ��,,���be��Z^Ō�7���R?>�R�uH���(凵y�C���O����L�1�/�&I�Y���]�uܶ�XZ�\ |������VJ�4@�� Չ�R;`��.sm��%� �P�ι��*o]z��ݮ=v���@�����g:]�x�=���,���E��|�àP��+,('	�$� `���gqA�h�� ��o�(F�.܈��C��%F����T�ѣ�Fп���M�i5���`Ak����f�va.h�F�-�M9�x^�䕦;,�D��6���m�_���J7���Y��\����Qo�#�%���Y������dQ�-NN�~�Nj�|Jɕ�"�pfዳ�}�b���QiFL�Yᐜ��\�z��]Ǻ��sPX|;��S�Ip����k2�6�(�8Q%����{ժS�m��u~B�n�I1�o5�®$)�Aj���)�6���R�-_� �.�J�}���QE����`��e�
��@ �O�O��Y�1��G��׻��HjM�٭�o5��P�_�F�_�(�,4�����~/�aeK�?����F���������sPsC�H�g@���"��|�yk��hN���>�����t�@�.�"b�rh��R6aª>T�R��#3SW�P$(�4u��1�īߕ+%��:�ۮ�R�eӴ��8<��;�6����\IM�H���Ж%�G�Z���T���b�7����5�qk�I�(�2Ca/צźVؚ�
��Ozl�O�/M��%��R+�,�S�[��:YE�D  ��J��[������{�S7=������$��D���d� ♳I�F&����9 w|hf0�~�D��}g8Ni|-��)gԢ�E \1��扠�p6^e��&ޫ���g�h��I	�󓰠�kT�����0O,����bȥ��.�|:=C�ǝ�u��~M�uo�s�X��x,L�M��8�J��G;MI����j�����v(j�HDQ�<�/�x�w	mL��9�˔�5�p��A%x�t���޾�`��	^=n
"W��A��=-{��e���Q�qº�ᓿ%���]&���?_y�d~|�y=�(jŃ9�� �h�s%��evJ�5�Q���/����[��|/rbq�F�f�$��U��^����&^�K��>�C��tv����A��J���E���prU�,��Y'lc.B�a��̂��>�,��R����e6�rGڧ_�����8ā����L�H��A\�.b�r��޸���C���㺗�s�s�#�Д2d��r5�՗^�O��S5j��]�j_�d�V��ء7+j�U�CIN)O��P��f��<������ ��~4hx�"�3�<���!���9�܀#��շ��{�������Y"�>:�0�;�������s��
�W�r_;��݁*���L�ȸޏ�ؐA��'��4u�(���C삝��EՓ�
��&Dn�x"�>�U�G"�ǜ?^�`��%�ӻ[�����!O킊�-�_����&"*���
�������E����b�yk:�?�����m�j(� ��0��Eː��!9V�$�hhS�����Ox��97��p��8�����G��O�f��`������@uˁXr��5�����n��3`��R�� `<���G�����������7F@J��t��9���:Of�n�x��~7�MӮOn�K�^u��L�D��:Ig�랿��
�楴�q�ye?�b?-Fv���C�z���E�<T���I�c�:����}q�_�4�0����0�HZ��V�+W����Om�Q_0b&�(��K,;pI�V �&|��9����G_8�%��gqeNf�`�6�&܊~4��J4U5��^�T
��la���RIޔ�Sqd+m3V�s��8�d��|�y�-x�������-;��SҨ(6�������2�L���ݵ�fP�rEe}'�3C�����p�wWYҋ���wg��l���Dx��1rN��ú��hh�9cJ����gȳ�F�ϷO��;�$��C�pbW1ۧ�тI)��.I-<��>���g�ي�M��Z�'�C�mna<�5`G�)ɷ�QY�!�ش2O�zO��2`��PprW��y�J_�)m+�22a�Q�4�ӰyN�� 5�\�y쯺gp:�grT���٠!EP"_��ȱ�rc�3��cx�u��'A�6����
O�ŗ��T��ѧ��$�rfN3	���
�5[}A�Kl�z��,&cS�2X�'�/BM�� V�;چ��@7f���>0]4E$��y(Nj�������:
�/@�<�i��O�
s�Ҳjp�S�I=@����u��+��Ǔ�L��Z4�*�|z�ש�TM��ӌB5y�P��&uk�_p��Z̤��}���Y��bf��$�E\W�9�L����LU,ʬB��S�ܶ�t7mѩ��=�Cx;�*�D����AHHY���~P�/���d�� [����FRA�rJ���i,��gr�}@�.��(ĄB���@�.��z�7�H{�3�8'���H]mx'S�8�z8%C/>b�F(v���A������ ��gR5P?�A-��K�;��4K� �Fzp�saT�2\��>�UUu'/��f��8P���]V��+�&��%s�Bg]�dܴOv�&�Rz��A�ģ_��.%f����-P<Ф&.8������K9�e	/:C<��dX�V	�S�8���t��h��6�̻�/���Z؜��1�1��X%a���|^E���$�W����[/RM��n��6@4?./p7�������ճ��/Ǳ:������nW�t)�g�2\�)y!�c��w�p�
�6��[����2d��(�6��hNȤO�*���*��XC�"�?�,C
��nL�W
qUϝ�?�r��>�I��i�y6sc�_g>K.��{�j<��GULd�˳��L�}��z��K��ؚ�4I^���[���>�������A.�^;�gc���}6L�5�-k'�(X�.����D�bx>��6���ad��K�o�8!�ŀ|,�Y��or�̸�a�h#�1��l���Q�W3p_>7��:ހ���k6�5���w�@�'e��
tǘX���x��K��Ie/�b} \���Z�H�������|�� ���3�\���K'�F\�胄xܓvYdN��y��w��$�ۨ/;�$�	�� ���{m_�nS(�����k���\�m"�8:�%�>dk����;�@Ɵ�2v���qI��pI�S|D�?8���Ȳ�`�<:�-�1��k��D�+`WM�&B�3u��gXU|�tԤ��A��p�*��{��,�d'�$�G��R���P:tF���#u�ޠ���T�_�h+iX*��0m��R�^�C:oQ�.F#e��1��$�vr�-i?J��>BIk�J��n�5q�#��tn�j˖U��̃9��h�u�����F%̾�4X��m~��{�Ǘ�c�7��Ƭ8C�;��/:77�~Ӡ�!qؑY�gT�9�P+��`&���Iӷ&��r-n�5-"e�g|S�ޒ����h��e�ǣVd��רu��Z0ŉ�Q-�խ[�78�F�,�f�p�_�5*�=�����k�O2aBIm)ȭAm��\��!�UcՒ�����>G�1�/��M���z�MՌK���A0�LNP�E���j%*W�/l�� 5�~g��hF�ڿ3!��
�l��J^/�H�A�E�G��֖O	��4�*��JP ��%g7��U=a����N���DG�ѻ�hГgz[\K��D����^V�# ���:K����d��}�*ɦ�7� �:�$[x��ֺ�M������z��3�$נ�T�YӚ�����n8U�޶�u�.'\�Ϻ�!�9Y:(z`E ��j�i�S����^�sW�-����lz,3��r���� H�Rzr}Lߔ���,���1���2�{L\�R���օ���i:1��E^CJ��sk=(���g��[8V����Ic�$D�����;w<��e�Bf�F-[d�E��8�B6q-\������!��Ɲ_�."&������~/�9	۰���%�te���#���B�p�%�����`�9���b��*ܹ��f��dd�0z{��M�"��@�Z}l�*������[�������ͅǑ~�#�#ٕB��Ec���@�H��fi-l�oR�xcQ��XrP~� �^�>�}��
�P U���)2��H�?���ݠ��v<<q�3�: �&�1*]����?��w��C�G����,�c��8L�O�g ��j�Y~m�&Zp�����hk��}~�8�yGtG����9�Gw�Dr��N's�]��%�Q?َ���%]��sʚ�~~�S��dVi�?D�n ��P8$� �CZ���� �k�k�@�"��̭��F0�xrPGW��͐�+��I� &��N���ԩcs�"����F`rXQ����U��.�E2�啺:M�Rux����V�G�+�ќN�0�sA�����?6��#����\9K8v���腊J�!P=���3g�&�$���ީ�{˴�-|���fF_S��{&�)��G��6'�ٯ�E��5cROz+*��mf��i��3�j���H>RGH�.[$��$c���K�>�`S�@��Se�ݖ�66j��YO���(xx�:�6�d6�Sw,N�m�E�{�D��������}�Ҹl� ��ˡM㖗}�[��XpB�ՂaZ�+7z�,;�n�#���z!����U��#�!0s�7��5���9 �:��#J�l�ް�7�@�������o'�g�E���[�8S+�M�	��hisd�_6��[���Jg��Λ�@�xf��j��LӠ-��:\�gD�4����X5�~�����5-�	�����t�±��]�KDn|�6J'P������LEvq��=�j�ل�"��Lg\ f���wZ4s$W��cV�tC���{� ���1E���Dƞm3D��N��n����w|�\` ����ԗ�X�/�ISfwF:����{�@�eVd�n�nEҹb|f�wu�A�U�K��#l�t3�ZׁML������޵�:�G�&���&%���ef�D��co^���WJ���<^��F(2y7'���RS�L6<�V@M��c�[Z]8��v@/G#��s�n���BSf颕������y�z�L������z_�[�����7�_�r.ߵ�g��-�=��k��t����Y@��8�3c_N2��o��m���H>�r9jmen!�ږ`H5֯~RJ���L�6��e)��Rd˗��p2��gS��'U�`�����ZB�0ԈZ�p�"l��z��"f�f�y~�ހ�Sãk�^K�?�L�����s��/8ǰ���:2�?���Z���!�A��ٟz��H�Tc��쇅�����;�yܭ�\�3u�k*���{c�ɱV=�G+.���ѩ�`��*���s����'EWL2f�9�`��\09Z���F��7�q�'����3
Ja��/�	\߄�9Ĝ!��$��2rx x��В%޺�A�>�$@FsT�^5�9�wN�M�z�,��S\�вo{O?�������W����O���r,�7�O-wW̾D�l�r�#���xR9�ԭ9 nt$ �͈���ĸ@b>!t��XD�Y�^��#t��i^2r��B����g6�)�0��� EAMHa��6eAL.Œk����R�����d��\Ӝ�;���_�s9�����/��/�$)
� �84��ra[��MXk56�!ds�W��_�Ǒq�x�u� {(��H+�.����MH�:�A�̛o��ǁ�O��8vM3z�l7b����s�����"0���C#���	�pz���_��ل�P��g��"$�E=SiyCd�[�C}�w��3�۬�I�ى�M�ѫ)��#���T%>Y~I��,Y
��G!����ĥ�ƌ�r��q��i����JT9V��H�]K3�aDF^��Dԧ;�gQE�JP9�g��P~�!߾x�\k>����#R�e�~d(�m�.��8���U7�����5�4�a�����Bw�O��4W]�ؠ��ۼ��j܅R�zDH����SZ�4Q��.]�F�_�#�̋�ڱq����)6n�lP.�o�Ge��;#�%6mgg�T�n%��r�e�)P<0��p��ʵ2v�t���E� ���~V[v6�O�Jr�)�é)AJcE�5v>��ʺ���B܊�|�r����i�ᆒ^M���!˫�e�����Mhz�A�Rv`�����CyPǖ0.Q7�0:�p��")��^�el��h � ��`Z�.�wQ���ƿ� t"Y�<p�=�,��& k��Y�7����'�Co���%��qdd+�&�
����~h����%l
� *ː���+p#��
�={��#*#�{��d�3�&뷧*��4ٌ����%Έ� QiUM�	ܽ5����?l�Q)��pX��M��a�a��V�WP��rӹ�����I���P�ѧֿ��=��d��Ѭ2d���:e��G�V~pɺIu�, s���y�YŶxAL:��J�Ee�n"� d���Ɗ�O�o���L��*U���h��!�e���*�9瘓l��"��g�>O���%O�[L�LT���w�7�)�1�3�����l�wg���)��9�2�b�(Na%s+[�Q��� �V��"ġ�"�������ZqQ�ܯy�#U�7��H���,O�J?����Qֿ9�]�B ��bQU?J&��C5�� ������f80����TU��g����_e�9���o6�͈�t���ļG� ��o�d�ZUc۷�z�\j�� >��o�{i^����bO]��a/W����Tto1��t��䘹�4��G�T�͙�/e4���?�]8Oj���g��H-�_2c���qK͚Ƅ�Z=�����m-I�``w���:��?s1�<��{�χf���ױl��x,��U�D�y�5SĪ�,���r�se��l����}�0��Y�b�<+V���VC��h��qR��C-��CB�V�>p�e���wt����3)�W/֟�^D�i_z8;�;U� ��zN�$�Dg�4�KS��B2ރw���U��&����	����W��Q��/���D٤��D]|��a�ˋ�5I�Q��C	��i���&]���_����l����oucE�}X���w��lE��
��� ���Zs��>D�ؖ.��N�d5ov���]��>�M�qƮ͂��?��K[K���w�ҽwU����1��o�:�|/�k����y3����F��rf��r��bu2���edJ�$�.�I�-����5����(�)�:�䌤ʬ[%���W�v���)Q^�r�av�z�1/��	\הqѤz�� }M�Ŷ�g�s�_�p����Y��