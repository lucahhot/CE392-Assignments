// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
nmg8wQRUUTnOQGzy7dGxy+5Xoc4lerg4HFJ3IkJ5SH175n5OXo5EDcIDp2Y9EUSB
uWatSLYNXk6/gLDTnduR/dSpoJmvehfbq1nf1TgQPkg8zFWDXf6x2RSgSWhmAVFe
awDblz9SG9dEvmiUT1uEGJPlwrjN9A6kIDe3lyzLLzKwbFpTJc9eLw==
//pragma protect end_key_block
//pragma protect digest_block
gzE9Ww/mt08YX9mS3cjdOl3VzEA=
//pragma protect end_digest_block
//pragma protect data_block
Wkys5SvzLdQD00Y6G/ciFRAC8EzhJK+Nh1WBT2devUP59Z/z96I/m4egZU/eLxXx
q9iLTf72vGBNegDvWD1ru1z9UxF0ZL1KvlM8H55kuTFTFLeKbcdMC2pP4pE4NG5G
gWZ0s9TetiRLvu57VWP7sMpLQeKS2vo2JyY4ydQBAOjgwKG7HXYdziYvV7MouLu8
i6BekdDQJaV5daeHo+3GHSi569MSrEiLee7pxZvkM+gyP+Cl9aLcp0sUnY4cGvlA
Q2RpjypyUKyi92s1CIoi7reXCHgDtzGhBpYgDmAbQMZJayhQCJSpaoH1GD411tqP
K0RnJOfopd+S8Vb7oWV53bAL5JHyIgVSlPHyP+AUOYAqdOro/ExWm8brSnMNuy3x
VvXZUvwqvzPDEN1Jj/QkPPu8Ai7/DKp27vS9dCG3cAAjlhJawarnFnrscWheNlvX
v2iIxxWs3kTvfwl5QNHrk/tuZfRUJXpiwn3hGxE0X6TxA7KQU4/9O26m2qMK89Iv
XzXQL9vi1RnHZnGmYHawehYc0vFg5x1skFi29hBxmiyCW4ctzIZC853ZO/GNBVN/
Aytqumb3c2ZFNEtadax3ScFmsh/pOFzEWeOMA0YNQCd3loEIl9eN2FE56wdgDhme
5X+JPNK5AE95gMe1IB+/zleSeOwP7rDAo3pu8bL6+AuEMr3OuHRILEFFuvyDpu87
AoaX8P3xtT4BBU5oUsR77KLJDKx6euecHeWOsjUB07Gp9S8gGT/knXopDcnf6y7Q
2ugVpXBzloe2WBGMKVoWRLE3RVdUf/ryyHKa2rfmSF3cZZUaVGMrKqPP1Bfwr89n
H0Y5OU1ttUxzirFyAwNjHk2dFiHqnZny1GsMc20DAP6vPQgRNtmTplQjEg5nfX+o
9Y+54ca1f/G4EslZspJjGv1CcHMGx2WDgA+S1bwiBzhMz9DVKwov+7kVPwhNFuAX
9+f3qi/svzYqDDVVHselYIcvQkhGlfzoa3aPu+ueA5OMAwaGla5xF+hUxhsjF0tw
K5t9CkT8pWsGQsi9R1ItKWXhZpzplX15K2PQ44J3gkzeN0bCOMJWO5MgudSnPwqh
DtWg0/XepMSn366tcDIPB2Cc6zOkWMDVL3p9tNhrOLZu8IVsAs+PlZgLqmZjknRy
gR51uU42gZmijk1V9Gor0pwfPI2ZH9dtJ5GbKBW08IycQ4geezD7JJZf4YV5P5Iw
BnicFfbEW/CAY+pfmvRdpRzCFOaBN5cpN4KDMOMe3bRpfGfCHbbNta+m7o+RK+59
SviM9OX3qiJJ+TUDAPe+Q1ZZQpuuv8IJyMZFydDBTJ28itq9UV7uhDaO3Aq5+Q3b
PAIS0RTn2ClTikpeW3zzk1QbAIcDCYde5V4eYqQ+h9dcpvDwRaXtwzpy15G7iRcw
qVS1j+5u42LmpIt7Uee5dOcF+Jmo9/EB77MLH0Yaix+0sxtez5GP9rlYMXg6vR1w
V3TmhJ1SwlBVI0XC38Q0XKzuiEnzC4ENzER3uKSrOaJWr6OzUoThaJ71GyFKtmXS
ty3UDm68oUBHLmkypnp/CxWYG6+j/V/GTXf+4mqOl7IrCTHanJll++ufbNgLzNdB
ji3mvYztdsdztMFDopH4P+2V/5yACpzHhjI3MUfvLBkyuTS4Tnr28kAh8ATxI4Sa
TDjU8Mc4It1xkidx/qOdvQfvQX8eDJND1aG7jGuVT6T9vI+QqDy1cPENXo/8yUa0
lq5yw8zqtLU9jqS5yVu68Zu/TCYdJ5DYDnwhjSJpyjmn7oilY4AcX0TVvwNCZasS
dG1mXow9qTGSuhj/W3pF5EIjxzM0JfXq7ipcL5yBr73Scwth3Xtxoa/TyH3oeHuM
cKEXq+T2AwRoc4zbZdXbuoNFGX+qWZp46/KxASylQ0+uTqLu5tKC7V5uP9F+RJ+4
V7kkV9j7d4QadXzc5JmJZScsgBtvMjgmWZdWtkOq8kLmYWqi3uTC+wuXxnzFp21P
8ZHuh++6ykhX3wt3MXHBzyAXRiSBeXdF0LZPtxDG4T9QQu/L7sHxNZkPbdqnFL3H
5T2F2x0H7GOqCc/NjhaSCTIOUMlpWLMz8gFNfSbzEv9BLVA3iLg78T+GUjbTFaAh
xTxDHBPLPg+I/DuPemnUGzcxUkIh3e++u4R33+ooXRO1mTfw9GlBQsIAMRYS4OGg
RkaXpRkmhJhtKY3ehBc6Gm3aDh9s4+yc2rDjxBQNxBo+kAWs+JtGQzD63JHBoT9b
yTeOF9g77IArT4Eh2fms+EYiK8JH+kFAxL7gsjSwpmewY4VR6Q8nwBwSmo/YZ4+P
NmDy7R+Q7lttY/S4bzSG6uyrkF9fafFTM9vA8s+CmGp2ogadkalBCWxmpmgcQ2GD
u+TQ8jvm/NGztZ0GM8MQURKqJI449yOkAFv9oI1oH4WpdjLWX1X1cXARuyjlvsVj
BiMZnilKzEZqftF9koOkrTrwiDfsYV78776lIn2N1HN8UJxTQYgBIaFCCf9Mwdvc
FXfoH1Cv241ciSK6I/7R1HfGurIpk/pnvi1haFPp0wlbb/Uscc2IdTrs2c8M9ASB
vnTXtQuNxpKORAIPOwjVbKRMiEd0WWuK5AaqTRaw+McatwJE5robvDjKnYgwxzkA
we3q2YZh4xaDjsquSGcTFFXfcs1o5Hc/7ml1VK9CSCNEKNSHnXcDMW64KhThNMDM
6JVXRXU243Q39fYH+VScZJoWG22LWxxndEPqqMcua7FPpmAdBu5wxgn8POMRAnrk
NXsaeRyYeFn1FO8eHxc/55I/debZct0oQuLaPTjzcgBjHXKu7xaigrEs3pnyJ9bV
Jy14FxbkGqg+es0evlyCXri2oKGLSh1l+2itwnMgkGx4M+8P+6wB0oXjLDtPe9+T
Oy0kIQ4epLiUKQhCjHjQ5cv9x4e6IwbmsjGS0yURP2GlcUqbeiPVS6XjOGbTOSJE
WgS5Ja9NG6hL2jNZk2VnKIAz4yJd+kVJd2PUIOO6nnZGoi1DWeu3ZHOhmvFeTO4i
pPNrVUhfhiYOOwzMarNWmFUlRidgBrmdxNmqG/AHu0498BxeifrtehRnu9z3Fjd4
aoC48WNUyODYh4gFJt9BxNzl5n6NKzbW5Ituk+ede2WRyIaLUZaDCDlb+7J90jOC
KQMv2PABkQk2rznxi9wTigCR2I7UygAxeiflXgZ6jTcakrEmbnoKon0w4z6iuCxH
6x5dIVtpql2ixSX6E6yYuF7re+zEEXEea4h7mOGi83Ejwe491fIqXpofrYRIRj59
U2e1rgYlu7Ks4F6MVvglEyASzg/GTos1+0KUxera4MiCA53h52gLm6hLULmxrRZy
7fzmhYAjRTr09QD6PE01lyL4b3/yBJ3hI7GPIrQIBl0OgPoXcZot0gws1nhPDzCp
WIMPnX5k4UPOD6ZTbRRwaAU/a1/g4izgyyyWWF2Ml0MQkopPchF51jYPzXZDQb+R
smnntJy/d3bd8MJPDoOF0eNUYMvBl72ONiT9H/UxnBWvLSjK0NHzh1h+ECqGrkIk
lRxjWZ5tT4WgeVuEQEFEGnWaDmgMXrCPZQAWuGsX4s9yEUIoBVF8DhXilkSlU1Ad
psMQPJ1/JT09Eo0brVZNo1em3IAhDT47MJARi5Ddjlj/93RoB8AY9yLcoHmxho94
O6gRkYmFS7BBARPMsjk4s0aFTtl/lc8SYCKC8Qn8c5dUM4oZSrWRpyP91K9W3Uxi
plUXZDvJr2hvDOb72FZF/3+xC2rav7lkALHb5POTbAt4mMbZiOYjJO1Hmupfwxw1
OLfuXZycKvVh3ugWD9hJ/w0bfHMg37v9Is3uJCxkaw7qPbo9rUdsLAAbIoVZAi0z
b/Vvwz0ZedahqV54mY0kmCKZR3YorUeH6Qf1N/wrw/JHPGxJvoV2YYyevjJXDrGl
8yzV9TJulkpdblMptvjtXHUVvz83bzGXsbOepd9FbwBCPOIAfOoDXz8oq2Usa706
j8TmEEulo5RXil4ye9nYKHSTinwueFDLKe2XEVcbuKluiWyPmMcXVRC3ixQkzV/E
ZW5sKiq/bgS71ll8bX46uYRadpVc6eJdGUor0TZJ9Oov2EIh/hPhbhNLshf2B1gz
6GRJnCnqvbhJHj0TvkYQ6EEW89PPcsqpxRiKaRMm1iX0b4Pai7n1kyxavIq39Lwt
vdgFMxojeNguWUY/bA9dQO5Ek60aNDzDsdCEywoKFb3aX76IfD9ZX0ljOiok+CNv
n6XtoMCFS41Ut+q6DRUIFQSh9lF+TpUOsi1BrAN5bc3+EnnhcQf4TGB71NSIjlSJ
L+94lEhJuX92QqHgLuP00Aa3VsGxpaYXAbilOI2ma/6GkK66TxKoY9Q0t/N/gC3+
YizRNev8eA8vaqhs++hOXUWwZZqVbu15jOQkh6npM5jfWDWyshEBoJCpWJ8s8Tq0
/RE0rSHbDgEn2t+Ff3b2mBWYsSoJNyiYXL3bLRpjXsaP59nThROB6AscSaMtUL/I
c0hQNwXnbtkdPhfcWJXUOLzJNTvFY6spgo2sV04nvr1IbcNsS8X5QJVvwnAzAuZY
3zGgwY4mWHrOPkpuGvIak/xpXs4PiY5hCde63nceIjDXwIOAe41YFVSyoEogqBNA
ozforjliFDadDFUlD4PFfHjPZ3m/PQWNGQh1iXeE/S3ridxjb2/u5Jsr1KxWK+Rx
3jV+OD3gRGWmfhJkQtxJNg6bDRpFdXS2seD9er8SLdtps3ICDk7zHgmCw4ahcNiF
377q1zYjVNx1gBigAdGSzR+71ljKDZhxIVeBd2BrtwElLf+LhVwpMVJZDQjgyw11
PF2xk/DUfZPIog6/yldbZO3rFAZC6cBoVRvMXR52rKRkBk6knuHQlS8ShO7wCoL5
si2mMPMb9+eLM5OZZB7bf1kBjF4MNLnsiKkLTLYMjN+b0Qy2SyGQN0uT2pV7hGkF
BjyW4/yXTLdD15meUSqX6J8PowAcy4c9uJ/u4SYu/hi12RrG6+GnSqc8QLqOEPfy
b6o0fGfa6U6SWQyE1OsP5h01CtiztwRcx+DBA16kUBF9lpkivp5P5hcaNg2/UX2v
rBlTbs2fzi1dn3IqeI/G4yGdAiiyqWPIKkycSq4Mmj0KtQYlOALVJyEn/tznrH07
dJwsYFjGal4WRjPJDzq+09IHh9md9P10c3CbUh1jzmfr6JTXkFg3Q0Z2ZLb2k/wh
AtTH39XB4AHBwaOkVGMalqL0DP3uXDArqFW8Zm//fn8LoZfW7SDD3UQOJVHR93EA
1wJiw0rGY0qx4tE7ZyRzA/7wQUhMYsJSfLXkmidQOilCG9oOeMXjCNppluK9XHjI
ZQbnc6NglwoQ5rQVzPML1iNop8cQjJTVI6JS//wPsRjtIweB42xrV2QpxM7KOBqj
eV1cCBAFLGBFMHpNBRcHispWD5WfFHonrFWvDfwQHws/dhTmjh4nBk/ssjvUpBPt
G/CwGmumAioWYGwKBNdC5FARxEoqwtFZgNLZ1xzh2NyjEw0lR0biqFGvVCPc98mx
dchFM/El7IYNMDVp5aFelNJi+AmZwYhI8c0rw3lNNXQSCtQLnR4qQvJG/IbisR7b
EHCxUcYRJvA1e0Yd732cELgHLCY4IavRxga91kvr3YSd19/KPq+Xh2BRrBXPxVz7
ha7xib+6K7/9K6INkLgIZ/LgjNGYkoWDFtWZ27FFAfYPEmW9melF9aI766OoN2V2
fTkiqCnxv5X70DCW62J6TexsjPiHKc0l8hnDgUVFRTSpJ837qodJbyuCpTBQU5At
/Dgc60TOYZFxgsCd4ae0HkxKNvEZFsJXYCLr4IXKM+9sQqOCbMwVNMcDGNnVXuM5
1LsnI0WNespwwxzfnin/TQGJT4lgCCaxQlavqx5x/NnswW0vWxWHGjfepih6CNpg
QAbJ1DR2WyWv2JD19SDctATczzbLu0EueoPVfmbrUwgEnxVKJhLw7IevYMWdUpCO
IbppCLs1MjnatClXKi+iLarsnRBuOtPEi7M3JUI8qLr5sVLeHsHz91qcpJtNmV3S
GLE1Zyxd1lbB1ix1Zvq0VPRRTsDyGB3cOlpvZaDU3kMFh1746b8yaS9brTW1GJas
s/b2z9MFlRM8JpdqgT+aakbex9eG38qk8zImnI4kzxQmbHnYk8EqbmK9DT3HI9z0
Ap7HUe6UQ3j+PNCEc3FkkO0tbYcYe7KbfI3NV5JFfOvme7NqtJz4iWnqKBVtUz/F
yo+uq4OviFQqHFR7XbnVQL5cF5cc+lRZ8gnsVG4SW7Xye3xt2QAWWH5elMLyk++s
DKO0eojV1OjphXTEXJs4qVDEIbJmZlNypigCt5dhlnA66yTvUQRC6QAwq8nqCPIP
6FaGwF09KtYpasgdm/2K1+IE9V7ny/dQpYIEmiBsbLUwd82F7mrZnVQ5hSNpzrMU
CA09ruXrEeKONA+DbW9Fw+aBG4jX7VTb/rZg8wGsVFEsL/oMFOYSvszY21h3BIf3
hY8xjsz1dCNoB7OraMM5rn8RHxtEMSB5FyENQVZqam8P7Bxm5NGEUoSivI1XEOgG
vDVqTJcooKk7tws/dUisqGVhYhiJPAGlXydwSYQgUQ4yCXqKtwGC/6XbGFgHDm5F
jL8fVIS3r9XUZV6/XmOQ2U4eOQlRtqVCWHVhNiWuCGvcTqHVmv0ZX+TiYON6+NuK
POUvvO/oXDhDxyKLBbc4ZpOWpg2+YKLDJxDQZc2B3DPI3ZO7QISw7trF8GmnVvbN
DVsDzLIDU6rbabwtu5QR/cdBugV0TNNKOmZ2zZFKOfp1ie3PgIRKiz+unNhpGdIg
9n9o1Kqsw/QwBSUHbeqMZZG9xqutgxEMTdAV96sJIMTD7KtjTEs8P5zkZZG3Wdhd
NCTMxV4+yTtyCBUUldVBPcF2TlBlOi16j+2w5kP4EogsOqjd6eKCFsvFzFf4g4IQ
08AcXTgvm1Kr4jkvPzquv4QrcBJa5EjYhNmowXeyC95LTQwV/mIaWx+px2kRpzwe
B8+dtm650U4+4lIUmFPgBlCCR4u3XWJrr/Qriouv00jESmdWtFIRQRoSQ37BIom3
QUWMzROrDGpVdukgkt6Lisc3th7IDkdx9t+oSa4XzvxrhJq1O5v/3hTFUS+rILdU
xyA90PRgAhiXclpAanx1hH1wClaJxa7j03/4Gp+PhAZhCexQIfGefpg4s2qosPGZ
lX8AXhyOst7wENyW3mU8YLwFG+tufZzxHatJ1jgzhCWSIvzr1Qiqk0AbAoWbrwVk
G3y+vCw9dIdAFBaYgDeB2eQHCpTbuMLCNtfWkCSIX4HajYJ7Is2ooLcRG9QDdIm6
6vtq7wpgt52cc4bJaLthSESW54jtGkQ7E0+L88sDEQXWNy8iiRYSy0t8Cc9A61k3
YDX0XaIK+Ubw5Byf2TSUTwK14C6Wde2qYjYvJpr0OCQ7RO/gJP4aiq3e94MApEM6
NJmlrHHU5MrOM6x0FGsRQx1J6YkPcDdHMadPb5j7AfgxHahLTjxswbQ1B0jVb7of
gNAScDznwlYKPhxSWyjoVf9tKST9nYxbTBRVrG6M9xIxD5ajod8BP/oBdISAgddb
Ft0gxqMXUbyISAfQKeATPrXOMsLOzYDT3Z3mhYUarzd20mW/YzLW7I0eQSneuuaq
/cC14WZmkuBpQoAhEW5SgYE310QNwAEscgarhdvvIACp1uBHrKbc+Ayadyd/Vq0s
kG288IFlKCJbbzaxxyMyzf9I9Qw61Y4kuv+kHIIHTZZLFcshia1/rmLOZ5l/vcDm
de0W6FND+kl0TY4L1lDmuMmsymH9uv+7iFK4rk5yPlLhQSVqUk5RDbCNDpCRaikm
cOtWNyIFL2D8weUUXb+t77lZVpEtlruF6ra2TTQk7B/yC0fj4wsk4mCyyQ5nLv/D
kVr6QjiegWJVv5CsgCNJca+osP9VqgYaIZnJz2Nb4sHOqZrVKt8bsQNXx/PoAeYW
hIugoRdxkCTk8NlkOeNe2eFrqcxqodN0FPgVsfyySsN7mrjQaG8+N/Aj+jBo7FDC
ByiUI/owMk3Xm99M15L2T87bIMFOmBLjtWK4D4ZWAOZnr14FKFWL8hKzkPuLJIct
trCZaPYKsUj1K6HSKrWUe7pLPuwa4Ajt6nXjOA61Z9VWbfSzsSlomOtyhNeJ8iNe
uOCGQltab7HfsMlDncsynmy++mEoPunifYlaqq+sPgJJsTijpiQjZjxIKvMrKR5L
HSfyhGytKgbUl9gcmRw52fj/sU6Zu4ipGgRyULJBWNIrMowe5SPmy9VeUpihuoM7
OphFo41NFdgUlrD88Mwkt2bdaaOPboDxJ79tzOaPbhB2KWW+VkvfC4w2I+nXGsR7
Y5Zy3AKXKXisHMryVo+J2oCthOc6s+C3R6NPG5Mag14ODQMXwznwVR02VD/oaN7i
FRiBlWZmktnp1iCbPfTBGg3qDMuIIWEx2UwRudFQIiUvsgvVjrQJ9UlVK2nuiM/g
+7byeAHk6iTdsx486QkcslL74FTlG/N8/9gGGSiffYMoEQOo8RWGoAsczKLmcuiS
bAXD3h73CbYeDJHLgUtbTmvI5xW9cOkILTfkf22inaFMqryE35JPsxLjtPI+vAtM
QOqPCK/5AyW4hCASy0WSWLiefAcqG5Ilt7xe81EBRQnFrQNpGW2m1dhcZ9Mz10Jw
QeJAkKrcG/Co86WVdr5vpzopaaTegC/6ebavvmPYC0MJ+m6OqMx1r0xdEBi3AxWI
hiKP8xi/DX+1/yS5xkFKbme40eCrVA5CMufFw966PzD9ieEiYSS1BY5KWgxAXp7M
+3nG7AHYvzb8jm3Dou18buwQM37iZxxFXqaPrW4GBR9dMXV1OnJK49tLbgqXtTyH
j4pp96wjsCU6ywGCghfWNEVge9qCwUPucaKUs45o6vx275hfEQxFd1WttRjqiIpI
whZljrAy9NYq0KVcRwrr/LgVDO0tkQ2ZUxbA3UHUg0k7KubvuCuW8gYfHY5XUQdV
svCadp6QuVVNkwiTEIPq3mnnY6u6U4Tt1MDwDbHFNeMCfHR6Rj2yQ3RqR3n89MHe
aEzhPyxcvsUW6H8qzhuW0qJl+c3RNdUf+IZbtX9dlU6C93bfTWYGuYXuUcc+zF1g
N7mGKyo1ajVz0Rs0PoFal4YxkCS+4RRrEhzijl02v4PbVjF8SkfQ0VCKcLWS8g/n
Ej/LxqT56w6y6Q6Zm+6n8zLZN5LzHRq3IupcEtEjV1dtqRrgINYzEMBah+FUarpD
DEGVWGqw36xvDv4nt2YROuncH+3WZDV+3qpLjS/U7UuMv/bg9traqMoZx6aw01Y7
a6pyerDpOqjyQZ4Nzfir/H/k7yebMHK0X7puFbtqwiyd36CIkssv+a4fm8Wwcgal
x1DUTireumPpflnCk8NLuqq06fZlpdOL9nRUeVlQZOsZePB1H148WUeoWzQ3tSII
1+r5l9m9qvkuCvsC+WEpvxwdl68QuwfG0ysM2V57fOgMDG7S00XjQ/lsQkuwmDJE
n+nMZPXNw1TDItjfrZW+GGU2QSAddzgDG++Lf+SJll3lZyjI0hirQKKOBH/JRY/X
4nNWwNTnDGNRvdtZj/hq5OYYnJ+HoCw/p8H8e81COB1VffhgqUimFYcfTajEquxf
EJfSfoQLLuvYqmGudXxAkn2JEhZpvVCvc+yv3x+wHKraloAfYcl9038qd/XD43C+
+cApjrAnZ4MTdQW86cqhbalK0fl5CVkzXtagKKYGNrSLVAtHGPXnNFBsLszLPGDc
MiQePjdqNhR9gPJVKwDU6eW10CJhzLeFaO6p+1Re3cN9+847B/M7oByx5pwon/Lu
6ecOJ/LaW7ZkzGJCMSeW9zYrNwSkuc7Fc264CbYaxjK7oFuRWLRdBBnmQ3F4B1mc
8zXpkugz1Zg74Sobu/whQryf+a/MdIz1HqLunowlq04MLI8Y3tM0cNYM86Q3AOyb
dvpg+995bYFkbrpiCnlpHFYsu9tSqPvG7Ly6JfLhCm995yRDTtfo2CsLN7zWg7l+
tYa2oDgFWUuvr+44xHUbPbym/TDeQV+JOTX0TfS5DC9jZPgYGIjAhdkr0bw7AvX2
Lj8pHZdUrBk3SLDoM2l7BKZ85R2XTW1i1dtUe+jtUE6MR0Tnw3fn5f/wCHPmjEia
PVA7ZDhZR2r9uUCIZfvZJ/FjQlrORJEtL5IhqokF2PdJvJV4EogDGrzloiZkt+h3
0DWPYyss/3NvWX3CZ9pmTLeujNQDZNQEUv3QN38ZrLJbF2XB1Q7vYoLOFIDevyP1
rK00wzEsIWHyjALcg1O/L8N8byMcWQBG95KSBQVMAt7HtEXqYLVJYiUrzt1CQdo4
plLA2oDh/C11ljH9e3aYE9LaqUfdZx+dtqSvr0ob4LhdrhvL5hn+UrF+kseaEYqA
sM65saMY+r9RegKt0eIrO+a5MQk7okh5SqO6nFsz2Hw0Mgcm6+nw8/SoH9txFPFS
6XDqAZ2wMnudhplnIzm+c0z8a/ElVKMDzm/8gjt/L0NtmYs1tKFSr77cG6cOEBaY
xFuMeHzy6cC/0uKxopNqdg5ZNt8aQzE+YIjPA5daF2Ju4j4QOB14n4AnVuKAAetY
w9OYaoWBVK6PIEm/ByiYslXWc56V6So78UatSMZSNEV/ws2iPgT4apw2xmsmyNiD
MdCBU+CV+q4N6rJ1gCLzToAvq33a+9oDxt8+j3ETmwQmGBJM2Ff9b2tikLzksF0G
A/yUeNEzIOQVAnE4gRvmGoAy98eRFuBUJgp+hnQZD5ek0EslPjGJfxg6ZcE721JI
zkLrPNYda0ox2ILBycxNw5F4IXgT3XbuCMFv4kCQ/nTrAEuO7L+fZFwQDAtWcTft
8Sd7D0q6NgRsdN3r1Ajw7FwidIgh+vXIe42CxyONF9FUZ5wAegnZZ7YAzEl1mHrL
UbkOPprXYCk+665G+7PkTZEXeaizM9almMo2mX3SaNJXiBB+hFqaov77tO46Ynu5
YN6CMZ8xAuc9Vmvks9Yaz9TIgABva8qpLmijCNSpD3gA6x++F7Mnsl/sZMX1IbAV
C2syZqV5P9NvHDfx5qydDkGeioFSP3to0Bhddshj71D7gITGMEsAQOwH435sAuZA
fprjJtnBGG30+YXwboXQeuos4lUO+KI+6Tz4gKM6EWlwMqutOSiVmOnRuIgd8IZo
xK5F4hbb7A19g1Gu8z+ULq2K780Pn5+CvyViS6hYbwkO9zlbXCgXSjbUtnKrg6NG
ucAgllBduLdmhgshH8Z9u6fGKx3zARDmDI4O2fJGbNQJ3S42wAPR6Hp5StFNVorg
kL+GeMszpSrOawxRKf51JIxnzEs7xEOW5aYMDyQ1odcAT4JWabu+/cbjy1bXF2QP
r1G+hXYyr+MK4TzeiH8O0QN600V9bMla/j2Cl4jsTTFaIY0QREs7CRVdPE3eYluz
lUFD9B4Cs0gXghLwVjunGZQhxEslajLDD8dzBFSPFa6nx8yoN/cph84gu44tUMzb
a2Oa05cDuQbxkcmiQoqZnin4E/kFWLiTiVDjjkKbVHaejp6wkORuzmCyu9pjnTw+
3vtd/oruDvdLtm5PHxMa4OGvYosfNYOikd9bS9I7YvvAHRX9sunFxyObhXyBxiL2
56gXIyLy/+h8HQnZkNllHakbA8gUXNeIOli8ceh9wYMh5PF6JpHl/KqHkdv7erDq
/M4BYfCUKWzVmaV7GU7kNKOeXEOPNuilyKbAM7oEz5SiGFV9+zIJLpkC/O6wtCDx
dSbDlSZjyHC/XPaly0AInZjjq1jX8/EUkdCSilgx/V4ltyM0WE3b/7FG0vwQgpne
e2wwCdGNzBRANJMOsh/DsKgyDR5y5qFKX7fZrK66a79QJwJjqtCLZxOmeOU2xUU5
/zgnMYNgEna4m8sM3u8y0ohQyXRHqtx3ntxj2VioIXTCnIeSp3mmOK8xvlygu8Vr
mkTNqLV8VwzlbvP+4O6vOsykcJhTp9JfZvROfd1h31eaplABll3TUa0aK8iVh2sZ
9+4EsLiKkYTKb3ngQkug5OeO5DCGFNm1AZudh4UHYyPdO4M+09uqNg0fl0uUToxo
SCOzAPI/tTvJOnwTLpALJpW4ewd2+v18gZf4/KeBDMNifA9ysCL5PawFWQ1i/oOZ
Jc6BjbYvAm/kp5KEgkeJWGriQzXWpWoPdQJx1irdHUXYj/Cm6VfYvCCmzzlx317R
lev+rYfLa9E0qfWfOcAm9qevLdjiAInKhGRfQmgElPzAFVEMtwedVU68/lXZaun9
GI/cmDCGKwnx5Ew0eECeCJp2ZIuB3Q3hBsA6huNGLcAeI9UXL4LpAEUZ0JgPxiYv
PzXdvFP/G3zFcNg0gGXTPkJxLObWBOtp+CE87m9GgVYdV8pQ4qjIVjSHxeBhkqDR
O1e0UaQhlF8TsNG2BV0HwN6gSYS1o2c8BNTMfjbr0oZxZvkMKwT5meQMfWTauLGl
XApMGOPveKMpkT6B8Gnw0MOv0QgzMKO5liJSeSL2OKehQPbold69QCjYI8/EO+hz
wT2SunhLYJCekvPNlSVEq/SygRhpdwaBpyMwxLEIsSE4FJyiLJMPKvsSq9Mc9Qu7
1DU/zOxgUr3AxGZEw0Sygs6DnuRE383tmmmxIEnHSmf1zCaFB2F7OfTxrNfv/4Wy
DGhP/a+qo9jaM4GRx6WRF5HrykgVfkcBH3P6KoQLdhcJEu6pWGy7oXByUoZ4UelB
GcTSzAsfiXEl1ttEpK2NhoqJZVGdAst6GOvLEy5hTzjlCsizA0+YC79SAb2Xvhiw
TeQFLgo9sPBurAg+gPsqBN4jvBehUXfqWdxULFYOdyKnu+LbOnaxK8AvYpX/Y/h2
XcIQw5iYr2WC9Qy6rlufMD2Vn21HsY0BO/Z6fLW1uvfMCc+a6l+ERS1QqtLXP1lB
cL9hmF0Ov3+P95F3v7A4ozMOW85n8U4FzitUg/h920MlFrLzoRlB3si+RUarB4VU
tligIJPiEwAIuwYbaU4wOhdVplmKSRL16qMlpTJ+9+S5bO6l3LyysA2r4j23uojT
8yxz/mDbL1xAPq/P/psVMHFWge24snmTPITn0RZNCAnnuVqbu7u6udoAGoIgkF/Q
R3uV9+y61eYLtGRGSqCVUyzyJ8Qsy2XlOMzq4BTqWelkUrXmJx8elRJW17BF6U4f
jwxivZduNxpnXaT20TYR/pm3vUfBaonrrEEStp3fey6hxp5uTX52uq1aGqmUWexL
ssh7gu2SZsRtMOUg7lC4xpyIqIOCoNpK8CjK+EBcQ4kte4gmpzSpSGnPXOjjVN/9
MgtXoZS0BYSETO8hKnhb48PpzhwKvnw0GNNqxJ5FaQiDTFUznXnMfb3FwYSYJw4P
ETPD2vJfXyzOQz3mgTcU8C1T3iylCeBXdexSZp31nWjPXU6kh0F3M9QzH8aIdiX2
eMs2+XYd/PeWcO4+itUiVzwVIhlTIVinqOOO0c4OJlFBoJYOnEJCKpYZaa9ZuRzu
TbsMyBg870xJy6YBVcCFr4ZK9fLuJWdqiAA/ViBt9k29MEzsFLsriS+7mu0tcBbM
TO4s9Dv/r6k54yol+Je4VkGkc8tSSXr7N3iZ8C1hSxHYC8KkWN/4OqJcWRoztKWY
dy1s40Ct5SJN5zBBR+n63lDt74EgDc4X0utZ+Vv46V1gjJzr96MTFinYi+cphff5
mP5nKZ9/uULsIdLeStqsvDhfsphrPXpra1pBIInjqwr+AmZ9Fl0fDH40SPsN/5PX
ONoJmSevjR+uOk+IqBeTUBegHJ9KRg9xEgfc2wQOQKjTfGIDaNQhU9RyIFsw9E5I
AxHcDExHTLBkSi/CVcsjufYK/D2VZmeUrUV11GYgdxqYBIScXyjHcdHzTHM03hjk
xGmTtfYsLX+cI5tjNxrw1VXma6QLrWkNja8cH3btt6bYuaxDlGklOFc54KCydwUr
Z2QsMXSfGl4bpjnTM6wF3CYbLX72wyqSpsI9po9IkAppnrYRgkPPR80OC0uv1Vt6
Fyh+PMBE5SUK8QNjx+92hTfBPdu4sQA1aZUepbFAMGsRsfeEZCfPiZJuuQ5gQNOR
jVpBZFBCmtx2JG3R/FAGivPZgclJPcRax0ni9px4v38pfmhHZswX13EG74iqJH84
g7ZlpzrYnt+tZuNX6fIWqtGpDtPySm5rgyjyZUbIkJp812RbMLnE6I2CROS3W1yW
TuMRLJHrZncRG4RSzaWwSMgJ18P8XDyC+mae6jHw4wmYx5LrhXsvIp+5W8WIVa5m
8vLSavo2CNzEDIUe5CFIF494HHz8fO5I9qPecYT2pM++DjUURNI9G27A0IfCTyWv
/RZvxCmig1r0ocLLH2cKRazfGWItPMLU4AZGpEba15RPJWtQQg3aPx+ZKlcA5452
nvsVByy9g2d26NAdA0YLednzqaCjbIHhR9vc9YVG6Wqo7wDK4i/h/aklvwkzuGRO
M8tV72IKJzkSrvmGItQaxRifomnIz+qVAFxaWCuoxg5eQL5KhUnMgpWZ6fzTx5dE
5Muw9aKYXGbWtmcXdbkBHhrB0XvTBgSk5Z9Dr0eYcqFZ0r1yLq5QRQm5SQiGsP5U
tSP+iw4q+NwrkvjbGGaqVPFxs6m4gXU+VPAPM9XIl8UD6DLeuMI1cm9xO7ieieiz
pOCgcBI11FPizxX15/hHPXuwOJVO6WXjuhB/HbUhcwdnGM34o02E1bov8h8c7mHt
HkBo3+XOR1cPuKicdGOcN4TCYyXhZmgzgwpVrI6SOF1okhkEhJO4p32V77PXZQvt
EqLhfBkkvCtW8VTwiSbn7AKCtBBDEB2U9kJjjplsUHkGf1448MIfZnxhZuvr8Bsu
zksd39VFjGShiwU+VkVG38WDDG4cu18qkSC1oR0Xwu0xSwwWDwetbkzGZhZU2paW
MjE/W9myvC+/GRyKrlTqlObOOC+Om8H/iE9nuUGjkJSLkqnJ2URd3SIwi7dxYk7+
eKl5Q4q1YytX2hrm4TMualocYsYqaW9HqUXIGxhtiUMRSjkLaUFApI4B6EiLkrwv
hFlsjSDYeoR6UVX04epFD+o/CVQxVfqGDCavV3i04lkbpa2kFprwXkyDH3uVcAMl
OqbSfkFFJnBCRKojcyOwWLSWxA+vdmks8nH/rTYnAU1GusA2tN/WdxEZUfru8SfC
lIiN0IBwq42IQTjurqnUJ1cj8bs8ky2SDDIoqTjJQk4fGf+R7NcndL9iVBxs4eE1
SHBG7CXlAv61Nu+uGLx6AFc2h9RbBuRgqy+5IpdkejzUPOnS5DGp9Y2MOHYIfQ+l
5MGOoLJTtAVV+T1QC9FzaCSiW4AUBOI2XWnWMh/0XwZe6a90TPGsmuG56XRVp1a6
h1KTKarqf0P4RTwDK9xUgHG2sUYhpo8voskAiVdXpT64D2T0O82gsZrj1FXhaGO5
9OLi8vY//pCEwRtuk/+rI1gzOdlEKQtgueK4Slj+0z2ykOmKfL57gCAN1+x8SrJ+
ENDpppEa76ygbbweZrJCXv81lL8DhpSeBesSRMshZv9OxYClUHvqcWarVhAkrvpC
cHuIMGSFR9wOwWNMwEj70ZdfeZFuBb7HkG0eU2AR2BEdSbFTqTSZhUIZK3c7Wb0w
IhD5u4PAez3Ev0YmFxVkI3Mw0WIVCuLW5RH6TwzU4SyWkJTjfwgj66ArYuSGfTXq
ckEZ5up4g3Wolo2/JfRmQjxSxR0dLnuXKZZDIhIfxXJTCPtkfC2s2odQKgRSpqEY
zm4YJ3KgLJOaUDPUbEdGp93Zvlb238RNIgttoDJC34TW5P2XLYVYkabxz7DZ0P0O
K6qLzKfboL8M1nyY4G6iupAuOLiagr9eQ9nZnJv37EMDXhOVS3t2xwQ1vA3qG76F
6uBIozZiFSydM4LRV/Pli4FxRpmS9kf3KZAam82KG2Z6T/Gm3U5auL8XW/gouLpo
z6SGBgKLi+nXo2l5kR0ITD7dQ+iJJKsC5WQ9k+9e3KFUW9tTJzK7XWmamzqiX2wb
02PzxcHU9SPDEwIhIXtS+4V2WVi4fPjPQ4Uyovp7Zo6MM3KePbQqUBbVOgBDYBgo
oPI/etaANmvGAeAuKCnI4y/t09+zlWOy4Qg64Xx/6Y0pi9E0LhB122UFUwJ6eGQk
ZnlShAaZZYDt3teBwJWbJAbeHysSi5CeqlYSAVDZW7Vu7RNlriH+uZzmIL9SF9qm
JFJgZgCymdA/dNewZBpCKcoDXnJoLhrB9JhKWUoxFVliJ3+P+fBEwjOZwIVgYZQ5
BivyYe8YnlQVXquwIWhKwt8Tnaq1dCPXnqUF4dkzUIAzZjVQsHeAmWgMsyyxBH2M
qGFh2j8OFVeqcZlxHFi8JjrPUWqsziAo+cMfr5c8gOHZIDj/YHgU4oNk/oMWgA2T
hcoTU4bU5fvVvqXPnvdQKaOUwa9o+XOHNEYlAtzEhJ4ZySG13WN6pJB8mNfK8lFr
O5hfqg5PeUAbHs77F04nX+MYi/QqedcOWzNiCdRhK85DQFeNZpch3tApJD0+zKho
ZUVtogscD3Oqb4pp0P1PBn9RRkyfWFvrozZd4PsIzRdbSjE0wPAPejEe+aXiqaoJ
lk3230A5L5w2XNLIToZoYw/AvdKQ2+Dedb9ZQH7VohNLWpYC6zISGxYFyvKkXj4b
1B77J/j7KdtT6q42imGJFf0zB8InG6ZkbKrmnB+Shb43MyqcsbMXi7gpQ9Q5UfvT
mTFu82GoTuZufqQrAYPF2hSFrjClKeJmkMduynQVdGtMjLz/u33aShgzCOjXL6n9
gBympIpVsjNpUcavSwn1LuFdVsYOe2xvoKySe2gLiQ7jzpDc+tnhb7oTb4HS5CRv
/dYJYzvhiHo+KoykjHuuKQB1c4H0vVb+5wUDbkqvxheOjYR8egBETsU9HxQmjuO3
COj7vWTFmdf88TBUYxsJDoRzq8Wj6Dp5zhLKe1VbmhDFD7CVHGrKphp4DTP511+d
z7xOVmEp7pxCN9ubk1S6l9pz6rgEqIREpMnoMjs0Kk7aETQj7AzXaQChfe0b2MEA
5eWedhZxDbrSci6WmUmySXwcL5RHnIWvEir3JK+3gFM6OZs0u0sJQgEYBpZ55a+m
XbWK4yqFfcoYAeWENAFs1sY5mwQIZ1wYqxM2FJLhYabym+iD8T4kVIqXtvMxu1a3
pDZ9d4XLyeC3dw02WFEHZUP1e8tvIYCd6W4koGRdkJk6iIaXXkJFlxSqHm3wpnwS
aguABKcy+AJ8qWb6ZTXeyyLQggFrPBvSDJJhx65HzJbyb8I7+dtJPa2QI2iFXFHw
tR126+9kJaJ4dGWkY3Z/qGTtyoqFBILkvi2IEZ9lvpIM9hfpjL1NXlj+cBM7CNah
jEymlPPt4y3J1U7G6vL1E3q4e7/onKHry0LaX8JtBS0P6/yVlqmV32+71f0aQFsJ
HCpuukhAT+dEnTCUGwhZk041jWPQUEjD1EbR1cKHnAYRqYD0FHi0LGdRz+kXhTTV
DW3KRnjgRr5NEFreW/5gZ5YGSKGCHTfQog6VFf0NfiC2H1h3OGJITn+HyWDkTPno
j5LBRut5BuGqgbcUfVDoWFGWDIPmDKuYDI9mqYLX3G4icynYU/jdKjHhi0ExKW/2
Y42OsR7tYI3aVWQCNDIGLkYs39qRCFuSBXKcsCsl7EojNHrKuWgz3NGBxNlBVk6t
FgSgH4U5sSJ8nHQ7MD34sho9T5DjJHBzOoMZVfxmeVkgj+NgtArl+QMEn+gEQo8H
qha5t3FD5Pr2AgQZjoDXB+l4BO3dr/nKOtYxp1LOAspsEhPS3vsnqKFsv9KJUQjc
onZcq8Rm9cvQda6H4yqpg+YFvj2J4O277BHcoqqjx3MqPzDAFOBwhoxn3citXYWk
0phhVJkHHFaa54tDO3d4ultPRUi1CIikNdl18OTRO6TLlc3QU+yPAHJUEVSFWkiX
EGbh4ATsGCn3GQNJC+Ft2AgS4yHcxLXuKOBqne/yGGKxJTVTDU9BqfkqwZbVbgwj
bCS3wMOeew9Caz6TJh6mQGXj7EmT4MtQ+TgoWasOnKHqqd4mKyX4+ZvR8TO0F2f7
s2ajQqb5CoTxdh+LYEhaPBHz2w8D6DCe+VAJi/X2BDoOXb6Us6HpPH81U7bjSc4h
zUmglD2njgJDxocwYANkNWavEtfY+j41tZw1bW/pCMOa2I//C+N3YMuvqiA1fnOU
JTxz6BFNliANY7b9vplOhy+hFs598g4PSGacfwslojI3CkxBhLkusrEhX/XakTa5
Bnd0BmGTA6qSY5YI4EektQk8dOiuM5aWEBHhkOlveAL2dMJk7irsgDKAOR8Ig8TO
GJSf1x0fkCYRWFl270k2O9++2fZUuzsLAmsPG8xNnFtpKcx7xo1V4OvKl6arG2Uv
ccW+ZqjkZE6C6pobZ4nc7zCZiWWolSwcxh4bYlY6PARP0dRVzVbtAFO8WtGhsa/N
YZl88+a/cRDVI5lSqlT8OeHIPhNnUc3gXlXGfgE1TbpbJk3LlV2vjyEGQNXw4cgC
LrKCCX69neyyVOlrC7Z+M+iIDYlwqMf5n9rSo3PkPYmvi80MCi+EC/NqBgTrQGgM
G7Rwh0UObJrR5ANmAaroPDk6Vaiek5Q75XC/VpQCYeNsoVNXMAlR6uOtAI9mmBmX
fkwg4xTFPgldAJIaUvyQl8Tsf9iArDgTi5SBwLdHYJUEe2emoON8xeZy0Ur7DZQy
pwkG/OyRE286E7Zs8ZyYxAZo6R6O5zPNV9a9eid7h4isMWks1CAkhY9tTDcEljPA
zexCG26aqLBwZ9ydB9e/gxzcFuXSWBwMqfVpQiA1458eIQlXLKsB4MUmJfPIcVlM
iKPUy+tZhnR/ia/hysydoZa59yE+3WSgIj1mCRZ2scLXi2/72TPztgpbmloer8zo
8+yuhmJihpkNXolFiR4FlA9QvpPzs7isv12m47FeL2S5Gay0I7jSm6wBt7Q2eEP0
TVgyjRyUzgTBhdTpK617ju0u9ydp9CkIBre0f0Rt8lxK8RevZUVKv4tR6lTl4BaT
7FVcXiPI+zg2O/Oxz2c4FmmANvpbZok5JxxaQ1awb4tSP5PgTWudSrB3iZ6xL0Wf
3hjBHy8WLIVFEDi5/5nhIyd/dO3Y4CmnRBzIHKHc4iC+xNze6k4KzPf6W4qZBDzD
KEMkXl1eSht0tgQfLDVLcjE9R2oZj/HWFVPaYTSCES+gc4IFGcg9rw/dEPAsJGf0
07EbZi33zJaUubB7hgfOmOrKbRWSdAS722qysXalaZHnNhYVwFr2rnI8nO7Ksqzc
LzijqTZ+fZMhMmRp6caFe/qedcjjPooL0IRvLcmqh1BfstxYIYR7wm4xvH+Wc+EJ
5Ad3pLCD1HUDK467TO/KQSzB2+WWq4D6/S95ImgFXMb9C56jHBBbQ4PRgN5TDGGC
iOdmdBX/WdWPbBRqAy+zE/8GKtHRMrWtxfHL2TlGGCrPwc8Qex4moEds91sFZadB
+MR9XNintLY6VpOAQyCLzvRsa5tjlVBt/NNDiqBkJ8GDzUOBcGHBBQE65p7ZP+ex
vUMF2D4QitqoE1JakY2aCpSCRN5z8vX15KqY5OdwF82d/DvTkMWwFHy4xuHYDPwc
vfekmY0O5ZDp+L1YbnWTnKSZJBcxQxcL2eyWSj013+0F20qviQnXgRamubxz+1pi
I1lKSH34Yl/2LLBq+98ImGsVjZo50/1Ksw1hh61/ndbBQbSLRwoAur+1CqnTs6tU
vM7jeeylEXtr06Sz30cJUt0d4+yRBROvO7nU54SlqSN7SrHimFlYuD5cRsuHFmJX
3IPj5T3eJFZtb6GaIz8r+0ZrBjfwtl26oMgL+JszhF3HlTauF4ue8CqWiLwJpa8t
oh/kav2/KNymoAjN/1avCLIqtfO3m/+FUHDcJ9aMGozfvyJ47LWNnCnt+46feiTi
ysSBgNrBUIA9Ed4ZAWNA01z04saTjTifADiyyWXsHXi8179POhkZo4hiDM65uSuF
W0PeQy5oyna3WLIWSjDxzRZasX1I6oCTstTgM+LTJbHXDebVwd2uHBokn79zFGAI
6qjUlEXgpXXgIpNSY4tt8sXsLPgioSAXHk5YsNIjJXqZolZn3bV5rFhFKAvnvc12
SsvFMoiS/gW4FpY5KBk4sR709bo/+vF/p9pRxCLggxdMeKIr+Gf9NIvAnPBm3Zzl
jliVle6xCmYEQjYRO8Gqe6kTNFRtkmcJIjGGkzjAXt5J/P42IMPZb0J2XU3iDSFF
X9UK06yaBzkUOSJCIPIPMfyV5TRwzyy1er9v7+yusX9k5wNXCg8vPZd88Clojur7
qujKqZET+KAE3xEvN1iBUOp/kX5bD7OeyMfkBwcO7HZ7rZaXaMjoZBjwjKDOoGd/
bkbVBYg9KunWeNIJ/h8axbHLLR3vivI8fgiIRN6JftLhb28hOz1c5Kqm6Bw7s4K0
jPR7oj9ekO7e1Y3Na2DlcY63dDPFmk2d7vr0NSs9BimTIyfAgVv4VZRW9KXAUUAe
57wZoB91B7DXHSyoXQa9LSuUIlJ9Swg9s1ShhoFTTo5q8hfUy366Iw75q0EZ8R1p
YEQ/uiZcItZdeQmPXwO6M7A7bZUHkMyBZsit6pAwyFc16kJa1DCuAc1xgoaYqK/X
DT+kilwEma6WLG0YulM8M0nGOlzSYxpPVEWck6GzTpbgIXGOUANBXXkWiY1qMVV4
1Fjlm4cED3S5DAgPWAxLycSY5zG00VBQUqbNHBxpgwBiQxoNe/kgCIHsLandJQyG
tK6EpZFAuoMewNU5xAOq61dt2/wzzlyjrVyg13ZGPq4jfDkx1/yvjCMHqvrQAbq5
6JWR1MR0TXJElP1ApJD1+c4d26Y/fUZ1bGJHWbs6sCuFLOhW7Ar9Q2UdeKK10LCA
koQC8oqB55jJBneWfbzdbal3F5v+wWtEEx5Yhs6xC01LswxlN+lCMZ3YfKAQbTiJ
E49O3w6QjLnhCuIOkdHvVf4mMb+8KhGt4rSuiCtIuwFN2F7OwfQDmC1JpvG1O/5G
JtGJJNBREUtLP2EaIb6NUlN1lock1S9ZF98FGd7PqKqaaBJC5iNnwJxjTabaSGVC
jw/4T12czCeetzdVaQMBa4ZusOWaLYhSFE+XC3Fhc+5LiZAwL7LUx2iIyJcIVSxe
4ZJfcevDyFvmyb6ya4RE+120OZoPoyTX4OUDzWNhcfJys29Y7COEaaRZlMbytpCf
L7qGlBC4ouBoy06NsLk10TULuPVRvYBx0vn9cKPGPNv9GDl9t5Wn7W4TOjibngAk
VWOaFL5HidjXXo8UOw4s9jxIIt3uWDmy+46SgDZMYBwljIPLmr0HsZnI4tgki/2a
24OFsST1NHOObobeNfm7xCirzKsP5C0XsUfcYkOG/yIk/0FVK8Y1swEp+izzVJ/Z
+JKEft0vBWBepNO0+mZsHu4MFAJ+c/4fB0QIejP4OvWGEDKWk66A4+3ZN/7ivRUj
P6qsTjc2VfSgA+vkngP/QWt12QhaNA7A7CaSa/ORo9IAfQA1cSMonPh1fqDMTNI7
U6PEiO/9TGTUqzIgRTBWPlmENExbtaonJ3wfqCZrYMYLrqHcBUJh8fzp4q63uJwa
APVwAKcf6dr2nMsbSf5Iw4RTazpbhT6rpZC+MjJai+csmc+NS2YlfzbgUlf+VyHK
/742gt7xhYBkBT8r8F6HZGXJL5AQif4P2FKX49SDQZP3+e+1eMhho+1SzXB0DxYp
YyNXKVmIlxbKmod4b71Wwl4rN+viGkv2Cckm7UO/hgo2PRlSJU/2LwjWbI/xKJPR
8dNeVaHApTRq7y+Y4sDx2jKQ3rgGnf3Imy1R9HsKNuEt8FEKYbbNqMcCcOeGjSu/
BhBpzMkJEy0gzs9x4dUp+nwkx74daVRSdVWSFt3HTTg2fSbub+pQCqK195DjrKur
jAhZpMosrWgYUzwNYdTXQE7JZDPLVfhXxBtVwhRDjSyVMp/Om0V6Pm88bSVw3V7/
ynaF6X4gpIJSNi0fp+Z8OtWPwwduGeyGKHAxbaDPa22UpLSWXwcPIdgMUngQ55Hj
oK0rK3d0RUejZ1Go0MoXt/ThH13wrWfmXTCXGA0lcMD/OT83c0WU7QRXXxcbwGkb
DkUyhu1mDg10LIOMXVN6nVuhdLKbzIF8udWob8p5Tp1DUGqvDg+4/1T5hc/aOPoC
GnrgGGquGnbSgNMpYnl+Csw4SvRCcwRLbQhAXE9nBDCqBGmbW75EZBDToy+I7UPj
hM7zXvFd+jQyCyjq+pUG9ju2lWt4cJxp7HkvNme6noQbT7GdRTj2YSnce9H0rXV4
H1w2Ch0kYC7LiL0d8W72wTwEehDfEnHPqLk/fN5ImcMQ239VKdr7Ixp2CEdG1AMu
lpdByvMOmoxy+w4/cz3do6ECz6ggjmQdHJcce8lWNw2/UwwgKQ6AIAG+bQyKYsQ8
xRBDZzXOEPAjjZFJh7uJAIkOM9soBLPLYCoWZvDhscVM2XSNCAx+fbONwR2cjkho
+kXpe2gSOD48VAt9jwSjGmaVzKEuAqKsxKKYRNOkvSTTZsKFc/EB9pPHjU5MffiU
jqvUXAeiJ9oVE8B3qqA1p1pHpJxt1tTc5UPjUbnboO0kftC5CLiBcs6dLlnpcopp
8hWiHt9CGvldBFb4D/3XJ/vyYyFFNo95+RmtgJ/qk1gMpnIUlLsU15sXaqL+QZhT
etzl4heX2a2tpRv2BRScK4zn3Ac8BzIy04Wfgik30AfLy583TARkI3y3on5HPZca
sq6cUuF4a1N3lgJCwsQ0zhakjJizHXWL85HoQAE4bk732VoQOyRkEQFWZUCaQPO6
EhfAcC3FBcrWU+UFxD7vNipATT4rdWBir8md6oEvMm4ov732/+0FG3B0vPx4W+zl
cHUlDLwPmkBigBc0RteqQ0PVCSdkM3TYmNSX7ssJmxi8077ReDAsR4WVzPTyN76k
XKFI+qETxINamCSdN3CxuH1CD/YEuwQA5FlGb/K/1eGyT74+eSdkkvNW4fp1tscZ
oUNiYF1MkWkDBA9JIhOjtkFSlFZAEvv3ooqU6SeSGgvFbBcqWYIbdrS8zhiGB5zY
nVKJRgmtO8/N03QkbOHDJlrVI4OE6IoR3l1WLwjjoOqJ5/gYtHNPwMXuguVdd0Tp
8aVm4SJnc/zpnSppZS5aAX+bTaRIROzjvVSJskLhWb6h4Z+Kw9j3q2OF/SnvkPqr
tuv8ceCms+mABjx99CVFtOxw3K3ruULhEezrMqqt2YWYBv3MLK1vld9F6byqIQAt
zvYj8zNMQ7m88r8uAK7JA3fSXmUcSRui/novtpDyqmW9oUO6uI2ZOd0WDt0B91Ij
WCe2HO+PGRtf6hfVMsG0blP1si8D4VDtwjLDUSEtr7if8We7Rd93KxiQcjyWsdcV
0a7x8xQyGtKU2AsmlRJSrZsJXOKhQsgzHVAA88PVEx6sNniN3/z+jK+89zD0zUjO
deLXCAfxww5pYY3x7niZMI9O+tPGrYFBr5d1c2l6rHSjNaOo+/jWTVnMCtmgGSoO
jHS97d2Ykeg1VrRfUH7shimgyOXGjJc+9ab8xsRB3UEZ4w3Be4Ue/ELDUqsqGv/c
2r4u/r+HXkHscSRnbm/qTZHMgMUxJy1VsycS1Sd669K6wepCdBsR5M+VhltFb8GX
cadoOW0dh92QHidN+YpzHw2tzeOcq/X09hvqrthqyQ0IDS0FJYime7WJa1TBhRSG
C6OJs5iPUX1JuzRPbMlIQ6kV5qfp4NNkiXHdzpvcvejqhrBxRrQBk3jznYYDFyR2
jHLQFnb3yQwEMl4h0nALyKMZpwDrrv25ntCDh+3ffP6iXpzMJcD2ZwPOT6pul7QD
5Vqy63Kz5ApQe6cwWbY0kZfw1Aojcl0TM+ia719nUCBo7ao8bAK8br3/pQlgiYZ+
acTP0T3PIqsNELe/GnJhMAXxF2FZ/lSQx6rUmRDwQ72UMrxQpUkQ28zHxn0KN5Av
CkpT+VFodaUp7tm6TGxARFgWU+Lxd745GTZsQfP3yNHQXAkBct2nAKVC6L03sUrt
Z4VxBt+u1MkUr2lzR1UM3+aDzqAXDe5u1iUj+WwsDpXva72ZCVgrbbiw/Qr4pLKF
9y/q1CqrdhHq9xp8XT37LMln6w74W40S2yHXgd1WuZPFpmRhQGcpRfQLpNCgN7c2
lGGW1BPO1CVOTlrk/qHBe2qq9kjbuo1svfJBSap2s5evUcBmutWCbej7Te10DXty
8OjF4eqTzjELY++WWEpZUEBLHXEW0NaLVNPfWZGxvJZE0kojjIPDsxmw8vfDNZGn
ZizOqYhn4JQSqBGncpj/eMlLgqxbrxgbeyqdZMdR3qp2DDmUKSPcgw4Ciuut8t09
ifgXewtpaJeSJLZ6ieMTVnot7VPEREbhtxMNiKj5UOEmPZytUBYI+/Cx2noSJv7B
JIjhgjRCliIr7SRc3YQ7qgRwk54n0cTvmBJ7m7Y1OzOeDTA3lW93V7MXjmIOSxuf
RJJBtxXJNJE+SkV3oggO/GyOkZf5tm9N0lgEJ2QWh2xbsTlA8ImhVLGrPnT0VdxG
OHbe7OUHaNeqODWxO6DSLJYQs6WrrEsPOSLOHJS/J8cqiyRpnrSMKPNyLPR2dBXk
5jYDmi6vCJKATUny96sAd2W1k22EFikMiSfXuKwXzElcGihJlb+/Lc8ivEIPY4EN
5iJ+bVAc6MFrFVMwKL+dTQoyAYn7ZLOLa95dLiz3j6yuElzMKXGdbdVGsgFpLcZQ
Y0/g2hNSQJ/cM5FvdNcQaKoBQoXhalmRNxH6+hZYVqysa4y8jAbYJELzlGryGoLF
uxeuF5aLO50fKi/w1g6bA0WHg1mX4i6nlY7rDn4XzhtXCIiocYgcwJ/xa62Jg3+0
bYBRrqoDhAXkpkqRKYIqdlBtQOeJtJ4hJsM2NerGqUm02cy9m5sAXh9uVtEFCb4Q
h3R065VN170qJegh49Ef5W/Lj/kxgDAG7B050woHXFj9FhRKmB8j3eKjZI1BSHq6
+ZxYXVCE8I5W5GheOo3Ok/E4KQVTC6CFhPKAeoubZ8CSnsh/A1ojJoSKerUiwYXT
kXwvzOtkjHA7QndZTT1zJnmmJRARNO6Im8JtpPIeiGeoKyMq14r19TAfykHra/3t
1mbL46k7tOfasmegQuNxQDWZ2K19ratdazymGt/6TVAChIpJ/6v2LM7hZK+uS6aV
CENeecGGOnEueZo7oK8AnSHAvTR2CGyodOrg0Rb+2gU/egvfCn/1ojD0rptZ8Hbt
YZ+l3/s4QxSj0rNY7IVTGf6Y91nQTt+lJ6G09b7B++MWeql+81oWw8QPGxuyHwra
/BwXcaadgz8Uncoak1CHi6V+N0CT7qPJ/ThXw/XJ/lDcMg3/793r5xumWdyP1inm
ZhW4qW7cgyNQGgA0vN/1L2GxXKuwZ2qTDp1Y9AsLjZYlEjklgoYeg3jRBlnlIgb3
JCzsa6l+0LW/G+7AIS1hIsVHAT1vMmuS6wU4v3J4O0cM+h9Qs5enkPn7E9XfIA7B
ZlDptHOqKuYj0MXm+rCICbWsozyyMcV96QfYWycq/l3kv3ucBsdbk2EZPWb6zwJP
geiz0aRJnUEbIvz28OaJWbkbkbVi+lIweHN18prVDQf9e1G6QSKMGgTl7bnGtMrl
DXdJUphlWBDy3UlsEWJd3dxWwko4F4Ai5wlTAATwXQRAKFshudqrkOYlZ62Bd43s
5cE623AbYr16IZ78CnmhOkhkBkzAs86ITiTxtr8oSzBUfA9Hyl/oAiLsLJ55YdbN
V+hj8hVG4Me4znqoMNYFVqHhj5d5DZ8NXj3gT0SSTrn/1WgeqS7kYXdXd6UmMRT/
1wKPHKTnm1dMyV8OhemuqwHhGONbyD5i7+ipLexn3zEpW44SKwKeoqabO1wBTpyt
Lg8J6jmR5E+Ic3YR0/IA4t7PdGcbOjLJt8xKHHuMQuGU2Gp4Fkp0gvFymMn/1OTJ
+Sf+Znl+Up2Y1NjFBAE1uD7mn36lIsGA4EmOLcXxVjSZ5ATAC1bHJfD0jtYk3k53
tERoKh5XxsPDrLZBiQP617zSv8qMUBO9zaIRrOlySVwNcDTIFsmV5b3BmFvmZVEJ
l7DrcYQFeal+VfmDquUcxFD7yyMGzz8wBM+Rhn8Zta+BX09/9zBMDQDJmt2kT+cz
cAVDGb/PrnfAxo6mGCpWts6df+SMj+QaSrszB6SFheF/SoWW7H6JVgnrvFcPLBgA
mqqi7bFFzV8ol32oRAS+IO5xjJ+XoeuTid4VX8tfEFrA6F3R2/KKJZ6tYw0HnCKF
HOzI496GztIZjRx5XpUueyrPsxtgLCPoH7PttXW1d1cQhtVonu9rseO84MoqcW5s
Lkst2Q2jXuOT8rFd3M4SNI1V97LiTjRwDO9xwPLy3K9WFUMuzMb7uYN+qG1xFUh4
uzVaxEky6lyyZLwFJ3TepH5eQr6EAwwrPR8jF1RgX8DPfK76tmlS6Y87+MZDutv0
CHre2cn8O0wGqjsZQjbzXKkam97dsXJnf2knzmNELR0uNPap0zkYkKlV58l1HVCd
7l7BOW500wKix85gZg0jdz28yD/LXrRSFez31qWZmjCRvkc9bIV1itjP+8pVquK4
RJs86XZ1msHDP1FfMYrsvL4aDkoj4e11UxIjVZXDrKFZ/Wy1zZMrOKZsvp97XVyw
4aIf/r7icqWXOp29Lsfl6loVdnbIy5jorROPKjoDxvL7PoQU9VEVT9Awx7AsCqKE
s3/NtPf5R7abA1KsNGm61sdiavbbFG8P+ZPzBLrQgU7wqOVNsQbBMwc/8z7KPwW1
yvBeDHLrvhhBkstf+wHtu6u4Qat58J/fzW23LInbvBwVwaOkIimUS8twPFYjLf6x
MOhSfFyMR/mGwFeEIztJaNC2M+ixOenDjTTIkkqzZbr6UmHVMcIEKUX4FShvTlql
ASiRwJnVfRmp7Ho9Su/iveB3fd8G6/BJzyEcD36IHGIIY2q3ST/ouH3HnTsHp9W/
L4KcJIIZ1D+O+wp370v5Cn9DbwYhpgfncvghLFuDNW9Pj9JzF11AHi8XwZeBEae6
UMjfqU4U1s4/Y6QKTX/1VmSPhp2lRMK1lfVho9rMIVjmVbgUrsUp+zsFNYRGMyp9
fDbqFji0ChAbvjbWHPV3+hQ79QAminsq4ve1fqbDypaBP3nIdOx+snCiTdPRKboD
4kgwBDrKLpHIFKYdBOS2N8UDD2A6CUsUjUaitI0WZrLF3ql8dYWcDAiLtvwqsw3I
Lx7GB7zUXj1s/Tlu5dtn6WTQvGsF3jnmrabVkK7XieRGqUV8tiv12Mr25Avnl+7a
TS4Q8RiVH7QY1wew0MQaKM0qiIJ7Y3bX0tHxbwuxQ4PiU2VMoCfvWpiul8co7bYA
BR61fe1hgTX7p+X2tMmq87zc8+ZPaXXVvTkAHZzGB/G1cWTcpfWpsjFNFygEbWi+
6gngdWUgRzIcaVIe0cQk3FVO+Q0YdsbCeuNPrgRR2YktwB+CuiHd/ZiXbHLI8t7Y
1gYjzVjgGyFFX4bQh2GWleBECJZHrjJZpuT/VpjRvLCo/wJqLQuN2zXhqhnMoC/5
tJzLyXv4eOCqgkDh3OW4+GGY/FUNBK4d7bYN9sXugvhwHgeerEuc+eesKASzdaQ4
sqgTOld32WbwAJljdI01b/J7xnhoWrJC8QHCT1J+gH/yM/Ur2LHNHchz32yoHaqL
vD8FvyVAfHVJA0Np804DzdzqYbZ1QpHXrxc8zUImUv5bhvur3uBj3sxOboMhMieH
s7+0r5iqMUyD9laMtyyZx0GaIS68V3APHbYh0R26HyqU8pnvJaD1K3KEMvoXTIlh
dgIuAUyZ+LoifW24VM/TlYsvHzgoELAJWFmXvrV63NezutUb2SCbwB0M2IfGJNmC
ezG5K6zELGNMasu1d5sh0GRuVAqsXuqyPLriG856Uk4FUXwQBPxU5ZCdBEXGtmBs
vNJpNApS2Wvn/c5pZ87pSoGgRBDccwx2QxUlUvts2pknxsLp+BcMt/cUlQ6/l3Zq
OttC5RmsqQhY2QY8IoKOl598yMq4b/bW0yBwn51hLEj3QIv6+6ox6kFVIqIcJdEk
Ye0T2SGpqsFPNRYcZHgMhGNHy2HNEAi+RIeZTDF8VjXTbePyOzY2lY7E5Orb23b6
1+NWyhW313YrOonHCvG/QyjRpVscHhXCbZCg2E12ru0LsBAsbzeAtOshcmCzxmnt
D9NFtc2bdvyCSfFibdra7RBOkozf0PTDq13Z/Rs3SZVglWbN9lFFZDJ8fM4LP8B1
qYRNZQ7p1joGxK5nAo/7kOf1NtmJcFltTKzsKwBbiNbQxMISEWSX4oGtqn3WDMqG
KlnetKHlkYyJAWQYpi/WLlCsSa+QCv1WtiNVnuXv6QZH1UFKy0IzT/jmTRVhCGL7
a8Fjez79o/DtBLSxDvY9vhvmAW3tLYxY/oMdghKKN88HD9Ey/QquCrd2fI0Gu9aw
bH2L8QCgblZ2FT+LK97zUlUyBLKFfN0ykAGgiFTw96wPD6Vov/Mwr859ERTMMNTc
dKTane3v2q+U5NZARRS5dNMsDxnl+4aRrqi5O5BXzZOfMYerbCzGXSRPFZgNDlKa
1gmeCcsnx0igOIHym77cEz8bDf2zdwc2Vd9T6YQtPya7FxWHqQCyD3kqbo8EIo0J
MCxqH8BnAyn2uFUzfaVvBvzuBC2kY3gNG0hd6ETobjytHwtO936AXDGTQ5YSlGTN
yDZQtd+rJPbrLGnl0d9kxL4sWnZI/dsI89oHyWyYaLxmFWbzbzVllYEZaHcVzBl/
qAI8u50GJcx/csy3Vt60CiIBfuD4j4EZCwx+65t4eElUtWTgEc0cEPBmbHu3CQt/
h5Wn60ytWHAmN2VLMYO8up6lJbidMtwvJ5BvWH5mb/eykqmLJU5GLJ9lC3qJainZ
NNbdq1bxgSu6ua6LC6ka1dGC1EEXXcCb1ezq9axfM1/Kl76HdY6nJOB080w14zJJ
bFWjB7pGrh2kemrDpUXyQwyQmNLM1jekByTuU9Q9OLYUAcPrzSi7fHoIkSVXmvtV
fsWxlcO2rt/cFJApwviyFnfQqLkYzHF48QfPMDoILN1paAwjeTv4TyBnOcKao6YK
UWu4IQ1SPa/S75JbpwK1yvKe3jk5gl1H+ncmE6FscchHt5JoO6SRzK+4wWOnshsK
4zRzQHX+/ejhAXSl8zTrq6NPnq89NOXXD6j6XAjt5QWteDfgBgkdQU215BpyVPue
SsraQnfSvr2iFyTGNZs2MXn6CA6PpVJ76Z02mhjovqREbwdwtGOQ+IcY62uR1D9p
UiviULmsCDWIP6cR2ammwHEmtJq2vFVeYCbpDXtCm7O+zKebxv4jXb+zStgs9lBV
77bGqXh55+sHktD8VPzCZn1HO6mbAwFyfq5+RTj9CVGocWbnTebZNp2EqWafPLe3
fryU0nV1l5FL8qD9ysR/m3wiCIv0tmNacxCczeRekrpRcIhQdUx3vK8RptDtBmBU
HsnLjWxygnWsG9BfQ6+VJOcuVMzNoaR3viiBvot3nsHhB8oeuCD3/l0AeHQ+PjPd
4TV7+d1mo6KSK/pDkd9OmXZT7V1yQSXxnsnwD8elHU5mGLRjw41j2l9sgpRLp8D/
vnzSfJPDhygZYOJ3KE0uNYtJNUVU8XYHaM+zFaLQMo6xAkB0Y5WedhKEykBeMctQ
hvJLRXSbGWShpkQD4NRYi+Ng0h7h7Vprph9F12B8MFifNPqZYWekwXR5FBJLa5yx
+4e93ezPN7Svm4x07THH0sCoQY9K9LuDHuxYmtvMkwvOr7CzLJyQrkZUbsVcGc6/
9lnLNOfW188c5KyhvcmnS4fTtpQlIxp+PIUI3WYCJ8MpkFjezggrkwTrSt3sf+T8
EL3F5tD1BH3QiXg6kU3MJarFDP4mzbxMhaqzIsqfHDsGPJFZdo1uYX7OOVLfSZdH
RJ+Y7eJEh0POIhDr1dJGMzpuH4luCfnG0w7bL8rKAh+uYkQsLODvG5RJgHxerQTq
m8SB4KYwcJQew/gS8lJyv7mli6JG0zvwX+FKyfn4fkl6+rkwK95paXw6D/3LTWuB
VyyTQ26lF+MEhE9pjrILM1+7wq/nfGB9pA0s7fLg2wX+/eTfdQKf+1J8ym2Ogs3j
AbueqAQXIIcpN0L6VJ714gVpsKMF6Cv5QWAU9t122vNtmJJwj4bt8kfT4d5yaTr2
6aO4YRTAqhpDqgjSD7Se4BtG5gWmuWyE8LOKklELDMWukM2sL+Xdt5NZY7nE1Ynk
Pb6gQDC2LtKIqiLp3NBlu7OSQAf33IT1ADBj3JBjQAuIE2nRVlAvn1umvLKEzLIe
RCxGXME1+3kCi+us5IJRxKrPLtOiiayBTTo3N4wAxG9twxbHlUmUvg6pIgeXwcF9
OX7kIHrXHP0+moZJIucZtzddgjPZQLIvT3T9WR1fhrASOuuaD09nUr2mivHnubdk
dTGnzUxJPMv2DqT8EAfPWBF5Tpk9bpy8CTwKsE3g1P2YpyqSjwha247ZIF6Ss1td
1CEHhnxIrS0hcOyfHs8K4QuQyCyy7FqwqNhG4XExhByd5MN3irMNmCHLHeA+jzz2
cAqURooJpV+1zMbOqfJlnj5artzkhVlFxm30J3Mi0jt+j8WJ/1JvWPuHXC/QvcnU
ypSzrcMjo7ykVqDZdL8nBP+d1OhtSqSC/L8J1Bn4UWDLURL0BNgNBZ6mpgUKPlMC
tOLu7HZbQ2+cXNAlHEQOJa25JpeO9YdtOxBsQljTqthXZjNjYqAoNCpT3zfRA2Df
3Prv4438u4vM+jAs1ktej31kbmkYjYbWDUcesHAmvPEZdJjOJ5fKxOZQijkb/cIG
I/I1i9CUq9wGErQyrEeNP7O5uakdVF03Bq3/32Yb2z3kVVuF1QNn0HuDspCMFA4l
iLDuWJpamOqI1FOTtpX8f+59wCwa0rhgWU7CaF3E+VwnzfxPzkJ/LuB6f7v1FG9l
YJcyzs4uqiVYUgKKU8uRURluj6zCAPWYkTs2t/c2iAJhnwQYwCc2vnMyahJPUM1C
Ij8sI2dGBbeP9uv19IGrZ2qWFO+45wnyw1izwH8gixQtg+U75xX8N3QSBrVYjCVE
PDeclLxUnTrmuzrw/6jPk405EdZaPDRLxdIS85ImvFjT+u8khEN9Ko7vUu80UgPy
1spXF/Oh1EiGNstswcbqRe4yIdIEWHjM7SWiHVK0cCXPK/p6dpnC9ZPvZ2GzTmMp
IjN57nrPpMmX2MnSaslXtDYYKoC34wKIm+AyX0TMN4fL8qEgYpe+ErrPd+kKbBha
dxa7vm6ClUfaxKYv4GJnd/NRQ8MCDcqG9LN1DZ1drpMcHgN1T+52pm3ejkhXVkGg
SaNepLox29DVyEWRrz13Hc81e6b7V0V6UdtQf6Bd7jiRCKEx/MZqrTrZmbbDZ1rI
umOI9u+MEEKWSYCoXV2bYHX5qQrUugVAhTjk/c5L7FzYjWflE/+h7RwRCbyW4NWv
P373eb7ox7QBTqHaTsV7+961NIbWjW6zk3CLBY0gURGtF0H1ajCN931Unm7lqnP1
OtIRwqZWEfL5S3L0YYnVXLRDtnEKCkBAITd9GjOLTRvOw5Ke1kNPf6yXReBAPJa2
pKO24xaW0nwtQcEFMgws4mzSAO/mUNAHSYhhdn3WPp9zWuZMlWbs4qmjOwdsCZ6k
Mjq5RV+4kncVryBQmHhwXLSC+GBnSuprqwyXQdiNJ4tfTIIFcMsWoq68dWVL1Tjn
Jr5vVCqVWHUrS0zRvR6NQdHoFugOLR7Ss3PoTTVbyj0s73sgTnLOIbV6rtMaCAxn
gTbq4OJpjoGAe80LwlI4QORiF16B+OI0n6wA9KwLiRZHjDc8fFRpKdDVmpDkMjTh
J78x378onlt9R3tMIvJuTfZnqQdDJJD4f5n3p23VE9W8RebNcjrpB2JG+xLQdFxW
iYbQbrsduBxcg+hBcWagK+raMUuaZx4WuM3KIhvn4FBfSMaczph4kcKwrVY3ACQu
uTTfrqlJKR6nax5IYmFa5uZ+fdqdTZjwTJXPzobTFtqGNECD0BAz587uNHGpVv6f
+C4i8yZ8h13tMSSbpX2CQG5ya6YJq+qKQ80yVfJLjeDFwTucDoDtNMlZqCf4qQ0f
HasCEy6nweCfRuFQxAlwJuR3avPZIwdrc09Ku0oy+UvZe2nCoTsIVfOErwNkYALw
GrONBMFO56fL1e3Asgz2FKh/3wR5/G00ttT7oMHm3B2Ir0UvO0Wp6vyr5bczEWmS
h/njLpb+TrRDc8OGD5RQ++11HuBFl59lH6h88le8FLPJCLJjhSh0ttnoLC9deW1c
2ifKRAYS9r87ffHf1XStV3g+T8iFKFgNHDBDpnCQXKmI85oRoocHlzi4ZS2eDP6m
q+OHfqjnTS7tb3hUHryTL0CDoEtyceuh/9FCTyj7peIO6KJCNK70n7eY8Qmg7QJE
2u/x1tUmgUHo9lAFzOJm95PJs+EWhrdNfAude8d4gxDdKP5g8M8nv9gxwprNVTpD
yiBi9xhUx7eAtMB4H1SBsy+diVODdZgvIJV2ARcXApLJHdZ+nIHAyRqceVvZOI/r
VUzmo1wqYT/u/HxjKkYwPcCyJiEXXWbd4NrB5Fo1LVat9ajQmBJTrKD215XqTe46
P7IEvxVzdX/tT0DetWd9It8zlBWz8wqx196wQ8AJyuuziBjHl8r4I6LqLQ/XvjO/
Wqju326ttM5ZIecK1NjiWuF5u0BMi0YTxbdr6wIJdSYZ5dXlkLLBmmHIJ7MElvMb
m0AnOBZRp67fdQoII1/p8Rw2smcxS5aHuR58IsJ766SldWQkbWfzhC6BbWxTkaA0
cwljrSDtFFWOEx1UbVuj5UxxzSH93u/xmAvqBRWlQwcimA2g1lIgpikc7LS8Mb9M
X6ECMrQXXx8DhIiLr7wNURfk4sBWG5le1kCjwXM7xrfn7CjgOQsea9TxQ/7A7oFd
1S0IycAMldoUERXusFPXcL2NuLvJmadJ1rmEZeFk3mkbrdBfw6c1dp7w4reu6Lgj
wRhe5sc7gL6UgkMRExkXxCjBTJCVSS4PdKQaqesH+j6FhR/lvHAmRA4Hs+Yp9+kn
kZFva1KPuHOdVxyLuMYekTqaDqF7jR+btpnEMydyEqkithxxb8NpFbvSiELDsNjJ
iv0/zHcXs3VS3yx/6PgMRwtOIp3MFDO3+B7jG+vejvt1fEdOhCeqsMY1oKwu7Ut3
XbbNVJE+JG+vwzoO3rWIozAnPRnsAAYkrtUbgdjT8LBPjh4xmK3QmLvpyDkp8Xr7
HtLjedAxl4jOMCotrAG9OfPau6ogtHv9aspi2kApIDuZ3ufS7OGlACq5vMNPlp4t
VfSb/qr7h/mCBGIFpvUOoGZYOnyGOKV+WtyDkiQ6rv1ShSabR6d0rU1nm5Jk2PtJ
9hVVykHCgPrFycLZLz/BO3wGOaMG+k8EMXnTJlSREd7lp7rvWgmcxYdDanlq7ZBG
LNG6Bo6oGwbYm7/BkKW99BZ5UvhUfQPodMEEyPaauw9j5gZ6cTcwLW9d/0iNw1S6
nfdiXhgKbo90mHrUETUxm+kCRUq6d/Io/ZqVcUQhrzAueNPpu+U1gpDk7rorTHsw
7ZFVcHPPcn9BU5Q+fnA1/A/pualJEQ5hCe2Jp/YxK5wgxY1NAmC4YuAakpuV3kkE
umMLPNUutF7xHpZ8FXUHBZyQkSBkrjQUp3SoRu1YMyTaTalt361yQTuDCU9IdYqy
Qu6AR+Gk+4dXt1gFnzTzzo2oH5yUHDUo/55z59o0kM7pB53mdlmYVBqDV2HlWUZm
3P8F1MoBi5ozwZUM/XfnPSjBpSDrhmtRK5gT54oON/IcN2bUso9VUBMyJo+D2Vua
hOnaZ7xonr5XSjTbbfndKSZYnWB5bfzuVglbyWCEisqht5qK4ndc/pEqOCOp0zQh
nQdP5Yo2AudllpwZKCKBQdAyXIF9YKXA2E6CCyBcPNA9T8gGLiHhNNoCVP0R+YqZ
BlSwslWq+21fIMjMfJl6K6bbA+oS3Hm5DpGSOAvTHR7Ls0YZ76+Svt34cZ9Q+w/s
EIyVRki8ANfpSavoYH5ERuhobTPXpHUlLmDrwOwlh+mKWUCO3orzAQluFjSTMMYZ
pMDBXWpHj/2Qy5WbIVcuZ06Z73uvzggd7mSmuDohnFj2zIRV+DxFOSAwgLQywruT
fUVG3UbUQ9g94iITSNKdnc0E5nLkdnCtyXhNVvl+/0DwNMHfgMM/vKxSqcThWMMG
WILdBBB6lbqrD1CdomRY6Ghv0MDhv6WQwTumMUxFM6RzJHECunaANwWKB7oIpOSN
IveS3eURfdKRnnfvjgdGvvdRaRVP0HbjDweAouq8LZI4KbW0FOztGkhT7AC5yvwG
k5wB+EFh2aS4frVIPKyO/q7SQMOq2Y0T+DUwmB7wDOCDf4Lkzl707Xmsx0/8mrwa
T0m3md8DKEWjQBkecLyK93PUN325QCnvSxA448h7GHehpVaXFat9Vgv5Zb3ag/w7
cXq5P1GNvpvctvj8DJ+lgM1jHD/hUBKc5OkcznpXDLRr+ywtqn3AEDkW9aLiR02a
wGCa84kU8FglE96xTszyiHKMrCPORBJ6XCRVfIGGF7lQhKg4FIeRC+Lr4bEEx6BI
bnUv9O6PyFWfLp+ty58Jngzfj72BtBrVJmkD7QDlH+bMvx4j8fp5ys7YKqnvQiZC
8xNcESVdGNYmzrmBZr96a4lG+8wsC/ItdbNB21UCZ5bsd4uu9glgPciuRH5D2bau
2mdchXmyVN+kLUQ5aTxd21KurQh8K4qE3cwhgJpjPSv4Rw1WibGioKM/NFMEbH7E
2Zm84MMJeOm8hfXGtHOxJCBvIHMLH6kMTp+7cJ8bHwy/pn9hKf0MOhfgORna6az8
6WVQufsyAUsI3svD7/e/OuBoh6Qq7Vqxq2oWAXQwwRlZj3JxMReDcmHtSvZmINVe
bYHTUxbVG3PSc2R6M+7tg0p4P5nShIyZLrA8VmfDetUnPSLUW5In6lY3uKNskVX4
Lfm9JqU5B2uERBjoGQ6GbhQvgnqJmuXs3ovg487Z3hwkQmiHYlUX54MeoIHy9wPI
qTiqQbmkqxDwDS3Ku2wysAaVTjiAxdJMO8xlWTIpETcT3wpD1MrTrq1po2AO12yn
B9giZJmAnMAcKZfqaYWMMNO71HQ7ZTl7I28CCJujXPFyV2nYU8jIX+9bGh4TGVn5
AYAWUO1NJvt5FxuU70kg4afWUhRBxFX1NefnJwKiZXDz5TZ1+GYf0J124XBx4r/J
zme+8h7Ry8xfNnilPDbwStrtxBVJZGiYhobu8uzEpbK3ILCKVz2V6IeuD08dKUWV
xtkQv2pS0aiCo8h282hgJQ+4cCwrmCm2pU/NBz1mgCBn5Tao1TpJ5k3e/rTPWIBG
8/6ymm+lgDi9HKZkYqyeng837FwgHUEi1++dwRS1r1QsER8+lxmZ5KOrxTegq2cs
NJVpf2VQd+JNsLTCkvv+Ffy7RmHQT7mq8Rt5xrtR8opDqgx3K64ImabCnyo39SX1
66OS2v2tbtWbDuFS4K03pLY9oYTU0YLYgpqNdJZBz+lVMf8DaYMVx4ksN0sFCBxF
3D+OTaZ0aZzLhdYvDpoZnzttRP0dofXEFvi7BUb0v1Zfxu7QGaNczXoaAmGSlzPu
l3p1c2Bkd9eJMGh5OE1sLJNX1Dmz3vpzVscPqj8wDVS0A++j8Fue/4uDTFakO91S
Zk6uFIElSuuC3CNA8NMewS8YeUnKLvBNr75+CzwUTcN18ZyWzPG6Xlp937b9LmAD
DRNh5K9NTf93n/zEN1s27mDfDDI5glSxyNeOocfXT7RCsyuLN0hEbLFiPXM6gL38
G+c0mkv3dflrDYCPIR5CmDkn9xeBEaPNZz2a3K2PKfK3b7hGdYz+Cz7OziS8UZs3
UQv8HOSLk5RLV4US/qac+6LSFmZHugaVSDiqe1/7qPRIETNMqIykPTfrCCY8cHMS
wPfRfZSbfccze6yUcrxtgiGFeR+iRMyRtYP3ZnWOcZBl2qK+VRk7Zl0pg/V2Dkk4
vxXHwwc8iyUsjNk3En2gXqZcZeiHHTrWltjiPZ+rfwMyNrDwvuO4yyGtVXioxmVD
EvND0ugNGSz9HXubV9yxKSvip6Sj9YTIeNJ7WZkxc63BIEDowAFjQ9Z/NNHknzf7
xA/QFfKRgmRbKlvEG7GiIXce+3rnbs6qm1W7y71TD6q16oAXNnt9bpOUlA/fpa7+
d8CcuX7CAMPB68i7SM+A/bZVOfp9pqAR73fON8MQFX4HoCFsc7YwhssZBo+zHWis
QjkTW6MLZGfmFGml0yPqJgaaMLGGZOi3GfKVZ2MN6ggzSeEsEIlhSlA7Wu64eCqO
C38QXn3q233KWSe0552j1Ukg30O8dYljU4w/rBiVZWiVoKLzUeY3NuFW8nZ93a+k
g+wdjkCY7GCTfpE1k9zVFsMoSgEekoGhsV98lbFG/94C1utlwE+TBVrlGmJimwZy
HOsUgj37EWvJOAkEoKzPQJRsaXf46jbEVd6Gr5ur7RnKb9FHKAuBNQCnk6zK/DSZ
4Z0fKZRYvc4+dAKJfbXkVNQegQYR59/PBO6/AX9WGjaUY0kGKrPizjMK9MBHrFy0
4Ckab427fTU6HEShd+msNVWzVQyV4Mmvu5KjQi2V1VcZ8O/n7CwCYHihuxSJySnH
F0BNuFUoxrnkRVqhfNmbJUw6xx1XDUFkjw6KqGEXzd2pS/hpjtHWogMeyF6sQqP2
/3vbqJTUNW+z2aAddgl0Zd4fI/4U6opgiER5fNmfyXzvqvc0MwjEVh9mmlA4vciP
LULugahAoWKoa0TzTC6w/EGhzRJRCWJ4vBpleM6cUY4Lb+g+MK90O1zny4PM/9bd
7FAiSYxDUQETIYbrRA+bIDVjDGuaeP6zmDE9/QLQUNCtaOUIjvCA4zGEwu9BFCSs
jbH6kCpJC7O5NXFnBejRoRt7+cgzlwYi+eo7GIS/y4cpF+JLWrWByHaN+lvIukRY
jbI7dE+RdSbG0DjPUcUqwVFYCcrTdxchBjqmd0EeTslwOJSYaDO3hjmdg/PZOL2y
3+P9Ts0YPFIkg70VuRdWSxhEXqEpnUk1Gp7oGRHHywF51m0hZBLC1c5RtBBIJsXY
CO/fpmYkQ1hlp2q5AbmZguKjUyxs8aMlp/7gsYTjM2+TpYfbKI3T1Z8OuCcXzjji
ujnX2q1yrLvzd0YUqcFMLfAyoMMEUXiVgREvJEWrZ0kNWFwpk0FAAclrbuJ7U7rA
8cwW4lajO/sUpBqRoVznjOtkhVN2gXFXWpQWTfhTnIHSubsyl0r06sU7a/4jJRY/
iVtBEhi9Ss3jwlJQCQNIAUdQNYTqaW9dXRn9jSwS7L2GCf+5X6s69qDOjA1EaTOD
8iHL8mTr/AFyMa2a4aNJsZvozyS1jP3fHYwzWtLu7mUe9S9NGK2V9dV6f+cXV8Zv
TSq/hqLdI8csFyP8O12V4Eo+liyMVkoCCsYg/PDjR1tBwt6SHX0KCr9doXKQ2PYA
UtJe0DlUM6JAlXxTZE0edIuzl/8kvt4RJHlkTAGGjAjBapFdUI+nYmFd/1rpgPhM
BK3AzMeHioKvhZMpsh+WmjFXCkF4eTYEvmcEG2a7nPjr415VIM+5Tr94Xy8hGHmB
mHcAZYClFX0uIyb5aXarLx2Wq4nrmxDLqIwuZJGJhaYU5NfHhYbi0X4oaBzT6B82
crEDSDFKMmeAhJkC4whVfbCEHMVR5L+Izi6LrZQEQabpJ76PCmgDdYehh/1U/X8i
2/RvA9fHHDx80aIxo02APJrQypp6U1RG92OAZslt+esvIbtfJ99GPRquISMk28LJ
xcBnzpk0jGneOy/ThvvNO6UJqT9Ixxe50akSmk3SivZfSOQS++b3cvNw4z2oRk5b
cZTOOpsuMXRHVtbki/jr1k66NBKZLjhCTP7jGQyTDjYLgUMtegbaE1FqcpADV5zF
rjJebY1+ujri+fftMAh8qn7TL4f/4Yk5xJlomTQBCcxQChNqK/roW+hXBpoyjJTK
TTYeesxog9TERV8qSED/Pn2zsY6o3dHAqy9M3Lun6oGT+8gFHdAMhiFmz2hjFO8y
Z8BEEF2vR1A87AJRr76xNatw66wSoyg4twgJN+3QMmPn0PQIjOLUq+YUKnJw+cOQ
j46JJ8k1feA10XR8ae8sN1XdasDTZNd8MgIdRRzb0fcRvECL8OdUyNYfZkl5AzbW
bl1pTZOCMYULpFBuqCOG+dtsFpxmLqVkcd+5orlzvW7yI4qIHbwm7zPv4sYMEtEE
MlCPatWhw+BP5paJEDX2OKLzfUUV839NHGT3h4vtd/iXLEa+tVvtqGF4yReggRxy
HRTfWLq3xsZG9yKZYoUhr7RNJ6GlkdYSUvjajAuYsJBqwRoPgPvitpoGWSB0s08C
vBW6f7vvfkwzzXqiDgsT1Rs/jdukHXCVVWU7nKMhkKtApx6ZkPitNd80YYyivzaR
xksw0a2fjocPSv1/bkU9Jvsgnobdx8/g6/4YgLSFRQF/spj8IP0DKIleJx6+tjTY
IvDluo7Cr2Hd1UZWNVv9BZNnUIdbBK3Y9YdIN+/DaxXoF2h+FIJPbsek8j8rD8gP
H7u0+Izb6a+OnqWFl/vi3bRNFwJjm1ZWEuwrerJRiViPzUVxgFechelxaUaoxjSz
mqeMpRNX546TILHx4vZEJ/ikg+TH2al93GOFeqGGOrhk4AyeoBpbt4icmNzOkMaZ
kKTPqYEGPVUjq17vinK2n24BWcCNaxilzh9Tfu74cgjZnXcq8f9fGE663F8LwPRy
KqYwygnPiIIzAJ5OMBvo4bEnG9zw+8Z77IF0RHiOfm2LMFmd39qbmdztxMbi9M/v
peaY9qF4zWaOpza+x8GmoAlkv8IEFon7zFO+F6/kt4cy1C0FwhTQv9Hv/mGkRvMU
AXDAsgpjUib7UovASBEhHusS44P6xeL+VW5y3FpJyTg2m6QI4D1kS1L1NHSH0fpV
r/MaLKltX0A2vZovNUCojfNeMD6PaX8cPTlLx4J1cq4FcbBkXNk4ck9A04PKLEsx
HACzi0ZlyVxaGJty0s22nxIyaH2XitrmxFJBsSu6a8Cm6Zcu6KFLwDMy1ea46HKW
yYH/xig/ymqX+A56cfFmhrcXN1zEOIuWNUXKTSZS8Q1NLbyvu8kB4KSp6CkdaUTI
b5QMzcF8y4vLc76aUKyeEvrPIFS0wY2zuYm4JynDN97NHzSC25N4IQVPDUdewFXo
Ra9xffvRyG6JEu9FPUWhP8RELRA5UQvPGacZVYq0glASjBg+Wo5kv50Gv41VliTo
aGQCPxBAA5aXen05wSBBN/igvHpUDa0NuQHT22nZaKy4ECofaN4L3VDJdIDHKDVi
sYKwj03+snsjdpr8oIv/r+PDU2DQ9dv+g4uC2YrncQRucLF4+zwE9S/S5Zxnsig3
0XXO71dQcA0zUGwOEwPstIHUHPLivwxNa8K3BQYgZbv2kyMj2nyBwso8LnXXnCoS
XohDcghQzWd7YWg4kTD20gl4INORZ+tkBvxQ4eWT+9fyo3it62nXYkIMNFllE6Qn
iyk88B6LoNeHhkjXISN2b08hiGe2BxrP1+J8JLL3lNxVFGTrCjnlTmLVdMQNJT4d
wmqDFm5ikkdHnDiYBOXCm6C2Mx2XVOMyFul5NnzR6X6lc4qQYvUK87Fm1Sk8GEHF
Favi9l3jFT75wkNqFKljq+/DnQuDaP3tgzmRJEIY/wkone+xdJTt1tqsPROC3nNY
+9w8hnUKKgVQ1oCZc9BjevnFTdKg8qhxpSryq9WgtqA42pp9AA0/WHAclZDhxXkq
AbLZkKStjxS4y+xzEqweIhykuRAeZVcKg+7J7Kc8KJPPMwuaMZIaiNIAHjWkbdbf
tcjR4IcxanMJzPEDiE6d/fLCKlmhKKddbTMI/d47GgXX06l9UWXu0SGG0VEMFgxS
GahcJs/T+icfnx1DgJ8gJnLW6eJhgLgqgsDjmbNbvV0FeIuH0yJztppeB5qxwg5u
ZKAgzNNgzDa9SV4BzSWpPEHfHMtuHZNezDapXNdHKHgvQCXOOw2fLPh8Hui/T0Aa
XhumSG6g5r205PKsIq1rDHqCCTpPDsxqNZhjyBxcQwO+pOJ6LD6+tKtds4VuFv9i
Y8kn0wBzla3BcqBmtlvB1Yqcfopz6KTOAGDLJ4H7NawiVn4WQtuynfKLvNvfB+nL
wncSe+o/eJDqusA8Ketts1us2WPmBvAGYP9GBRFofisv1DqITFpu7uNzzfW7UNLe
G5m5gO75fNj5D+6VTh+dPulScvQ6+GVcomcEJG9L+Cv8x0ItzsKmLwj7j1shn8ua
1NxDN3HFsX/1lYpq/TSEmayTjnDcYHkHKAmoyFJ13dj0saJXdKWPCRcgJWPrE7P6
ufjszbK4wE8Fm6vAoLJlqa8bgSFT8f/08+Nc0GqrI9bkVYdsE9d63xzXeaZ9yRWc
OPxLD6p5iFpBz1XTMu7Eav1SqSbxhCJie15ZTS1U4Lgr4QloYN5dFO7REO6jSsq9
xNpGJa5gwYQsmHxWWWdCbbEoYVLsVgW8cZ7x1QG1JsvWHaiNXs6ZksM7Tz0zLazg
Uox2YUFQwgdekrgYj8VEDtxlcQSs8+BdaBmGS6XqXzpa+Q/g1ucfHeFH27HSa+qj
RsmfMHwt414onGLV7iwWHiJsG0jdZ4hg80RCdWPI2MVCSVBS7jQuwZx8gAAUXA3Z
AUw1vQCDZPcM2znvEw3h/nanSonph2CaFHBQNOuq/T+OtQH7xch/zJMUdPEgVa6o
ksnecNX3I/ujpMjRK4BPKSiq894rlUNPH1fpmpH+KIXkpDB1cSTQHS/4YoD3Oq8L
jB0aIHw8kdbos6sx3RSU5siosRFgZSJUwIhC41mqmogmNRcreigdPY17Y+GnGJZ2
QY5F8H3rnPopCaMgSYUTQUWbJ/QiUOlQQt7fPndInhuxwF18fbmYL2ZbZdik3wzA
lCOfESn9Tycerkj7TBSsQxMOB8+BpMV7/kjTys5GVe17G1plapwM3h6lREh7h0wb
/NAgAN4sp4Oa7plEaefl3SzT00ToJXiv4ZI4RE3sosXguDIl2eE6lppxBvsCTxzq
grJUBx8S6juTYKmaJi2T0QBGPoiNfiu/HHuk3+eav+knm9wYOlGWTSzoORjjhg0x
VJBcCZHrnaYC8Zl3p4Hm3wMsYRojIRseOaQukHKugsPPAlGPUTT06ynBcXYC3Fwo
W759/UZYpz0zcSIYh+UQNhOlodowHQnnbQJyvOOqrgRZQVE9vSxXaMhQVIU4gwy2
3Oef6AQ71xpjrUGhnpcn6TQhcAlhXl5pBwW1OoGptI6D0O+N57gEHIOEjC9Smisn
Of+PuOApwxxLZ3HZ5hTODEKQUFdFrXjPRIfmUCw7OILXHDLw2NRwFcBObfSQbqEG
qTRtnRl60WIUdaThbDDxxbNjz4gK1qFzIDlD0FSNLt36xwBzKiiyUa2R8opONerG
ldaym5upRW54kKZNUdy+DZRQ4s+ppdUdbAM15VQxv5R4srJT0mRVE7EhEyfbw1n/
o1BCNQ0BlP/77SmZ31l1HU1x4LNPGGhGD3SkQ+usAeqbY3NjRN4JjbwxRsuIN/RO
YGcShS23qJgJFcQAeQEaYVsrN+iRmMnjjiKNTLj/I4aAkpARfqnZ6nktBuB0gDIs
fJW/KdaVVQNPPllDqptE757d8nRxwvx2M8R9/J86NF3PSvO4mzAJZ3WA9Lmk88Hp
SZCMpQ1lM6TfBTOA0aloMIxB1bx7uLiMsfDD+gOiO9rHl8nuHRuZ5tqPeDVhy/py
Q+BCUUCZUilsncDq80SbVjyjlL/jJqq4YTvCbebmPCW0RgjebxhQiHix3Sipqw2M
TlzuWjoEu6FHApxDa674qv0Wl9FoLOkX7CvVeh3X2qEVwyJybGmp/tXin2nAcRDe
1mPzSCPCtkj8l9gVQrHlXQa1CizewJWYGewTkZrAVh3+ELsj2NTUaqt4Z1gBCJ/G
gtZXkrgr6sUlc1IE4aJ9bVQZP7zsKR81bU7OVeNS7NxloUP6fCGqNb6tQHMWiJqK
kNuGnZCyt90cDDN/VoV3ESc+ISvEJtxaiFk5aQuG9KwObuAEGLxk4137YPaBc6p6
5Mqcx9C8x2uWmAaVYyTikKolrC2kCNXLa+tHTaBzIDJhMIsAkxRwc535Cf2IfzZl
Bx1EGOa5yBne8fTinmqMPpwq+kj9e2WFeK3gDEgTq2nu5eis6KH3DVGqivsdQHIb
uO8iJh99XKzWyE3qnFLuh51erOMVGM7TPOH+WwLUgx1TtEplWS19LPS5ngQTChOn
ThQ+RvVB1NiNkWLpLTnjt6kZSwJIMQ2PuyVETXZB8VsY0s1s0F7BBiJ02haqDazx
gq1nDAMXSewklWvg5Mnn7zQrn1jI8DX6if3CkirH/q2OHjGN9y/QKujkE39Y6/z2
vwt0vUPzuMelbwUQd8oq5YPDPpH3mOpcUQTBog+1dAFhg86jCXqQsEK5tZwIt7va
CJCKkUWyP/8iFDu3aUL4W8RweiaSqT5RjQJKaxBIWhf+NtjOQcQbAARBnv9eCdST
Td/axcO3eAnmARhTxVX3Qd/fz6Oyk3BXfsWZoOBgKjtLxPAbJ1Mlm7ySRbdjeYa5
SoJFENSgNbXpmb3O7dakAyqMHy3pZ6tkss+gEE5CA+7Fi/YwjZmLIRUQ+eg9caDN
xRsRlvM1ttnZ9wNbL24QoqZVZSQl+XElLfhO4TLrjYNAqB3jGs+4qC4UiSfnB4P2
0uPUYKcJMKL2uLAOlaMxtFyW7+HmGcdhLJWO/odI+f11IPJNR1NysG/viGbnnTWw
TFACL7Zcp96gQUwg7DUi1l4QsiXnffIqzhbLoAfJTuEmpTVMAoVuKY1AFRj8O3RS
qtFz3gsAbCea8m/phnUxXuXnBw2QbpPqlIG0tlGKtM9Q9UswOEXbIFTnkkaI9XKX
ATGTs5mqq9TNIVn6PxjoPp2iXx5Dh+nDZlaf18E/xwjcZxLH7An+mFghfX09co/U
VAekFNQne4G3cwMnGD88joE6EfQabq4IDP5cmCYqawWmM9Wq+PfVD/hrCltP2cZr
s0euJ4/KOzO/5cHJh0CSLfMEJTNR2MbSEk03+0WikDbijq9rmIoBmM9dZgSbNCL7
bTlQpswwnLDX0hWW4uPNM26mfIMARSxk9NLyct4V9RnxGNL7CqO07mA3RsOSSm8l
Z/yj7GR5Ayp33xF0B2ecDLQzsZPlsFgPeKCfA3ztm8xwF9U+FZ0gVRi/4sWR0HMI
/22mpEwPExrAdBcFRKraKL+76iJdlv7vAbilsG/ppzX9JJuKaoa6rt1fZoiA4u0D
OHlNSiykM8mDM9z4y3xSel15HK9b3S3Dy/mIkvlQXGAZEhqo6c/8IQKzvs8Nxx1V
mg9WscIQ9wXCijv225ZhG9i7jzD9+t1ha8ka5FTIOuKwyw79ll75aHnhKBtfxl6O
UVR5epYQS5pTt4yO998pN+EEVhmzr7WQS/R8svk/RK5754avrgkd0vIZNMgjFH3v
E1wcmyt+eMfS8DJNsW1OVOcauy3NvW1XPrtMD6C/PTBOoTPhUc5DEAgC1LoIJcRd
b+3e2EGj0fJZ70k7R7H5ZYpyZKI8Of48gj1wLqPpVMYYV3FQ4hbuOiEg6uDY5a4A
xqytHKD2XmRIc/MxFaLF1hGvQhfzHmmpSV4kSnOC6oB9zRBM/KF3dg96oertbqal
Z9vbfdVtX1BqrY72HsTRbqYv/4w9/1CnOYKCnPkf0mWX2by8oEXLq7Wf/Jl4Qbeh
Jv/zLWuU0zvdl/OPFg+SbCpkW8XZJJAV69pVS9BeO6C5Y83RYhoCdsdwKverZMKC
vDSQrX8p9cuig0EK7FH1qyjTDnzD/DEQ1auO/4vipnlEYRLpEm9lQk8Y0RFQty/L
EUUiE+Fnn7osjGquNnccqzxhGFgdHWfOSC126kq4HpS+j0DdnpNyjnS6sW42Uec3
gV/IuA2JE+VHi9LPJRmNSv0SPZN05RAiSstREdqwphC0dYPxrx27Xd53Tq9/NHeW
Ar8VSmRVCur1sAv0xkXG/tBn4UMWfCT2HUNrqdMuGN7L7T0kIKP5D4aG+88FT3e+
pvsZ2w8f3zuMCiaekbHnggfQIVw63TpVukrvRsJ1EMd7V+Ls6i26qUl/rvAQ/uIF
R/aBalX0J8tYrHLujjLsr66kuQ9mfpOqplptV82BNu2wVGInoNgPZn9GIad7Q7sD
xbImG1TC2DWshkZfe5ME60jIDtswmxHqdb6vrRKTvfRtU14f1/19qisjpPFVRGZu
/cQEfmTzkw8xYrWTwwefqw8Cy+VQolDeI377YxwNaCRPK/2oL9ag0XveQiguu87b
aW3aQir8Qwp0r7TaMTRunavuL2+JSanuNLWxekvlIlmyDIcbtGrKZygqs2C2fq58
mNUsQgMHRkGzVVHq1MFncbLJtq/cZQq2jGLxaPRv4PXHkUyd0EpPGoBrfOQVZV0v
+TDQPh/7b5bic8htf5DB/aqiBZ+93G3UO2xZPbSEUSZjSjKHQUN0fPWEGa5YagK+
inEPtmKUu0FbA1COj+KkTZbxMJgDx1PoiNQcPZVlP4jPnf4KlREChwTW6GQBYJed
UT/UURpk0oxU6ZrOebqHHnmBU2ur6b0lkjro1G7BOPs9dEWSHnvWTVbGy+G+uTwG
2X/kw5MQrEuF/SlcRZHu+3khaBn5jhWt504TUCSscF8onxAHRT2bOJ/bTH209qq4
Xt2vIKnJldHYqhoeQy6ezZXfqpsPe/9QeEXMXphIi1mE8nF1F0umZOLnI6cQ2vRV
yNHp/X3LzbgUR+WofJWjdIk4/uiVqSEiPiQ49ed6Mg+XRm3v+m/yzSWOdML3N/uP
/Y3Zv3EZC92MqDHWDZstpus3DY/eiiZRkD6JxKyO+Qb8pUvuPKlykOVYaMFnWRiR
S9crhNzEkJKMXZ1MEoWZLKZbC9PT2umodQjm0x7ONXvy1u2bJ6Paz799TPf6PqYS
yeGPD6Isd5g3eJkstCA/j2akWrQxu/11/CsQj2u8wI/7jRxvrIawXqqRu8n3W2dC
5lOMA5uwOU6danS298D07rmdXWxXsNdnEwDdYYi44Lm3hUHvnUJ+3j0+rEfwVwGJ
fun24V6R4WyMn7CXPqGzHYOrMw2AFoDllemjJzeiupz/pNI4756gRnVGFp0fEtEh
A9ejfXo3GlWLAfKy5mN7SLkxshPrs+pcxsOTVmimOFLd9R8a7cqsX5UlyUzLc3t9
S69G/kEWBnoJ51tnwIiAW0CmRmL4eG0H9jFkkd54Pg/Q/EYHP5spIjChr8Q1aay8
uw8TuVuMuKipbZtfUq7xosUtoyt+gaiKwcvkR69NTK6v3Nf3zTNXhQaCwPpxysec
t6JN6nK0pO/zO/Plzomlj0gcDzjuX903cG0bhS4BqNf1jHsgDbUFYSATmANgk9Hh
aVdZiy/SUxmtoH1gzKuKjTJ+X0J6q6d9n7XzqcdJKm9VjpUDfetJd/9L3dpvVQw3
2/CQ+d2wcOPSigTbUuxSADznQ3o5fPtFgQ+kUh67tNFtP26zDh41kuYvrVuIiq7U
Wv+8c9kSEq4m28LGEYkF/Bg2NtEou5vwepIBDzeQufnJE4f5ISYcUvnRD3ziGtgs
6FeS8zMjDTOcrofZJAsBYwBg6AI4pcEuesAh3U5GmPDofmGVTUvfrv4ZtRDYjxdA
CnVXc9SETXJ27xHZOvlGr196NSFz6TcDKK7qkslRGIwXEA5hgT5Jb2YglTfgA74w
pspFj+axG/1q+Zz+STkpaD2iQnslcMIJ6I/ShOgvH58bEFvErvxi0Sd755Jn8v2n
1mHcNN06IYosgfzq8GKkPFSHx91tCp11XiT/v7pbzvJlwd1s6bKKuTQniU98BQEd
RT2A1488HE0vuCdvD4pTOno2JfG9d0Jl9Tj9Eud4e59Vx5uj3OqdavaJaAT4ESBn
XpIvB1+z6M2Js29ReXV/nTanEMX4oTVZg+Mbm5sfEA9WjEBB6klIjSs3e2yR2e7t
zCe3BjEHyY95rUtmhMz9MhXYbv2Ru/g+mKbDM3/L6C1R71LYLK81KiSgtW9oWtHp
XU/8Oexb06Eg88GpNRcnqU6EReVT/2q3dKFrurU5vW7+dQjNXhJqWPLZawiyOkrk
oOHEtTSNf9QQf9ujS7b8OraKTlbPDyKPz6qHHkQn2npoCpJj/4bCnZJlT76j0MYI
JauAof7edBCl3v74g4GZqaG6mVxQZ091nauAUU8/950=
//pragma protect end_data_block
//pragma protect digest_block
e7fp14+QVGyotz0RpP7YK7L9n+c=
//pragma protect end_digest_block
//pragma protect end_protected
