// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
fbimcccxgDFS1pkPRGAKZI69V2+bScuZhFPS4F6KXrHHGbD6yM5qZHahRRZmfNi5
mfhEuljBfltRWDK973JOcHsmDLaEQWNluHKezntKScb83ounuZNCH43gAwQr5xSD
fV3QgS1/k2LservQ1dTxEW1UzlJLzU+lex2XYW3NuzQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8384 )
`pragma protect data_block
EvlQaFKA4NDllFHj9uY1hggVHy5CYdDkZU56pi3Zqm32ME0f6WtzXVBuYMiQR3L4
a3NKMSOFMlaKOV25HE9RBsEjC4x+5jUva9tlUaz0P9ALk8OoYfemMenw03ckUzuI
jYnIcbLC7rnXLu0EmureFierMk1qrT3lPYHICU24eUcXPL6bAsTdm8rDbW6n3aZz
K/g7isQzhw6TKfSfwPRb+yZCCDunAJNtxIdbEIhZvKCvOImSRL9EIO6ys5mWz6FR
/Lds+0xkbU+kcfqS6KV2roPLEwAm3AnWMwgOTzNraXGQWMN1txkib/8AI1L0klKi
BjRArzXsL9QNIt2oaJz6Sr2TmhmaSv+YUApOtVP1ywEIteSdaExQPK8Z/XuZ/v1y
MBsqlfWh6HJG79/j7k1NaLfLsnDQn0S9561EL5mXacpOk6/Mk20zGyzVfUZKesZb
Ca8pCpp7D+jkV02dvPEaPYzqMMfbCk/TJPvEB3PZ1w1NEje4r7W18+8z3I/ypQmI
+7A1Mc13qRrXPPJPysp1YeDL8HJ/gk+kqzxW5ziDzMXlKqLxL+ostSQshJXhjmMb
nANtwmQmiY+Nybfr2hiSkeFBA5RvLQENmkDdkt1PWEPWhO/oLBtxrGSiBhC3YZfw
6r/hQgE/NglPwMtVpm4e8NQHnvmxd+IMVxS2FFYZqevvUZRP7wwlFWkX3v6yXsRl
P5bSrYxh40a5M70aVk1eJ6RUH5W1GJndNUAahag7czCH/N4GodTvG1GyNG3hQ1H8
9Xoa1dIDoRbWzDZkOCbXLFl9nr1949cZqpOKd9QbosIvUTFlkJagdVf/McD2fp+U
mIilgEv0A8YWeS9/HQmbW4ftaNY7X+N0JGe97hEQ+wn6XwsXQ5z0WvLVSnL9Qfyt
oYAQ+DZzbm1oanbg2GwpuyA3SzfKO85afLxKQsxEpO2s3y9xSa41wdzBdX4dem3/
PRk9k8DUB0R+FautKt0NnoZR/2FYSatGEyw/NPz2szFGrvFH19ulU7Rggmk6norI
SF4kQ6WjA0AkRtzEr75SZU3NrFA44ibUKVovz7NZcgf4c0yMHdMZahiSh5uQKssz
4sNnh7h7i+pLivKhL8+T4ZG1+/33HY7PlFEsc1hxhePOH6vsSweeb0KOxO4pjKSS
6sbsbI6t+HvTlINOMtp2orb4VIJgdas9iNeSktn8rnTfbnBsHkDXiUwJc/VwvyLk
N2dU4aT2G/yktG/im58krqp2SGe0RvmlVHmiHRk0HLfYYyCbxxRluclYKhbV9Oin
2lzScZ0jRCGYpHYl8yiV+l/goxvgbjbeyuJw3K8+W8iVguUXA82V5hqzIlmU8CSv
YTffI+yLuYgjZqwePhkoD3jB0dqZKy2w+MvtYh6jrGt4RJ0kgI1goco5kRZn5a8s
mllwcTHcdCKVSzVNT+7NoCqoKYg1UN8BO6FeYJUt1vzj47q49UJUBNghjq/PHsUb
HTnr0MJyzpRCMO0rdWvxqfFqzfRV2hIV5VUhwbr0LVgYiRUlm8WHaa+/SvAGgDyn
0Q6afQUWzMHKqozyO0zQCinf76/sAgALhZa0/FGvxLMi7jXh8iw9WqwnYOhVLxlj
ycfnI04FJHvJGkbpfdGu6xLN6YaICXTAPh2FgsUHaN4AZ++Ri6d00yI2fK+w5NJh
cv/7jS1qwpIXbM/NheYArWBe0CDVUJXFzira4FEWvhuEaTZ9Gom4Hw3pBVgiriDx
gfNOmc2Ljr3DZXkXIG+ey8FgTt+OPA4s0eCGOJcWvbQl87E/aY/8ZR360NIx9qwx
Q025R1CxMEfO+AGFmIID4mbuJkzh0TL9+8NT+bcrjimWsTQxbs/NY3CIeCKhcW6C
eXPncaNGWGxQ62mH6bsF0cy9dLRHgUG7PZ3foS27yNGEj8H4pnM8yXFvO5AcfWvk
TzNdYOk2OZg8ff9DWnSQZhgMkcMhCml25YRVtyjQv8nVS7NqxD9PEgbWMvYvYsmj
ru0wBz9y8KtybU5jvqnnSnK/JdeWxT1wqCehC2rL0b+bFy5uySGf36Z6R/5hpRD8
6FbItoHH66XY+PfU+Ovt7no6cxXRsrXNAJGwkFrzXDStEWsaqyw4AJruTg6rqjf6
lS5HE4WhTdKo3rnO3ruLzEkaGoyo1qeCYq6okWftrT5dYj2YcgkylPfEvTAVaa08
MeRAL/4m+Mww0bBECvnBV/6VbtAaScHLW43exLSEyuJqdTpr3KY4eZhulY7rbfpi
iXgsof++6KTE6ZZuO4qUYM8Pys/OGVr4Ppjin+MxJkWhvWvrj6Lw/+wZqb903o+0
hbG7WMAqIeVhg4L0T1BfjWPkNcea9yVfN1ZR977RX9b7IXd5gDfm07mht5y2l9g4
+qIaHFYSCWw0vB/LavNxyoVtE82oNW95hDxnk0UG1SpFkmIOTZ6Q5yyOHM+YoRMc
qu+iCrHjWZrz2a4x96puS5rUaxFpiKeYJYKTdK0AZfRdyxFNLN3Rn7r3pT9s1/8v
5rCRkV0m6nvyol1/jodL7SZnWamf6bskBy3ZCkOoVeby1XqaDPfV7wxzQGVpDbHz
K+GpQJTsEYopPFXfRh4qnwjoCvsbQaExGFMgqmMP+fGp31NnWFYURytFK6ATLVIA
dhJyPPzh0G1KnKhlAXERsudGa112Vb6PWBSqVqKoV9peIh3+0K/uxrYqenNgU1rp
TnKl7JsqTg5vhfXtQNSENn/8u1xQy2DWql+xoXsuvXOVcgtY7FWOFGiu3d/5erE0
SB8Mbkxl8GgTWKPlOnue9ZaJfSEMyAbUNKr+0cr3IW3G/BAQj+pS/EWCXZDjJNSd
w+l86W6YlcQcJxRCDjqiK/Btq2FEOao2hzlLwY7LsX0wpe2x/fohwTZE+CpG2//h
ExBC1bS9eswjvRhk6E74P4CiBpXbwWx+P+1Y4pIjQCdyVNryHlPbFp2qr/mA7O09
axd/U/R5Qh8p21v2SYLzq2+w1ZgzKXXqZfI5cKHX87j+/UdofjUVDjL25BUjTFzc
Tw1Gl54P9tBw4ku50dJpj0Ftye6F7JdT1qodZ4TepCHMbedudMXpIKTGAxF2NH8o
eDrAEDvthYvoqQeuZoD9cTo4DZ1/a/h1rYRnEve11M19wRxGrtoK3bebHxuNmKvz
iznMVgv4wJI/5R4RdRMgTjbLONIbQkacW3Ruv324I+kM7lYg9jwBGyDXwoVVjQKY
HqixIqfq6HE/B1yvMlU0XhUXvAGjimrbsFmQZ4/lUD26m56I42MYs+zu9v3G8Sxq
jF0RTH26zGQV0/6K6i830jEuUEVK0/oOq0S5Mz67WVhGCAXOK9Lq3icZJ1eGCvRz
ph/LCF4FDW1n2PQABLwocR51qs1IJ50sg2r3weT+Zh4LYcJS8L851u2cXL7IZsOB
Z91xbCofhGCRIq3K2jXO5lmR+5UsO/5PAGMk1+T+G5eBq93PA5QKrYwBEYxb4S05
avudgIPlotxWCqTc6UoL7X+kZbvKx7DKoz8Yhj69+BA8Zm6ygwA/c+ZoDESFVzVo
eJ7Q2HVO186hl1j3/dqMQX/4t/Zc+9W+9qJYWH8cqYsTgYEYP8qeqAaxLeyol+Gv
wF20yjbAW0QUO8qpmQoaKnVYYGCXSdhRICYacA0xetIk49/8adhA9n0X7vHpl3Pv
tv1Vqb0nnaioTYjGNwUH0KQd32+BO/LMYlAHW/sEPFgMpJJaC/BG7sQfQEggyeat
I1IKvqIubax9XehHyjHXEFI2LrzpP0Dpi6ORjV4z64y9GupbkZqNQWr6jxhswFHx
BU+43FQK//41gRv7OoCRYrse6D0mcjg5fkS3sDA6KOX1pQ9HKCcNF7Vrqy1zsiZt
tFkhHUnHg95o7owtNmMZldU24BlFjJYyp3SsnFVBq8DVuAFY/O/gbS+Gkz6aGdD+
3AzPSSEQW5GiCKl3gW70dBoHdLygCtrUtSrHDUOV2IZc182J0xShKNwTZJ4e++HB
w5yaMSXFGZ0sl02jgcOfdIHInK14+rBlcdKl/uSB2JlzNAvFwIhG6jABioNBHluE
gH1VVYlqeZUlGVueU6oQqDUY03lAVOywzRRZvsRvRtMa/qMqK4Lk6MfgKa93iZLG
xRkKR2hN2fyTRBgY0sS0rNiBxE11fh1CwRn/k0wRy4CxZFHxgLZnorhquN7yt7Yk
PBfTSskUPkjbJiMfyga4Gic7E9VZ83RERh1aegqcsfV9709pvG9tUFNMQcaixL/g
KK/YM4pkZaQYWM7Mw+gYnExVZ6cDhL54h8FeibNsw8VFkqmTRUPPc689w8osZRew
tCfWXHvqvz5Sb1HQMTF5Ho8/x9oLS51tvw+/SQ8rgOxVyciQ8N9i3dRNNgmbg+YY
rSneNqx1A+rEXZPNoOiZMN+BiAKvGIWEVLH99yHpFHvXeDuZMxuEkmGmwtIhY2Js
Sfa9p/MCq64S5VN6TcLEVRLDAcwLDiw8SVj0UGRxMYDgzrL0ZV0bZlkB8j8FLM1Y
JpegDFAwmpgzB1hediPNa8z9F7L+/K/PD2yszOC0HF+fJKK6lv7TLbMmSzuR7vPi
3rEDpJCWAqZsBNKqPIiJaRdJXkz9sPGg7n8dtbJ0YAHs/ZhF8ap9ZxcOaPZd7Qbi
eW88JPwNqblZrYwMi2qkd3QMUxz5QUtf3de1rZ/BoVr/h032UU6qvx4WBeWMEAuM
vkyUoAifOGOTJ6BoV5iY3IN65kind26OVFwz9VCRU/R7+Yxam5if7yIsnFS9RFhe
xo1xNcCX188MZ6YB7b04tISVz1rklkkWN6WJM5hOr3wcbkkjxfd9Erm9Q9EzIpVz
Yat6H3i1f26O61JbvxmqySfbMO3DedbU1w0qcaNE9s1443x33y2h7J9X8kAqsDMu
FTcABkPubLA12dNnWSYQQUXj/2C4A+TsSevKWzBSreFF0+fOS6MB6VvKsmR0/+sx
sbVkNeWiw/pjz81Bkd7toWkedzZ7cVaVoPAxlv7arVa2F/YP/jvIpwsMznrE47CT
4kmHlBLiDItXJ1yjoZb46rFs7cN0CFmy2GCIlAotfqIbcYIn1pZM2x3U9AuGK3mz
r+jSLXucPNLy0iqStAD5SSkH1Iir5aoFOmMX2Z5DXdNQfMPADa7qSXMr4Xm7B1XK
9NimSt5D6QuNhpdj8G5XcPzkR2xq9oYSnjKlB00TQtM3A29hDeSwWRAQMq0CvIaC
U9t/sFfcOvGJ45haoVlLDMs3Xdaq69K/M82qpnkHWZptvJGE3zdwqVDEx/zn78sk
RaINvRuetyoyKrOnrTW4SdHjnvvus0h3oOf06qGhIs5hYx7r1SxSayCcQCzvYe+8
o+ua9V8TBOC4e0sAsw8IyiArUeOkDWBCwsxdzcKiUBia9eGeU/H66GTpf50RI0gt
bwYzWfwJ6KNhEECLcGAEGpyeOsLUcB21AfB7F6ZJr362vtU9xEMHLf4jEVH3ulyB
+JBndm8fSKoDfzG7t/AMurRrLHJrv5Tu9QEFG3gI26Oq7bhaoY3UXQIkyPaz+fo1
+TAzIduVyi+S6MyYYPqP7D1u8kjXbGKjcxpv37TPcr3wzjPs4TPNTI51KHzq1DfJ
aalQUsgHusj/f1Kf2qSQIv743bPClqMcayRu9rFd1PW0JqlQmwS+DZLOBaarmpXz
PIKUrxJw+3PmwI2KYmwgW7hSrEpTDCY4IbJM61/RpZLbGboYbXiWf6HD1t8Ux+tL
sNM1GiTiiYCc284IItfMqFnJYI0YWoGLJdGJDgr1qk3ENCi4hxDZu8SB6uBKE+1R
FhAVX/B9anmS5GzUFbYoprcGYDSqJiOfNcRokYQ7I8AcZ6PxBmJhFoZgatzwWNhO
xn3/EIajTnE+L1yzAJ8fJYC7XWHpAJhOnM6nHT2uHzJGOm/OarviKnwp0X/WKmjj
gr9M0mhXCQ1xU0XL7KT3KxFoTcKuEiXnDfEOjCPiHtNH1VHu0JXplzyaetywaOCb
nWRbysqSP0aUFBMtfqIeD3xSwyc2ApXdbmYaVTiFj2LWKKJGiHjvl0Yqful+Pzgm
MbmOjMRxYZk9bL3DoD/judgCuDgShAA0+H7cEtuPSl5deEqnEpcZjfhN19QPpcBK
X6q2ZaPE+UChgwsZYaLvV7cYrP3YSVsMk6qLREg6ECB7Snpa9vfbyr4GYNv118tm
H+kD8nm/gLCbcjlQzfYPNm2lRumzEIlrS9M/6Y2fvq4noxh08vLmXQv5DcBunXXn
4BLS0+XZeAdXhMX2qhxLjMhhbtRuK9XrvT9I9V92z5smYJUrFbXX0bOC8Xrvyw7u
r3o03HzJWHNhVdHTF5StzAlBxpshe+c77yGp6AKC/krqaq3Li5d37gmFX2zjKtVR
vCpusRytOQnO2YXw38IQ5SKBDcYUT6IMAkhC7mD4zCRSlVZ881d0Hh6WU/tpd/r1
pK6iBsb73GxwxLXPJj9YKq0F9l4qDl90C6F1bweOxiFO2OMYh4DX4rm2eAOLwqSk
9LbRTwyZq+E29lfV+Zr4BKYAKPGZylQYFM40srpHjO07UFZUdvouDZKmIqoc+Txv
5qDBbekasOh4Z1So5rGZwCRVIbnuRkPZ2WN+nBueC4gdhd1MiwiivIyZ4JQBVUFS
dtt945+lBjpWaG9zX7dcpcxMJAEvMmZ72ioDTQXWUJBrwKtDjoPVgjEvu7DWBqgB
89kXmBeoyE1JuK/FS9IVI83CHfaseHX30Py+1SspzS3PivUBl2lF3FpVwgJMDtD4
E0l1KIj2W2eyfdhKu5oDc8k8nwTA9qXaGwAtawK95fi3RpaCM3EQ+Eb7jKouX0/W
6/5B4guG6qlwO+g84xs2Uko7XHUGZaHNx235/Rq5b7DiT9q3a7u3Kj6skg8R/z/6
ODbaobPqmzWLtdfE7eQf65LpR5e9Ipzn5gYr3m4GpKCOLO+DiJ23hfnoTFZuctRG
Loei6w7OTc15Lwj64aAiZ5imx/KEVxev+OGjwbIhS8XLJbYhLZMO4PkrLbRBAddb
QmnHXccHW0TTBsrdatsr487fTWuxfSpCY65IyMwuCeGS3cJqzcBEmEpO+ur/dVBu
DrBr7WBs/Gptp8+csxciXhUUR84Q2yWja++fzQfmSOueTiLFZVMF85CwpZ1dCuMC
VvLWXfxerF3hAfuT5ycMO7SrEzWeRADaIArklFobw9o4TqP6Vqzq4aZySV/NK+zp
O02PfFZL04s0G0ksBRpdCuZKHDjzrG61oddiUN0odM9QcATwjudMUO1WHDWdsEPq
qdC1J7+KIGC2Zrx2xAZEJVqElK4G7CLT0R2xYBmqIAePS210/ccNgLo0iv3tFI/0
rxjYWv+vp8nqIDqoE6yUzXxaN5jrY+Q7eUTrjNZ9t52trgq9VfLSsBS9lOWG/Ojc
dPSxzcJJ+eUb8z8McUS/oalcTf1xdygut4x8HiOcM080fvc3hjj91V8qHM2WzT3A
DGGQHeeoX3KDkGOvokb7ZfIgYwaIsWfgsKJxgtU1nAQIhPH6+6kRH3H7MVAhzGxm
3khWJ2IMjk2l/v43KcBbMCrtY7AIaSe9XsHCqfg5up40ngPG51FR8ldTadLlv/dE
nnhB20t63VMiAxXnUjr69oo94JlzJz9wMAfqSEjix/lA9mAFVxM+bE7JbQasRX3E
bDycrBU3aXOa3ZHlTvDL4aNZ6+oKHA31c7Je/U0fIVKeBAVAPlsKvp6DPqTWCX+X
m4V4cPcmn8BxtACdFXDFPMTYBbNWi0KBSUOJd4PJqynPJ5MTH4HYho/9OQ69R1Up
KOAZ2baBHwYe/E3gUddBWMCOc3AlngPQ9e0gkrttouPGpT6onKrmicrJDvfZJ4SU
rhxc0aEpqJ6wWsiLvaPymk/Wxr/Ef2BoyuokEdrsJPY9vn3XlbzSr40SjZ+zGIzw
9YFDJPs18aWZ9KUYFKJpfXGTGoYBRRmfzGXaYhldAnGbc8oSA8A8dIcmYWDIX8qT
bRMwNNk/zeyYSV1OpLxxYg8urDJN9mN8LAv/iSL9MMmQyjApsE5LrldGfHJmNQPM
OZEjzSMQZV3FQsewJVliUwB3UwB6HI6uedwQsrsvbZGyWGA2baa4rb7cvRiPVbfu
14H3z+MBBS4iLUMOOu10VyqqxISS6NWt4rK0/u5ATtmxwdUtohWySDNPZl7Z8JEG
4CtZzcawWtpExSLRzq6IUaVZlpREXW5UL9VRGPhu8s92AhUakX/iW64F7fGc47Oy
Tzdmw628ZLERhL3kO85n0HuDrhXLoXEjcZa49boYOkRGmqb5xyfrTAcsF78NrLZ1
qu7TRVUcDIaQ3uuRmTIWgKMmhFpDRbxxSwZY7466IH9AwRa9lsRbLfYlQzvUqOqq
KXH6fXuaeKMquSU/CJZb2FctjgUxYtj0Z0iteVJyiZpXcTXPbZbs5FidnrWzeuXU
cOjMJhZAOWoPQA+ZECRg4zz/A0sbOvABDFpkIoAzzQ1MOh/XhqaSTtyrm7MaLort
z8NXX7PbL+wmMkoJbWqaiAFtIc4inOJO+GUWkwYTaE48p5k+3nbhIMDVSnmJCHTH
Kh1Xd+ppUX+kwXH95L6K8WG84gJhu4xtcoZDQU0SJ0wg7Bi91cysIaFeyr7N9UjY
ZMzemJiX6rH4vpPp2uP/Ezn3LRQVkvYCMkP9yJYkBDPZt5FfeOZlQb4YavbBVQ2f
mNvo7I8loGcAFxG38xBabQaVIdjrWWzxYSKonbmmg38K7CWcWSjyNMEO2lou3h8s
1e1TW7mnYL8p3dJvTRDhbe3A4C+3IRA13KQddhKhYB3AU1/M8dLWjjkOG2yy6K+S
K/Ir5u8EnK1oVKGp6+AFnhJ8O1SaOb1XRkkRahgrnPUrdR9jg/2d0G+X+/NfChI7
B2X4bSNlEQTNIJzxblqivfXF4lgjF4dmcTpBDfdciZGTBjqvJoxYCVClDw4d4Wl5
Fr/+yn/MmCcbFJwzdEgDtXerrNy+m+0JNu8OMpn0ViqzTs+Rr1LB0765XZyNHZy+
s8woSGA2+GSSMb+klDgcd62eJbddbsdhMtlh5yaYzy3zNvJ/ofiR4tVjoIuYsR3m
DiuT94hhkCvX6lbuRKhtTfs/n5mN57Y9aRJ9eKrQwxkP/z4YSSnKsmfMwTCmeIMX
PAO2FNjRAxoFLLEqqL2MekF2aWI6Tz+18dcJqC0gX969QHpSiACiw5EVzpyEe6Xa
kElikeNM7uYq1DlctwvXhSPSvWZcEyG6rlYQ105LUspkzjG4+sxUNO1YV4bbwyXz
a58XeuSniK6JqbMWA3QUX0mVPR53z9ZgPEh7MbHpNtIQokQMkOtu6AHtRGU0U7OH
5NGMUp2kWoAMtSwQ9Pgj1u8cuzKtigQ4mBDw431/aQZN6yE3uCov/W/tv0B8DPYz
6PX8XUlAyrrtatg4Acf+d9uWV0YtCzchqP4caFC6xhSRci/pNrkQW+O2FM3vMlPA
PgOaQG+DlpE+k/3y4fVNEbmGowIZwWuOnqRHKBr+ZqCpwmq7h2IAS3bNRHaDWdZ9
pOepAgOXvZF4HHu0LEhgYFAZO/7zzIK5tcPf+xdQfGg/IRrn5psUt2PYCPdOTFua
7JyjE5BWBwsUuZ4Kh1I7qr5bnbUCpGasNgATCc5isWMtNoHlCV9v4/Z9X3kBFY2L
y3YEJUUU6ZOC30VXMh1SRICB1BKbc/7IupaGMmtOY11osPnoPBNmcqapsAItz5Pv
5qJ6CQCqt9upoTKj+4sY/+lN7gqwYqnaW0LylLxrR1UHQxR+RUOqwyTVdN+moUZT
rU8poMfKgGXPGnS4itHGncjRaocKumzfKj55+hyPg1YqsU9It2/uaTi6/J8n3jXa
zNfATB67q1I+6bjQr4dBBhclh1xvVeCDFLBGfuaGGok7Dkvb8ntidOJnuvnE55pH
Y6/K+lG7j8mQfwZoTUgVWZr5g4bGTfK8q3XAWme71DQniC3KBmyd6vWOgz8/EzKZ
y5B4pkuN4gKjNjUewWWv2FktYpPYABq64bN90whQnS77Ok8C3ENK5V69ZAmwtWaB
OJwBCI3lJk6BeTQx2h4FITuwQWJy5KUHUPj2reyCnWFoeZOsxVOqvf5PyFhsxaKC
HVugLIi6gaPWnPwjYpXia97RFMI7xv6hy6l+SrIfbGR2eC9FWxDVQMAi2M102PL1
5kSIJRI8mVKiNfshf4usnfOGJT2k3AdC84+z/IOfD5WqHbfG9SBxNF3ZNJMBZvMq
9dCxPDHIWfZiXmIHg2GGuxr0T00ZZPZT9BVwegFOq8PRDWRuVut0329UKItosIaa
1hjdvzL9+XMObwraFjozgJYxKHgXPhmZ7L0OasrVYyv5npfhq+c/jkjgFfet/3Kf
HSx5iheyVspAIwvr1hZVJr0xPKAj1/v1zezi0GwkvRa2NdBfA+Kv/BdEZPaNobaE
g7Wx2vu6trK/Q/f4yMt0Mp2RYz89n6FGHAqYk5mgqdCrOdg/6Hpwzw8xNgvmUUHA
NwhAv7NJ7hEp4Jcy3AuESDbVo1qZc/8XewSyplESw2Yybg1pB3G0IiYT22pMogoG
vrViR3T1F9D6hdVZwwBQypiwnVXb/v/qLs8D9C/RU+lTfaJsC6xsRsTqke+ds6CM
fa1k4HZEUQmrgrz9WVDrZ/lRYS4QQsfYFh/kiZGXmXWaSq1938sakyefN4z0HeJh
wis6VNFLZQz0ucn3NR+avd79FkZkggONrsv6y89Z6Ul53XLx3sua4MJzRnZ+N468
TQsZYTVr5uLUGqLZ3SWaAy53Xojesmi2B6Q1I9z2R9QEMg4mxkmd5eQPxLbl7seH
/xdjBNV6LFLsx2sBbvKlOoff0oyCGMAjY29eZDpZz+aPg8349H+5npg8ZW+rn1IU
CWLm0PvwqPbYaM1pk1Q9o7mpUZvmq5BuWzs9c4KW5KpvjzINHpmRp+veVcu46W+o
wBERMTEPzZGAo8nzCH4LlLUMvtJqmugeMrKHhGn5rOdQbOiO77dfXbkfkmXgHGCj
vl8UcmV6T65ytol/+eTFtVV2YNNp+omdfXwREg/4L4hgAVaPR56kZBE1XnLZOwYD
AdpRYPLf4ErioSd+f7jqHZclBnyNAnuZFZx1T0ho3iOb03E2OSMFCWdK6iEIvavb
CMtkGAJAV0sD3ualFBQ79jbHiwJVzEW2MatvRp/XYIwHAOJbbDS0/6l+HwKkb/0C
r6kcXbJnrFmtQRu6Llv0Dv5jCJc/n86Vb3DA2B+YLTY=

`pragma protect end_protected
