��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�a�ȝ��j��^5O�w?�cF�9}�ʢ]��� ���?0��k��j��c������������	yna�Z�1���������}}Ci�^E��Cd'>���$>^,�dζR�Y��k
Og3u�&�x���PЬJ����/m4����0��e�[�c@�a,B�8��?#	�+�:B�mh��2"�϶�k]���l����u	<�P��>��b!b5��%Ə>��n�ȉ���x&�r�
a"Ί[~�"0��]Ri�`��_��Qe�"^]i0�N��b������]�@��),o��RR�4�H�z���o����'��� ) �՜WII�6ʥj�U��7�&��߽��ɣu�!����6�H��B:��^�<��p�b$ 掖�R���(��a$NDd7�D��z�8g[^���]�\rT�O�?��v{&L�0k����;�T6o�S�(_�D�׼Kzf:���U�Üͨ��ς�`��b����ū��D�\�)���)h���J�����ꤖCS:R�GK;��\jw��uXO���q)����vA�7��zCq��@@� ����7�� ���>�Ҭ��4��@�����$d2��r�8����s�����4�%��l��C��&5F�YV}S�Ő��B�T���\�Dk!���A~�����&��<9�}܁P�Q�*m��kj60����+�tM\�vf��@j�`����X���'h~n�!�2�����kC�'�|���9�l_�-2��Gk��
�ٚ
�،�֠-�?X&ICr}$����yFi�ʩ
�y}�տz�5��:�XxC�*Z'���A���f�����ium�5q��<G��0��+?~�rJ ��\C�2�Ii�����IB��~_X�ģ�I�^s��
���D5�DP��S�<!�4q��ة�F:���z�;&�!��ƍ�1y"���VO脔�vw��ҹ�a��`k�zJE�����~����b�K}Z%��6�p�Y�L�SG *!�?�:�Q*���T�4e�\8��D��t�.+�Stp����h�ۚ1�&�՛ʃ@-�h��N�{i"R��܏ ���yף�ɚg,���w`��M!�D�s�a�wO7�����=m�h���~P��s -R�!�upu�`�w�J ��:���4�(��e%����@���DR��G��T��ND�M=.S=U�06�F����j�em]mI����F@�LN�w�����^9x{H�$������R�z�i���.�l^3�P�z{'ƊcE"QTS-����9���d�{����>)� ~���q���FZ�
o���ܴ�7�@�|P�$������<��S!�{�Ƽ��ƒ��`6�� ���c�碔�HW�q�wιŚ%�X�fPHbYʉ��S��9[k�Dy�a8͗�%��3�u^;^�W�dna�l�|��|�Ym`����n���	W�S�w�`�S��PX�h����"r1v&H�\
����3�r7�SA� �B��kԝ-�B�݌������P��B]�_�Vs�{��̰� E�������P[�Io6�4�[Hd��?�	�ѢR^8����|��(+�+D���)(U�
�Z�f�W��M<9h	��sz��a��rN`	�-�$�\'���
zROq?/��g�w<�V9<W$��u�2�s��Q��Em$��'D�߈�s��H�*
ꅟ-1�����z�A��S|����%g�tIhzQ�2�Q�ܹt !7�
����:r�����+<KuW΍aɕ�����P�\���o�g~eW�&ؕ3i@pLI.wV�����ζ�ߥ�Z�e�K0�����g>�n<��p�F�!�!J�Qs�zv��w��w�Ӕ^����S_K'uTǆ�T�7��@I����/���#ي��a��BH�q6"�t��XFHA�IK!^wj
�vB@�h��$r�2�Zdh��;8.�j�,>~����Q��t�;�Y�cA�&$���y����ղ󾳢F1D�~���A�2�����N�Ά:��Q�~/�rr啈�BYt�
�5�}�I�I��⤾�`�o�dd1���� `f	���?H���X#(�q8����.
T��t��.��.}vM��ul#PBe�fZeO����K6�K�c����N��Sl�,�
]�*+����?z�7�}Umu���4d�Mp����I�H@�*۸�#�Z�b;� }AE۠߯��ΈB��E�R8zR[f�O%��N,b��ޥ���%�[q��Tʻ��$��T�X��4��&��&4	�@���S��f�� �\�OY,��]��<�>�G%��a�p�+j���S��dy(�D��5�g7AVJ;���H,�bVH�~�Hy"�Vr���r�E�l��u�B��x���N�zo�^�Ihy�AX��n����#��l>��#0僙�����R�i �:z�Dz�I��&� ̙��eK~��	oPKA�4˞�n���uF���	2ݿמ�ܪM�e��D��	#3��>Du�N�q4��a#�]�+I�U��~�g��%����4���/F����������L��G����
"��:�y/���R�ҧ���K�˖�p�������O���ˈ��Nx��y�uX5*��(���A���D�G�m��ݍ�Ԏx������|���p!��oU@؅G$����9�}�Cp�S�t'#Je�QyN*�yJj���N\��!X\~�#��\MŘQZ�.Nx�Hh��m+�p=5~G����q��K~9�tcj
�����0T��(#%�d1G�Dؒ��ҝr۟�4�FT��7�$C���~s�8�H2,D��ktl�&�4m��%��<��ۃ�2���AJ�(�Q�+,��u��=Y��@��Bb�~����C�o���� �C���mK��d���q����V�e��N���z�"��
e�	�,1Mg�W�R�VV�y�V�%$�tǓlQJfDư�o@Ąͻ�p٤:�[8���c�w?�b"��_ ����_�C�_zԆݛ�r-�5V���P���8q�Ay�?C��똂'���`�OD�C!\o���lzuK:�SA�� 恷�l�?�G��~�1���5��Ų����Z`po�N�h�8�G���z?Oe3�&j͙�5���ڹ��ޭU\ˁ�����h����ø�RZ]�/WBxd�b���~HPG����� ��-�x"�n1�f~��`U���O>$?���n���R;�)�B�#�4he�PN����[Md{g�~n?������8�h�MwA�q��\+���ϭ2�p!� ��'��õ�
���?`6�iM��L����Z�~ѫo{�[�x�?!�K����w��n&W��_�l�qr�d�������XuS�ry#�)����=���x�Y�U+yH������Оvf�rO�U4t9�$j�'M�\Xe�S7V9���px�yԄKx��g��ʇ3�#�,@[~X3e����}�8��s[ps4�r�����$P����5ˮ��v.IE巘14��j��9��])�WS�_��._ʕ��8�ow���2K�c����g�U=��s�?�����7�Ȼ�?���N�%���l�]���E59�X��Sa��_o�|^%��9� e>8�N�J�!�l�*�)عN^55S٧�5��@d��K���ܹس�I�1t�q�4�
qKf+��`���B�����;�v�Li>��<I�t�9��,R��<���D���C������j,���Zf3��_�[�*0��m�3UwW��9:6UXB@�P�P��s��W������pT9d�a5T�ݑ�x�D�����s��ZN'�4��G�i��v[E�	Ј;��<nWr�X�#��b�	������twBQ�B��]�Ʃ�h�MeB���_��Q#�N�����1F��l��vS���������\��kk�rKq~L�RC�K*؜'�F�j�p̠����syzȃ�j�����v��M�F�F��W?�v����F��{�;�ׁj�ZX��;Y8�=���-��SR����}b#�� ��sС���RL �f�(n&�x �@dD��\�� � ���m���u�^,�n�G0�vy��x^,~������T;��։t��V�_/�뉯������#�I�]x�P�EU֕�ѽ6���N���%X'�ȐG�*�̏H#w�1ՠ���.|͘���~�f���+�u�ջ��3)�tAݱp�j��(��w\2q�(H�k�'_|��ᥦ<�)d��F^��A�B�h� �d�-P���X'�e{h��÷������WunӾA�\�F��G�+6�����ҟ_	]C�%E��k�A�V��`�y�h��te�G�P�=d��C��G�Ƀ���d�#�^hx�4V��'4?c�x�\?>b���n��S��L�iX��Y�D�����$��1�|'q{2���2��h�ת��95G9f��LbII��Զ%KwX\G�N��:�!����_�Em21e]&���Y��v������bKJ���#����@��]�$.���0���z�ߌ����iN>eyP��wZխ�2aUp�E�$����~�AI�����'H"�$��#.��|Lt<CFxV;��@Tn��[�x1�86N�Ai�������7�1O�gd�XRv2���~�^���a-$t7�q�{��p�;L�"*~��wnK/'����ʨa�p��D��;Ă�PL�a��Z#O�oO���(*��ݘte�m��oC���@�)�;�R��	9�l��8�@;C�g����k�{+!�c�fGbq�w���(� K_Mu��oŶd޴$ߢ/�lA�&�f��18ڔ������}�r i��V�[���{�HuH����ֲf�W��eayW�{u�]��eV�7���	,�l;��$�?:zɀ��&������aW�4,+Ŏ1=M��ϒ�9Ld�~�©��/��1�6 ������8aa���|��"�c/I�:�g���:����xY��e���R���H�&���Դ<Q�9��J��{�>��;��	`�lWB��e�m��G��)���A{�Դ�_|F
k���\>+�uKQq�!赖G���iu
��8��ߑd\r����_��t�yS� =���JM]���%����ı"��0cu#i�#��&�@#�����ߧ�]��aazhU�艵P����|�u~��)\V���n�Wx�\��h�Wo��0�R�s�Z{;�������Y���x���<�ΪKU�C�Ƶ��uJ_����:�B���v���8�����#M-��F����@�*꤅L�oKؗ�ǅ-g��ņ���+���r�$�p1L���{Y�y�tX�{2%�����S/5�'�xkɗ �p��`�Y���|�m����������#ߘ��Xb��%�1�#���UE��/�'�XXE�u���h�M��Ճ�t<hL�h.������%{b� \L2�����/��9O��b��X�!�:���@h����n�!�5��n#�^��O�Qc��_�{�������rd��V$��8�<	���VG�/bG�.l�K���{v��&��!����4��!b~�6m
�r�M,y/Ty
 :��1������L�+�M��O��5�Q�hh0�tSX0o.��8�0� �}��g	���~3�<�T�Ha�����=K҃���Z�t"�*}mcoʑ���������Y!7C�b���a�7���<H>y�*��XD����d���0_l
�;���e��-e�G��B�U���M�)�ƅ�l����O��zQ����R�V\:���9�%�[O?��6�u�GXYm�����n�phs�}l���DS����7L�/��W�mW��{����sEyA�xl����2��K�G����i7gCz��6V��"��B�/yM�f��E��?uA<Qo�C76�X��~eT���ilgIQ���7w��u�C����o�Tx��|�?�NA)�1�6G���EVe��t؟���x+"��/��t���;�����ޮ�7.�C����Y8�1������֧����G�	�v]���,�,8A�0�o0�Nk�MyOx������b��
T���{@�J�<�oڹ��n�c.��n �pO���SN6LѠ�q��Ky��q��}3a(Pz�bċ�	K(�:�ﻃ������O�bAc���:�bMh����Wvv��-O)%)%�����Q�g:򮏈Jk* �
j����6**U���z6L=́�e;X�X'�Ay�4�3Em����������Ed��kH����I.�����u:4C��G�"s�0��|ޅML�w���Ш1W��go�ɰ���/�0\���SEN0>wg�wu��	SrWH$�m�)F��F��w�I]�y��-]�yS�N(�!�"՝*:�6�8���_�C�!���W�z��~�p��n�o���2R�Y0�n���P�E}��2��E��w�r��_�cM����Ғt��tny=@L$�Q��JXu���o���n�ea��)9M����\U���H�c�l��O@��nr�D�6�|��W�¡El@f��aCj����X7r��Gl�m�Q�G|W� wD�⌲Ft�n�4��%�=Y�[����K�Z�!�q��n�ig,U�]vɲ`y/���A9�����F�� _7̆My���Sh4T�n��ќ��C�ˑ8���q����q?7X��#��� ��ͩ�٢*$a�b��e�����ۨ��t��)#1U,D5:�JbO�Z\
�O*�4����Z�8�d����%��Ʈ�]�
%����|t~æGV<P�Q�bPQ�))��h7�)�C&=�#��,�i����Yaя��v[�=T)��L��D��w֫�ǘ'���鳗2{Zh7�u��q�޿��a���Ұ�$��nAًa�x�Ï�J"�l�R�C�~){��@����4�1K#;���}�Y��Z[��u�k�����ڨ�c�~ ��q]�����O7u�B�T��"�$��noe/�B����Ђ����hd���l����<�Y�߸�3Wy�K+zo[k���g#���ј�.��KU�\�e8{���v���){���U���qGTyT�2����ژ��y0�sp��1�+�uO��M��w��ꌑU�E�@�}
t�J4*<Q#j ���Dl��?c>?��m��`�<X����Sr e֣a�Y���^ʊ�������*P�����V�V�2 #<������v�s��g<8*Ǹ��C���L�i\�`	�e��rJ�i/�!2iőz��8L�*�ikeDϐ���ĕ��H�i�ҝ����ܙA��C�>9nBVH��O�J�l\���=�LF����D����
�VƔJ�9VI�4*ˮ=�v�nY��w��R��ȏ�zۦ�`  ����t#��ٛ0��3q$�� �q��h�u�g&�K�Y�h-K��sX�C_1��1�+%� MT����o��=����J5�{%[+��!���Au������T�A1����ߎ�Ul�IڮlK��/Ӿ�0�?�Aڑ�� f�)��nFB���|̩�LH<��}&��3�1S5>�ul� 1�L��:]	7��$<���]�LI{^�;�8c%��2�mw������
�#!� �>I����T�����_��!�h�W~\���X2���&�8�4���F5l.z�7���Vx�9y��{��o�i�����H8eѩ����W-�m*5%��%��e��!�+������w�"	�h��/���(�^i�ZM�,r
i��[ꚝ8����_	)�+����܅����܅��C����������w��� �	th<a7[ ��?��#(h�C��\V|u�9�å$�Q=f�jw�������i�#e�7t�l�t! �2Lн�m�Ѝ��؆)���Y��Bá/��JE
�cQMo��݋h�4!:G:Z 
P�x��ёg6eެ�����T2�I^�=}�f�$� �
sx>Lcny.�ד��������sg!	��%	K���Z߿`с� f�����7��c^�)�Ž/�i<g�.��O��ؤ����oj����@�H?��#����1K�
�|L*��թ�u��	� �+g�|��?�c���
�<�r^�������ޗ�!alƻ��7Q���)�)����9�L!����Z]q�.��7�+B!;�E�%9S9>j�|���y��e�OK�����k�!�&G}A��٫�m�wb��!�1*sd�˧	��&���qͤ�]�qY�cS�b��eF~@�E�Y.����A���a�	����*#/�D��qtM�ɜ.y,�9O@s�6P��'lQY �s��3�d��� ��>�į�E����ܼ�^s��&�ٸ.��tf��#^��\�������y]^�ӆ�g�����S*C�/C�v%�g�~��r�����D�r-��]
>+�;�,b��H�*�?W[�����Sv��BC�pN�;ii����nކ�uG�nZ�h5��k��[�K.���`6�9~��)��.Ve2M�^YY��dX���K$<N��`y�
|�(Y<ۍKz�����碬F�ۺ<���SG5+\������ܓ�O��?�k��}K0ط�I�U�|��*�?�P�����e�@��0bh��lW�煉^�xE�u���>��o{����lTGcC���`?��>�?bz�T��eLƋE4i=���{�+f�.��:/�PX��g������-_iU)��P��>�� �-��U?h=�S��,*̥ ؖ���C�����yj�CD3�g��I*H�q2F&�h�wFw�	Tα�n�k0)�❞:�'�~F�5A���lּ'5�W�F?V�-����ߨ:����IXZg�"e��j��?Ƽ�a�|\}JQ+�m����P�"~��X y}�M#�ݲb����o̹:E3�G�R��ەun�!E����y^������x�W��&p�#�������T֌��:ԫ�X��l#�53ׯX��:��#\q��"�~�˖����Jt�
�[j���7�ZDo_ب��EH!�¼܊%�������:���Rez�2Z���k�6v��f��#x��b�$�WcP���<tTPUU�jz�h1��86����S�I���F�i�~䎈>�z�Zw6 �j��"Y�*I"~�n�@�S�
�č��a�@H��ԧ�����"��>]b~��Ҽ)n}�$� cpX��Ƅ��}��:���S_}�ﶆB�wc�y�^p����Nҷ$�.M�"���:a9� �Vt�'3���G+�"��*&�Y�щ�@{�Y >)ĕ	�%�J�\'Ε!��V���6kr9�|so�ݡl�3��h�Q2W�U
`N#���On�W��WN�6a2��ƶ8o�2�rE����n*ԝ�OZ��I���6M	|��N
�@�a685�6�Yn=�%���R�> ����v�"gⶒ�%:���|���Y��x�Dv&	���FK/Λ%��cŀƼa.�Xq_�k�Bd@p@v�>@rJ�3`p:A��uЦ�Z��Dҽ"[rl3�'�XU�[����q��>��.�)9G�ބu�BA���9q���P�İ;ۍ��g�>�d�˻��G�i#�G�m�Ɠ�G�[&#�`R�MK��!��� ˣ�jwM}��1כEe���Rr�P]	�m֝�FJ���
��EV��"?IM�\�օ쭃�;w�Sp���j�}M����e
s�u8G�/~���;�=1�d<w��G���I) ���L�Fި!A�m͈���-W�`��a���y�U2�#�a�6�4���>��i6�No�pÛ�i�� �[�<ͨs�4�����dg�F7p�v�*�J����c���7H�Z���h}�<i/{�� �V���&�5�=��q����-�N�v�x�V垳p��E���$Ǔ��
ot@V��o6���Zˑ��$�C�����D��P��Ի�N�n�V�$ˠ��(f%���B�*&��œu�p�
9��������Hʸې������:���b�vk-���O|�]Hc#
\U��[0u|{�k!
&P�j�-�=����"r���:-�((6��Bx�I�c�ms�:Yd�&�L�p�&}���Sh���c@��""`� ���@�7� ����~'��M�;��=�xzԓ�0�׉`_����RM19�����NJ�a�{�V�@fڗ����^a����ZTUڸ<&w[C���1Ǧ�v1�.b5�[�d�IP��$,$=@<�T ����b��s����K�x�Φbx�u�-U*������9xM�Dh��;P��&~�����6�P�# h�kV6�G=ږu<ew?�*\p9���W��)�`J����>��DQk�m����U��� �Q�J�]%*����@�T`)f�\";"�t��Y�����=�UN���,��5�;�yL*T��1��*?rZ]�R"Lrs~�Y���J���i��)�9�ez�������yC�-jd�ső�|ymp 
k��	F�~b#�͂��p�1쯌fJk���VT�4�m�q
��h&h�^���wp��dc�~J_�y��*
Lau�֜Y.��u\�Xȓ��P>P��9�K*"��t�(�@�+�6=s�e����l��<)�D��\�*�2���a����� �����U+�M�"�v�x�@jz���������P�N+�g!�+Ur9APw2u�f�2g �����I�a���{�ӥ�-����F�߃��m�bD�� ��1@�t��5�������BI�I�	ݫ)�`��n�q[}7pQ�7��Ҧ`�=�ʖI0�(����*q1�f��d�)�h��N��4��甍��疤���0��B��'��b��ǫ��u~��_� �<��+�P/4�9oZ� �mf��٫�������H��������.5�:�Vh��f�q=>���{ ���Q��\�M)<M��K��HX`�ieeS{����fz��9م�[8-�*�E;�>]߯���K��[�z&��T
��ږl�k�h�
����^��/�\{A�1�̃��c�͑�׀���o����\�~
�Psv�r�N�w�����RM���^'v�F#�GXA1�c��"���{�l���s������a�g,a�R/A�&8��5��G�:K7�z��u�;/ ǈ_b/���{nR�&L`�����&�#�v�]{��ܮ�AI���x���)W͔I���>z+�B/U� hC�X7�^���ĹS���B�'�/��.�ۋ��G"��?xXN��2�nZ�[��/w�2�be�9��E������l���g|�M�:�W��HkG{OnB,7���}�e�^�)��:Y�������?!EA ������b� ��@��B�y��@�M'�a�n�v����YX2O�c�^�"�ƒ �GdGv/�gA�ん`\�,tQ���u���%T[<^E�A��XK�PI�u��5 �B�����9�%����D8��(&�
����.�a���Q���G$m8��:=�?�3e���:�b�\L��� |�nd��fTK`�1��g3 �iaW�sۥl��lzn�Fpu��f7���/Ņ�H��{�Rqy�A�ҳY.���Y�a
�L����Lﱲ���C2��cI��N �f��y�����{�SӜ���KGe���Ugi���њ'�L]C5�ͣ�c�����S/!�m�?k��΂Kt��5�u`v�㖭�`Z�d��/�y_F� ���(�6�}�|��;���>��(T�X~F?Р�7�m]b��'A�.�?<A��M�P�72v����u�T�$���l�ץ�!nY!�|���`ý֓���z�tY���<�L���ZT�����
��o�ɡ|�HʖA5����[M�THBb���J!�/��-H2��5x(����������N�-�I���i�[i"�����HH�hg��dǭ�Q�p �f��0by>q�����@MO�0K$����� {�)�j1
��Ѳ�1dI����3�&�=�p�pI&���UM������qq�4����{��Vh�[�93gL,��5&��~�y6���IT�߃Z����n�dV��P�]����D��i���s
o]p�~��a��J�L����*�Ȏ7����`k0�	�K��,��Z�3��U�7~��ͮI�,����@�0Ļ��[IJ3	��	�Z}8��A3��:�|�X�C�����Ķ��p��'��P�T�4���"�i�	gY��;	TLn;���=��Kv�Ѩ]�!Y3�bW��vM��:�~��@1�
��+`��ue�P؁��U�F"	?�7�@2��I,�!E��
��D黬����
����%H<��OA(x�����1F��Y�!��y�z8���).)��`Ї�_�sE�3rT��0y�#�Y ����U����\E�Y���Hf�,H��!p�F<�k�ޜ��?n�ˣ�Y�U>�Y1_�d�oJf
�VC�݉A��PH�ƳuG2��k�f�M�?�͇g�k���o��ƌ�a�K+�8�j��A��'V��Ry�[]�D̶P9-M*o��Fܐ�z�8|�����40�|�N�'ˢ�`~��Th�ړ`90�)?;ڳ��UCi�&w�Ҧ08���bh�k	���p���`_W�?��J��8��/3Qh&��9������c�N^���E��Qm�FF?IP�F̛o���B�K�e�G�߻�o��g|c�G&e��,��֤�U"�wlb�6I�$f���_��r9]��֥�B5i��'0��n�u�e�����5W����u���*��4���K��pK�9�����!�ҳbj�*c,��s�r����y�ǻSO�z����u�+��Z����� (���U�@=���bz�ջ����Z���5vwy��l�� ���	�[�����¢B�n�g4�<K�YZsç��=hxz/�Tj��~���f�Q<�:�0��$'�-g��&=bνc�$�O���z�|�@��]
�Fd0/��n��\N�'K'7��*�����LC�gt`)�S�ڜ���棤����\���:�D�w(3�A[V����PR��b�Ä�E�(tn��6e]|k���tF����Q�ݗ�fHz�@S�D9��I�ƥ̯��s=��[��f��Dg&!���1�s��=�����c�Uݼ?$L�x"EŜ���/]1*Xo���IJ\T�D�L|�~����Q�ڀ�1�md�F+���/��C�0��%��\XGb�}�S�;�ʐ-���"��dX�� ��Q�G���-��m���?8o�25P���]�F�,�6n����-�U*\IT?6^�2�N~x�j8V�r�>�L1~��󂄛�6�����X���xj�l��8U>��c�z$t����Ġ����K����]���p�l\��kn=�կ37"��:	�E9�Cg� @�x���Vw�6�[��$����P'L�BE�"{n��V��F���O*����4���k�<QgoD��. �����ۂ�e���.;�������KabE_�1��3�Q:�G����V�頫�pY���/�Wp�����ѽ�������CK�\� �A���ɨ�'��!0�X�{�J �U�qϣ�'L�p��LE=_���9p�4�\?�i � Y��k��Xf�Z��y[�]��6�b?Q����[3�㍉rS�)6x���>#�czM���A�c����m�����Ra�*ݸ��������nm�o;p��όb���C[�3z�L� ��7�����3�`����p��ύ��O'(�|���o1,�9��ʳd{ �h�}��F�4�ڗ��EBर��Z�v�#��Y�gDM�ʌ��x�nek4��H�F_j�K�A���SiW����a�#��n�[r���{{_m����o���;�F�������jz� w1>R/�:X ����
(�|����nQ���D��Ulmw>�|cp%�os6yG�Y�.�y�͆��˿��ӮD~�g��8_�[�XAqc�o�A6@�tǴ���٧+m�F^�h��)�CH���{��z�A�3z��y� ~�ߍ�,Q{�F��]�y��Ɇ�ɬ����}ݱ��;H��=���T�e��誓G3�	�b9 ����eLM�{	�H�j���F�ɂ��#n➺}X ���|6B ��4n�[����4CR�����P�GwMXhG�'�I���3>u���a��`�פW?"E�����i�T� �c�FY�~��δI��cN���}��~o�T�Ն��@]�FP��=�(�@���9�mۈ�Lw�?���vBo4���z�xn".�E�� ��Pn�.\�M�Iâ��Օ+�ɩ� U���ʩ�����Q��F0]������17c�����)����뭭�#�?0tr�.w����+K��f����ܫo�<z,оss�,��@% ��FK�	���ҵal�i�$����@���qk�Q���Vi�PƘ��e��x���D��T4?e�;����1/���!�_oՃ)���x��iL%��b�ĝ>�x��tx�$Q��bl�&�#8ศ�}ws7��=?�zD��z�8;3`�E�~	~�-or����o��oO�$o-����S�ه5B�Rv[x�BN��AO�=B	��ϸ���խ��Ѥ�Y{nq5o{�]^\�
��[�I��9���D�8[y<\OFe�	�Ć�{�N-<�p��2�+�w�?)ż'Q�T��2��8�'�.i��T�����èS�6j��5qɊ#WD�t��Y�TiH�!�)���A�:�p��͛�GwG��/{2�*��]�Z`�xz�0I���[𧬪(3����g�6d�)�M�q����p#µO���侠�$�eW�=�?Tb%��U&�	l&����f^V`�%e�F�>0
b?�®� �K��~���{����Jg��P�����T&?y(�-ŭ��Cke�Ed�����/M��8�JҜY�i��sSĪ�EJz���0�j�X�7���_�l61�;&��]9f5�YC����I��0����
�A)���ϹU�x�(�b.�Zܘ�r3�Y�b�8g��^���5C�/b%1y*W1��*�s�Uz*��P��ȃr�WGa(si
�4��k�o��-zV�Z�O������4S
�� ��~�����u�����w~,K���@w�k�ɯ����e�k���.�d͚yp7�u������xL���1�E��p�� �:V�/`܇�ƙ؜�م3�mJ�S��s�/���7�Dhb�R��O�P� c'��d`-�/���=�6���'���;@�¬��X�M��ۢҳ�a�
���/�3?��v��Q� ��4��b�?��qFgrЮ3��g%~�f�� QY�o}��	mn�{����o	�c�����F��|��gE����-�c+d9&:0�9�i
%J��q����� �c��)��+�������Ƌ��Q�e�6c^���姈0YB8���9�d �ɡb��u8�\�ȟI8C�Y��g̙��jB��&ɷ�R��'�!�y����bV�(��#A4�~���N�z��zd9�m�0s��r+Qy7IE�I�Q���P�׮��@C�·\jħ\�I�iϒj?�"=9���*X�N��5]y�{XIs�Zc�T�jM�K�s)��g�:y�o
�SRq��Y��nϓNg���;T��3��d���m�7�=��0g�_W7�.�SOmͯ9H�ɠ�����h{�*���C��p)Gh����A���#Q:�FpD�XyFd������R�����DىeG�1K�H�Q*�t���5=�ߚ��ą�DB�Ԁ�������P���Ԑ�!ΟT�����Y^5RS�b8n>��g����O	����*T=�c�Mv�q%pV���9�ⰼh/�)�v��v��!}�(��U2䠃�����U�)R�X�n]fJ����&�U�F���t��"e��c6�̛-{�S��]�[�ΌJxgNr+�ꨦ�Mb��:-%����uDҺ}�B��Œ�*2 t��W��׆������S/[�
��� B����0��p|lͱ5�6�'�^m�7:�sb�u��.�ha�1����K�Ym
��o���?5��e��:.]rЁ�	��%����!����9Y�]}9rc�. � -fq})�\s��g�d&�D񞾛���7���J���?Q>����ƣz�k��PM��>�C���aҫI��#��6������nc�=���v��2�z=���_�Ӕ�{]_�lZ�;���A:�z��lՠX�
u4�E��$�0C����/7
(�h�� �;��Vf�� �u8>�-� 塱��y���W$5Aw�'^N���՝w�NFvB�� ��Wlm���W�`�.S�w-|��0>	S�����