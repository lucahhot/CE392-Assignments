��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�a�ȝ��M�(�A@�=u�R�%�0ŋ �/(������'���2ǽ�{c�ke���ml]��$C�w�=:�n�����P[O#JB&txq38k��r���#D>)����FQ���u�z�&�_(�Ί�`���L�qR(潍D�ܔ�G*���=)�O]�M\��y%FI���hlԆ���QE\�{���5gGuC;��ԓ��)�����Ab�U����U1F�Y��zki-j�����)�֗uҰ�+���v�YQ�1���\�G޼��<4���q��~�}5�~(U_�X�@Z�'�h�8�tvS�R
�]�{�)�	��U�Z�Å���j�orT��K�cH+�V�gXч)�A~C#]�;9̴�;��T��M	w�;��?������
+!*�&?�ژ;i�h��WHS/�^�������Hvai�c�Cm�Ӵ�eT��ʵ��/��+�������{>�KZH; O���:jt�QB)}��
��T��n%���HmF�%�G滀v��w2�{�.=�R��q<p��b9�?�J��Q��f�k �;oK�B1��U���z���W�t==�����Tj�����L}��h�Z����vg%������W=��ʚ���d����`�Y}�~��q�8����@'
v�S�gԤ�+kh-�︓�����脻�#T�7�ͽV[�]p�_v���5��;�âS��b(U֬-(�=|�?eg�K�2����ϥ�"�>S�G�@ 
�]�i`��*/�F��@���9|��71
�Q|m��'3x�d�&���ܱ')�hŌC�A�FE���+_�z�O��ijY@UZ�3����9�����6W��)O�ۍ��M��d���u�8�J@Ľx�WC����HV�l>�2Ē���%��\x�?�,k�
��p�j�t&b2�7-[K�@�Z�da>#�s��6���%�ǲ���__�'�}3�W�c�'fex�7Q���e�k-I�3>�>m��k2��2"�7�Fi��㯻���GJ��lE�k/�,�˄�!Cc�'�����Bm%���򞃌Ǧ�ϖ�3ȫ����s`*��l��N��-w6J�����f��_׿mr@��W,?��B=���tS�D��5&�R�쫥Pd~"���Z�����#mK��������[e7�ϡ5x:w��H�]�%@� �5}�Z�`	d�؏�[�4�#?�[:�C��QTZ&��\�\2�����RO��@�0�lV�0e��t�R2���G	��Ra�����a��i)�����&�#$?\Q�����.����kU�a9�\��4��B8��D��s�
��:��d�2�+2h̸CዜNED�x7��ƟtU�\��Ϻ�R"���+"�����h*݃��]�;�*~�C��W߾�n�n�3r���9�͚ݢ�[�˼I-���@���%�é䗨`P��׳���q�~�ܦ����qq�v֍�#�)Oqzŧŝ���[���o_T�%�
y���
�:�'��YeX[X2��h�ξJ*R"���!ǒ��g�(B8w�5,���aٲ��]�` 7eN	'�ώ�2�{H���I��&��nD���Z�5Q�+��ؚ<�~�N����H֞��`J��gە�n^B�r�|�>5��<���_�+/�F-�N��R^k��!Ǜ����}z˙����Z�~�����*�%�<="m.�s���H��U����cʴ�0�c8��*CD}@M�vL�L6�����d�i��=�`bGG�3v�/?򠮗�_�����!V
@�)���2���������.o�蚑�zK*z�r�=<��1,;���'��T9����M�#�x�kT7��:d�f��'�`�*s��a����[G4-(':A��@����7#o�
�v�����W-\�0�/�t�����mo7O����� �J�{�>h�#pf,�nɬ�ߚ|����]זd���tF!��X��S����\Lc��>���M�i�A��LԼ^b�"�����b�5�S�9(�W$;	/Î@�!n��ȗՓg�(�Pٞ밖�/H2��3퍴�0�먃c���^]�����s�*g��Dmf��8�;_x����d]���Bs�*�]��\ Sk�þ(�=��t��PR8����غ2#�ɎD�������k��;ȕ���f����޲�8���'�F��w?��Ij��{�e)�a��� 7{x��^Թ��~�)���ЛNJ;=�+"c8�:���@�^���Q�{�[p�wwv� �����o���!�Z{��Ћ�o�Ig�u�x�f�r ��pm��F�r�K�`��l����Ū��_���$�4t t�$A��Ƈ�~�SN���:%����EOB#�W����3f�����$�������9��1�_)p��L9t̅��K|��h�{6���]z� Ӭ<q�P�c_ c��I��1�����$���Atm'��}֚����K��4$x����O�Ԓ�~fE�Ěۭ���ѓ�ElL��U5����[R�:��ԉ�D˯_[��Z�с9zX�Y�W;�����>w9jK'񐌒$N�) {�-1pb>Z��uksV��)iW�X���#����0���@����'�U��ܢ��B�1�ۂ~3X�(���L/��1�
�B�p�P�$���ʺ[��hK>/�4�!;t!��:����M�@�s���������� �g�Ƞ�V�F�؝6�5_�m���y �UML�Y�Z���Q � r��/��]#D0�-d�E�fAGAG�@��44��y��-���T�8~�*4�~�]Ė�ZÎU���<��ȫ�~17�6�Y��o���'f0�VR.}�4Q�y�}'UV�� �B�/;������z�(�R���]��&���{[;e*��F�>���ῥW�f{0[puvE��f\�L갴�>�gYY���HM݌ZN��-4�YW��ڏ-�[?����{c�(
��Ht�ҭ������}������6@�3�o��M�g�K��6�G���-�7��c��-�)�;o@���c�H����YQ��;D%c;Τ��,�jP�u�#�PFڳ}ɑ>���|AB��F^pxLkmy�B_z��n�nܳZ��R�Jn��0����5]G��c���:<�E;D�"�ma��oE�W���b���ݰ�,p=i�3��%&p��S'��B:�=�5G�^.Qs	�n3D8�A�}�g�:�AL Q*t�������A������Tx��]!�L�\��=S�����������㊓e��k�����@�&��ݟ������� ~��T���K�g�+���=�S?~�N�&Ŕ��.�%H�\�3���8\�+��ˢ,���)A�z%D��[����jҪ8,O� ��Jzbtv�c�<�y��%5a�"�Jӿ�7���hQ�ta�c�h��e�jF\LnUxR��`*G��A�H �,m��%L���J��/�'(G�X�{�g�!s�!���~�(+z�
��R#��T�5�lFy����{��3�Ox"1�Q͟k�/�,�V-�]o�p��+M}nu��>�8G�N�Ё]K�"�a�߳t�{<1������Fk�
��C2��>������*(�p1K�{��#���7�F�b1`_�dv�õ'��&󁀃�7�Z�#$�ͳ�u=�g#_=��i6l�6��Og��>t��o�U�{>'�s>^�N�g1���D��V�O'��|��z7��F�ÿ猗) G�U1�I����j=GPQ�m�^�lZ� 6����w����0y���YQ�l�h)t3 GB�έ�Ew��R��1�{��$�y�)���s;Pvr��c��O�{�%=~7��G�[H��Qׁ��|?Y��{斶EX��x:NɈMU��U&�x��[�R��獢c*[��6���2xHѴ`�K�w��{n�E}w����TISe �[<�gĥ^p��6���B �{��!�y\��`�8�p��_A�Q�º�˯4koz'��X��_��^]�3��#t\V�}�5:#́��K�S�I�M~�e�z��W��U��1��Ę�1��l�1��3wE�݀&hB8f$�����U��f�o0�`�[:�����|�o,�VcԱ�e�l��A�� �ol�I����-���p��R��5��c�I��.m�0o�m��/
�y�Cŧ�"�.	;ͣ�����ÛgD�ѪU��Xܵf��RrtoM�/u��ʛ�(E��d<�j֚-.y8����#��$�*�xpt�.W��#�J�*0&U&��H�;Xt�c���S(����՟ʃe����F���t(��-���ݰ#�(���1�Lf����z;:���֪1���J��T}���������`�`�����:�+�vb��χ�fdg��t�+M�̓c�J-��&�35"xe��{`UeEF�ի�y��V������g(z/�:�~��q���9`6߽�j�>���@�pp}�������,,��S��"�X��g��8�$��u�E��dam*tǎ[�!w,�7�W~�\b�+:��e�2��R�grF��G�Ȏ�apRO��	#�Nn�)
��{K=7i4�!|z8T�@�)%R*N�]��� �n(�SOa�z"�;�e�E���2��h+���ؙ���b M�a_����S�Z�:q��Os 6�"�h��r��&0�7ӻI�Β(x,6�8��m�Y�5)���L�{^����p�;Qk�( �t�e�����+Ac�2֤[�	���n<Ք�l�FA��14�Cd��8>O\�e?�&x�3�o^��+#�Ƈ�
����K5���2\z	z�����&ŽhQ�F��F����9[�F�J��=\��(�Ay���z�+���0���#Ci1�J����G�r6}�v��p��q�@r$�
Xr��v'ݷ�y
�y�1��[�Yܟ�( uJzEeU�(�K<Yr��u�Ɛ	S��0��<n;T�����^q��R����d�����yrk	�s��~�I�>�R�i
��\��'u`�Kd P���M��g��)��߫	���C��0&�.�M�T�wc	D��)|�Py���%�n��Td.^ߟ\�a��S����v�ӯ�r��G���M;Ur�5�V����km��iJaU��|�4�mT~��Fѝd�In2��m���J52(g6�����@�� ���J��by5�Π�.�&��p�t�WO+?<�8&�P�m"� �ʯY�Vީ�x���Zp�ڔ�IH�
}��{�|s����]��t�WK��p�!	PXM,����p&Qi%y�8#�dy�4�	�ưKe݂C�����*}��I�%~�q�(�
̸��;9o-%����%6Y�֯��8��3!�ۆTEe$C}���{���t�]sCiY|=��:���Y�8�z����vj��%�^�����L�L
��(�����!�g"�s�6u;vJ�^��MǍ8gWv:u��;G��m��JfB�r��0Ӣh�>YӺ�޽��������"527(�:�q��w��zJx��� �
v�K8;��L�v="Ҹ�X+j�|��;d<v��0�nEm"�z�=��Lp7.z����0M#������rkCL�/��Y��Wov��f~{H� 4'����H�]L��ǩ�l��#�B5��>A\�����t 1�zC�9yD6xM$vi`Ƽ]���#z���e.1"�]K�ư�+�G �c�R*�LrB��k��*����,KГ'�w���Xέ��ދ���2`l��_M���'�0�D�5��jd}Q����~=�No8�J�p������ʥTs9�9S��>�w�� �w#\M^�ޞ9F��t�S16l��E2+��j4�� !3.'��Źץ���"��]��Ŗ��5xg���V�B��͜�p�����_���t��2t�k�.ya
����E��x0x*�X�گ��k7�V����8�u�OG�дOH���F*��L�ej-�lĤ��aeKj�+�3��	~k˖�s�Ӌ���!�:Z��y4[C�/K�oP���Hji;=���9���|��[�>C�6���͠�O�RlɄ.'l�X����U7T�X!m),�[�@
��-km�02��CfY�����o&���,䓟�J� g��"V\��Db��Lw���>�H�|��ʔ��`\ZK��Q�>��j�.�V>A��$�/�˳ �Of{d�����	��\8M�T��q�ph5�E\��\A��܍�V�m�W��Z,0�Z3�\��r6���p�����x#�$O#���o���n �Y�g�p?�Vg��F��<��6-�lN%e�l�Qe� �o~" ���%b�<խ�H�`j3u3�|,��lB5dt~M]z��o!옗3h��2k�!�";r{���o6u4�`��J��/��U�A�U�hU�r
�������H@v}�S������}��ݯ=Q��%Ut
�J�P$Z���	",��
���H����B�}�|��"��M6襣�+�W9z��#�E�1�|�`J�ۍ�;��Z!�/����r����@�mo*)ҧţ�X>��q�^��8o�-�	���ŝ�i��n��搄�q����_��6���O�j!S����sf�)g���l��W��"�T��VObD�;����qo���������A�Y=q�s��l�>�@{�A����Y���p�Ơߵ�D� Mf���N��4~u�Gh"��w�$d��1����������ɓ$��h+��)Y@d@4�)?i\��5ZNCP��׍럍�=%|�f@���Mυ��R�������I���
�Vь��JC�.�	������g�W@��mf���<y `cgE=z�nEUe��5�y8Ɛ��b ��W�D5�:�.˘���օ���^!�?ׅ��H�z���A�⽴��k��H��(U��Z���"Y
��HS6f��ʗ\5��J�O��:8�#]��˃��{"�P])J�Yi-r�4�e� �Z�i2��P }�.ha+pfE�6�#�c��B�h����9�� u�z��KXk	�ds�I�`.0�����jǱͅ��و��G�uE�>{s��W��+�cr:�:�	��y4ȑG���1S�t�)��y��U�ε�:B5"I�`%Ƿ�5��3p�&���0�	dr��S����9E����m�ao��p#�?�ؒ�ꖕA`h�0��t�P��-F����̌yT6�Jlw-U"�G��4��c7��p�?�UL x3�p���f*9�Z�����E`�
3���K�'��>��l"�$��&��{���ݨWp�p+����CUW���df��iYvߙ�b6~�����$�/����OG�ի�|�}���V��0��������f *rc|�f��˳j�P�
�i/�}=-L�RG��ϰ�@��54'z����C���c�-[�9f=�G��;��M4o
:r�Pf5x��g\��`5�$v(,�e��B���Q�1��i�F+���h&�Qs6�c�\���K���('dZ�)5f�;'�>}Q1ΐ�$0o���8I���$yRX�'\��Ã��Կ������z�1\W�U��"y;�1��eC&�l||c#��{�M�{�,��5�-��hQ�£G����$V���f^�
"�<K�"���ȁ��l�����a���Ȇ�<��0���`)��=�@�#/��V��Д���F�Ȝ�����^���k`]�[�7�HF׀�P�Bmw�|���v�.#�#)B�[��Fz��>!��S��Sg�#l59�Hl8?�I��a������F4#��ߡ/�,p�޵O�_�,�-E���loB-��m6t�������[cR{���������3ڛ�Eň�q�E��i"K�[�
RWԷR�>��W���w�h�:7ӛ�R�"S\�9�O?��Jr��'�?d����oL���:�K5'������J'��vo�/�h5!:�&�o	�k��U�m#� 	\�[����%{X�������PN�Ⱦ4�eMA��Ǭ�W��Zmya�֖���Z���x�+�w�][�t�:Mi���K7�I��j��=�\��N^����1��Ϛ�O�'L7{��/���ԐiC�_A��Y��ݑ���e�Oa�}�*�����.HD�A�&M����!6`��UuooA��{�*��%�X�)~���~��ݡ�%���@�0���ݾ��Z�@�����AbD�:�҈��˴j�&?r�������K��R�K���@�4����g-�<mF��8V'�Q���9f��/�Jܗ+�^�T����x9�1\Y���T�����Y�>M�E�	l��ME�	�ҡ=W}�����'�����9j!��:�8bZ!�`2]�cx~��������P�ˬ�
��K�7�N��J�x��I�|dԈwݫ�Y�|Ŵ�8T���v��{����s+I���I�� ���J�|�TL*gV��e����=�x���waB�k�/d��1{�O̩�NG��#���6��ޔ��/�=bu$b����3�)������^�߽�I�7@�69ο%�$���&�$B�1�\E����4F�`����8�I>bʵ��/-����g���pN���3�����h�6,u��6��л�sK�9��!��0�t�d]Z߶N�k}�����>�rY@4���䂤P��9S;`�=���q�v\�����	��ɯƛz�����U�.s�5�y	����VO$�^�DbM.xH�-�)�PV����XX�GH�'t�0��Zk��z��c�yc �y�q�~Z;[^�g��+*���#��'�e���D^.E������v kz氫,�����%?9Q ��k|��H�1�b�]4%��J�?����d����^�/�����2:k�	��Y4[�*M���F����둫������}"Ɖf�we���{�,)�pBSIT~��:���Ч`A�L��Ւ�`��8�*�<�ںB,��~5:ttq�=Q�z }	��R,�.7yCZ"�\�K���sma��#(��(��JFo�P�x@�Z��(�q�\�c�t�$\�Ƌ��t����W�}u������R{��G�ͦc+�]�H��H����!���l͋Q��p��f�YAq���m�P��3D7�3�|��q�)'�SN��J�5���E�ɔ��d����d���W�M��W���獄/���I��G�+�Յ����E�_��V�]�����o���F
0D�k�')Yo�شe��p�G!��"��]~CL�"m3_M��e��L��d���X.���(+�t G4�g�S/��;i�'����&h,u��u�&�!@�XS=�z�cw�I�%��݀����Aẋ��U�֑�J�8s����@;n�O�#P��h�~�{;`Y���\^`�j��(,oEz�0�+T�+���O��#�6#�P]���o`�{�,��'�j�SPi�/i��s혗2�f`O��Ð]����Ʒ̪���]�K���`:	� `7�P#���Ab����5R�t41Beg�����5W�c���r&��mM���Ƨ��!#����p��}'�G #�:��W���:v�SPX��3+c??#A���>U	�� �6ʆ���|�g+f$�G'e}�1���YA�S��'c�HNƃHϰ�tݦ˅!&l���TLPx���3v�|��r,��Ǣ��a���\A��I��o`_���/�:��"s��^���~pgEt?Ҫ ��pk���?�Pv�âU�-"��T��ϟ��ߔ�����?�6���^��#��h؇M�?rhR�����8d
J_"�j�ڤ�����Y��6m8&l����t�Lb$^p}���S�UsS�7��D�B�������:�F�f8:�Z�:��W��6��}��=�y�ҧ��i)A�]�(M����� (�1/qp!�uFʜ�;��} ��aܝ�99��Q�[��O���'(�6~ڴ]�UK}z��@�W��c����=�}D�eG?��q�g����@����!�"U�[N	ծ�i&�x��vL�83������S�}��*�fp�ͬ���<�Z��a�8�66ײ�5ޛq���8������B���:���;ݘ#&wGh�vo���m��F5_��!b���/ċ](�sm�:È��M9��E��Q����){X��������&�Кa���6����
�a�:�**g4)����� !�a��,L�#w�9I���a���BZ�d=BP�f�4_X�eNO;/ģ�7��.�}�Ԝ_�DU+#�w;{��Z������k�J�O�gg�a�d��a�|���r��<��&�h�l�nR���a�?�w��*��gZ|�&</>l;�ő�,�,S�ۖi��+�y���c@��>CZr��F�Qw`����!}h+Zq��^k6��!J-:��;��l����W���Eyq]���	��o��
�]6��(麮XE��%�ML�Q�r��g�1v/T�5LFɫ8�.��z����u��7�wC�,x�bFe5֦q��3>�a�Dܤ/�-"=߽JZ���>��%��C��bC]��5����y[H�t6� JC׭�Œ�^��w�_�[��~�@�G�:�m��,���4ϳF�%hfQ#{5��=QM
����~�(�q���
�#�,"��V����q`uSyO�Z�lnʨ���%����ދ	n���E�װ�Q�z�+2��dR���4B�j@��b�w����n�c�8�x�5lB����,\t��9v�~��Ɛ�#���P"���1��.or�J�̎����}��k*Kg���8[����f�j�Yy�dkw�4Uh��iN����,�R���!^��/�x� �Q��-D5b�Z�ɣ�9������6������M0L�ȵ^�Xn�X�Yei9�e̊�ޛ�H���Z���|(���&�[cU,�en� �"�mnB�1���:~�r��J�<�J���6r�I9�(~�o�L�=",�n��`�zdS3ѦH������BPe� Q6�z��K���3��`7������U�dр��U�&>a;�p��av&n��y5���t�m6G�N?��*���^��5�AX,cyV�KjN'2T���9_1���>��N��\&Ga����p�R
l*̄K��R��7���0�;���hu;�4�t����C��͹7��Im7� �����!敕q�ôވBs�Ò�Z�1U
.RH?.�'$Z�(zI�N�_�TC��W�גvm�G��ZDT|v�nE:ԅ�6DM�@�F�h�ٓ�LG�'����u�q�tx�3���c�j+���y��Z���>
CUl���l�\s9��w���NK�����c'�s�Ƃ�d��
ǵ�Y�P�2í�;@���`��}������j�J���H�����ދ��t�Ӯ�{��$
�A�J�F�*_}/E!��pѱ�$�Fiɤ7V��i*{ڳ�s�'�G{i�e]v�ŵvxzM��.�h�h���T0��UI���keʯ�����4F@J���4�Zuj��a.\.�k+�4�D����h��Ka=��'Gp��X�|(U�`�m�M���UL���+(���"�pS8]��#7Fk��n��K�A8�jP^����uԼ�)!M^���*�sEW�
���T<C��eg�y)d�������қ�Sl :����*�y_�;�Un�>si�bncX1M��J�en8�E��ǽ&IC��l�&� �̞y�6�%,]1��?�/l��z�}�����tR�Կ�vuT�f7T��;2���!��%��r�nb��[����x�U�)8�/嘎@�+��0C}��QEl���e�c�q�+����[Gn����SsX�p�$�����Ks�ﮨ#�]�.C�w-�,�����#�cByN� b�c�@��N���P/kE��r�RM��o�<�`��q&�d��Ƈ)�)�X���c�_�o�n�v��*�<���[�\c�f�#��K�H�yȆ&%��bW�)�,_\Z�]��������l+Tk ,g�-͙���m9�[�{Dϓl��`/M1(�Q���>^���21���(��]�WԸ������(��+�H�`'�)�����tb�r���&$�
,�d�����6��5PVW�����N�O�.ҽ.���N$����m��Ap��|gk�z�+羭���Ku�>�i)L�N3��� i�,��/N}p��r'��oL�����BJ�q2k�yF��H"�m�J���l�8t|=&�YyW���/���j&�F#��²+K��6Us�����5{�����ɦ��#�U,���s7t��J�(Ȇ{�D����xd���H��w��)��
��]�1�FD���A'"���g;@��O�}�H/�9�LLx��i�C����������:4#n2�];���Di]l} O��3#��^��!����غ]�r��-R�<�!��3H�����-���2�d]Mz��0*��XSS�OZo�k�e{�b���X+�µfh��Ü3v�s���-�+,������|�[�A\c? V�_�ۓ=�tLN���D�A�����g:E�3$�����}� e3�J�ȶ�7`<]��?�6�a%�ܟFc��A�#KM������*pT�x��T)��7��u��l3#��Y!Yq�׵�bO=O��.1ރh���?6-f����a����)M��I<���hE/�v��) mU����HŁ��Fo��5KrSM2�N�,�i��N�;m^��N2'�C��̍-Q8�`��'~�DY�B���Ұ��)���� mG����(�An�E���� r_@���X���'�l�p�^���q�%N��D���U��L��gp�11����V�EJoX,9Yŵ��m'7�#26�bm��_�j���q���u|嫿��#ca�C�?D,_t֍� �*5�К��H�.)�O����qP��og����bXח^�M����tŘ���9=���c)���_;�՟�;l���O�ڎ�v����Gi��ē�g��XNf�p�̽1��ac�`�	���D�C��u���*��껲�yb^AϠP�ךޡ��ak�L��|[�s�?��|��� ���*����{�x����Z���#�+4pb��'e�t`��f��?��b�����VΕ���L��W��V;Gz�E'�><�ԪQi�|t3��Fb�4ঋb�t��6F����<�@��0ZeX�?�t�?���]���%�:��mg�*�t���Q0n��������B�KۖfpZ����Q�{Ue�%�������Xִ�6n� �x�S�b?V�(�s�I�=�0�|�͠�ʐru=*�x�L����N�\_J�H,	�����ds����Y|5z`^Ph�mM��|R�v����|�ѰL���%�f��I)٘`���ϊa)u(��E|G�:�5�o�
M��%�ʾ��&�Dp!�)��e�-�&=�o���R8���x����ϔ�>�n��5km}�^FJ"W:�,b(P;��7��}H66���v�`�0��3a�x Q���C���V�����"�"q��3�p��8���[�_nE�NO��� ����t����^��$h�e�e��Tz��DI�2̋Hzw�`���r�I�_փ�4J䔳��#6^��}�E�1���5��(ZIq�5n�2~�ٌ$��T�e�G<��'���:�̪Ԏr�VV�В�����Ne'���S�7���j&R��6����ͥ%����s�IBL��d{��K,Ym��NV�0� }�m��B���6�)KEF43)��UZ���n�"El�<�+c���U�yN�Fh�s���K��'�gI�aM"��P�&�~��6B�T7\N*�0z�]��7����՜[��+D��bV-�L�'J/.�W�N�X0b�|5�+�M��Pl��*t�\��nQZ��.�I�n��3;�HIk����������$�"l��ľE͍}Z��hc�،��w��o���fi�U����	1 ��FX��-]=�C�`�?�L�`2�w]IP���W�>�;{�, �ؤ�{r؅�4
�`�<p�n��C@�ZM ��V�A�� M�ļ���ǲ��)�*�F��v�;�D�Y����ߨţ�K���?  ��j��2A�n��i����%0JWا�9��y�v��������9d_ɤ��b]������g� ��������47�[h4����1�`�w�-��Qjn�1��ĳ��q����|�σ�c�P�vh�H7��Ӱ3�7�ee��_Ԭ�y�'Y��G� �d������4�&�79�s�!R���g�n�W\4��������W^�q.!���p�-mN�B�1�u�H��F�D<�}$(4!>~�����	 ����F����B����ko=E�'���<���a��s1o��RR���˙uK׭�/���1G����K>��dބ���B�ex-�<�$Zy��T�n_��ٱ�����V�=�V��{�哘,����*3K�qE��T��7������Fp�*��9������t�ݬ!E8tgC������?���5>W��{�\��ٝ��EVH6~N��eЪ1$ w�T�H�h�Y�y�`7NϏ�\�:<l�}m	+n�X���G7�0#�r��a@�<M��$��7�gK�u��ބjN���_����r�e�h]���Lm��$�7S�<#�O�N��Jp�	�UG�q�_/��3~����8}����,�(a[�P�3X2}U�Ѣu�H�YR7-Xƾ��'�}eV��oln�ʍV��.Ւ�s�1����8��A��3�W
��W3��m���9>M��'�ѝ��Xz��X����\4���W4�L�I6z�E�YI��n�hl��&�˗�t�Q�uW�ޜ$蚷�8�w¹v�,���-N*@�:y� X��`H����_�l;+��	]忋V��Q��S��+M�����p�6O$�;�=��ҍ�]����)�Œ�k?��F|��	�4��@��T[Jyr��o�0�l��>0KP��%g���P:#L���,5��<@�;ߟlx�."܃Iل��#���4ۮ@s��.ﯳY@���*��!BT�GI;K.�99��뎝�����xt��X���8�Q��ã���1� �j{	M Fr���E�����t�?�������K�嬚�P%��N0;|�?�j�:M�"<1���9Z�Åu��5���W�ɧ\�	����/g1J��Q[O�x�˷�\��a#�����ޔ�=�/�x�c#���G�����Y
"��/�|��ۏm��|��r��^��]��Q�k�����E��٧1*�+C�4��N eK�˞���o~�D�?�0E�m'�d�����xK\[
gݐ���W���M��O�ӄ����A��ޣn��M��
�˪�߁mJ��������!��;͖�r`�.%���kc/���k�Rk�F�Lk���� ��L*T�ط�)!e7���B�֟��3Ɓ��2�~�3/����`�d�Ay$Q\�}P�#F��#6�������.����"�]_���{'�h1�r��4��O���"X:��3��KuI㉕�0��5;�����3�LԢ��FL�l�����F�Ċ~�����Ot�5�l)}��������D60�n����1B]��z�i�I~�B����f�%�I��(ڏC�Du7���� �s���F�S���aS�^�m��G�
���5�R���CE�F�3�-��t�O�x_hU惔Xb�j'�����8�D�0�J�31�R�v���A�ݭ2y��v\��S��/.1}� Ke����>�1�$���k�6�}�!��Ͷ�6���TQ)��/�Ѣ�L���aҷ�:Eگ�4��3�H��s�YN9�}i
)�# `��bH��O��&UHTol�}:� F=w�9RZ������~P���G�>:����L��3j�w�fF0���#Xb�x�j�n��j�5GS��n��Ń�8��e�E�����Nd��s�i��h�W��7�dJw���y8�DP���9l[�l!#����/�g-���!����{�iڙ�� � (���b��:^�/��AH�D�^2�À_*PfsT{��!�[36�`�N���͠)^�D4���7:�e4�7� VVaN��\S�}�ܒk���(ˠ����F���^f�g8Z���9����5�02f�")Ӝ�nd�<�}�	D~�%�sKh���Vt����m�#ν�_�J�G�\�}����S��8<(��cDoFe2���Zl�؈ ��:���pt��4�îzӔ�@��R#���SM?
�Xy��%A.j�R7T3�J�����eA�Ħ�e66F2dƾ��s��u�$t�ʥr�ѵe�D��)u����ȋP#�Q��:�������3�:܇C��@I~��,�B�� w�C���D�v���������"+�f�'�n��ŝ�W�{AJ2g.7���H��c�ث?)sNVz:t%�<�gcc`���fU�?��(�(|r�C-%݂� ���RK_��m����bwGAf�xʍ+��q�2��6�/8��i�l�\dAS�	4���燫<�q�c��]�����sp��\}�Z�vb��c��T��L�?a���@ �2(CO)6k��$j�֕'ry�E�$A�6�����Ht{'6�A���Q���z�B�z�����������
��d��j[����M_.ji�c�d
�7̎o>�9�I���\�>"��y,f$D���'^�H��fфT&�$���7<揤{�c�:�'�1����vcS��a�V�c`{�q>2�	<3��8I+nO�`��vr �	����N�UX�AL��;���/�����>��$����n�#\�}���B������5�^�8����/ t�A]`������EAt窕�mH���TQ]����U����9{ƀM����+���OD\U����֛�p���'S4�k��Y�op=�|�4�!�Q��҇��}Rz�K���Րƴ��6��]a�-��..�lS��H�T���w�tX�DJ*#��i��4�	Ϩ$�s���p{ �t�@e����^�Z�R���<��7�+4�
����_Ŭ��G�gx�4�oD�J&�ӉYdKj �[�d��F�(�u7�����7Yk!�]���Q�;��i�v�C���(K[���a8�afɯ�b����q����$�����Q�n�9��v��7T�0̚��56�+�}h��Tn;�j��wIܧ�J�~��MO��Fl� ��!'џXʛ~5���	�
Og߉�)Dt"�t��vǅi�7�S'�}x��L���&�f����R��� ���J�Ή|�M
�N���hQ@���k{��<�]ؑb��u5I����p$@���9���O�!G̉<ʁ�\D-�Ɋ� ���u����I�06�ݹ����]dW,�ӡY!�,ndv�M@fV�j���6(�|k��J�����+se�f}h���T$�J��]�}ψ.gH�Mu�@��P�9��[r���1	%�cmk�+b���	�8��d[�L;UU�6یG$���`:�s	ˏ��5��`��PWN!��t�� ���ԛ`)=�0�@�����<Vz�����M��	!!��� Ҷ�dN��,��Գ5F@1l�����`���������n^����X<y}j�I�y܃�)0��xu�#��#>m]ጥ
=�����:i�:qm��J�]0/�����Y��.[/�jײ�H��=�Sy�`�N (z31���6�y�9���S�$>��sg0���[���f����w�}�i0P�[�h�"�F�������8�8��\ɧe\(�%�	����NQ��߈���o
�s)����v�礬Q)ė�x��s���o��*�[�HZT�k�:@�Z=����m=3�t?�H�L�ׇXC�g���3�"$���<L�F��@��#�{_��o��r�Pm۶�-����O��ǲӐeq���8��uMU6��y�fV(6Ճ��pC�6�n��u�q��D��cU-s���N�Ӽm�2���������P�jm
�-�F�]N�*�m `5�+����[����0��P�d���\^���z�~!1��{�94ED�˦����K��]��G>�%��8ɋRX��	�I��{j̓�b{��M H�KȰ6�p~�w��a[�š)>��O�����9��x��b}6��>hzF�<VA����붞�3"��g	S9~��o��s�H�����T������Iz��
sG�mV���2����x�H�j���C('(f-d���5�v:�e�C���0~-�[y���bOo�����s��*����1K4�y3(F���}���h-�d����"f�b1��d�m�d����_Q؉ 3�r��U�0���**o���^��#��]F� Č+kWؐ��G@6�:�sўd�x>�,cd�ظ�ż�4x�l���[��Ґ���:�J ����*�L)~M�ň-ZN�$����5���A��RHI�	������'��:�Avf��X���P��;0�����Q�1����ډ��mb����\�F0�Ϡ�u��d 
�!Z0dg?s�.����x��ֽ�!r�sj]a����v�W��H1e��p�zo����A�p�>߯@���mypB�����G�WQE��h�,�F��%3����y�9�u����FcNul�lHx��Jf���%��Q1Gx���j��fޣ2q)��������t�d��>l�V4��*{�x��Y�.a�DF(�@��
;�%0u��hj�w���yۦq�*�f>�g2r��P��Vf��E3[�Q^V�k��	���:Un�]����t�bQ����g`�`x�^��d�;��K�֞����qoS�<�6��L<T���s_�m��%�M娔g�~՟�BOC���z����iʸ(���J�W��C=Q��V^/�J����k��K���fv������r/�!�;=C.���RB�r�K�d"x��B�D�|}�Ӌ�3���#9��J�ňZ65�-�yR�qj�E\;��[R��b�O���0f�n���[��׬G7�i$-)&�"�=_�u�b�#&.����:,��ڡ�[�*��:�2��`<�	X�Asus8�v{�g�������|\��y��.�3�T��6���r4<�ӻO'܌���g�wc��@�\u��;�ѧ%�3U����ڔ�3����<��psޢ����S*m��rty9C��=ߧ�s�b�.���E��`u�8W:V!��-4��B���=)`@�� ����w�ۜ�6��rI#Ō��n!.�z�+�Y_nk4%咧!9����)����#�J�`k<
/�8���
�t^oTO4��8����M�4E��$^��ҴYO���'��=�A�Aң��i�c}�t(n�b��4�~�;BпR��L��zш��8r�R�XdL�����1m�?A2�B*���3�
�8S#rLcB�u�$��SՐ���*�ԞɺWL�&40h��o.�I��-�Y����Ao��>H�_��V7�~���v�n��Yf��!!���C$���2�}�\[�+�CKD-�,��rC�S3���(� k�46�n��P�i1�t)S��F�J��.��$�qn���b�!�+�g|��*û�c�	���.�į��72>�`�������Tg��	=-��K�F7Q��X�r��E�-��&EB��/"�&�C�5��4��{'���?^��-��'��9L�~0��Tɔ���r�Tn~��s��Ɨ'��u�AB�s0/��u�O)Z��N#�v!�)�/��t4x_#�x��<I�8@x��ɻ�+ �xrٖfQw�7ێ0p�����_�J&��x�Uߌ��9�L�|��X���
]�O#�3����x��,/,ו���g��DJ5؆�h]͓_�\�1Y����3{뒋�]a��j�=@��>S��6�?Y)��ʰd2�*�,�ƥ�	=d4�/�����1���W�U��P��RV�v��;����(�$A{�L �8G���4ֿU���ZT���Ci���|i��w��V�Os�>C���?f�Ķ�|��)�J����{����cK�D�S�S��w���~�s��ɦ-m��p�/�c�L�ˈl&���;2��Y��zȷU�����I��V��S��ߘ�ݻ���c�ő���#���Ǟ�`6'��-��9�E��^l�j'H��@�r�5*θWN�D���Li�E��7��IoL��������Gxrp�81�J*�/Ý~ [����gk�F�+J�)��°�
�v������a	��t�������[ka^�@k����Rȉ���]��D K:���h%tK�7=]�w�2S���Bye(<��B������� ��*tO̚#��g�����E���d ������b\�E��Pz^��g�������umYs�Fa����,����Dv�x�n��E�%�ƙ-�j[�"r$��>7���`cZ �>ə�6L��E��)9�����(�F�qXQ�-��,c��(6�YV�Ū�v#�u��R}��`����CD�M��ɅW�)W�_�+����G�S�f��V$lD�;�A���*�2m;��9��n�o�����|i�����*���w�L��6�T��+w\u{�S�U{D�V�ۄ*9��%0-�.���W9P2.�y2�[
�y��2�*F���~�v__�;���tB��?緡�?�43ӽ�-N�Z�<�x�]wv{��Ӈ�
�
d��zӵ�k��;\权@�AcU�L�ȨIn�)�"�ٻ���������ucV�����k|s��h�����uf�>�k%��͗"�u���!1ޤ?�7:��*�l�o�,P	�*��힉�3�d�>���^Ʈ�?�L���腬%�~JޒJ�m�/��*��������ޏ~�P�k"��pH��������ד�����:u�B\B��w��~�j���;����p���� ږ\��'V�2�Np�n�'��_�K������^H�A������	��`��$��t�ե����En���I^�q��aʀju�����8��755ē�\
N�X\v2�E���|��@�Wq�X��bŚuJE������ye�$������d��Z�~�2^y��ktf���45iO�=�'����ᓱ�W�|�XV¾N�����.�m*Na\4b����و��L@C��f&��(L�P
���㷏��K���*���SzS �o'hk>讱��7���	�zEzQ�}�(��Iw���*��Ld2(�.*i�,��ܠ;�]|T����NQWf8��gA@:����۶-`6��z� 2����WZJ��p��➱%;s"�%�,�?��kY<�S��vU1Xx�A� �@m@q���ѓ���^L:�kn��%4����)���Gj8w�Q5����a��&�ڰyj\�X93���L��N�lH�_Q�g�}�Ҝ��4�CD�����Q<�yAzݤYC,b��cR;d�;k�Y��˷�r����o�me"Aՠz�	]9�/W\d����f5E�}���Ek��D y4��(����%�CJ��G�ՙ'�ln./�;�㙔lՃ{_o���ܖ��԰��Z��]�y�z���t���ط�+�������^���qrϸ��N5I����>�߶i�j��O�K3����^�������.�Q�i���h�2'XAc��߈X�I�8J�2@�k���"��{L���g���m��;����]����Q�!���4�T�:,�x9f4GtM�^�2��r� ��i_x����je��c��Q���&ٷ*��k�Z�'�D�(�I�ﺮ���G�G��gS��� ���>5�ؑ9�o���ڽ���E�¨�؛/S_w*g����S����{����]�\/E��d�ҧ���p��F�uR�ջK�K<�=�� ���Ǿ�:XRb�,�����r��
��>5u�������&L���GM��?��"�ME��Yu?���e-�&��n���cn`>w˰<䩡���(�ߝ�α��9�6��X�[��C�W֒��L���ryO^���-�� L���/�s�ꩍ:��E=j�?t.�|���-|�
���9�7�|ʳ��Ezm%��7�g�]��S��������vF�Qg#+�'���lo�+44i�}��C{Z.��ڡM��r{;3?���Gn%�+��`���ڢR�o>�lFH�}^����`a�t�)�2�2�qCT1/����<�	#=�~N����6:�i	��j?�����'x��&7�Űy�&��H�P?�\Q��Y�&"3={�]�ڴc�RL&"L�����z3���������.���`���D5G�U<��NM�뇙ΟU� ��S�Te�68�Qx��{��fD�xˇ[��WY(*��R��N�P����Dt���^͵��~�
L��Q�$��n���`F�w�����4Dy� �!_�7a;<�K<�\����^�.m��o���j~�7�.��D�F��\(4�j��@��lx��?|v�d�W'7z	y�_V%�-���>�,z�(���}�,��k��\|R*��pa��>��^��ƶ��'B�@!>����$����2Vإ�7ꤴ�����I�	?����mc��.O�����#$�=�;���������N(n+׻ ų��oʘ1&�A�`�RېU�:���{�l_E���3$�U�K�%W 2=�V��ڟ�4(M�>e�@º߲��d�s�zѴʻ����\�W�Ɗ�����{5�m�+�-���@��b�C�j�z�L�����!&g�U�@WD\�ǫ��dw�C.u��x  �V�U��}I�J�CG��a���{9��{��+tE �4�?������v�x�+S ���W�B!H������3N-�J�۸ēR��f;�N]�E�Ŀ��/pk�o=1�s���e�t���L�7�U�M��b�����7��,��+���i;�|��0Y�y�a7D�q>W�c��oU���K WI����0Kn@m�u�l6s�@������s��]�PR�4_Q�5�V�Le�6��'��Z,No�d}1�NĽ�d����'�!���\c��<[�����I�C�W}��L~i�K�vf�[�-$�����;�+��3���`�i���͹_�	�U�2�Mb����fσu$#su�C��N�I���ە�h��sk͡x�������!ǣ[�1M>�Q�|}��`�K� v7P�N��%厜%�d��E�(0�aǏ�ӟ�*->;�x�ň~�^�׍��tf���J�1Ѷu73��M8�3�=Հ��Э_&��*&5����*�@�mW� ���Ef�d����'S��k����XM����'tL�a��f�����F�lv?R.�����S+i��P�:��Y]�[��Q��
3�~��?�DZ�����ǝ�i��^\]K6�q걍���$>w�\�H��8/�-�n|f߲قY��	���r7��ʋdXX �dO�N'+�$���L���X2��*�~�2��.B�r���
�J���?�$E"��n�$��&dʪ K�ixu�n� A�<�?Tt��K'�b�V����QM3����^/w�{v����s�?D�Go����K��%�[I�#m)��R4)Y��Q�,���Tf�C�ލ ����A.��-��
�]��eAX�-�Wr@�"��A�g�����D�c�� ��U�Q�k��`z[�yšr�[�j����*�NvS8u�!�~`E��C���\�	1_�L���$s~�8V�-�"��bS-�|p3�-y]5�b�]�l�(m�X��E6H4�j-}�D�k�5q�`�H��U��7��v��%�LQ5��3~p�j��.�8�A�]Bޠ.��R���_>k��W��#9c��m�E�0v9#%������ ��d�%��9K���<��
�ݺ��>�싟��f��w��!p��~�g�ڣ�8��yR�܊����a�7a�ᕳ�����Bi��c��'XMmP�4��,_�$�"��D���X�f}�����o�j��\Z��x�sAq�jή�؟6�Eo-���{�[~��C�z�E��<�tLNr�.����7�M�!I�t�Ԗ��x�5%2���`њ�\��|�3Q޳ cՅ��D��@�+b�C������ݎN%�2�*b�u������>����c ����R��:��Jn��w���}?M$�q�UOL��垇w̄�(5�#1&ϖ��8d�?I�Å�t������~��!>�!� ��J��2����>��dj�F�����ɬξ�	���F|�[��%ǥ�]�*�/�=��t#����g��%(L�$(�ے�w���2�;a�_F��cǑ�;�x�a��[\���ó��؎	ۇ�d�JO\��Gq�[��E���Y�x���C�Iw����[��l��H��|A~j�;��$�g(ڟ��O�Ӄϲ�S2��TP�&��L?������j ೯����S'�o0��><�C#�i;�V4˨�e+�&fp��Ę�4j�G1���*,k�q�*Gk��uV��I��	����P�>x�*B���;���:hF�K	N���'��Fp_P��m�6܇�ȏ5Y��Q�����B�ʰ����3��WZ������K%��S��f;V�L�Ʉ�} �������r�,Rl��G�=5�%)l�~��TѠ!�K�,��!;D�}��\0|k��j7����$L'
���X��d�<��+xSo��Z�m�1�yĸ���t� ���Lj�r7� ��l�7�����e�;�����Ś+f1�d�7K`� �E�EF>p��eB Ꚍ��>V��~x�3L{����܂�����Q���1�l�54�>�Vy�g��isp_��G�SJ�J�0��۹-�$n��dprѣ�1�4�v�������h�^c�V�aB�/H:!4��s�Q��Y�?��Y]=B�脂��I���,(�%|�L��98C��mu��t�n�Yxw�7�>�dnCUd�%�F�4���K�4x��[%x���x���mTz=� ��L5x�� ~��9��݊s���@z,6L`-�D,��A���pe�1�����Yfc�zw��[e�̨�����c��~�R2;�0u����-��s���v#�g(�G��B�{����)�fU�}��ϑ���5Q�6�M2D|W�.�V�V�!*7�e�29��W�Ӿ���/�2\��� gK��4̳]��t@�(/]�&��/�*�0@�S=�\O�Ʉ-RzD ����2Κ�YD���R���_2w�r;;�j�j&�wΚ�O�R��k؎ǃ�I&7���7���Tk=�gM����S�}