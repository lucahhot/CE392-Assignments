// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
tnQIaRm/rPTZDB8bOtmXa5o9p0AVNbuXCGDPTaEWRopkCJhHbDudGFpfIpqrMEsl
ERnwFq1Zvw1Vt8rC0GisedieRJy1n5N+p2Qc1COkYe2uHN7+++mLAQWnkq/sKOuE
GKdtvfy3wwM9Ix6ckArCbmcdJuSh/wFCLRH6pYPtFz+REWfAIuU4oQ==
//pragma protect end_key_block
//pragma protect digest_block
70M0FBVh4M9Z0+E8rBD04N1+HQ0=
//pragma protect end_digest_block
//pragma protect data_block
5fzq+7fU6o82Pj/VkTwhmoIy7Lk4oHUq57pyalXe5ThaUXKhOCXAHGvWPHlG4Nlq
rNLaK28/zrCkUAMEPfmpqHZfDAjDW6IS0Qms9WH13YaBUx/+1Fj7JwzCXtsqQwiC
q+swNF4rMufJFzc6Nf+ZvBjjXIM0FYEMwdtPyGWGPNQq9AG4MgCY6X4AqUM+4KjA
dkOhgCCcr59Wd0vKtx4tZtycsbC7DoWZpDfE3uoaakknRoeYmUp9twRQWAQx5XKF
bLRRC+aP7T3TGpt+Pt4qHH2qukNE77+0vh8oNgiSkBUZbBo749QwbtWJfqRHoVV5
OexoopON50/RUFxxDJ8arycUDTUoTOdDzf4uLr7k+34NdXpKoDTjEDK8IVBbijrh
2Nare5m1xw0P7FGY+Nkn7VyPhk12haRL1MnzIiwMaFM7KQ4UOt3UJ0T95LRRRbHu
vrrnAoPIVdbXmqewbuMGSzO2CS+rHK/mWEx1MAPk5oCBaUUyM1OkPU89mepOt0dy
JPR8Qp/uLETiYah+AmO9eV5ckabOZXIZvw7un5J7sI4ACtc4ZXmfrVoPXrtApsum
YA2VM7THwuXYaZLDH4E6CIOUbsEa2uI24VOCaAqcbfNYUs71tcbzWP3KYJbeORaC
7SgXVc7pCMtfKUNj8vpfJ8SbYLUT5tUgDcLW5TRbUxXhDHvXkOPbb28GTgXxoANc
vrS5RQtZtLsvnp7deVdia9GV6nRb20GJz8Y/GFB1hhQQIku46KJu4ca4YePYBnM4
uiQ+ADw/ni50o9kO52HnbLFN3WKCzY7Z6gCgDrtfxM53B+/Sww+R6DrPiGVYA0Zs
8ti5ibRBuRHM4SgUc+cMVYcq38GlRNLvL1VIFMphDrdq4XIensMoQal95HHqyfKL
G/57CRuSM1/hAYbHI67xGcZYNt6DrCJFhU1ZnIDbhkry6rcNrM78tPY3076r8cmf
qZNRXyAuD1H0M98ehMMYfXfCqdI7mFvvbx8I9B/4slXD7Om3IPtXtN2hwoupWsga
JzJp//XU+RblFBmSdGfoH+jEjT6BKbq2Uza/oH0goDpXJ9kpkOrORe6h96kJSxt0
Cv/EIr/wxccYRrIWg77Q2L678s9B0RJM9rIXwn4AJ4jmdyk9esmaceXm6c29iDiQ
fU4QhCOsDuFjo6c2XlqwUz6Yjjwmspw/b1ZG1PdnBcBDGtixAj2qnlRT5OYgHtkh
JXWccAOeIvfFeeb0l0xQMTa+1TIIxhPNK4ImjNZsb2zMPzj1OiKdgWyFzzzhTKOo
nCV2dXz/+rVfgmWgAJeQ1UBrdaRN3xs9mf4QRbuX+VkhpROFHuShMbVrCAH2odAU
7GIjHHUobqxZbPao6/yVdqO+PyVAk+iXne9VbZbe82MkAXSRfs4jz6pmVNdBffCZ
KwnWpnz1rZPmKTaWz31jQ4DbL+yNj0S9hAWCmaAhJzBMLw3keJqEGvN1nvBxXk4Q
shfxFjsN0lIgOn2HVwq7PhU7GVoZ7BEfml67IyOZJOiLRPI5XIXKiEzRpYBIfyYa
ZPSgZRoBEz8Fy3fKCgMIu8F31OdqmHm8pTNYkRVdn4uj0tTX7uBAWQPlVlSvz4hX
RGwV/0oM76JyyrAiiCF2U9CI/0bMP7A7w75dpKBRAaYMvAM2LxJ/wbc8VaicObkS
/OlY5ihukiTiCG4Uwpk03/7gXeQfPEGsEZKzQ7Bw7dVHnwuDTpJQkuDJ5WfQ+Nn/
zlpUNvgzI8cI5W8TxBiEIPYhKX2nqoTgblk9hswILk+6DmCDm4sZeyL/hsRLwwRi
RNFyby/ZHkyrj6s1yH/tBMyNVnvY3c+6kjyaD6dO503cOUGRMTJKBjPb7OEhhHGJ
4/tBu3bMLEXIIWsXNNjizVPdEsfNB2vBQlsbZfBKerCCfe/a5JMZtpszTtmP7KIO
jEE0ibkCsOQw1uuI4J0lj6j8y7O1YAbTWPAgbcBeOTYWco4GZnHWHMgnxGUmSrqP
xSEqMC/ug31N1gdRXBPRrtzrTxjlErsabIgZEc6r7j0yp9TX+ATdoFZJJ9OwAobF
u3QTy4HHPxM7akTsRDIuewm7IZce+EK1ufheTuYUuGhbnrJVJOXgg83BBav+exei
c77pkYSS9+DO3DPvDj89uFfzcFq9G7+JMdndutWLMPmDNLFMdE7OMVenptaEU8XM
pinY6w1W0EIUAtl4Tsz83t8XjO6id7mFdc8kpoJkhztReSDjOe4Hq7WoqhxVvRoX
RyKYFtIOvL9t2sZBv1jWpFitBZwCIdPc3lSKriHcWN9edbD/OMqe65J+bOW+WLDL
IWNG2HDYC2IwajbD6pssZAHV3qNiXgwdr3TyL+Xv1iowY2iMHGsZjskT6jsrxX5G
iuucjJDTQ57aVz7v1oEvuaCLt1Yn0kF4ZepwGcu+dtT1VlZYPZKI5VLqkUzeeOoz
aCT6bIG1qs4M/W+gg3uaki8BggLXaPrhX0PyqRUcuzWO5sKlh7iFqNwl8fbNSZ6l
auX8KZTUXK/VxbCA/vS3wdIwn8M4oKoTeWzNEM9Kz7Vl0s5HW3RlljEoL1ZGNlPJ
W3Q8wGB4nB5PLMYkK5JDFyQP6rK/L9l15g/LIlZNEb8lnZ+RanNr20sq0EyDHtnE
dj9/XKaADqTTnvimxVHtizr3qHKpj06JvgC0bUA/g1zJI4z+0qJvwC47a+x5yBaR
+/p7xGMYO14Dmx0t/qkmC61daWbQbcMgNXVX7M02AA892vT/5pmguJi2Ao4zfsVb
J1+PfBSmtLBlRkSSeYgB/kXFAFe929v4ZmO0HdxNEHN1sUaUTUrx23FTsMrJJUUF
2rh1tbu2jObhikSojRddQ/XVu0UOnPig9CwClTpEIQu0WhLyDs3HEL17b3GBmKdE
WafIGh/Qo7o+DgQ+BkoOlBeRxjS2BbQU41MRLp/gi76uqukEJtWqytOqHatMrm70
hjGWWqk1nTuWrUeVZy9f/6BSx3DEJ57sy/s0pubQpGA3cnc900fw/jtTrd4lZ115
DqYJPpSOu3sEC8HYGVmajtMu6shbi/TTPhkuoZbXpcZ9uun5m3U9YyH9GQWI9yhf
ylGKoTPVyDWwQ3+z//TGni33l4G76GvalAT/0nz/nOAwBhe9sKgD9xjcNiqVSEJc
uOFhUqN99Due2doJqqQpJPEriBOEG187DOH+AYwxyQNcSIfN3Z4gTqVDJw/L4tuG
omDVjGshqGywax43SIQ5g+x4S73Da+7zubiL3aZGrDtmSPCd67agp38R2o91B6Ic
CgQUHgShFX701QIlPdqR3zJaP5daLIU8Y5xxrEk+pAQXBP6q4U//lONXXbt9SGaN
Fth/ExFmuFNG9+t0zPqM2YFALoH5JYpNZOBh15rkz3l9WF8TP0SDvVM4oOGJBapQ
mfdzawg5dh3fLLM7ARifcCqPVjkBaWfp6SYdMTTd3p9wsMjZ3LubBQbJeVuy44hz
WDmPBDTJcYU4rKliJNuB4j1vjXphlroILIy4rsbKoVEIJ8ER5NauHZM+GBxfj2XM
Jei1f727+hNMv6wlNiEFNIgJTRxQG5EaoPQTeRuJGLeGDrKJqWHs3uTLCRxQ5HyF
baeVaXXU1qQGa6OwLegqSwYcBU95NLaLvSLk1Oldl/69Y3G0zOep5yUFHfH2Crv4
dAsEig4+MDw+VvISehRIuoe4ibsQL7uoE9+xxNKaAr8HJ2cJyBfn2jzu1tx3OPr6
edZ5EuUHyblS3VmFmsW/x6CZPd+Q7DpU+jqldQtxrHA1YgoO/YgUA1lpj8sA/+C7
Pnsxd2VLcMxSxR68ja9/WOoc9u8CihIFVDUI1LyClcfDVSzc7TW6krFWwz3TPto7
PBuS8nokj07Nx7QtXeqjsVBVwTLFvn2kiynLmAH6x0Rp5UHkNlpANjXdImzcrYRb
FEpIg4PSrm5iFJgrF3ffiNZUA2TWEqJjowjRUjdHxY+3YWUv1g1FDIJ728v/ef1O
m4l0F+B5pAnvlwyJFFyUG0BqYTfv5aCzBS4w3syDu4YQ3n1Fhf8xpFep8C4z6Hwv
WGfJBrTGR2z8k13WjxZDvz6BjYNdbYRJgB5b8CXUcX0aR4eUixvabDkjgbl2P8cH
lKuflIzZhFrdhgkdQIkVb3aEFPHJfNGqXvVBueNIKzJFPTl5I96hunej41xDe1MA
DQGGu9PcFbP8TK4sqUEZp4ArSRzFgsKE4Y3TH2u22H+yMHeahYaeWYSF2+ECgQvY
KgvhHDcAWO5nMzNfYX0ZP4NkW8jFZB40qbBT8KIwY5m8aA8LkNT9W+OFbu1z79F5
sc6KHqDaFnBN8rZv0ScDNbV+f/KsrQvWWjZk3ARBCzwL6anc4poIWXHzTGlaHgeH
lS59/yDrsN27Ep/hh1tOuE3jPb+6ojjC2whYl7rlkzP8OX1DJfGjCDdzpSvyk7K6
J6+s48p/u9t19vsLDa6jY7GzPugG5PItrk0u+uckv3chGsc2zia/teUCh0KvcF1x
0mKi+DBZlc+tPfdj/BlM7CbptZavRwBqxKKZXWrul3MSVJJfEIebHIe4ZdrSqquO
wx9W1GP5VfhMjTmrYfxM9V+/tnl4yfOa4mWb7CaB04FpbykELDj3I9btfJhVzohT
ytJQugBMQwy+FToKhw2SqaqkmH9aZU0BFUjbLmCL80wFLutZGVLSwvOLTizg1X18
ANkhlv7YSObxbctsD90q+ZhLEFsGtiSej7veQp8ZNBGi4G1ATOlbuFzjFFdGue+c
9+ZhzDVFVC/htrvQpW6Uw/2GYr5qSAGLNjxQe2badswIM+OjkuiTpujwfoZDn0Gk
k/jHC3UwmnD9K95hHBhrq7fr6HWuOs30wLW1nrRmRIGzQM/Q9+V9pJOTyjruB3Oh
qozQIlh2ltm2MYHTmBbuUhmXTX5nAECR2U9FG3EKx/+SLKBVaKaX8vePnNfClvXI
younWAL5bRbgfIzHNYus1lZozTBdzwE0u88rR2hmW5bx/cxTjQch9saDszuoqd7Z
g5bXfndEZ8P/q2hgW7R4C9PZE0YwOzoh8s8QIS9NLwOLyq7sO9hDdnldviAioffV
p8yBtTAKgEsVrRArJYRgAtdqtLYgplKh97OTFut+7YE96UYlqYOibPpjlQohohj1
9J+XQEitS/jnXL7cqU+Khn19jYmdtPDsB1swBlZQu5DxZ4X27QfXFlO8IpzCLVn6
Hg35NaUaTysUXWuWg7jDY/76uYCJH+V+saDg7yiTHvAU4FdL1EzBBwChUR0bhK1I
D77oiAD5GBJHhbsw//zrdWhNFY/g6aTxdY0FUK2eBRdJLWUDdgStnkl6k8ZNtWwg
IRqoCeb1wgK/8MCOd/6EFO2Ey4UH0p06u+l3+gQJV2QuV4zxpf3bgOZpDaGRZ5Z3
VOPg/divKsASy/YQNnen+/1GA9oPfvIcPkFS9G4/b/VVD2ma0Rm+XCSeBu3RJ0Bx
/yZTfcMDIP2FXHEKE41jzOC59hqIURMBKVUqvWF/Vo4ucdwBZcUo08mw8/Q231Z3
8uM+TWf/woAmSS0JH+jt2xlvi9MNFU7UD9nfewc33F/S2hkiMy8UW4Jozt488yp5
PoC3RJYprtU5Nj0MFGsyyRCRqIx0/LdXClG/swmxmZjwsOJL8aOLBnFfaX5flRp4
sXWHX/5hbGBjfTEIkss2owMTA1WkMrn1NYOAGbDGpg4QW2vMJK7GkBvkEQT6RX8A
RxPchJVqUyrBJeqNkavPPTVlYVxiquoDbvpxKvIsxLpk/8xVBiqENArRQPNWmmvE
kZn0QevJE9YvPq6bPIQd+gxkG+xNmU0T16v4AsB6VDHbq0aypI1nkCPWkg9l7Kgn
3AFXJyAxXbMXSCLl0uHhw2msCc2C6luuH+GV+0By9zGaBNbnXxRZs1j8G015nvMC
aKLtl5uF7cXmQPewDAOvdJGgQOauQhjcgU7SSxQq1tsIGgY8uUEMYh3GisFIVjAf
2Aein3xtOPoqXifF/PqikN7hisvK4w9irvnYZf1HnF7vjEwEAgYlSJg9DGKjCYvI
ofYJvzWMjfAE2ELV+0npOlHG+VlUPn65qfvJiU2qp3nHxvJF7JfzUAyExvV+hVHd
vxT3cdt2885y/yulVhaCr7ZJF1s433C7QanIttroq/V/bmL2MCVG483ltegs0oUR
xjdpAWI9mOUJYBA5cZPffsXQoRiKDgK/H32ExJgR/bM12kbxR8vjCOhAm5QUB7Aq
cG/2ryLCWBfgGx2y/scQnqdA6NUCkvaUr0M70U8s9gaLMQTe31VpNGKi4+nabIhD
MO4FNu53UZqZsAH6CRFxj5v5BQ1twfw5YFXo0I0N0Wbfv46RqwWo08VCASsfCV0t
R6bJcBte4elCvRnzmaa7ntNi2pBPZAkiZ4v4fkvbi/Wami0kGRRnriar7vy1AB43
64Swf14VPafeiCGwhWrFM0v2j0V4TnXFnEMj/b+eoMIkoMWKvJvkDlba4GfWQtMv
jxcb/nzYC78LaqIDvxt0x0QkiZIgvP2cTHpPS5oMnhZ3/gb7sqU6WW/aUHyDyXes
w/Sm/XK2zlP3pbZn/YLUncIP5xGKrt9RCr0oPm9lcxFjjnpNiyWyRTxt+DPvHnU4
PPDUBY8MAvqxPTDJ+yqLDlCSEtOeS/NN+rZgyKAyL7L0d01GJR6vCt9XQsTNFyLS
nbuzdpQpp6uDIwrPZOU1e+UZrSwnDwbUQMOF0Ldr1rjIaxByZ39BrXL43Bu5zvHv
vsT9XQcQBH4trl3yIvftwB/TAth+2Var1b+5qOf4YlDZI8fSCIVNvG3aKj2fb8KC
JDynQP+cR43S+a3mRw6J53qrJguwAr81beoMW2dDU/fK6FC3OWYOWaj3M4MmeeX0
E2orYSr8umPuGBMF50h+dksbYtVPvUGwolVqhvXXtz8A+NlmMUb/ZGAh6ecabX5b
Pw7CbU4yK68wHq+bSBXOY65OGPlk6qzjjPNUBj6IGOc1qqx8WjrdbaiyxPbCCU30
YCYQiNU4bsiPwyYVuaV8ilF+k/Y38eV0CLdvMS0AY+ePvVCQWZkK6gLy1KV1QizQ
OyyUtmEGU8g5kWTqb8cv+wrtR4T+MxZyoglZ+7AZ4Lcj5P7/yCeBvLNcfzJqfEkA
9ajyDgrovS9Knmm1KzZ0kx3eLSVojO55P9t7FnMhF6i9pyYN/Gm4leoW1znhhPpp
hEqpuAbVydJGHejngN0WfRo0l/2O5BjQWy/iUrEiNMAWYakFXZct2Vf500XdvxQ5
Wl5Jmlwjw7M4hb2ZxFsUKoz5JnQAQcEGjqiN11DguKGHVoM3wDkdlkTij8GAMCoQ
fER5qHGCfKYYMrxrSD/HbCgVUAg7f0b+TrE/uAOjepfHmHFacP8fT2WCHWetL70w
NiWofrtMZkFvQeWMQ7tnKkbHaVBE90T2r9SV2XNkJm0R8z9VEdUeTTTl1mj9/5rb
/Lf7f3/kfuMDWpQhjHp4a9IYakO/VCbtTNrTrGchaV+w2k2Zfpya+oAn43J4Yx1l
1jqwJKZQ8RJxGv0oGtJCq/WZOLdfIpa0pcktZY6i0T+7fVYfiHkvOeHLB/oBNazX
eF4QJkv2g3oVlDoQUh3FvAko/hbN9gHV+nX7m/KUoihZ1kdFIO2C35cz2vQJpFLx
cjEN3gosx1zDZkK0i5tmpghYIwVg5ATrmlSyf6Bbw33yMwSK4362GqRbL/YOqZf/
olEdTmss1BM+X3jebXl+4DEOZSF3/j13VgR9n6vdO2bTA7rBuFZ57uCoNmUnlUp2
3ZJY9NEdBPRSTLf8V9zXaMFCvXmert0uCUF/Y5wPyt9dJHHgzZA8kwD3+G3f+Wrg
V8w05348LhX/irXUdcl+5HwfnZwrcPjvmH7ipGi92ugbHoQFXH/j9ViEuLlzMD8J
wtRBWm7GQ36rGt8AT+wYcPuIXoHzo06/MR6NB1nRC5CQAuFprkrh9YHNb6GaJBOc
WnSdUCzwpKFWV5HbfjrxfigpWu8CeT/cYN+02tjE2ywMPM+ubN4QLcsDvmwRGdjG
GWPXwrjIv5VhIL9EcD+m4utIdPlwpU+fpGgAd7v+yDYAnf3vfSbQY6swtFsvr9XH
I00ECuBHe52D97paf3jUphvGRneDlct/mzdtPi9mcCLSO42cK73/+ZozItwGbBjN
lofSs55f0ut9q+dqDB/qRtljWifG/EbGvcsiwlndqTKsJDhIv3iZymN2+JPYPPGd
wtegoT0X2wJdwIXdqwKCdFVo3Jd+nMT1X4Ub4NrwllDufozpfYzxhSEWl1RCsu98
JWykXs5idFupHH2XAlc0gOB7RLAy0p0AIdCswnr0ltjsCLZwEce/nlq+Q8eslaes
EcHCSBMTftjvVH0hDZAAiWNoRJOcDAiTuE6HnI4z99BS7ldmIcMw/zdnEb4imP4i
9/GxDn7MXNxdYiIRcIQsODUFxopustcocFa28iyeUicq98JqOTOt0EKtfZc1oFIX
+DICR7bgOjQp+FaK44r7M2bXcNx7Mz+V8dD4gFHypcnR+kbL4TIAeUv6PFH+Bq7I
4mlwWH4hTGuDgqP3Sn9bg9yU1+l5577bMilJr/MebFHSZJgkUm43v4mSkzTUVoVW
9SgMEnOtxcE7EONEgMjU0QHRvlTcWT95WwKXIoBMKngw+7CYGKQpMnIYdOC4xquH
0DcQjF0lBAILnuwK9YrcRlYwIoZx4dGVNAcPIsWa9ob/VsjBGWSHnRJV9m5S/UpH
To2uRQ/gR4i3CBLzxUCx6pcHabQK5sdKnnQCEN93tch1GGrTHoNAEKBCwjY8oOu/
cdZHyWxpMoJ6cm5ndaroibnZM97UWUiCt0JOQugwd928nSVB6oVQmGKONIIVhYSG
zc7PBl0RyNGgMDqsmRGstG0d7vcLhlF20hUQuaixe3fD9lJoOMFyyv6M0a3GOEGm
5Q8LqFOxP24kfqkIkHxMfWiyrjsZFIJLub9wT1dM0CjtTF9Q1gnJnXVKwdQx2+hm
PtJBUlhpQ0P3j+1wYxGyFwgWhwDZwagX+fyPYobZPtaeBFMzcjjFIlqAXhCQXZ6U
FtppkPjmU7s0u9WT5prsI3kKlGu7fqvJy0YDaGn7C6gXSCyUez9wvYeGwRWMZPP7
FTiyFIw/xROf9YgZ24jRPMG4o+mawrNvEhY9LW/GvuGlvWHzbAGX/Ubvkq+IMzus
5y2J1qBeA0nZiLkRHP1IgFKBru6wg2BBoIlyASd+H4FTyZOQ2dpPsjngnv3nn4H0
spo6NY+r+jAp8JYJOxSDcbNaF1B2tadzdX8Q/UOfbmb2i84hmeAL3neo0VvGnbQv
3nbQ4WTQNHat2o2FejWsDyNLEbRuJ2w8vBbafojs2nkEkmLVZwmMqER1fUy0msDk
rXw6n80rQ9wMXHnu+037sPknA5+LB9YddAmoj0KNaLxDk/lD2g/aLup/03EtxYN4
1kFx0QjnirbbGHFcg6pi5NPJcxqelihDlrqEEjnFpwLkc4vKTT8gY9EXUNEex0w3
J8j/3oA0JDCL6PbtyZG+DMFg16paEhSsAbQjuadvSczebcTZIPntEqd8uniwQ6JD
oBSZCsgDmLKz3I+l/zbbixVxJNkOLESFqgMndOxceDcnkR5waFUcOnul+gi7mxap
hMB8LeiMknV4Yj3ghXI9DGX0FQwMsnc2sho40P3l4y8Hk6w0tI76djsaKdpF523k
PScGlNtItPdPNj7E9DziTxE4zOhmXImQLYZMHfSmRdQJmhRcs8d6YPz7D+JYmzRj
N+uN3+WSNjbqn8LOt/W1zFdtDZSyIf4WsMjz5biGvwNcxiCbDNi76HwjrjQBhwxI
MjGWYw1ZUsnpQjAzupJuvYAy+eE+N6HMspCA+YI0QNujULhpXyv9HYwC/5zBeJ+a
vFwYxidZ93U1+lhQmKmQZgn3OYr+DzDdWPpWdERyG/GmJZBebk6wN5GmoJ1feFj1
7/fbSP5VaRyq604hGjx57hWNp0aVjqdugrPmdimsOtcBhNzSyLQycrJ75gF9OV5e
ZCKvX1aI2X0PXHam7OHves7uWgbFnS6n/ZXzoZRHi+qRyGxb+I+Pmr+w+RI2i61T
LAQwJMSl+2sdynzfp+YtYiRqDL1aPEgH1vFBEzIvKfBKyeMAmiwrtZC8dqD/IsM9
crBaH2Gnpxf/OGkNIaexe6aNub9D6soSuAbLQe6f30g/Amu+CO/FiW5T6QGqunQW
IrtVCafXopwX74J6SCpffZwzmkJWJsWPDEPro3lN9xld8ll3kw5pHz9GC6NTvzvy
AOS37oSsduBKu8B5ssBRZjEXBdVVDeG7ZVhhy7b5ranjxupgitdy9OXkveXDBpiT
6J4L8Z80qiiCWYxjBD+BYZaygPVZWS6qXt4XhUSOYItyA9liLjM0ItgXv7PPEtTV
sNEEfCh6NTA9D/RcG0Uwx5zcZGto3hNSyu73DBpryB7oKs7DtDxB8gZy0WwufqKy
7U34s54n6WADiknLYXtpUJeioD5BIIct+AQEigI9TejL+liI8QYm9c6tqJS0TT3b
MlZAK0Dc+IxzMD1pAACswm5uJmxmvPIuVaHN9KwmhKQkqtA2t1d8xdHvzD8ZICmx
aW5n7dEQ+YHsiNtNphfhbox3FKVAdwErM/WSqFKU/Rll5/m0wNld0Hh1ccQBGWXn
SEvvBw1G0DV0F5SDGoPo/k/JPLgYH+noxagmRqc55FDToJ9pO52M2cUGX3MTouBB
gv8UunlCDLQgeD03nywOw4Vsq1E0jW1xgbtbrDiYgIU0cHlAJXCCn0Cqm83JARQ1
nPVlSrWjgI/2PEo1fh1Oo3CCo4RMBoujLlfm0Vmf97T4OveE1HOCO7D/dt3C/0eB
k5IVXCwXysrOzk0moQw6iDOsr7KtZ8pOuDNKeUE0dxyfXUEhILI7GWoWPowRqyn+
L2YfE3lxslgTLUS8suiEmZ7ssR4pvLSzRLMip4gNAPwse+72QB2ilx1MO3ThK79z
LdMtYqPe4AHVi9eWvLA8dicyYBF5eOwHy9OD09DQYvw05DH0I/2daGVTTfrDV78i
V7UpoMxqemefffQVvrL79uB2AUGN6dKMh/I4Q9FOakjIJ4MBtt2ftGstHLYBQnjm
XOfAWaB6a/4JsXrCj2rJuy8WzzcxPceEh6TRPJVVwS4foAbW/V8stwmaFLiXs3H/
FBMLUlz08YINC08gmJYKFNSww0uwHWn4yMyICsIdMaAag21voJiY1HlEAxU7bmhj
7tQs3cxibDdu6xdKLayNZwFZ6iCsAzFpg4oubn9eAQlPgn5ub35L/Dm9O9AyiYbi
99/M4PjLimKetwDMbVbFZp1BI5brPJS0NOn4WUJGtlGyEP5Ii/r3c9Zq5zetFH0F
ONj4IOFiDZIJvqWOVUye/LhEGhyBOwawiMgW46otQ8oH99rtlGw4DRBkgl/LMVNd
8ue4z7qyXmeEBfr5zrIjBC9sdx5aSuLw6gSwPZeP/avhru1dHP1k2ToxGOCD4uGN
je33bdaxBBenUxiZ1XuZkuP0TrROulcDBW1gOcMQVwAW8p02QN5gSjH1YjdACRMl
i+SivW08L141pU/EWGGUcpfLDXHb0F0EKaxg9bIw9KjRWySXvwP9eVbuPh4Qjm2f
xChI6GSadaRDGIZpTMAfVK38zcMECsE5ozWOz5Rr2pZLk7ANeAXAClCZJ7fwHPZ7
riOH9WjOTPjkJDBKCC5nOv4gg5WHyUyJFAW8D5u7YTpG7LpeC/Bw3Ij9lLADyiG7
Bqqob2fc3mIYSjA5ch8wR9XCju5npjUFmwLMb5FMwdzH/Um8G3BGJszLd19OHZsL
2/e7X8IfKpOlmDZoGNxPUbT5dzzhouMCexLQp5sjftwl2S7ONCkLm2JSDtyI9NO7
Mz2mIB6F+kkRt/e31WmrNpdYs8tm+6+aPwuEAd0Aqv5TbI4xbTWmnnHzLWwUzGp5
4y3d72qWyQ2PcWipOQOzlrOK51gyVYxkVG44V1pTU5h3GRowkqigqMIeRBJc2iHX
GUMyqXCgp59oNK2RULyUGQc5rgqS33jhvVXyMKdvaXdn+qJjh0xVzf8rGM3HUjRA
qRpGAIojLtczWcZH3EeV55UTLBiR8Lqe1C3w6q0UhBYEIF0egYfx+xKttvQryRu3
3mnltXVo0ckZh/16sAyL8KsNTheMkiJNGyBwROz6m49l29/7o7j4hdeaXVoiaa55
e40mPSKogzjNiO0OuwWAAayEFueX0YARC8dartxkwDcaRE/VFgsowvFO5be+FZCe
r8QAdPZaiqv9lGKJyqtEtFYPhh9csgcBKgMqe3XAccHeP6KsI9QAVcmQflCrZJXe
xtRgNf+DEcI3OgfmiwGS1SGmPomfa9gNiXID4JkKDeGvcdVzHZfofGrQiNffvCVq
zCZP59ACqAi/wDKefzv8nZTq1VYOpCO27DlrwZ8LiZv+PHWekbj3h2NIHfekfPat
+KYAhFVmKgTaeD1OtU3WpNUo80SMtMKhVucbiDJOKruxpommBXU4uhdi5+U7otW/
8K9A//smiCL0MAqggQGa+ZRKvv3gjwe/dY6nZ2vNycicpZj0lVyA1pnF8bfhomfZ
xt5UpprBmJoHIQ+jNu/iywwnVDIgsSDVDJCqTJxEmGPMKNB5xz657auhsnm0lsan
bP4CddpH/5IMMLSp6mLwS1Zx4xa2XUE2i8nKgaTl0EuObgVu89nXdeDHYLcgrFHq
kwzzJwMxh2ix7/XU8oCrtlQbx/oAn4bmsSccE28Tady3eZebj5xpomdD6V0hAeHu
q8Dv8Kawk7qlEo01gXuZW5lDTLYbn+wZkzPq1LRERKFbmtsUySqj+3DUUi9yBq3D
UWZJAjIU8opVctDVJrydQm7oMyqRPuhjFbeIjKJFez2wSqdvUJMNGNIGztpZIEhU
vnFeGXGSpI2KCdWO1PwjMWrd43CRQhMP999b2qXwL4R4wDdOUR6LLUrPwUSey5Wz
9BvO2zr50kM5s3ZM8aGIYBCotXtr5uyBS+ASXYqyM9YAeYq0nn5TREqzaOLWuEEm
bJXAAQOBq/iF5BhXtEsmWSr7ylHD2Ttlg44wdTJY6dL0j9MFjAI6aKctn2J22Joj
b/AuaayRtUvkkhpQ1UP3NT4LS2XW9AjafCZjKsIkZnod1w/LYuWWj8TO3XMxPKQT
SJ/hxr5SjQ6sZaZRLdDoQK2+GGYIVVNAE62YuKBDgpaJGcyUXIrAJaMC8GQHPkZh
x98DamoHgmKEXg5K7KCLi7U2Quk/GKEEOybDGMI+q0TJPo8T2SlUhx8BdbUi7EV2
rJKxpJ/F/tXk/Cq694e/rMzua/dxTPhHynDkKbGDKlozsyMAkkwUgQej6p/X6XEL
Q2WD+5zOxlOf3JAqEl3cljDqgfglb4VuRk0S6JrjcQzIzHMq0Fn0benEYVE+LVv+
vpZCkYh4jnA/mmgkyMktFL4E8TinkuXv5T/LCQjiKyLAylIcwQcWHXPq92OlChGL
Z1tt6efBTWbDyjdceXqxBCj2FbB9RiZWhebhxFp+dQLuDpmYgiYDhyZdgWUitP/R
CMfZTcRs4qychQfzv46U35H6+kla3UZQjW0QgFOfFXVeLWFxQwAHlP3iSghJ+0y8
FYnoWTqvrYO5iUCJXzQUF2gGKiZHBJJog+vWodSW2lHNqXYKyLfqhXHMw4E+dIgF
2BLjlSb8uCxFqTiuhRkuCIbgMSkCow/K5SoSrtQDrVmelFcxYaJQWFaNIt104vXi
mW2OEY3UfqiO+Aan4XAzYfG9jzpMpsr3iAgnTHIdvxv8XRa/mChJ52jSRdV6jCZY
3igdx1NtpLsK1ijybrwbyE9iWAqWgs3IqcYDuF5Dip0Ceu0FYpv5qmj/ucCWfT6R
+2xvfRfo60aiRQxta2CW0ytFbiwhFZOiT8Z4KtbPlrkXMEt+XSEA3fm+rjdnipnm
3KBTzv+pDigTWE3bkwhA+X2cembnpcVrAVN7MZ93wCWJy0vQa4OBPOMUqQdUH7IM
RPIpGjD70UnjG2wwd6alFGChz78sUhrMUwiT78Qlb4B5/vsrjDaE/uJD2XfL4aiZ
zNp8NPjeuK5Ng3jexaoiUa7OTC9BUuHhqcRqbijtFoH351iPzr8syK/2uFlGWU6P
IriEj+SPKZMP18fwHNZBCtXoV+IGtmAg30eWg5QWbtXz3cygQbtlpnsXVdTPGz+I
lLdaEoJRTiTAy6vt9I7/pXmA2HEfsspPAY1QL95AWcsZDXv21qb2BXjKFFEYiCXw
mAhdUEt71le3c/mD31Y8grAKxdowSz4hVA+2vSRettq1Qc8dTbqvFF96NudFbmim
Hn6jaQ9AUO0ewi+2mdbYdB/n3y/Q9iut7nVKHZ0cCM15QhxZH6qatQdUzbYTOnjX
m7k/B3oHw4Ju2pkS1KdTId+6wYt5VG7LjZY7teOMWSs9FSY06viTKP3gvNiMyRuk
N5V6EyTbFGP+sRLSKy+cuKf8pQ1MKxqeiSrXCpEfjeRju1rv8r3u3htfLyNw1RpN
n3fVGxE/gD4dkMROv+v9vb0pEB2enctGi8qLmXGtjWrTH0R2kjOxyFWBHBjPurv8
nhAQIbZtESwJXId5UbI2AlwpqZrW5XNtgRqvC+2g/1glH2r/DOYAzIapBy66cHcu
ooyB3eDxJ0axnwVjvy/I2i1ZaGylds83SCweMnMc+EnRBgm8+DTy1d8puYMDSx+u
NRz0oCsg2qKTMMWRu8TGA6m2G6OHGoQwRpf8QSUME7shOWCRaGwdmI6j9opIi1Uw
mJhQpApG9A5y18wsRiA/WnUKl2AqzuzkDjJXw90OsRP+wTVSMsVcsvkwHZY2HmN5
Oh5fMHte/vSAYzlhQ+um6t2Dh0UzWY3ayZLs+VV7Uf2477EGK2KrRW6quiX6967m
mnGwTmWJ9/lIVvaC5ir7t5M3kuSlskTtdSTaBJOTTGdZXVnHspfJOZ9LpMGQ2prv
Nay2jjCwtTGzxTwmwqw19yRlA3Vrn8p2ZZYMQVSMEi//iD7/1GR/38krveSpAHvS
Nwv/lmJesHzTxuTZs7RmjCqhmrtrD69M8CRo6Bc/4GQVtAvK+cRxCfpmIoxhmRYC
qCn8IVsLtkEKhwtgv8iKz9Tm7XrR7VBNCYcXOA0zBk5ut2ovuxEfm081BTG2r3ZZ
HFCTi//x2WI48/+1ywvw2juqre1D+trFeN69aTynbU9ziJefdoz/bUshwa8+q90W
6saMi5OxzOdHkgEh33RTKKsoXqbFc+IdN/gqAp7rI3ABAqNbvEJEue/oc44tfpcE
zs2aqHdKGhpqcUKTsdgJxw2uC6ttUPG2SOXI2cM1f+0AecyHZU0Mrbyd0iOHL5qe
mqjOAQoLPXiXjEiGBGPCgoKtbogHmY+6v/XeGcSoQFy3l05RXizVQeGCSjHnbtnv
kJ4iUjnnmmcvr4SoRGSKwv5pZKACwGN4nKTAtKgMfgTFRRoaP/e1W6lzZmP9XzOA
3S9X2lYiPmHZFkknp8jjP0DHHVDCLjlac5RVa892ONjuk6FAStUXWGM7CeivLpCh
cBJLWHdtzLRi2u8DqufdmAWJc594Wk3lUFAA2HfXnvdAVbPAg4JyGGaExGRSfefg
jO3OmllZN618R3eaI7Feky824adnDQ9cGhw0nLc94Hnpure8tpLXW1LgDr7fcoq6
HhBGwWOorgyHn3Nyd8wsZEYWZ0ZZQ0t3xUt1biJwjfchy1ee7doj03fHdQeOAuMH
Z1nlrNmKiRDUSDnvfiSqSgIWH8ovMYamjyEHyDrYa/phIrxdHJrztJOELGgw2RTQ
nUwb2XNegEODIaOPHyD9tDxfcuFMpBAp6Um160gD/ThmI3Eo9V8CbPIr376Bg/qW
mQdT1jS6Or9kLN6LCQFypZ15tks3xz45OlzbUMH3ieHZHhyyAapA9vOLeH9ze9FD
U7UpkrIMDVVb/lvcoDWbMOUNXHGhl2Y7r1MdFjSiZo3Uq9VSnDT2K/ztwUpZnXFr
tKXOSLf38NcHEKrjRO65QKjShFLxEm20WHUaPYtyKiX+ns2aKlARY5Y24wKhE1y7
wh7R2PizBl9JmNW6lGvK/uzO7ATX19bqoNyrgAolRiJjNGVpSnw4rWFzj3wN9C2I
zPeG1o7KhMXiMC0KYC4Q+9k6GHCT4sROC3lBOHz+xqlYpMOw7ny/xZ0Eo2GIrFT1
vGsOsVaXMHVEkspV+dwqJC6ljgikQ5KT1avGD2pHm/d85YG4p0RRee+ygL+gy2w5
K8FcSl2Ju735rmhQH2l13EE6Ob0irmp6gYET08/SvZ6S++eVJhvGrk4lJc/E6NhT
HQs9kmxIIfO2a9JTreIvj445I3pB59UYuWIB0Rf/km7RQazG0jkZs08yQ54+hRzg
VfvEOhP7gFI18jCj+3aTb/FyOq9twFXIOMkv4RTLeEOkR07RPG3TW6IOTA6T1OS2
fKF3rgV1vFO5dU71d3+8OEaEfA08JdcHiCrUjTGDbC0MDmtBJlqpNahZZ241N68V
n90cllYhuxLjowTNf8Fx8SOEsYdoB3kuDQ9GbUT6AWNCEi4MXbEgnjwERscfpYqm
+4+oc3RcCupiRSFsCxMXl2C/8hkIg3DFI+zUvs9okLhW1bQwg/3zJkQPMuwC+a9A
YUgDFyhht6C3vWNtIIzeiY4uO8iDJNu4/Z3jke9bAuay52OECLNlHuu4lZm/+ZyE
aJvj+c47GlvpMTrXZ6qpKc6zMnsiB/PxdTat6MB1XfOzL47kqFnBg3/IbO/Lf1fM
bUuVjLOnhszJnNjDQsGwuBAXfzeBqBC9oQKLZAS/6QJ/NWBFPGOW2DFGkArhZJLc
9ofIHkGQgC14KieZbCFI3hjoJIl3lvSZemN11Co9o9EO0dzW2zzM8L3y+ZoVB6c7
W6Xtn8TCxd2gHE5kTIJUE3X2Q3TqG3P/Sj5XZVo+TUjS+0GIeNLjZzz3h99ekgU0
OMkMoGCayF+/E7RPOoDClXkxGBiTBA8lVGqIoVgfLgSQF4rrcp6DGj1H1PVVhydl
x+OxsaEd1S7rAhuE4rxIFnPvb3nGoUatAATa/gz8wHP5XLkKMTgK75sckmyzjptK
9N2MqzXDEvyOba+8sGeVVoz0wYFZ4B0zYp4I9jYjqvcLYqHt9AM4HpH0AiQPMzPf
F7w+RRu32CJnxNqgBf4Fj3tKMHmjhXPFFeV88vFGFgw+wXRJj3DSm+S3lQwwSth9
LI+uIVn1+CFaV2c8wx4gfc1l/ARnYvt9/+aEQ53HG5aj17E8QHbjvFByh0XY1C8G
tk+To/C1Wy6+jYpsu/9qpGdZvCjs5Cg869blJkmXeBlRcCBTiS569+8XUyPDJs97
CR9EcIR/GztIUdzpOxRIEjrFd0DpgQx1E92ANf4Zw/aY+T3lcI18w/L3OLcWul0E
AHaAcJh1dMT6abxpUKN7thQyqC4VIGAraRDCrteksDK77btWoW+fSCkTXMwxJE0C
bpEBSDZhc+p8vrKo5j4XqDju41OoTPjS1twR+QF0V6VDBGAUjmouMUYwXs/5uwvZ
UwBDR53ZquU1RINvtlR54DS+LInIPIdoI0MLvjM3o8wI/2M3VXQmn/d/6P9ccEBi
Kd6JjOSKuuzjefrj98ffC09MCVwFKhBmWJT/IWbDedNyiyG0eTjcB7fy2mhVaI3d
0Um9sBiAKDg7Tf2cF2noc+xRyWnJ4QKGhIXvNCCMyXVHeviH9OxYBNrbCDwteyBt
TGIri9W1BOns0MntdFKJRTTsZXLLNMj9bz8WaZMXWStiIh3Og5ArmXT0lxJxsd22
Ixrb5BtB0MDbEnQE+RCyRwvgzRIzz0Tzu1ySvu/FE58J6m+sCb4Y80pYNzsXYFaz
CeJ13vXjqd3LswsIkZ3RQ9lXpNA8hYFkvGoQJjPrYglM+dC2EB+dCIDaBppoPjav
06NMeLW3Is69spDj0y94vbKwD7DFArwQbbKEq+xrc8IKz44msyFbb0v4NMQreaol
X9WHX0yFb+P3aT1llnIWn2wuJiI/DSkRMR0mzjDUV06ubeCV3fz4DJZIyKBTxGR2
c0YSeD3T5StrxFN6cJ1m6p8LhUQGIIw78vIcT65BqgpH7WrkvcVFDPZ8wKdzSfjN
N+LVWrEYFeibhR28uUcF8TeItgdvf9r05yAIMO1pM8deyDTxE6WhaHywF+x9qy6B
I/b1iilA6x9P5TdCutAYSIV5aQa3FxyLZa+32FVGY7zUKT5IRMlJMyjImmue+s3l
zEAjl1E4mhNbGq9ItQ5IABslwzN9ay97oMvzwEpgmilij7UZvBNvHzIWtTphCIbz
IVrNylRp84YgmDvIHl9mkMgmD7kuyUoCX/pwacanB6qkb0iukSoGE8QW5Y5IoROf
PD/Nb2HAyaTtuYZcFgzETDO7Zg3g/oH108VubVOhMEMZWjS/qB0rbdlYhEqepl9x
I61YIpf0OHNMofkE0zNgSZcU4t4M5T/g6VHI4oktGDzRAp8oezcVT+x6PMzpqMzg
PicOscQcjPcAow+mJBT5OI0ZcYOZwujbiWu9xBdIqQjJpg/mDH9OVCr3xKcPaLGQ
XHyTGZ4BmKTnBI/7A/eewcWASs/deokML1LkXCKHFqFGzQCJXYonF5hB/ReW1Xh1
fk/m9tcMx9Bgpo6XdSf/Pwz/ryfSFZ0e7uROzbr3dIjRTD47u8Ggf+f3gG6PhF//
xPiRFQE/iTcWfBpagjvp/fcDd1PpxNrvtG66A6ZtDwhHBdbmJIY7nmQ0nduzrkNH
6JsJp+XcOswpzSnwjZiGCqi+m+UvuIhSrV9uPcYOVmqNDyMgt36BmPdB76MhFzp3
w59G4V8MTX8Ki5rxSQmCyqh3O5HkvqQF1iULF7Bryw75qWw8/BTlRA3AQK2dbAfn
rjO/AIkkSuRsyAQQj9Tt5mYDQcME8BQIEkn3BBJ7HhDZAYO6Efc+MfJLQnDdwZ9u
d2g+sf2x43p/azzYD2UIc8p/Eq9QzWSBv8JdykKnlBxmE35MTE5/EAlPGFNIVZDw
hAJ8VPdwDYC/FCrjpt/P6MsEZH6B7zbepAgWSDQClQJ43cdxOqEhKC6vljmR4Gz+
Xu6GfwiA4WkME9Z3cO3hWycfG5QCmVR7s4SUr7WycBG1/CKq+ikDO/19VvGOOQhO
2j40Mo193sTD/VTBRfioGlzFYVLurS688Mz1ZXhqgw1R4fku1guptUeObFyEUlzZ
b89WebJpC9V3tbVm6ZFhknJYaqQXHPyI7Y2pSIK+jIU5skmfNTkG+X4iqyoeQOwa
BFQcPrP5cOE8jcjIhBse2mqOhOq4zwoSx0XPyXzMghRAk17fEd8f5k8AOxESmUb6
FYmnT8S2+nofg4yb0JrHcwRo6pIrgH1trFWKVt+3UJAN2F3iEaWRuOOsZm4UQ0mN
twuIeJTzspWcU/wmk5rIFw3a6KCh6MY2YtkbnU1wWb2IbdlqN69ff2KX72OFi5C9
tXJqAVGb1ldDIgTJcN6mv/K8+TkVTd95E1J3q5UUJ+daWMGcSwf/NaQVIDyvHZAX
v9VqZpCs/IIUBx0Nj1r6e1O4tDNxwoYe3FfqkxZqQinZX36RlNtf5UNCBRvPaJ50
M9szIyIeUsYUQkaME0pOBWSzHOfQuVarHHDdXDpmqHdaVTz9zbp081aOdcJjtrH+
aJaCWPFXpdnqbfzamHR6OHXPpe/dsBRCSI4UOr27sW0DrRXTtPGsuyZOxYcv4MBO
WayKH13YkoeBZwDDhIPtcqR/TXp5xQS57uDvgyn64YOdRgt2TR/GWA8Z/GBUq6EK
cAS8PH5F9DFvO5Y7GoS2wmrL9tHyxUBkdwK6k3QmGVvk8cfww0e4TZlSNOBLcyz9
WwjPHLV3Eq8Cv194DRFVAXli7/Bw6fx76CtSfSXkNGmdGYKukLlIIM2F4474+Qj0
H2yND3P3PvNoKatYHWzJfMJ7T3/CgQPrLAKy+EK5+RzIcp7XWBHm7zPUdv/wwr/C
hsotQVQfrFe8EBr9JUwBHkc0VBn9KMsiANrieYw45jHOSXIX1ru6ZHX94cLrWAh0
uLctyvJVyvF42388rc19HXG62oKexKDdkvtxSJZgQ4J+dX6Q2DOLiR0/UqToWIYn
08zZUai6v2I8rvNad7gTXGWBy9N0Qv8iAne/ICdtGWlca+xS9vFSGcoFXr6/7IAu
++ICS9HEHA6NXHcBTRdeWI1dumGRRyAhHZSMbtqytz349iVFjEMh0qi+lYtjnNP2
QB+yFmmoFctBcCSaSse38C9Lyb1FK1ZMZ/tW7appbo4JTJqs8HebfIFafc3mbI2I
gNlbg+BuQtIFQBZmE4VAVsFWeLXDvC8Ayp43/YToZOG65EoSGKqtsoUdVrYZxw9r
9llfj2cHSlXdY/b+6vyRpYxgNIiwBD3d5eGYAufa2p9D8R+WxIyojaXKsMK0KHn4
P7ZHo2ErlRKaSmRNO4PxjEUp2vbefrA1VMMGYOBvw8QqQdTmRMqVGDSyjlVnN7xO
LY95FfOL26LSTdaWWD6ECWQJPNeWT9w8oZaxKcVjHCEG1JIfo3ca4f9LMbb9LxFi
mAWoPSy/rCkLc1pGOM9aPxZCudBOq1/+3Ti8jiiW0cgzQl4qjefPNdcoVR34W706
VAWV+cT2xmV/6ysInxDUfSMDAdeLbsVUzELSF9yUdSLyVoNv5tiqLlBbF/tZ7Ofk
knezBPeILWpnV5gLFYPDhhSUiuV/xUCBPhhaYcfiIzMQc31e5vwHyMqNu4cspqA/
GQj3fN+wsGzo48N+TcswvYbvv+yp9oqkPQqy8ut0W5laEw7Ng5orjVjiVk+5vRDX
ipERGQ9at2P0cpzqQ31DlI2l9TA/e183vkN46FMpOqc5+TvUKmwQWe33zE3pc1ir
hzThriceknIwzRcJOinFgWd1DgPbIGgK3tu9OxqC2kNYyxIfEl0C7UN/6Bii2qGj
2YNHbRkSbaKlIv5kJ02aBRV961p4MP/u4nRXAqcjp//S4UUlqUaQ4iMTG4MN01qe
3w1j4qmZrOE+Zx1j60TnnfI6YUtAGhAjXiJz0Rc32Vw22xFdylpJacRk/GqifSv7
XOrFde97Kz1B7WDKyg3Lb1p291zBgIhw817RtOC9OqCGbcvog/acDEoD0X5Fv2Jy
LvPsE+pySs5vTEuc3T0i/cR6esu9Rd6ForF6YhzFPBH/tyi/Aw8K58eAxEsSHkqW
aptDvTnULKV5AJrGJP7lalHrpbMCyo2h5mjtm/AusnS4zBgU5PfDaocsd+LuRznM
aYU8nw0aw2F7WhAT7aXjVCL02ZEF6qgrBMxJ4w67M5OmGV+g1JyiqOOQ2uVjvE5s
PpHd/N0M+6CxorwKiQWB0m620tMiQyxEW4b7PhD07lKoWbVDArqShT+w1UyaDXAt
CZFTVjFjyZEjPQTZO84Y1qwoX/8yJDta0SvpDyADDhb976ChHbx4xWA0wieXe5xq
cCBPu98Qoig7csA7j0fr3ep8N5+6tsJQT4/aJJtz4yI2NrbMetYpPHHY9gfYpLJf
qqetKjuant1xbrRifSb+Ip5ddt6GKeATvup0u/ITj0gYG53t3ERxJELcp1OFN7rW
W1gzXEox7tUmSO6q1jsRVgUxrT+acc9PIvGA1/b6y2kxDWqBsG7pQivCcVxl9cJ/
grabF7qPL9W/40DQ8eaJArsouXbYeL2mQix1AtoexK6EPTe3dFbSpFbuvo20ZDN+
YXlPA/IrafEpeDd1RS2FRCkPXATexTQHJ6iMUllEINqLT7Fg1DjJpdOIUcKYnHDu
yMuvI0uRhzirboh5SeV9OjwWa/wgyRZ/miMAkBRGLGcOfOFTmGnou4zyUdgCpN4x
1lUeRDT1TTPVy9FloYX6Fkad3jWTUiDlCoXKp37tQgPcO6CO4aqCc+JPpmHEODUt
E4B1PUFg3o3tDXCh5yPEo+Pf/UqyX1fYjWwEc8oMptgN/MvnjSU5OPeRlQTdA/5w
vMb5bOJrTSMZ+PhounoRke+rU7+A/OlvLvmgzbGi0tRa/Qd6b5B870FhanoYcJ3Z
DoqB7FqBp2FC8RmPEvv7C6ik5CgsLGRYAYN/lswFn/4PpeUuDz+wBDElFyrhxT3F
8gwxs7MRC3Y/NRq4RwMd2J9er1OtjFOoFu4YsiXYFvBopRdGjcjoffnAkYCSJeZL
IbqbywrUiyBBHGndpBq4sJXUf78V74UwaKj/Iav7LKwhMgoDdnFQsSL3H62bU7H8
ULWiVQ70iJ3BBarkykYKHR8QNjQxqjKZUiYENoxCdumxz3QIQnBgPsb9Jl2Y+bVM
8HhiLxnuhiA/P3H6L1UXkRClQC4jhf7cGTqQ0fkRk+47N4EpcERA8ExkbEVQ9MN6
gC226Dr2XnSkaxNCl09uBe9pKPVWrOKLTuqv7DA1eCh0+fL4SYH9BWuXfwGKUucV
l58pRtgerQthymeDJlsBJkYs3cf58A+zHUYf2SgS4KfLbkeF5xOf5kRc7SBiK8L7
cjb/nqrF4iaxSUYmd88KEUR0/WD6tf2NeU4+s5TcOIMd4Fw9MRSFGoIesZp4K0uS
Lw7Gg9SLUPBQu1SvnR5tk3t3Flo+Nq1SWREmemLzBXCXkx+TsT5QWgru+1vWbZjZ
WgVO0v9XFh3yytXXGey1uvGhyqX53TC/Cccim7Qh9QE+DhD6EW/Kd+A8td+3/yAO
u31rG+pg8EGl7IAuDnI2THb+rhYsAIFCnKu9jExMcmae1CwUQHZZ/BNJ2STMhOn5
xwuYLH3Sns5DW6pnDTX9Wwnc7UYVvJRJxY9Bp0S4MZ/jGLQY7CXZSA2XN1ZAm1v5
vDLFBNf5md6BsDfvBL+bJVTfR0HorgpNByl/1DwU2Jl8rfwbMzTpeOcru+rGIWgg
hOWp+vOFkhTuHuN2Ep0xlE+P7cgCtQXJsNgj4Msuu5qAu+q0TWmqXT+I4W4VLP8K
/zUONQ26i/VPl5fa2xviCc6jHueo2oYQOOew+RExlz4uUSg27qi4BXhYF922wfr6
zIJ2W8dr9ezjeXweOMS/LAlGseaunolWB/u+sNiee55Key5gB8Y3OPmdHAq7c0Pn
x5v9RY0jfDIMviGjvLPVONpMKksAqyNraoXQDncchI01UfHrs5OqaghkZz8bzqs5
X1Ld1NxZzUDbVYaa2VKhZt0sz7Rzco4ZGM5CcRNXSyfPf6PLEMZ8yz2Ek6Pq7R5j
rH46KGJue6z7nh5Xx5xHq7vzy7thJ4mvhrdDshHCI9V+olAC5ur/6PpKO5RD1z5z
xxU6vZdqXl1Wa6NlE4defDSofYMwPFrR9zNlPSQb0nzqoYKzpXjmoBRTgE3z+aq8
9btB5nO2pguEk+q5Fp+DiBgNlf7NQ4RsFMpfiRNyxh7IcNSlrLeUtHjEP+q//bx4
/TRSOeRuekNfmqRcuy2o1WYg6/cVXzTjR1dhZ6UX+6edfrNiT/EXFJAV0RmlI+Ck
oMrQJGpWIrWH9wGqQ3s8eD2sKXonZYymIij8de+qnQUQMIGyBTfaA/zpbsNdO6ZE
SH2+iHd2nyYGYMYghjDNcPwdtV+DbkcVZ0U7lt3JNCqYYERHcRUwc9VfsaAh4Pgv
s1YmgAWdwzSDfbbl02kTHk+pCGrfM8hP5vOF6BfwHLkKXDo0jbCUB86si1Msec21
jd3HjtG+eamNwSeYqWh3cxC3/nffV3vWSOmyAQufZryoCeFhw0Cq6y2FrEPt4QPE
QS4ZEKezHMnQhHODSS7irjuxSWN3oMZ4UmIyLs0GpaLUCK1UFzTcbCgsdALPrcf3
WNzs4CuhXrnt9HltFianTFvTc7H2ZO8fhZYT3IwF8n/ygXqh+AIG/Aq+z/yhEDEd
v6hFby/JsrVfUZiYIpBDM/iD0wxBvrzG1+meRS4Whqm0PbNbhegLLplyZ+yiCHEw
bbfllGX25/1p9UmoUACIt44WVBNEiW8Y9DrzggyZCnTTNp5Da83uo3rSjrpWX274
crCEgSu49QeFgJlotmFeRXKIf+FAVxGaJx1yt51/9FQcLs3aFWg2m/Fh3NiMDmbh
Eq4Sf8PV1sgiD1OhyfrM2ju9tWEyjRxXElJGkg47MCV17T7JovMOCKmW26LWJ1EQ
0Avip6u1uMTXH6Z5gThJugdaWqGXmJCTVmjhB4OI8aVFCyQIJ37gLZejMNybeHO2
5o2L6NEl/MIXZGmqNK3vKpI/BtbZN5prdPNELpYia4MB6E3zx7Jj2ueRTLLWmS09
IBidiTfJm90hYVfPp7an+Ek6T2VWIRepFkpNHwC9KUkgkZ8QOLPZN0YmKvGe3Rkc
HzvzH8Fm6DIala9aSlSJOv0lF1X9DbOZSXStRFlPJb6cG6gxMyI4XMx5gFye4X63
JV1gHdtaef00A/I0waLbeNb6J2BNRFn+wm1pvjEnIAnPV92K48EWjsixlfPN52u9
bOjjeAhHXhuimypZ2UXqzAPkkEVBNhjdDQVAiipmLTxHYnvW/dJCV2QCLHcFPZcb
x+Wd0ej8yzj2c2Ytx3nKuiLoaNTXnsUHi5j8HRfKXI2TIv5jjqY5dpoiyU6IGFat
/UXMD2YV/Pc8eJlJk5+fPUIyNkJHZiS1TfmvWDqRs0juAcP4p2Ycz21fyxG8h3JQ
tvLqOkbqoUc5Tdb7myHMsrXbiReXwY/rW2VOyYnIvjBoo8s40SZRwBH/pDvA27y4
exUIl7Ay/UhWyZrJ0+MjGZXz/SDTdbY3I9DHojw3dLBYyZXPb7QNLfJ5dchdu7RY
Agow3x80bkuBOlZfXtQCvf8b22fmdnjvrApURMVbVfK1XSXWzdW+znX10nNHbLOI
gtNlKuVo7+ut7wStBHtzDTJVUDNDjYR7aXM8K/9ICAWHR8TZwknyaDe0X9aHVBGH
4ZHrT80eyIkLZswp4v4U7zaB0l7prQCnzrBld3grussUMzFkwNmQHrmp2Cig62bI
wdtcawUqa+85hG/ZW3zRVDaNG+/p8RdVE17nM8MEdkb4f36alyRZyZmZiSpYZ+6m
EU7wHeiAM4A1sL/Dfs79vumO4BUGsn/jTl0nh5L1GyFHszGBvmiOX1mfyzt1MuUS
4xzvmdW31EDLdEN+nlXT52zf5stpJfbhLjHRNl/TG18xjdOxq4nBucpVa0tawZIJ
hFhyGq9yI9JhUJ14HiUJrPYfUjCqw0qQGjuAo279YfuVEcan5kFIdkuQwDPM+f0r
VExdN3d0nHUJDNf6uBinsMeDJGyofL/c86MtFPhh7daWeaGRtebnD8d7272Uba0l
303f7cVy4UrXuYW1pMo6MotRadCwstRbx6+4dAGv109U4g2XT4wTDcEvK/s2Dpi8
lO/8ERLHwCZ3TW/YeHAYqg7GwNeGNE1AEJjXFWkZEUTl5EjRLgVgao4IVyfWHPkG
bDIuuX0bboa+M+dzrJiXZOh/dKiYaByXpBtb9lthaKbp4mFZq2asRGCMt6551Zmj
S2CDeAv53YCARtzbRxj01xcODkeSzP5cdE7Dsj5CibDdv0FP6ODrr6D8cNcl2v8L
kqcP38q/I9ORmt8gOEVUuGO/5ylNgr5lopsBshqdXWqMkymDoqoavhBe/gnDwkMM
VTHuKMCZIgo0VLe+hAukFwRFjJcwuESc7BQUD9TER/d10AsPCpYwTwLrUjBLhXnk
mETSSNKzUa12WwhdEdw7hK8Gj13mEGIJgjftsngqdUezTzMCSKO1YyioVh59ZWs4
u7mtuoy9NqiPbWBrZV9livO+nvdrHb0Mnvk6mWQ47QfOyLMiBM8fUy933h4amMnJ
dEAonTuxETF/1BKvwMo+65Y/CETRDaDuy1waosqfnoZu7V1HOCBOgt0/E5zwPOiu
TPtSQTDBnacNu/Wf7jDbUQeIUSsysDDE9PG9wj9l6lXIUddQ8yevy00wdpBHGk/g
OpO43J0rqZjUl5x2U7sa95CXxxFDLO4/ceBxkv4jL46dhpPIxuEP2VqxKAyHLCyu
mFacUiqLRcnTMg/aatmgp7MvuTQT36TcOmYzv+STzqs606VCh8OdI91SBSCFlj8O
qVBgeOobeI+DAtjMn//9T5TKM6z9OeZZuPTnh4t4FqxZ+3H+Fb6UvdiMe0lGZLSx
zAvMMMZd8IqoV8+H0aGJZYwkUJf+3M1Dft/3MMb9dSO6fmdddZY5tseeDYt5OcSR
0UdhPl4I0DarSy0xFP873Z7c5p5GQeNH0DXcCqqIcWvQtzndyqyep2oKcH2TW7Bv
PXmAMu9XZwVdKmgA+zNswLGdCumOBMeaaQSK703jgJscmW5y7Hzth+vFnWCzD+5t
lh1P5y1nzJriZHbRcFzoHvf+7bWgY11W/eqcXc1wqIO+d8qAlFoBx4FJkmEt6ma+
E6CvtvB3FnKFALSGpegEmodtQWAQWFlzYMud4FRik15hMIk3RxZ5s1Zg9U8a/jrg
DH2XzVJ0c5mQxiXxPFPddtjtPZtTsFrKzEepPK1m+yqKNlMRjedAtvRGYFCkifRF
BQHyGrlQzY/poYN2t+SrFrrZ/hQaGX9oyK2EsGNYtH3x/7dMMFLpQz2KYYJB6GFE
H6Pg7mJBw32ISEG25BWiD1KsZtX+ZNafU2KayPj8oV7MWI6gBjsE2D/fi+nQ0Y2t
NPpgWHcBqyJlt4K9blBaYSqoMeFIK0ftJwr1m2jR51U3BO1Q8ZXOgCpV44aQ1qoW
dbX0qcIC1ycLCOqiAo4dfBicatQUG9Lu92Ey9JkjFiGnkAtZZOqbaZmG1xQusoMV
OWJnUahk/nX5sCJhPWGdvQFIRQcU0ZlYZ1m1AytPMJsaCxoi2KUcbTx2Eq41ZwuI
GtDObH276rIcR1P6jRemVyb6jluphsV+rcw6wuBnVPcAXBV5Re2RJieMjKk84k5k
IUMA4rarm84rAdqooreZl5UC2Cb3TGJQwZbnlOPYBFQIpn0yCpTcy11bI+UuvEeq
x5ieK0puARkvVKsedhx1dUezc4yzQDpMmKmLXfef458o1gg3pxZbXwE7zEv2vBmZ
IwCbSHaih0rjKKDTr1JSw3EHkexMb6CzFpEzB6+tczcxho30JUOc0/UA9WEreVIF
PZTjhwR2dg4fJdjBjzDcK8Nka5r3RaQ8UEOrzChjHMJk68qnHUXo+C+0Cj1uXrm5
WH4t3CxFBeieaktyS3jS+fJvZF+WiZPgEPGP2qsFSPRY0mAFeivCxe9cfV4nSUTh
UOQ4ZZ2kybb5gC9YdsQfSlrXu+8Aq3dYbZOX8KzTxc3ydmvDMQ8Qz2qEWriM1l0Z
J73/Ewoigp7q71eKWIxtABt5pvxTeMQGlbuXqLADMFcHzb7QeSxAi7r4D8eJdh5I
0RWNAC0QI805N8ILiO3IaoBtYcwtKY022nc+SnM4HeTujwRkai19mUwvPND6+Cvl
irtRe8x/SiHe4h6BoMiXdbZ7bFtyEUX67+SHqhK7CtO932KjP0RzSAsVOFWLbyvv
6UWiGn3bjJo6PJbXnSoVqPL1Vkimp9Guixl+J0MdhGFh3Hxn075+AVRL1DNNBlNp
yX6Y4EKyrsLvvHF0GiWMnm8OL2/bruDATePb3HmLiQeIybo/b1cJfls8VCDHuPrj
Fzg9Xzasuot8hOYTnw0Y7KFZ9movwsThfTcvv66tWMOJckEvsgUWRZsyg4eEOJMw
1+p39UtvES/ROkpP5uP0wDWqJhlv3pVMCLDsQr9UmMcHYyZ9jeRHZyQszHuiKUd2
abs9CmCqWBNMg0hPR8WrpYvTL5XGTbgj79s22UZsFf9NuQtEf9DEoWLuWQT4jlxd
0hnOzM+Ou3NEenzpCXlAgeVDJkhRdsw2x4vPlw5+ydKYY9F3Kp8PKmHtNhv8UNFi
8FzZHxnv4/WJxynsNf+dwhqkMxIlZzq65+byrHK79nu2aX/p35Ut7XPr7KxTVXKJ
ufObwey13OuaHvWoS2l4N2hA2V+xs0lb4ul8jF4Oizi7uUdz9trvcloVYK1c8z7t
FADH3wVgNWAgQEwLvi4cFQA3UFLAP4fXn+XdO/CgUPMnJ3H+J4W9VXc2EgI4t1jW
dTs50oEqFMBzOhrlrh0GSxdWW0c2sjU8+/54zaYLDH1ji9/VAFkafcSJ5yLMJiB1
QVXdOT1aecCHvFKsrbzgwRAE68ofqwwWJSeQQZhNLhcV0a2Ew8vCJsxZVfkOjrTP
/t3BlP5c1Wfs6U3Bh/+4nXxymrmlonHxgh1pAbMA5BXYkmo2FxhmQ6YE9KNIrr90
mZLboIk6g2K6/aCBQo6Ykf20iKuPPDQ6BNoqtUZG5Cs6sIsrKhX61CLwOJWBilzn
apqEY02HmunqNUXjl4bZMuwCffK5cTnLBN5z59qtuhcmY5o52JABjNmW/xZA0qHD
EVuHRNyuJCeiBs9tuUiPzlGsdfwqsJ8U3XUQehk40sWOrpGWDi1Rs3P59QKwf2zT
jWD4UGnkXPdQiFbjnJqVK6ZdcygkD3PP8+mSZzR+q6GAvonWg/EX0zIUTQPfJoch
8IgtMN6/oq1mx85pscfViRO20D9T8q5wC+VAHw7AOcnaUw+tNmlNcYRaWH/8Thbz
wOJLglUT1D/zyg9og3YBO1vI1ZiXCvkQ2P0TFNZm7qRk3yUPfLHZyXX58oFo1qwj
aCZ9m9SAy3qmobLw/35NzEa+b/N591VM9altjNrOA5rkmueszh6H8k8XXRPeoB4r
wNHH+1OVMYMNiaWnmhRerKeM/0zo67wxQk4Al2B2yDIT34VrWFM6+eGX7yr+/G++
J0q/HGbVqkRfFkoYWnL8FEMLKC+GuBCQCie6vNSIwG2hWQqUgztjWBwNHpcmsYnq
WvTX6rDwmoRXig0dnW2dL9R8TcouU+14yDVaNHIv0XJ+5InQzZ3CNHIVtZIUHBuN
ZcxJVQ6km8jlRom8VDMFKq8Xk1/v/+rp00MiYlKxWBWeAop29wJhI3cmih9e2Vp9
JF3MBklHthPondq2+MkIGt1o8sdomqc5jjjULL18Zvhqb1pEZbLEfYx74n9kfVee
uTuqeRL4xYqFGCo6wlmCWUQjt4Uxomf/AN4ouep8Iv1iaOhj0XjUiEQz7UlT9bq8
4YYSHfzdJA8pv4Odez86Rxl191RSGrlMF0KiWvYMFZfO0rZMg53+vxk8Ayu+MOIO
Efwu6G7IVylQ1JCoTOJslXF74DLxW3qOliaqaWqZro6uEn5bk6H4LyVyiPADO51F
RXEw9Xt0ToHv+Zm7oJoF+SD3/LDYUX9i2B9Vm4ZJWLaTKH9Vq1zdW4sT7VwEj0Ze
6iaGEEsp1GXxk5/C3WCT40SPkO17cY3xPmF3c8fs6CSlB2Sq3HhLfpYTxhT8rTMS
D6lNSVMi0KTwLTXwkEAfTQRKXlUOxWm8UG1im5VgDR+gyJcfolERzt54W7ziQiC8
V640dlQdfC5091F9ZiiV/VIgla9ZNILHC386ydLMHA8XcBIEAyz9KteWIfNbs+1z
BERI205aLq1hDtZd7rNid+jR4V/c/seNuZujK0ZCB2uwKW70/I7GkfAgTUnEVhfd
/CPfAwXd03lTkqkzbnbJvnyTfAnCGgn101e00IpXd4hH0Dk9zBMnxxcVHpL5kU/C
potJO2VCQJlvS5IuT8/4k2dZxdFDt6oAJuy8mIYVct1497zn0cQMomrTRUcx68SX
AsDJBKj2zoT9nXvlxK2boILro8E049gaxbGHBq8hD6oBFw2Xvb2wYBfnlqyTQXx8
dJF7PcTVhIB0x3UIGFaDdpwgVXrUZ/TzZLEX5BKyliX8JkwHpgTOI/WDvq8l/8Jt
TkASbjJRLs/dljxXmphL6w+gXpndUHuh82c6qX4vVUecI8ILyGhKnVa14vlb5ctq
+wq02/Yl4ZMnmoxVtcFZUeLuvPsyWKBmeylxKZGi3Zp9GACfDNHiL9s48Ej94pW0
XzVcKKgiscH6Vbq4rmr6hgUkniw/gvORUJiP1YzbJufzbur2t+F//iZwIfOtZUEn
Rt+K2xMLRwHgnAgpiqN9GQe+Efd9s5MVcApILDh1RCZlWEbGhsrEODND9G4nbhf/
gTRKdXIbUKKpyQcthp8ZyMR02Qk4r7CiRjEUG0sTh0Iv4Wi4rohrbvsT3jYwkome
fj97c13QNjPZ5GkTXM1gB+feFSCBeWK78ltmmsjhqv3KiheMaEtgOSbfga7ztxzG
ezP0ZIjZe724GXC0FvD145vJcdKT419OKiJgq3FGTdkmYbKxgecpGuBaGh627DVw
66A9vSPRcbDRRgTngET8h4yOoK5vnkwTPeiZjIL5jM+3d6hEIl2etxxSih1ZwR+4
Gzm60FklTK/fgetEL38QS8dKnvqjHeWrozqDqdr8zF9Y+IXGVdAlkQVWHVOlwpGy
8IdIave7Vvu7+Hmph6hr2F8bMS67hdRF5GiPpez3nkc8jJZfZLUST+9Qrtvzr4au
GzVuRhxHw+NV0v2L/4W6+9SE52cnkzTAD95lN+ILCzxwdfsui9h4HplKGN6kC59d
t6N//dvhohmaSKtTbSBV51UhW1U5sQRDRCz8fLQvj43aJH8BlQUEiD3c/4FDfMg3
zIe+C74ctSYrn4S3QHJRfI49Lm7AkWRXlNwb5piDo3MuJ8lgqaItB/TIcUPeTuUp
xc0dE1gZkYLMrlWCANxECeJGvpjZfbitNG06y0w7tYTjy6hxF/l1GYWULd52h5R7
mxlbGcVyshtjuPWTlVrq9RnHWs3VlxIyYCQ8gY5t4OvpSPxtCiKE2yhexk/XV6mz
Fg3URVUzUpJfnhHaqiNGwLHGGd9wY2Lu0zCW8+82uP9zj8egLr/ZMPKQuwkOMqHl
VYZ9qiCBrmt494La+efvSaiWeKsWAx4PXT4DILMdrp9Q/VvIzojd4qucD3L5Y5qB
tLNkOM5Yx9APivz8H1GhdmkwE7b5ZENE9xnUYLKFxUoF8Lv8JnsTO+44cByzrbyf
igQjN12UHtfh98qq1w0RmGXZZQ/AHkxO/RBnuCR1/XWftCSi4ikFwAlrXh7kw+7g
0+xk2He6zYyUfnoxWS8gS/BKv7wXhwWtlAYEPAmXy/6Y7/Hshvf+XbaEHQssOEit
6YWNnD6MJ9EvgatVZGDtkxppd1i/8adqqQkCbwuPO2Br7dj7jbZHbljv3eSvLn4w
vaK7S4lJtzyegG5ltKAQ5t99c7XSosF8TCw/ybSiHJf8Ix6dWrjktwfPM+NynYyS
IKkvPTT8EmjLxzdnMAOItIgyaik2FVZh+UPjMeuh7Wwc9j2CjFXSBLRFpum/04Ge
DwQr2TqfDLgZgSYLavo+pzXI8fm8IldmtO8KnCmaeIscvH1GGM75SrQVoVOOX0Fk
69LvMDIZseq6NCbdXLD+kZscx8LHM5BAqCNv9UPqXN/8A/dE22uFwmMqfNnObxtU
fM3hbB20644afYqD6BQlnuQAqdHZlZ5B8/vFxLz3+LAv/+2EYoV5k3hdCc75IFqn
aegcv7xe6VrcDKTmwR5+/nfwjeQJzuSlWIpPJWVnzzY3tVK50Ezp5k5UQ+Y2z12o
7QDikrVzzOdkKx/7+f3MCnlEwBGss3yZ3Arr0HYtxoj00DKXUXtM22zawbQAlMNg
7S5P/5LEc5inqWEhfGmvPxouDyw0INd22QWRhKYs3CKs/6RY9aOPoCVoZJmtYiEu
HO8kJBNl2ac5pQc1CIciFz+G8RBIZIaauuxFhKZnHmPX0tCEdMJYrbRn1Yi9apRR
LbLBiVOCtXUex+4fGA4N23odw2R25k/V6ARzSYUS3duXAjXxuH8XijjQ4aYnRbCJ
wNzpHtZWL/LGixroTepcAGJVJwuJO9Qb/VRZ4VjBArOyBZWQHrfkc4UNfo/QdedG
aCcF5sH/5a0fwMPYfbLZPsWTA3q7FXBL75M0D3UYKzBgCthDvqTzvhIpvqgaE/b1
GMI8DYH2nz2RoaDMcZlgNrqJLQkoX9btAZQ8/GUgxCYePb69MjrM5vD+2z80j0ki
bqIFb+GZMw5kOHFiwiHpzn1u6AFnyoLZLo76AWgZ3dacCR4tPpGAAbng5MkjiZG5
+8TxFgSIN0iXb+3YtcxhxXOtKbeGk0EOiPrSbfVbYw3cGjhy2ZOThGOeeIpl7/p9
snIVFMKTQgpWDL1+1k5AOcYnODd5CpypJ1sctt2dIncwrIMqvY3d9iJiqJ2PrcJX
39U1M8zuZqc89q+JMCRa5BMC9A/2bl3EuxB58XfgS3IXB2OOvMpSUcNO8PFSBSnl
umV6G02b5xVBcUyNZSnR0NndrShChUJHP+sr76ltBFKC5fQ/O7ijLGX9lv+/SFls
o7nO8UK6DssLfiXQl/9F5h6pDqLeHkFI0A+71QMCNGCPqn6QOxX79cE0WEfJlCKb
Y3F4BCA76DwWOeEJNsiACXoQOnvpO9OqF883pjBJzt6M506l3zQ1p+oiWAeDD3KW
W03lrnSzs7WAkfvABot1W3Gspvp2F0AsOHEWYQLtMk2OVeKUYKxpy1CZJbIumsTh
U4mkzgZm7jDpHxzs8JiRteAoqpSI+fxejqG0bfnDtp7HRSBgwHyfeP0XO3i4NUmm
TrrlCr1sWMZ6zKNYVCFRl3BfvGtOcsL2sCvsbPc/pmi2f3Erx7Tec5zB5cjWmEk7
nSv6Zxl8wls6RLplp+rW8mPh1o50fy790Tfy3OXZbL0kVmOYgD3COz4iwC2VLtXX
uAwxHS8NntDvWf8iULcoYy4Jgh1W7BnpixeZ9wPYEg66felSe6Tb76B8TJXY5De+
jA9RNruEnXYYmN/VJKDrvMNxCVKIkGyPeTT6RTcKaz7DrnfWNeOxFAaQLfzPV2lh
Kzirfob8jPiQDJHhbAKHL6BCVP5slf8Mkeui0Dmgfd8M0RFIspiYGds9mo+Uki91
VopyjnI8qKuJX2nKSCdmniMbzeKpTdCzLISbdNqfME8sbrnNr0ChIlbNk+1Vv+KY
MT/WMOZp+6jSZS61fA6KNXbIOZGiOZIaOC/UNnWmYa5zHDx9sIWTtmwZNiuvb5pb
7QrkCrQkhwNSVYjZ7ybeVAzaDMVvgvOFZMGv+tWm3unPadxb9SW0IHuKPjlnJXE5
xhju9n9szUzrwEO3B6s2PIBiihT1ocTwtZgtOpGDInafWXvUHxvDldnd1cb+1y6/
K5ZrebxzCetK+SiPnVPNWW9QvvVqHV/nuG0VmdYaGX9vxJ8o3XlJOxv0NVoBLiDE
81KPphKwB7R/+9ky167uKtG6izc7ZGufQFL2X1F+VucsB6CUrl0O4Mh6mKCmQp1+
kxONl854FxvoVuu9668lk0PPGM0Go8WYyJVq9Ja3z0Nx0pvoBbPjvMRR5q48K8i7
pHhu4EffO5kWlufcrYRshf6NP8Ng/fVksJiONqJ0F/6ApXLMBEXP/SCBnkIWjWJN
Jsk0mW1BK3YfZIuk9lvf+0GOyVsgSw25yoQI0B9qOV8I0VJdeMnHccALuyXPCQDM
Ud6uk9Txp1vnQWpCUE5znMEt6pP9V7MN0MRZGmJmO+ikeAYz7odULT9vGDHozwzc
a3Ds7E+rsoIesIwSZiJC3zeUYDb3GTs06ECpdc2WxHw79w5AxJejh2fCUZ1+/Pi6
uYY9b3fRFIuWl8xmdfSZiD5oGuxV/1V0CHlbN5STlljotqdExUFhL6b1SHReFjug
i5yaY7apfo90DDk5p3SQXIkzhKSdUWKZ90z7r9U6kuxILoKAwOFJlBz1eYTNzOJY
y9HHBHnIxXSJ9fE5uBaJoJX1XiW8Bq2w9q9W7qL9/4RB2gjCyTsv2j9D26ruljM7
9Gp1IfqhRl/kEmAprwIdCfzEEJWga0GcxdIvpPEKkQL5+T9CjzlXnjC6HXUZ7Fpj
raKnTQhEO2LEsGdk+gD6gKhJq2jiBaHsbkUjIT+PBu9dY+UCLbs4/l3cX+lkQtTM
LTQlX0ObgMuFOUtt19vzltKM/1zeKDMvJg9sPMMx4mZrchbYCmDtz8t/RF/uXJPO
G183UR1/WOy4EB7toLeJ10OD4HO8byrzK1vbadss/E3Lmkb4XpCG4jpvTsqSBTe4
GrIjbwVDIdxQ7bU62G1k1tf+c1zuVd1Ig84kHowutuvYgMPc1qvvxCQK1FIMa8/t
nmGXiCj+cHBnZppvepJ64Q7lm+dDEo7YrSuBFQ4WSPEKunsxW9GqDtwXyIo8QXoW
fe9x7w/213XqRr9pQ6Kn2btRThSwb+SRkMvewZbdGFZanqQVE77LvUQ/2t/qESjO
C5nzbcUf0eCAzQNfh0T3FFk1V7wlSSmbl6bFA2U2uKmqZfZyUpDVCQuj7Oe66Bg0
olAvcpngWUqkQEcIb6XLtOkIlq2q7tzEDl6YoVUDNAw4y0ZOFDEMo86Hw1QaYYgi
CmLBRot8TOZtstvY1AUdwYejFuD7ciTT02h6v4Fw5H7E+QuLaqs45E/YKFNvhQ9p
7Jf2j2dkfMCKDEjCnmCbFyt9yZYFg+e1L+NGd+m8J2zQTvIvqUDtumrq6TSsl0g3
GJEdqt+5gKKLo2/usGwWfIBimnWQ1BrhRZhAg/hov23ZQbrif3qBmS5bPEvgYhSO
+68zxKVsGZblp2UrCtTG3mXe83Rri8khHXojdK1jw5X5EhYXe8hVBfUKH7IjMWCq
X98BT+/bIj/yt0askXVO+M6sDFyfqzLpOem7oi4faMIcW9ZVQRu4FoYYC8ajpwhE
669LFwZauivOIqTRuFvzQCu4niPgSdB47mNstBVevuZR4NUVSwPU/4A3pteSRuDp
oZUOfMObAGlN1QEzMXh28VTJdIo14Wsf8iITwmiUmkVr3zKFQbYkjdgRr3aKlrhK
VxohGGhkDZ9EtKRhg7bteleowCz8PD/Of2Gpt87QvQ1mBy8V6gkXfY3z/m2Z44Fb
7eNSTXdf7PSNlPRzVxRvy9GE8I8Yy3orSOxg3hyaoiXF3yNCtBWGNaMmR0IAVxPq
IGpzS7UG13UCjmiu+RqFXspbr/Q9pwiMk1lkyQw9AEymMR6lStIlum8rcyyRiWJD
AOf55k22oMzhsfKxPiIvj3/hSKFvE/gpDi+NLrvCCCAQTsrWnya7CkZravTHC4hj
dy5GiSQ+1cnPIB3fMXgRKpqr4csFGKAO+y+f63wGD1hEYhfR/6B0UkEHTMABMmtC
hkTl+G3hEmevtwW2lLDSpiSTK5Nx+6Yq0WvlOaPM1Cv3J3U4JwJxTe07gQSBHJ9n
8/oJqrhvWoTxOZOKi+l+oozqIP0E65xTT53hnT5/zMoky68P7Vypn4CZi4G5kOzm
j1VulO7EQcLEV+FClqwfZvHUHDFizXJmTgMcz81HwVy8tePpkH2//v2S5/lYLhtk
nFUbMQ/sKG8pzG3Jh1bg/Qjk7rc3Rd8nRSBZhKSKx2uw5LfIRkrPsAEQom+HpFcS
rOOadN9zD+j91RsrIx3tMlMkbdm+fgKP37NZTPMDlWY8mcw5X6DnjWrVro7OjLeH
kfoMCnX86PCMOo/oV2OYVgQIDwX2TmYHSE5KdFQCAnKT2kBt4evIJ6C7YIHDPMLt
bAWZ4fcgqB6MiKDObH/rJVsp9gbSR/W0O9w8dcGlBUGoysMI8ApCz0dVHqSXlWy/
ysihccSRBbvbo3KJesBInN2f6gSQUHlKqnlVJpDU+Mf+g7L9LLRYBa0JSC4iE6X0
v71W5XSPAHozpvpHYR9dZ/e1gW85I3yanZ7JxaIOQ+kVVSPb5A4lssOkqmod8o7W
5wC7tyVPKKxSY02KqU78ORbhwoV9cPqhaPgKl75KenqhWX4pa6Xa12LdeHRf4wto
otcuOG4amrvmzsqEKei34vHizU7+J4uAVRCLr4ZsMbNgTnXDfh1OIvWgkEFzcCiS
iaOz7UDK0qqOYR7F90kpe6srTXr7RSzEWt/qJjK/rMc6oqcpw6uDFRTO7i7zsRQz
QezdTo8yNZXtYI17WCLqxHCEqIqIXFWMRdAQfICgxfA6CArX59m+ozX3E/szoDlo
XXAOZPsLR9noOFc0QI4g8xe62ULZzBQeUb61ETi9idPaw29XA6APRyY/N0/YD/0B
R0/zz6Cd6A1q+KVybDkl+i/LRttCBFqoiFbWWImVfg7ZQOVktpt1KyearQeOrVY3
dx4KyVNOymqf50TBuQkg8d2w3hl2amI+iBAmtZwpSWdMWINcRCMNh5uCqEWOUna2
d/9BIjmFbP/VAOKx52HqyVBr4ZiuxTA8dk5zoFe16ceggkb6WjTRxOjDa+hqJR5d
txJ+JsBEacm6NiZMKCfnsHExNHjx1FCSDRN1uS29LqiCV4vmF8I3dRC4YKOC2eBF
/uAeMGHlbWUVZ6ypWbVN+DmB0SqQ7arHZc22wZIP/hQ1+d2oOV7b0uEsm3vukQ3R
XnHZtByjtX4rG47H9hZujCwwHov55pV4mo1UCI1tSvyjoac4PLDxdSMM1aqYIKHT
dePoqbUdTjv9Nmhe175Nl+OEeItYc4eVkCOt3jRZXsJU1nYL1Ygj9UaRQsZg6u56
dr79l4tDHujgP8R766expmY4/89o0siLPdi1nwA0dkjjnJ69KEjjZUShdA72fakJ
zbug9h9kxfoOHDZXvVbIuQJtyag8DYamWBCJLXChRH4CJLo36rlshGE+RR/Jo+9A
hu/EMCv949ILmoOWeIL+UPhshz7byKPNH5haRU+uAF3l477myiO76yn6q4PXo1Kv
rXKNS7YhmBWSMPlW+Oq/K8P4mOyAwmcWkvZ9N7noNMWW5GKQkwgUoJm4/4LmHeSR
OBSUpXThIcCFPHq7sjDG8SZYYNWQI+HyX2oej5WpVOGGVTDolNY/QAMKrSXQoTVE
o9ZsDDFwhFuw1IHjHadPIDtusQ5egg6G6gc7mhSjDJjiiDliDqK8b9LBeyzxqGph
YL+P4D0lqZOpBZN+6xrgo+DIHiSm17Y/ImYxT7F5G4IyZ+oHmBPcHwOY79mLFwFZ
cL3wCE0i+x6FerorIligAUgEDdnvpXXn60k0Zi2Yx/NRaeAV4QYJD3SiEI64PAnQ
XYCxsOUK+YA+lwJm+64Px3if1O3YyDG9TOAYQa3yRai7ZfZahV+DaU/025jMtx8g
7Xa0gdtk/AUcgswFLEx9EWWA6ws6ZRu7bv89hfyUrvA7nYM7xZmhdcjTNRVmpMma
7nVcyI3aFK5SL9J6rWThT6G0OkV9kwz3ugYdX6GFaVX2pqU0+a8TWjWfs691JzkN
2FpxwwU6a8eDdi+YqYvbe7eL2ycDoF47Uew/xsUvNgjHfEVoWXTSorKYnPAfHVSu
SKq8CC54B4H1V0v3//t42+EVRa9N1T9rwevqHANgxHmUI2yxQokJGqWpUCevNcFw
evVLFSzpkPEXS218E3/XZjbAnjTJhGgjR1KdyfzC7ebgFWfP8SVq6vzImc4ksJh3
XmGwr1HuvgpaXHE1OYpgHeDkZmiB8JXZF/xVP633+8LRN4XYhMCo5zPU51q8JENw
puhq5lXu+u88G7cIv3tv9DV14v+vbjCpd2jvki+8YZh/+m/POvMc8Spplo3H1G8k
5IRXQG1RUImrCsDHTs4xQysdRLKn/Xhr6F4cQK2nrX1t97RF6kRjpF99eqJ1slcw
TQrEdtA1va/hHmOkhrAae4L/owgPAT8uf5p+h4FM3WPHRjXaO3sb3iv+aBUqMHU1
eg40QCnB6AqwiXiKjKSaeSPCRf0uSdsDF9LS3xRiYghV4+JRrl0/HtUplK7kkLmf
SIevvhPafg90nu6DTGJPAtU8Rqc0pLVl3bwvcf36P3j3kWggG3N069JMQnyFi5uy
m77vDQxxwJx3ymZmZAudD2tHHnwhy5e0R8k8lRqMKMeEmIxk0FU20hR44FmQYcAT
SammXjhilxHnjADBDeZLjHmdYhQIPvL82RtsbIxEIOeVib3tm5XTikNmoklSotVU
jkUqEn0wB38esJMyVVbpVx6w/msOGX9zrNZk9+Ix8PRSHCUx+QXlwxEVy7D5/Bdn
cnoylTLbWDJt0A1aZzWxxcRKNkWr6584NCynBqQ6h3M155LUpXNr4tDtQBLNdh0Q
H4jow+1sCyAV5d03KgfLtxFWGynv0ssXMwhUndEKqTOL0it7k2YtPyWSn876t/ij
gj+PE2pecJsrBoVtLObeJnlq+dfwtiTDf1QZK39Bd1qGr1OTm1dZYjbkRpIQY9m6
9ftkVfWSzrQGCREcwkMPBVEL7LrAOG5aeLH8ieYIhdvT1VAZtCx4oG5kg4fAs2zR
kVqh8jyy6cqaXnVNkPh7wvO1yMA7R32f0Fdiy3gxN0IiOMXuIHnjxrOLOyYJ2ioF
q8p7rsOmOfbtMq8bb7S4tCP+SJGqQI2t5t6DoXuJZu7P7hxDG76eUz9ii40JWwjg
fZM4N9jelCATADG1BEfgf1L1CuDlZ4EsWG2wFiAXdx85y1tKC5RSBuZXNUNpk9kD
WUbMSsChUEVnMJwXGAVedUsIu1rVD9h0z8r8lk1qWE8CkbpgfF4Fcgtb168lH/pj
GVPAOLOkOY8a5Y+UVfz2NK8TovMZwAUea/r88VEUTCYSJk+xiRKhsZVVswnJPOB2
MMQGOaFr/3ZWX6e9Elzv5w/RUsxsJn+4FBlTFTrrWcVlKBckOobbqSW9RHsx/Hbi
x9Bfi+7yoyoop9UZDYWl640JaPOA9Is9B0TocjrDGfrLuf3HKeemINu4kVSnhaIk
WMxDjjUSv/uR/qO53uNQVWtBCbvLfFAg+1JlFvnFbGsh0c3VlTnLC5qm4D9Xr+bq
52lYKB1DaArvC62G3k/2eyGk7MTP29vVFjuCgpYwgYDyKLAr8tRoT0sKkxNiedHA
07ufHMVO56Ud3bxUCpPonidTDEXcX2vqDVKyUaFwaPvaYF9TVwFfHDJIoiUbpv6T
hGvIddLRvwpW6QiGKEy7OcPHbkckLxD/E78C2JBabvlwil7DX+zSTx7BYMOyWxAx
lNjyoiQFHtT/57XljJpf7t9bWRHVDCH/KRihnGzoRJgE7/pVCSnZRgysKKWrAl/s
iiYklpHdz97HjPPlWu19Mpl+t4e7z4g8cq7ZmR245OcfzpCJPvUT5d6ZkLYAZaCy
ilcE9yaHGMNmlPNWIvHJRh9qCp6flj24n4OXLtXUFNEJtGQQ3ozyGhE44SEsc/xJ
2tp24napvHehzE0sQNlA2yPXhQDVAXBYOk8BMx7ZHFf2KPDN61jnsH8x9LzdIbgj
tqgEs/ZCXPDb5/rbOXQWq/4iIIwDhbGU3LfPvThVDPTUWyLMYnX3oK9PAxkBZxY8
A3XFY65Qvwyw7eDyno6ZJ3H7s2D5/kZRRF+a0U1Y3nNvyqPWEot9cKXaHzWvz2Gq
xoVspuAT1sZ4hILeT6yFQtFEemEI8f6tUtymTUbun9tp4lb9ju3+A/N2jWOIBMMU
JQC5apl6YvmIv6XdU/rvVaCgzZ5W8uTiuQjBE/Y2I/UJzLEMZaHzmStkGRdOBgRl
YCSK8pElEAEi89xT7H63lIGcOEXwu0VLMUFO5caRzNKnMN8DXinKUbBeiLo+xGbN
Qd6GnvSdBB9jUbKAls5FEvHZwFVDr/m7ac7Lvx9EXU+xP6siIxLerk4kcSDJ+lDY
KreUSrb7D+SOoPh+/0YLc7Zxg8rqX3pky0LJTuu1EAsrY+relhNs2bptCsc1Ut9Y
XotAUkG9l50+yAgiTX/sMN+dxUpoLXDhmacbfp0zTpjpbepjHjhOlArjuHEt6eHk
RCH+7s1DW0ilxWI2nfZ2b9Dj+TZkwm+QFIMsC1vyIh/Z13m9uGY2L4sZlCdSYHuQ
dh2xnzBASAvHnWpiclgaoswrJZhPWt8f/s+DC7udpxetT6aJ206JPDu55jX5tAIC
5Esru+9co4fMLFPM5qUCKSLXmThduJJVl+YslxD6XenJNH7J8fblJ96aZ30R85kS
X0m3ks2V+zf/nFyMdfsQM1CpkXDUdg6HPqJQyCYzC51+yMWikafTV6ISeuiCUPsc
gnPkcYb/Dpc9ETQJqxO/fyD93r/KZOzhxBh/Eubs4Vr9dzhF71YoN78vJpBAGHg9
gcgA6W5HhCna++01lcxoswqj0HnmilpLJlr2PUvv/jQmNi4SHYRixcMG+K7wbL76
tPaK4WpIbMEzqO2HvVCIiYqSzTjpZjrtHJteTTZfCDjV6/U5c6tKkUe+0tvGwwZ/
VORG94y1v/Z48kw73EKdddu4qARzeaY5I4R4QgZxvZxvpQVCcLBf0bu9zRJJokIn
XGK4Cwh2nCJso5ls1iXCZlEP9y38TdKGlc9C4Hun1KJtt03M3gquItcINuQ+SCrE
5hyGbKA5mW2Lvp+SWmu4Xc8afO08xo/ylLFiRL1Jv6cmpYoVURQj+Kc5CQPTmXbh
b0fxVo9gD9cN1AC21SxDmgMnswdj/clB5mC0wu5O/yZmXaXln5mt/Mpr3kb4O17U
lkheWV/RNF+j7xb+DbYRDXUBROt2iB6R/EGewIxBpSPUjK2xOJGIOOg6tkEgdTw5
3CRbW5J1WaCykC/6fvHQ2jeyr1R+gdHI7toTpS6Fxx0OQM5vL0UekeqGRtKmrclZ
TZGxVfJzHNLURTbno2nYHLIyAfF0tDqBwlyj2pb2Au6Y2zP9saBEB8tIGT8AIKXe
1+aa7HyDU1oL85sDsGhz8ZGsGQchdpqra/wgrE18268VabXJ6Hv6aVd+R8mEyJ1K
UHsARDz1JPvxPAyYULXJWFEvuuJ5fhHzcmMPU/bkoWP96uwhRQzFWONjUFzLCAHk
8+5PfcFcB6B4bLhcrUJhqJDtftxCyS4/4ABzl1rnbh04gzH0T2lytQ55FV/V6/Ho
aA2x4k3f7LqUEwT8eCupE7U511MO3s/xXzoXj4YTi/BkZEzxlNJjJ1J6d5YfUlcY
hz3ZHCQM0TQstfpsv4/56Wa8TppAQOHEO8/PXvDoAR9Yl8oQ/BaWMe2irH5EwWWe
eGGfteg3E2kOTOL7LKaZicgEYC740tth7fg4ZWm/OlGMPj5V3JiKtJ50aUW2oqbZ
k4QAQMAdo7Ox/OEoISJHiscpUZb623/eOu3Dj5Sk3RvmeLnQmoI7P/XlJwRk2PqW
TN+wza+WD7AXs1LIv7IrDndEi3inIpAeapderOs3L60gHlKle0AU7DfG/PPdA1CU
GxdNKMgoKGJi7Wp9UV7UY/93mk323UTBElJiOvbOTRUEWWYKEn5TVOw0Wx5PcByw
e0FKI9SdMW26Q6hGwtSL3c6hGqrD01bpEhvK7SbY1aWyd7CvRm60MR63mKJvRcL+
DfEruqXo9N3HNP/hvYjqhb58BEghP39tjKsXJNGuA6RVjDy/5F1sVnrZDR9DYtHJ
0n/0XiEpQT+eH8dH4jIlPCQphXR38PIxJnACLHLzvcdZvPv4pk6RFsXO8k5VFVvJ
WkDBDq9XWxOEILOYU6zHypxeg7/byWKkhasfGQN2fdwHBjdJNxuwITK9ZLhNmko8
Y0du14CqeK7IQ9UHfPeDLnE7jGSbZzPbJvLTXKyzKLRWqXxdT2JC9Epp38s0rKtU
Dk2eldFx4PSGKFF9caHh2C457R14MQ5BEc+Igx5vLtNfTtNTasBj7J6Mu+ivft8J
ULb0fPyKcqqL0VuAVoK8KOanPA1UTcH09KlN+SXFIzu+C3YOIZj3kAmrE7CDnLzQ
7ekXxfh40omBdDDLcW9fbMjkNhX8Uh5R8euexPeWPeXNXADtoHV+PvXILVgm74Xd
SqDI5OEin6vyQbkS7rAvPe+sZzNK6xTOz1nIIP9YyB5hXLLVTL+PAD1Z0N/Qyz9u
wpvJPiZ/ZF3AgMwezDngA0PEYHBgQB5aINzRTmbibXNuavFMKHmOCgQhkN0hPDr7
6c0w9CKmNnjHnFK/SZWikYUVjfJcRHLbeWKzGWOhjt7JNCJqfYVkenV03mjQ4UHb
x9RAq1YZRr6WW/fMvFgVmw6YbV0Rj9vvxHypdb3ycAH8RV8qXmL6wmBFAii91ueH
Lv97VHpWi90UXTZsEPfACO7B1IdMA+siyOAc9hvz4T3+QENPoZbvwv8W4s1rhfwy
fTuJFNJxPLCQYHy/8kl8sdDBniC891qvKrjNIGJ1KKSqFo40cM3dYIJRhLHlTDpa
lEZsYnYyHaldufTLfAmELKU+vzaXz0PRlJH8mQJAoUQtxfQRMChnzZdPZRFpZ26o
e2z1Ocr4yPRmEPv7ONGtqFiaHVlnXJkNwbt5nU0BM4VGUze1l6a4Hkqf+9q1/zfY
cO9yxmmvByuvI7wvvFtDSwhn+5JTRT4AG6WmEfpC8zf35OaBTeJNH2gf/F9YsCmh
Jx7S7P/HYbM+uq6qzl5BfufTfH8OipZ8n0uzxPOHVwjE4rbi8Rc7M+0tzXP7rle/
P1fo1ryXhq5skAi1ZZVR7BWJYMEo0uJE5AJiIyfg59uxkbqYcLfJE4xVd3wP0+lt
SYRqZLO9lbVrOuE4wkNI8H763+u2UmXJYasasboSnYIjtjzjV9RpcT8OLHBy2xvH
/9gFZ0hJe1zVZyFosKFGty9fCXl/emmj57vzGgpv5YpXp/gDJd1c4MgaBHTJxa8k
c6uOy+8QnU4v/Z5G0Xj5mZGK42BKlLYuQPlNed0ShxOcsB8tJqnjjRI8rholcI1e
IGDhPHubn0ySjweJLrG7o6+yzxCGfZ7Pn3Oigm3MyZDuOh3gGPgubWSdc7EIatzs
ohL/qjsKVgEE9+lIy6M33G9f4fVt2nrhqrOT07P83co1hMgxhGOKCmTuVijMyIHb
/6w8rHPpJsldNRy2FvkmWkcg9pRBQNfmtSah7lfgKdpenqiTNTy8y/C1jwCkntQK
8CddiHF3lBA3dtgxsDsmhtdzhVIqzAy2jfThi5IL5wRASD5dm5jxd1hor7NfEEjK
Or3gEM6kgScS6atiTedox9CcHTm3lNAF1eeWLXQEghI9idJfc5HhSXpePT4QGaxe
/hqgLf+P3SB6MGe8/bcV0IYrZWj/ZXbWLoOvRE0PBVy2wGwbcJekrrUCgDyp9RBC
7/X/VaTS1+OrVxTuxmvZddN68Kl0W7oQSgwYXTVs4dQq3i/ojUmmMID35+XB2mwk
+3Q2OZok9lK+tLG//iPp66ORjh+gH8mezKZ00Hl0MgVxqPgEprzKLD1DoMjeMPWG
EACinVwIhBOUqCYt6DA5u3Hh74GJNTPgncenSAO398HGk6epNCECjNG/wrUsOVH/
z0BHzh95nQRn4bOxPqjVfp4OPPWZnYnajIvPN6wo7Lz5l4HtkquphkdguSQd/S9l
0JCZUptBzccDnM1diGUaOiN9Dg2+dWIMZEnhLCzrnovdaXYADCCFeRx3HFX+AVeX
iiv8Y+brc5XZ/mCTOOxZ26kMbsPqSu2RZaaF5ZY4b9yf2Q2D4H9M8IJjOY+1TaP6
aC1gTZRsHsz1CgAguOTHZWo/d64goQgfGwUuLT9Pzl2oWbjADitmwmUqXjtIuqGb
qGDx6Oib4ZmH5X3n5F6BcWcVanPd837RdJgfAuwFo3BvrVFya9TyCfnBJPPWeswZ
SO1HZy/o4S2m+lUPDKphT9jak2+BaaX59a6/d/ZWuW8LTVJkcbA38lrnqhKgtW5i
Keuq7z0kNHt1Sx42A9IUyBhF2umyLhFmgOZcKnResJGkXafkn9AfdecZnc02vv5F
SXWtBGwHkPdjpVbygTQsrv0e6uWGgs9CQI3IF13NR1+PCRkZjzHXgC7Jw9RfE/Uv
DNHge2eWJ9wmGyQFkPjpoWo1SOk/4nfndBWAEK6qsmlALLPSA5yWyQpC5aF4d4s6
PhOAIkAy/teJdp6BTFL5iI1CtO2jjCl6R9EyRYMKNLiMc3a92UJvZYVUv6iN5gHv
JDnnqtyM4fG24gV0MQLkmVLYGizo/oFhZOcX/PM7oOynJkF1DERWBJXgquiwIiRB
LbeU8kz8czazrTLRyqXx8WyC7UtDaWWcDA80cV9teQQFd6pUbHooBaG5mscqKVrg
HyPq/YBnDvE53C/HuOLWxTKABw0pzSF2SaJYLG01Nhb1Zh4ipJt6xA/++lTahfNn
IiX+MbLEGHMGlgdVF1rKYk5CfnNYaiRjZ8M4hDzci5clCt8cSlSK1EHpo+vl2saD
bHreOJVQs+5XxhFbmrC12eE0VITc3ZrUhpqVeWR4ykyR1n+jT2kLevNvs0PqKvNo
kwLln7kocQN/DzvlCJb5OTG2BD3Sn552wj9wqkYJ8QbVOhItJqm4YWhApkAtpI90
+p2Hs3uzynTT2Y1yK0g+a/6IF6cjPDbDNpMEfdmv56+CBzPOhQSm3dGArnMkj1Jw
O0aoLVKC6g9vBZsmlfj/+53rnrclk5dR6P0GJhmhU+U0wSeGmx8W+gS7wH+PQRYE
K/GF7CQ/D1ca1MKSPFzE3Rq/ZOzXbcbCPe2EWOPI+D6lVC72QR14IRk+FIILhWE4
ZRDI4ytJAQqKeu0D8VqSnxwfUoClWlq5Bwiip1FN7i7+v1gELQAFzWmYdMNv4nou
DizIPVZNUEZ3IA1rnATlZPQ5Wbhp6/rrBD7Vf3QX5on+m8X/u3yJEgy6JPHZvKVX
8XZb10QACRVLxsEctPx8Qn7G3ALdN/a88f6VaPMm7Z2+i9eQjj0hxah28r7kbtdD
16xvKzn/2jEnaPfE4KT1C06aYOZzStcsTsy3R5MZiCGyWJngurqXS3AK30wSCfpe
2J2BQVcoX1WnS6QODjYymHal8Sj5j6Yh4vMqA3tTiSvo8StLQDC5MimCAY/gDLfz
nRqfbDjA4aOWaHt8RY6Z7oOND80qzx+dozxtQhU8KLxW4CHs3PM4BWbe3DWsprhv
rOJ7txm1+NQpBhufDAsiNW+e9BYTTUjbWyGUUUY2911iMcJQvc/pp0+3yk3+ynvr
cJPfqY59Rt0b36VUHOQuPVplZy91d3nxvGyB6CQS5lE6gUYzkCBGzfx/JLSm5BjX
hlrX1mn0m5elE7xUzmbKcm4aZGaCpUbRyzQeQMysPDLtv4hgnONMVHzxmgS2x+2Z
a8+xfsWhkjnQb25aOcVcpMFz7YvYVAwSbV9oylkQTyDKwsoPDYmT/44/vZ99h04S
3OP38NBD/QadwN5Vvc0trN3d881TcgEL2xzaZ76q9ptKqLx3Vhq2ZvEekz31gynM
avIMqR7NUHXTvXQjQvc98FeumpmFgOzwTUR/u3ruwEfD0cET2b84nW3vfXAz7U9i
Di5lLIB9KvqbJwC80eUxfFuOjPP51ZucmL/PF55+jFadOU//JyFSADOn+y5q2otd
ShY4GggNEhHBDK28WlukDovDOdemEIgvNbA6jTCsgTzyh963D2PNSZFtCNRFVV4b
mfTa5vCkMKzQ9bcEPYWT66/s2kmSrcY1f+3PLStu//ETnbYswb4lMK24kReGX7Ii
AxAznSs2BoSWP4lx8UNCXhaO51vXlADZXRO9b0TG4klix8TXd71lynU2y44NBDqG
XXWaamsESILM9SEn2NdCHagITNjd8v5Q0vfRKX3N0oKOQ0CSzSQkgHZFbz4qi4pe
agm9EqjgryFoN603V3NSkCXQ1axu0ImcxX+/P6A1c66WvISlDbLOKgjsmBTN/86Q
1FnGRPwhAebskzxy59BJ6zoBE2tpgPLMt0OODQfm/aNYrijyP3mrz5DW0VsvCJRD
CXpruer8+8uQipwSpUlIingjeuy5f9IrNsiUc+/Yw6I9MBNNMofxtLg/wXNAZAVF
hBvwZP8sWYStDpWRYQtD6vpSieh5aDvJFH2ENyTqg9YG2L2rJjJZMCgv/EYU/A08
Fvj95fM0KbrxRuiNifS+qFUwP/e2MQneDSKx95qdcKn6wPSLALOI+3VIlMVE1OzU
U8GhxEomtqOGHkooh2fhRUIRKDWm9PUq3m7BHTzDsG9RMenKDPwqUMRhw6yXSELu
mXiWJ+v9C+NhfTuncu/MxaKv9bi8tv3+ymjiudXK1pgJUWch9K72RfWfHAHM6+6d
6XE+LiGpBhvsKqcFFUWG9g9NU1yPIIDtuPx8FGXFAMTPQ9c2a8nTraohsJVV12Tu
c9cKYJwG042FP27cjdUsCSMs10ZrMrs1MVISSdVYoVrLBdOAVA2MAUfW1uktqi3V
L+GHJQ5ertmNSBrWsPn5xbSprxDrZZM5z4XK+MWq+YXUSFQWZr6Ad8+WDKzkKxeV
hZXHjUgBmR0fZNh+BvaUTIs/AG7PMw898HQQSC99ATJqoQXhaZ9e20BLFAfWFR9c
kNaR5ecUE4aOkiwR7p2cdjcNBKSnRsStQBzGzS1ZglM6b2Blh8M5DofaTdubMTdQ
M0QV7pU6cNffJXQAtriE/a38pZEWOUmJep4wouNbCxjczxzmUaiOeyvm6ZjhTM/Y
9nwuVwTshZ1FqCa3TFSiQUAp3VL70DrWhhi5+++YHRFR8l4x6+CCCB2xOSe42FNX
ErGhmNLuKS4RzMv9jbev1DIrc9dc9TLfcFC1Ct61Dy1scCEYPCYjeG50huT3D/Ob
9mZS4ZcZ81AGKsOh6zj7YqQO7NuRMAxe+BH+9f4QOQFmD868d2mGDcLYZ+IUuSFf
QmaQfOY7DqaMgoQ2Ht4WtKVYSf/fma94QBuYV1WDL7ZUL8xO/8Ujc40cbrzPClHu
+I3VcIz1ewM8XrVwZtTUrDE7b45dpHo7hD5N7QP9x1CqgafI92+03bcm7PeUXHZL
VUhqHZYh0DDKLlgScBucH9VpbeKatP/A01WS9H8eMzxxHutLqaTxNLKiRrqjiwV2
7fMtDG6Zv2JIsaHTf9GJzF0WZqUFaUHNtX1Viyeo4N6wDxss0BFcIuY158dWwtwH
GXjecglP1W3RHySVC7AZZVgXZNtqRRcN8iNcXxDtctcviPlO7B19MCabCjEDh+8T
7jqksh4g19Mum9bDhGLIFIX3pswbuLN/o6Dy8GIYUrTGeDQskLh92SLj6nIxRC5D
d+MwpDGmGdl0tAeGTymM20bJdJrzxwy+F/0khuPJ4wOjB0NTFWYUxPNMgd4vJypt
crbQACvu/1xBEi02RReAg19FHf1BI1IOUt+Z/96Xw2mXIgYISaPy07F9eefQ8j3Z
c5XS/NtudbvbUETZ0QBnOeME90pDmpVtuffWzIrtjrMpDwYMNIhFkcTfG3eThZsB
U5JDnlpXzdwPcxXSEjzdHMzWYuj29Mjmyr9jJbrCskB8yi2blCCnzfjENXDEi6VT
wn2hXyikQWWBDRi0sKflM6fAFtKXvsAppWBHhQkypbsALAh2c1kBjxiadgj79Tru
Kf/b2H3S4dOqhR8jNOMrPZLi1RsKVoEDYTG1u7Lf+JRecYaxgGZP4Ep6EpE0lDDD
emqep2ZyMyWyJLwvl+8xEKqxEhNBEGPMjWiJD9o5ddv6XnRvPu+W8QpMW+1Q1bkQ
IBrBRnqE9oDJx++kl39FoJvDLFCH/YrMgLSYz2PJpb/FLHPNERnN1wTEVx/MaGYM
C16SX+i8Imnz5UdaFW71XAwrafnR6/ISSL4kx+qT7lTdzfaJfC/jKJ9J4QrbVU9z
tMC6umtRJc6sbbRzDxPWax8ny6rmc6SqDS/OrHPCqUQ+10Lo5RQh7xbmB6nwy3lG
T6YC50cTQOlwksGODXGC17Xv/iBU/1aS7iQTPzg1bvpvavs5ZEM6zuxI5HvAVMkl
0fi5nNFNb4jhq41PWLsnJu1/5IDPhxyVN5JXGB9dyjwpGO0SVUvw4+qhDOE26VN8
rgEK1OsQxeAjjMEqPNyAW7PuTmabat12BMVhZDv2foVQXch083qqu7IbJxyGauks
zdsaCDxQKOXeMQQZQ8qNO92UY9tfmqxhQtn4WY+uQTw1VJvwO1zbgyr9dbutybtB
okDm7EEusrJG6CtWHn6KTDYQiVain7z5HyGUD4YKZcLrFqZqJZmoZseKb1FFq45d
oKrX2LHeI8oMYbboNcJv1vV5k1ZwOMXaIjiJq+YEtrC2nugTrmwJs7spOCP2rswa
Fdmhwlanan8IljhdRiXLmmpMQsXPfg4q6HeVe5Wy0CkXsoOPa+0xGnqCfqnp4nf/
FuAc6bfSol2gQRz43Hj1ljOMRf0QmQNnMQqgKCKRKgnBnWEMOOLa6P05PNXZN298
3exdgTmZg/1snL+86pQh8fxtHjDLhEcbXYJXUDOcAtqTpJ49LDG0tAVOW770T+Yx
x+Qg1EtcdSGNUTNkDvO41xzuqj9WmWNaBuLDzxrgwalfwgOYPmfefbTA3305QpIj
rqd6oBzeP/pE8KxNL83SfyEWGFFiMq+xtFzL/zIspH84D3VzavgelJ27uBnWFx2W
08viSPp4AWUgs36zLNZrvyB16TfvCHESiPAm9KMD5OHj1Y3V9YU4l1GxaV95hStD
N20Rii4Sijph3zBCBc+If5GYpDITC7G52CqEmEiLIlaoNocVwkG0o2dSYGH10blw
Xu0pz7wuZv5tO5dwjXXYNeSH4mqIdZVX/9GYEwmWQtm+N41/xujsCymT/NEIKkut
TuAJBjsDt4YXHJKuoy1sfq5JoWE1alj/YMxRxwA4rE9qCv/9zb0QNCDiVCqHSBwm
b4gA4JI/9PgOongU4iJ1JU2qQ7T8Xm8U6wQP0BQ5lbbwBUkNBR73GhkXHngnmcy4
rtFLOy0TAXWhUNbcRoFx6LY5IDb8FjRXzRqMpEhQk40f4WDfm9tCKTjsmNlpwPY4
eFo5Dq3ljXObMkSaweo9yoo+pOZNFFkvrt8FSnvb5HDoarBCdEJvLuRzjoi7Lmhb
oXtb6QiW0BjlQSVkFbax8m2aCMKpRqYh91vuSprdz0myPGoIqTSHcCNlhghy8Dfu
VXNMRJjMREzNdvlTtcN9kEm2KwFwrzNXwCSrgC5/zX6e0KSkPEDZncQLDop/IiRr
OSv3sgU4NrOXBRpJumjgH96AgXbwxW3aPc1asn289HD3ofNAPLGZtE4PjeFHamvu
3xDpgjNgKt+CCAFHou7qMvd5m6TtWMRUUmZMb7HRSiXa8mQM9VhE1iTDKSnHFOg/
htONYhJrtKm76Gtcp0qO+n13aWwIfn+TrRrNq4LiVys++SpkS4UkxxR5L+clUSce
VBu+O5SQeR+yvuM5Jk+Ux8KCs3pBGzdqwv1zJN9wJDKO7jnaPZQPT7t5KuBqwL7o
IhmJGnXbyyZS1Sr4yltikzAaWdJp1TkwGX8+0D9fcjb5vH3/r16Q0lDrVubHsCSK
tIdnrkr72anQeJpiY/KrAEpdQmkouZxCGvSOsykChuBgIyJG/9ProeqohJK4aU4M
FEztvF6S4etoJL+XllF3FtjGH1GffyyPmKLQasZiVMbAGKfZB9k8LtuZUMx6v9C5
w2qBrpZZxGPl0zCyCCo4uHneTwYWuX9kD33k/TJdq5dJoKCvUCG99jKOG9t1uYMy
1ghBEBJMSGeSBszAQCDLNSwz8G/zTwWbkr9AFB4DTl9zvFvrO7od66+GDFHX1WgO
H1wZ5RG3w4K4Kxfm0xsgfModcuPIgsBTkZXi+bYVrUIF6r5bX4ddvnnzQefvVtUa
NFZvTaxtI78FXFbGsdZ6Stfw3+7oGtSBN/cmPUrtQhPEZPIyhNB+7moQ+7vvGzKm
23OSmQO1CyeVHZt9/alPhUeQjrhYjYImrCkWuu1NtH818Cg0Xmq23vvty73nDb+e
w0GJjiEdWMG2eivXav3HykLlKoZqIKR9oRu3DDCb8tdyUuoy1WzUUUFQd47a848r
gRxQmRjzYxWbGySK3Q5YpKKaLJlKLNM5Bru2pB8ZcoSReqYI6cdJv33Dilp+LnoO
JnzeBaqZNVYq+1fY6jbDhS+33MuwxLxGlxCENPPMMGMI/Q1vsFYfn+WarEin+jRe
D36qVYxkzSgLgBjkaYBCYQRTLACWyKPLQnYRiSiEq2YaYdsuhb5jqt+n8whwYKdl
d40cf4v9LnGhtWZYBVNr1x/hbCXW7pr0t6mnvYJVjS83P1v6Jig7BnZV8/V5GJCd
xSDkPUhERYc1nCTdnHgjJthQoKOpZMFQbTzqr75sKpe0M/6RGx+Sck/AsjzQUZuh
dsidLVkSTIHhfN64jgvN/5DXyJBUKTL45b8JuovNqk979ZVAbUmZi/m8K7JPg3vw
kbCZiMcYk3oL6Yeuz7VVcEQd01vMiYA38QfwZHxjqil63NWyHPS+BGVE27MaSnxa
bfNkWUM3R9jaPsyQDW+zQiVZQ0zyQKFns2CiRSRfWaKNjyD8wxiK9wpfm+nuM0JR
m7bi+0KPmRi6Kg+u7zYU0HC0tqxAvcxE5DvzCthLsp3kkQfJI35Nrv6jYK4vqbEd
w74khJhh8E7z6ndOQTUUlKgOLLJ0+1zJWpboZemATokhq16xp0zN0GnRB3mc8xFP
to2zAZbkn7wfuPqCWMEMz4jNeNlzc348oPY+fRSQI8o50Wb004r2emG9kxb5G8WH
B/ZgbzXcjXhHuXwUGdOvZMOzbUM3YCqvPViRG2B9ut0oRE8RCPIlUzaPTcEDoUa5
NA4AJJNPBPht+IDWgX3lPHCy564tFD+vX26yTKE1sq1bhRMTafjF1cD42Etd1/os
cURy4+b4ufnbx3ryBuBTSIBKcbx1AFFP3V3sl9xLzZaazUDkBnLjpY3DVdjNH3OU
qHUvkl/WG7Mu9Qn61DEyQ4TYUwKuT+JctLOQbD/BPGGle4iK0cq3SjM5u7/+mOPe
utX0/D2np4RTDftP3U2/hYyR7BLnmiS1vAT5gLEIdidBnijw4Bm0P4MTNDyOiwiS
q6c+sJcStCF7/IQf7+c1Dy9YbuK3HTtIVlCrd2ud0hAPS+zs4Hpzz+r5/9obC3p2
pp8IaP13G+NILq/WNUATgg2hp4Qzb/NN9W9duVEH4iRp60jufk9J75c9kEL7F0Zx
NiC8gdzwR6s4Nmg1K8BgkOdPYGF8aAjbBmSV09iI2RcKxERjfZeiHOtkcTU+Eb2M
WAmiw9n3WH+dcCokFMM9GQyoYMEJVDRRwFRuESU8E3ol4A5GvqHiqfTUDmYYRXk3
IgDd/aLGD3nCmZbEKRuvl/9WGrmxJnfUqOwgmhekmo9bKRgqIO5rzH1/UijNe1wO
xCdfWbG3Al/GjBivJGvdL7Vc2nqsYNIdqYwe/D8hEbRcMf+EKqyjZXzk7Tflq1sr
e47FGj0a56mv+4P7/1lgnC9PtMC3c5itf89QDO9DW8/JFT7ataa0BzAAUyrGGiuW
wlfwDq4CuFvexDugkDVLOYtmg6oimdpZ7ZUlOUXl4OcZQg5OdBrvqxhGEnNzUh50
Rg0LZqQzWUrp0LhsHJwmnsfPBULyGYYh97jeQTGQvKSmukudKRIhMrOZbpTjEEU7
lJkNIlBx/z6hQHC/V2Tw6G4CBC1B0jsBD7+Eim4D4xuc7qWTQjCSGPrY7pmMt8o1
lxWp8zxsvnZCVBpifnWDjJyqc+/W79ZpriUoPx2LntqjFCQT969OWzSAJ7+66f8v
Mr+EdYOiQEZi0fO/PMZDnLx55YfJpDhFJWUVCNBCsN1xTOelVpayLcdqia21CbrT
sWdBen20iLYrvwSLHGnX1W6mFjbhQJwjZEIa7pSRhldySTfS8F0QgFiKD6hYPPFu
/eN3M3ci1Ao0M6OG2v6i2RwmDBB4exwbOfCAQsqLIQWbnzoLXuqYvrSGb12qRoHr
I/bKU645Mv+ZfAMduzVFBKDBm4uufT0B0obyNAAjuP8K6d6THl8WKqoPrJKNwdUk
9QDtgegT2sS249VX8oSNmck/W4hCdJVvufw5iwdxULLT4xRksCNBLeOLbkGN7sLV
1xrFHBjgaEE1JDGiJhOmUXxTMFFsywR038hCDKZSTFZmSkOlUUAMuxypklyjLzvN
BPrDboq5Qvx93fzYxT+cBC9neZ5fP5fU9rhMOSXoG9G+HuWHerC0CISX4YYgAq2c
p1Sitd2cu0WOTr5wWB/X6gaSeR9rk6LXLraUOZQsw8IdCakmx3Z3cvpcFZNlCqTU
7ys8X1UkXOV4Eeogg12jGhrToEIMJaGE7/vFiUm53g2kewGo4NfYSpFfkyClOI5v
O7WlxcVPip5HwAaggZtfeT3YCrI6jIob5twnwkPT5ft0CYaj8YWz6+ce/u+0Vc8i
eltjbvFim9HDJVG10mEc1RT0l7gFOEkgAwqyP1k0lq0MZqb0hIULMiwHJf3TSACy
N1g3eNWn+Rp88HGS4azHCc+VBEmphTjq2ybPebWhIZn5WsY1Qu7QG0hV7Ol6+n3n
QhrrQ2wmmY5qDeShYoyhoe1ZyU57Qx0at3SxB7w8G3K7NS7X8fT0gXtoghOYcptB
3J7jkX7Pi59x89oV+okSArRa790lt8uH65JZ2ubdXPBoN3muad7Naz7yYfx6xCFq
YVw/L8oWqbdHPyEoJ36xbzUtOJhi+9WWj+j/Uh6f31uplG/4DIFZFgs010wmr2MX
Rd467n2oWmyzBMLYypoKDD+DiwzqqOH1IRyyaMuJHejY4p6qvKHazPMW29PWaBI9
KTuIIivbqwHSQtgtegHEB1Jm6DpAwZSrAb11OJhr9WHlOP6Z196ca1QRNidyjZLI
lhEAXEzt3ib59cBB7wdqAyUDuOGiiLXMfL6L0HZ/sVw5hzKe+Ezi4u78Auk304vY
AkbRLAzL14u7lQfc3aVXtXKLQp+MvqTZ8QCzP7YrqlUXPgFihBO6Z6YMD6bjL59K
wvUltllaYNufQ2yEMSZuSlSQtuG1On3T1uG98ADfZ7GvmRLt4NpnIRt/xaESNyB0
1tC1CUJkCAjnTUrJbnhKSJ7V0aAD4Wtc7d5iNgqtcv0vehZN3UIDi0g73IXPqapt
Cnyyqq3/GVSc/Cx8kBzb5mDxkkG+pAaFV6g7YbpF0MNZyLRioUgRnj0vZfMPcn3A
quiTjKzTqJuQKl3qeq6nX+onXIckKp9xxhxztMiSnUizWtKv9mtLUP7TxO6YAz65
EykIDBpl3Y7gfHuVILqkTkC/g0UucvTI78Y2XfszhifUTtHrW2fJO1MNbJ+eLyvt
xLHx9cKp67C2SSYwP4EkOtjWj4PUTl2TAKAWmnxKfGMt251cNtu7bfbYxrNMW5ze
djNeD9lxIAjhClacBs+d0XR1s207MCS2XOtWVO8Mpp7Op/wlDclRCMpjUrKaq6SY
yLcleeTMoT3REFRuqLnwn2AH1TWhw441XcsnQMhJLVZ+iVtNQVcd58xvwNYPPWFs
aVL6ttqiqjsJSvbK4L3m3DBgu23t64e1tEJkIDa8fkdhSDmBMNZIRFLQvoU5oPEH
TfnzzhFC1woCYu2NpCM0mwGgmVGYJJIal23N2KaNsvk3Rj+sky9Fz/c3if5p54xz
YOXEnm5uZuog2iBTl6kJrNoEdAgOJlx5xHWxTesz4CRUIvJ2mosNnVVZxdEKVEE2
WfWPV5LAS2YbFPcmCGAzoWxnhfgiMVp12z2u7XZeSoMFPh7OY6O4+PGoX+/0yQ5Q
A8hw2H1S3+ParYPTC7YmYJdlL4aQil9/Gri10PtZnhhk/hsBVg6ylRaKOJ1eUcbF
XmuVjA9HFsJsEqtpFr1T1kit2hhNVEU94WdQ6LEjYkU3fgC31vK/kGJdSZC0XKI1
1WsGYeluNhwVG2uhKbMCygQuSHhptxGedrFQ5aLM5a+FvIlDQsHztlOHAGMo3xuv
pC+W2435qBRe8LA1mD8OvHNQK9ipobB5hZrVe6JuGBW0rzVTRLu58SNBQTbviB94
WIO/gO8nu8BFphXelb3aERqNt54ctAst1atIapPDo98TjA9L39Ov2EcmLEbwQZ/c
xO6pWnryQlRv6Xf7+DdPA9ZfU126SBg8YuK65cBLSsjMgin74Il6U6yGI2K4rByc
wy+YfzJfibz7sp8IgGDfmqjmqFWRvnXPm/15DgLxcxD1cFbeBmzpRPsWZF253slm
KtXSzRDQdo2z6RcryEnyiYtUAENId30dV/xqpG0l3q29XfyDYFAbj+t74SuLeWhu
06JYY/eOE1QRbPExINgMjUHWYuc6b13S81QQ5YeAuqFUz0RYDPlj9sSLP+ugZrmg
OQLmFUpTEK1k9IxseIo6FfJu0Yv5glEHoIhwhypFQM4TvU9ut64s03U/vJ4MW/9L
wHHZZwdhIw3glsA5IL8H+s4sRcC1BgMO7SFxoPVueFGiggLviwVVUowjZuju3UVK
UxUIPCYeHRfrj4rXz1FfDLAyx4iLvaSUxacFSCwqPr47sWyRXyhmPRbXdDKDaDzN
xSQDyzqq4hZyw26SHK9a3+Dyu3abyrDBBbPZwBjeem00X37EhS35Nz73XGc2PrgW
QtuFo914xadeL5TCed3l4QNe5i2miaIFCOCUCzksEb5iOK3pJizdzLQar12EsXP8
+z2/gQOLZ/0WrckkU3ii/jX0ta/64ADYaDt/vKneq83Rs84ziPITbG0zFBDz6xyk
jgafVk6oASaWTUm2IrtLcH0V7C2qh0Y+35f6ZwFdKTjMu9xx4IrO/S/XVI1AUssN
a49+hZseRa0KB9pp94Dagw2AJPZM9WFCZHnwGAxalkA/FJRKzQV0ktKabDOtNgzd
u2hRGDFTwQJchsRQKpfgcgYLOWR93tGRsFlPbX8LYRaO81ytaJ3r6hkUhPT/Bv2k
xmon4OVZIK6E5Cin3tR7/uPt2CyhsPD8MdRe17T+ANMQ/bu0qdBXnYts24HBKqOf
3XXYYXJ618d/RO7yrWHFnraZ7rMqnUEKJ7+szOigtJfKBm51ykGvPhkjR4bkFquH
mw1RPWsYzC+KV/3w1osAlg1Usq6fH+Com9DULDxh1F+9QF9jNW/UbysKzwcAN5IR
uSeciFmSPpkW/8jQ/jfFcRVf88ged1XAE1Or0AUYwbYHcrMrYjELA/PeXNHEnqtk
5mS5NUbRpxJfE0NqJsvp8uYkgT6zRLuDDmTcajGvnAOdJWZyEmDjYK88f6/ttF7M
PFjiwCMIllHhmks3hu9m2PXerQpTSq048ml94qsUcPAyQEbEOqR79n2ZnbE+TCvJ
LaZ3t+aExl7k02OhnfiEddM8ZvG68Mdmv7aQuexTps9ozyQw66/GFXO9bFuWfkha
8PwTRCtIkK8Q0AJAUiBNybDykDj6Xj6mdvwF3EcZvyvbwxzM/mkN37jSyooroOO4
os68rgk1ym6GqEhMqV0LBBUT9vuXUNtIeiCtJ8gFgUZqwv51LnknTjAKDR6GAhQO
WDXRQ/81N8g/SuCGwB7UjbPtYlnflfyNj9otLAcGg9uLMz2Pm6sGnEIXvqlOzNex
zdOGv94CLS9cjOLDDneTQ+R3jSoa+Fs7+c7faCbXEBtdyiGjhw40WNUAqkJf/Guy
lvEIvqxY3XviZjjHZHc5Pa0/i4+sdRBmMYY4J9WuucAY8Qe3FllNBTCrnpcBDG+4
jkRSeQX374sx2pHCj1kBcbQbxgpVqkaU+Ry1ASG0mFXWCHa2xrhmkAt2KnXSlqbL
3frvWvGSPlj6q1EGNH3qnAxXH89OsjqFJ0IjTZxtIFYIQvbbz9NI+BgPUV9p+iG3
dyLmtiVWh0RKutcU6j3zTQKfWTbDjAuTtYIAszfSaunxaVqTxDmZPkbC6Zsi6vce
saRsDvQIEXJQ3fW0r6c5vTkU8ieyIFQRzxpVOTmJdVg1efER2gJBAkEmcZeamNTt
CfCjSn41H1Xa9Cz9BOZzGfH4/4mGaSQXrqG7R1E1Sp6BFcfOhx0FgpAnxdHyYAjk
FSdRQDyvliD3QI818qU5eX6jfRWOP5cP3R3Emg7APLR+4UFT8I8NV/lE9Z49EdJ7
K9PPTOU1/x8nRwWFg4nUFusi7T8/bokuLrMW6crJ4M5NzpgrKg5XNEoQk/VjlSEF
Hiy0hCS1M3yJv0ohPcWwQIXlgbkm6VTpIyHG5FYi/N0mWzPsednYZyxqxHZGROwM
wrmeajJ0U0FWe5jIJOP+l7a2sHanRDafI/4C/GMYKhElWMCqWkHui+nJLJrpiI/O
iy7ljm1YXhYDhljVHC6dOsEDeKiwAYJcY44MYlPY6tn0c8xAPPrYpGmJ/aoZULam
awJzvQAzwfKATmrp959bNxNlhqcC6KhSY1K7azefO26v81y6pUodXPkN4EwA9Ib+
VCoie/7+Ocb8Y2NhHCart/TdU2VrqWckejJ+SZoovbe519cvK8L4QpRAqqqeLUhf
A//y5iXUY2x6AltVY1wYklvxc51+YBqFJQcy1MJEz60Yot5xTZbc90dP6H/j1mCA
qZQ8xeKUdPzExJwkA38BigrvJfxG+NcXovmHoNwkIbYtTnSV8FyEP5kAeXHGeG/q
U04wi9OcKtks8mf7Lbl4eVfkNvTYNn6cjtbfeqTBd71przv5GBvcFQ9bn128q851
5HZf+otmd7o8lrazbX+TaMFtzA8cWgQMRYZz7ftI+9uHm+lkaJeze68oGlH2SOil
GP58+5gqus3zV9LoSqk6k1fxvWG1JoDfIzWSbCP8+XpVrJ7S7ADaRS7xOf1BcLaj
3gFVL7sKWFA7dQoW2IutHfLo2YcSWntM9QOLAxvFFQEUQun9EAAgGb+YW32aT3I0
kkhNE1DA4TJsiaunWPTURwaCzaAh7Ei+FL1aOryM/XDdRBDHv4R6qh0epq5kmrVf
kQCai/4NIMg2XXZH/6uR2zYhenlJk1Uwznj8Yo6NG4eh/cl4SqkmiO8SgtFZIGDb
mCjAqSUY92bhgAjmBm9ICgXtHXXEmVZxMXPe69PKbuxreAzDOZ4+wqD0cQfRuxCg
BtShKmrknOet3eMflRlZloFCEmRO6EidyCczwgsIev3Qoa2L3VHwOVnhx9t0W0ku
BEMshxqW7UMELfJ305Sk8YQx9a2xwFt9ynUiR6qdwCfPUFWQkFHw2QK1GpLrTTOD
xb9jGMRHNKVnVFLb5sDz0FpwpIOvNjolHGZB4G8pUqzXpp9ADRNr2GaUeoOzU6OP
IOV382VtJnVCTfp69IsQo/O1rXtBKZVW8mkmaAm7UOsziLwVrfE0LbQl03ov/R5R
ukQvljD8tbxLK1b4OLH+dFcH1OydyuBFRXFmVZ4zTNpzB90CRA0DOAvA0EeN6jKj
vFS1fBMnHDq+4r/Qwpbsr5h5uOAqw0h3tYa20pnu5J+rk2s+QjeWnIsLIRJykach
BOOXB9ObcbDenwXaq0NMLKrcWsuWPSNmn9OOzRnrgY0huj3kl0OHgsf8X0okO5ov
lRx0cF5bhmNZhIqyacG6ASFPUX+kSROc5BpilwOavMVExldRZ6EpoHXpkQ6SfTla
tPCzNvJDTXLhhbxQ6dvV2Mgr/WkVHTuaotc+RhocoUoePAe3p1Y7jtQfkUW4Ljbe
l3YuEi0689uFaCHD93qJFvhXCsAldJWjS3WaSrfb6gZhY3a10g+jc5DdYQpE33e+
q2BUfSNj45AP3aUeZUy4AqqevbafE4pPjwmDDvcXrDaKz6TmuQErldF+fmV5n+fR
ftBijJJa5Cg6uKlSfiNOC/Lhgn7gVKZZKWEj3IGEALMDVHrna7mzR9YBzxfAZ7tV
mnrcgKfTafn/Lq1r5iyWP9zhy6K0JQ36y6qKsrLoe8/6UT3Mj3ORN/a2s3k+tfPy
QZYQAFAHrOB299PcPDhXg+FcUfOPPCEXMFDxPjBiQLHNNkQU8bTg1IVYa0bpm4DB
tC7OoVpJk2mJjb2XoxOEYuY4CGWvsdaSb7eu9sbgAhdR7V5tq9AszJunexp1xyKo
kZzpmBOoupUMTKd0kFmCFvm7z19NRpu50IEAHxjVxgXF5G3TtySF04gz1Uaa7+bS
y9WFbGYsyAvkvTV9J5q9obXmpIHxeJoSHaSNgvv/2AILeU3QRxeT9GIiqcdcsyFl
ap8O5zdXaTQtFtmN8/hvlSk3WccTAIV43tasuALC28QWu73ukkpbIhqkWsUANOgy
mu+D/DsZQOv6ZvhfaeXYogxLsmI84EyWDFMvKVftNOE3O2liNa0Qs2G3PYwLBtlO
l8EcRlSabck1L5DV0gkQMV9D/8K38mSRLn0M+tF6y+kon/CgvV2lb558R6+j5dE7
tWr1u+QvynKUgPfrhrX6vjWXijwwrVursqEmE3rs78LqA1eHQVbdbE31d9Ocoevg
QPjzMQoYbN6D12yw7FXYDvcn/c22slA0Par9O4bCWsOXZdW/qMSnsJW8l8fVz7HT
sFRyXqiy943Nz3v/a50xYMoW7nxJQbsHSi7VYfu3GRj8PRYUCQ0YDLFJNg+75Uc+
X944HDqpWXAjTzNNzgATRjEBZLCLSNPC6jMdq+RbeazhYpluK+URATUfMwVonCxx
OtA52UFi7TFeqQtXR2qWa8Z6DCfyqjrViLlx+hrN9RmWLleePlHGP4SDvVWWoRLs
64xTjW5Gkz/bpCx52DXrPnm0T4RoaQKe8KWfgKK+kX2H9+RPBF+9Ptxpz+o7F8zF
oaxYOBNkMvnaURDry7mv0d49C+Sg/5dWhlrpEioT85ekIAi1UH5ZjaQMIqt0GyFB
oRehGerkG25/WhQjpl4zreBoIVminR2gjaBjgPpl7f1R0TYW6+/9sxC49fe9i8i5
LW8++RXRn7oWF/MVtlmoPuB2yazBTvwTx1gr8EJWhxF0A6m3rOGxxAEkVOfFsMZ2
vHLVWdOeUYEbaMm/E6bbqnUbsd9Y1/GGmsFlGHXuXEd1WnXHlsrNXAB2B2xsaHpg
MpewbT0hCRPS/6pXJk62Rzl03Jw5A6hF9Lr5Vc2SbH5H7j7arlzbjjIDswBsJuyY
sesi25HRJOxw0rPzEwvkvBGyrDS9jb2pz2XdCSZPjptZ9U6XBf0FMJfqFhliSk2z
XcoBUeUu/1VjmCSNIROQ5aiYTpow1Kg3BzVQe/lLP/S12DqfyJjvx7RR4FdLleAc
LT/T1NstLJ45ovhRa996iGElNU8ADvUIP+uoStE+UDNDpESXr6yQGNLx5szika8T
xSImp/p9Rsdzexn91QO2DqYvtvzTLGFdGDOgoFefXY9QtqHNb95paViYdIBP2iHH
n5J+I90QSUtWtRBeLcLga3XW7f5lfmOcpaoFzPg784tfkSYK0t4O1kssx+tHEpec
SmQdW0djVFCOUTS2TfSnDGvwpRDnl6LGZ8mzldh4wVmSBJGCf9HdVBwDuhRrNNg4
c3vHTAajXOqzXq57kmu46XlITD4pkqxFJRRooRwtcW/tQaOUDEP/Bftj40rAUDah
fUXVMqxDWvFxpYZtD9xYOHexeEPVvs4MclSJtU1aKW+dnTTls0pr4lWPvf/3t6JA
KcEbGSrj1et/GV8xfQoM+P2iNDYNtlf7gWeIC7IypFY9jFP4UfhdfCuJ5ioA+2Ap
nAGWQ6It4xJyA+J2tt856R5FinmV/znBrFrhobPHw5fYgwyTLvy2AHk+FMNBbo6p
imCq7Gwbeo0Kl9Za/Ii6MvkS7FP3V92ajXF1UnDKe8111EdD3M4KiaBdtBHQczxY
pg2Flbz789iVtjrUcAG5nNmFKXyHEUqjSxBWwp84qCVikuHE0PGBF25TVj3XBVm/
5Du1qA03CSM2IaVL+G6KmGR6nBFy/sNtwPW5PJcYwCu+/NAmxqblGzoRlj+K0q5U
esngWtSa4PcQiXHxnAt+8jqnT9B+ym1C/Ze2HcbCqFY4QcrKOx0YSeekt804KPMB
5tMf5MSfyugilB5Pb/LJpNgWi+IEd6t0EVyZYiVTHPMdv//Vcv4RgfLC2fbUGzHw
YNEIAE73Pnz4Rb4Vfiy0RrjHyx30U4G550xjFHqrGQQjKppeAWvJKQ9tMuRz+4Nf
7rYG3WTmxIHJnd+WHEmQuleoqVOswKzhs7Fn9cErbXH21FfSQR0bBt4qUcx226Sa
cxgFlyLdlSe6u0U8kIGOs4DNoE80Q6PoAGARQyOgh2A+IK9+t21730d4RfJ2LcSy
qsnJKJZF0LzBdHnR2qIxnjjZYdspFfgOh58pgx62fxpjoIumC9ihZQUXiHev07Rd
qNSH5wRbOA1YzU2oKcNRrSSOWjQ9x4QtCqX5YCRVrjoEOax5XOuyecGegC/N64ic
AYNz0B+KnAemwz/qw9om1aUrXFDz3DSR9HNo2QeqMkXABnAOavF9NXbQwLJq7K2j
AQuFn3lyYPkNjnzto1g5DLG8u8UZhulK27Gg1ruN1wes/xemsAysyNeDVCJ12aqz
txKa9BsDKcoYh+qx2I8LgaoLmeRNis1KzTKCtli2sbBH21RVHfPbMobw7WhpCvzv
A2OljiK7l86wnFUwPxh0hzlL/zAnnA2LT3eM4oT5GadPwe4f7wo4rIsmPs8cm/CM
pOF2SDlJDUzoIbaNdKvnxWDuSh98rZJIgAXrbERAWigbWGUbA3ZX9SFsB76ZWb+8
zGUMET8/iRW4kkq0RpNoiAWK0Sn6TTw+j7piyeNhNViFA6VFQHmctaeVOhA/3gU1
GAlB5g8pVWjFJyUUU2rAYQcpaKOX+WxVMMkDG1QEu+RmZFiznsgX9/fyqKz8p8Jr
bHzIVa/i2CMiFD9Bha0/DV2LnsOeyCUUYrGWaCBdmX5VFSw9iesmNl46a20yLLge
54zYynsC/Ge7AO8fZQKtYrvRHFq8lOiHiO9WxBQrR0Ev+EzgezMOf8E3NPUbQvPI
rvu2vh4v8mdzqy+zAGcjYjdv5dc/dSb8oRHocPY9/Wz9CvBeLbIaKqRJ0/wwWV3z
HYbwJ0iEugSugSxwIjXWlISjPx9AUXVp/06jBRWpDACXD7XOGalKqPLiN/nFrDpg
2PLCbBcZqVqK/FKJFqL8/IY6mzSwQE/gi4btmxFAsdukt14g6WSSxJ2FuTFMN59x
weCLtOYJ1yBlGqRXDfVWNIO251ZmFiK/LKfVm++VenuGoOs/d7DP9Jp8n8UmzNxk
1vBR1xp/HBjVNTIZPN0SG8S5ANs+2/PcH3Q1NMVekDob58vgh+nCinmDGhSsUWYl
uEjJ1QPk4EFNAQkOmP3WHMK8Jbhk0xyNb4D8d/gOEgxYrZVGAc5I9qiAnZ6/JzLt
v+EM5olf9gHQootdhTNYNhRffK7R5i2IjiLkAh39VCGIEQ/JHNvsQVv1QjbAlZNp
tVFU5nsLmgFy6DxHn5XCETQv2l4Qyw23uoCLywpfotFAEYfCYh1z0K4o8X5pNjba
x24FChuvkn1mKj1qCdfY4vOiXKMbIMcRdyPP4xH37NvmfdrQFvdLXZ/24w8Z/e+A
kQwwLnyGIbMOHgz4Xem5RBENBKS4EdTYgp3Y6UfuUYCygI2it4DMwyZ23z3XZuao
4MRQW6VDJcCpx0rh9e7Y6FwdA5Zko3ls6QdUEbaxeNUMB2ujJisJ7ST9Q4l2WU6j
3GMrIq1/XdDlgmDi6jOKvPpim8T617K2iXoacs+1Ma9BlOZjHlW42++sb/zFirFr
To4B8Ay4f7xEGVdKTGMFA6pX7yD/+y85KGR9obqTAr6Botf0eBuQK8ZoVWvE5hWH
LhiWWws0kuX/ez+1v3EOgmjwLa/9pm3LgS4bsEcMlLJvboMVaduBoVThVcJ/rl8M
6qE5paHK6cVJlsx2kC+tIrpkNjyk1LdCDaeJ+ZHiVcdP9l1d+wuqNFMHWjHEr/Ma
6sKa0w618dFau7gmtzmGVwZwNxdYMdOPIn0EnEYKm6W/qceloNKQRSLCXC+dl7NE
cgMWw5w2RXCZO28sUvMy0+ti30WVcQUycTjJ0bUPBVEdLzdvOKf/op1LA1ylUfUc
OgH/TgLx2mFRio2AP29y+5oqT7EOJ17RjjgxOPk4YLZhkHBSBP/8MdxqutZi9YqO
DgR0dtAf9WsjzN7n0vXm0m4QVEVUGsitbIupHS1z/m7FCloaCa8+M8gxrdRg8/5E
eNRm+2NJHG+Rsa7sjh/XrCnuQoum4FBmuepRSmms0V3c74aQb5xOKQA+2SH/SA0L
4EN6vCK5TLwjDxO3tperhlYwLzYvU4y5mspT51ELF+piuQIrEYATqEsfWbB94+94
RCLQMYKj32tkCRaCnMgr5jOAlIS/2iilliBrAcriBqCJQ9FqXHM2LwnP6ZjJYXRE
ROoQE5wm2x2+XnF9AnRgC9ecEk2qph82nC9vsU+j5A7keE/63+ZUKOhfBLBQ9JIm
3oYIYfj3y047ez0GTqg4NBkfSxAfY0souB8HGjwcjBvGqVzQRKy3IhNONd/V6zds
DMoYO2OWNKQtxBnbeQbu8OER6O8wFIZa9jPdTHWD4Tpy/LIezwatv1JM7RQDQ3YW
r4BPuxe/khYt1q/80cqI2axmOvSHp+9fTTqLDDojLAXcuujXC1SaM4V3pOVD/uJo
McsfWW2gUo/5uJZwOpfktOKtjEGTrkc2PnKHRv2vBLOR4BzmaqiMKkkX54qgyCQH
eQzjXvlQcPH3IjZQKDqHdQfKFDfiWAjEno1uCsNmD/1c6I2a1s3MQri4ONSNqDlY
5AP9mrJ6FChSkWl91nu7l2A9f5inVIzdsUMP9njCK5L0MiHnIxldF0KhDgwT+whi
CDxLWGAlUWqJFDZqHawVmJor6R32rN9bhpwaEEjcwYGCaAvizRWJDtITJ9gzBoBF
TJ/puuhJxtQ0BDA8ZHR5kyn1WfzuLQGRVFF7g2CBoOdkGbyS5YDtKYsunlhNPDjr
iSg471nqlgo5nuNkYp0IGVh0CqsEoOjT3TEgSuIX4nd3JIkUB2+U0yy8OoEaDYBr
1w8+UANE8qN/AtKAF5vqh/NfX/OuBfyYkP90MT9H+HAKVkW3D+pVkIPtx19tw7BN
Wv8tZj4orNavw1jt9j7aGz7MSTTEYZh15aAaTqBs0CFdpSfpDF0bjb7XNL4tkXWm
e4Un0Lnk3HE6nzZ5DFlqYA+xQfsY94A3c+rkIc0MZoesTmfbQMz+m7hPhTnIPJjP
yfGyBJbleBdNKe2CWg8SN4ghoaXLLl1bFAbY0z/qf5fE7F0Z3I7sigzPqHZ2d4rm
rG3OXZ9r0BDTXkCwrqhxuHKc0Lq1T1VtErQtK3TLM0PWaqRsijRr7PHTjClZwPX6
bdPgo1dCD/zP0vtPz4YeSX0nu9dXdROZHgn+u13yozVhGcpnHHadMTJe5F8oEdEu
CnKx5gQ8IFlrSe5jGGAEt5sz+kPtgn0hdCxFDXQrzkEDFQBPviZ+t5e3p7xDPenn
+I+V87xq3hELxdTjuBdelRNfuz0Wgh2PFU3qgZIxzT3Q8uUbsm2znEUnqnPrF11i
7afp3qf4WyRlQluCxjjTP+IDlCjGMqnxG+NxRqfX6iCe7UOm3QCiL88ch9Y6sp42
0vjKftdMngOkFYObyeHCAKE8uVDsSeooUxZLc5BjrJQMQDTGqRHMcOaJjY6OG3ar
GubrE37rU8o+06UBVrqwseHnxjPgAYh/UWkYxOFgJYLoqIXi6e96GapukJTv1Ipz
1J1XMkfC+CsYIk/fI2vgzQhaDe/hIrd/plrJV9/CWTs0mGbNgyzYuSYMbFB4Pk+S
uWuagp3ebqBTo1JACPNw7/mO8ZP7j9k+CmA4xoXWjkJzSGk0gLLdlYsa84frhGac
gCgvFYtBxHmycBEzCEbM533gRnb4pMTrOGpEapa85W0LYzIsjEQ6XOsvw4pIstzG
FXZIKyabaktFqArxtPoA/pxSEyGK+9rQN/x+Ir3I9GNitcQeziT1GD+ej52PIVbJ
/A6O8KJa8vq1VqbjysObuECIKamqyco1cvbFRXovHqWX1yLV/epr0ceTslp5zfuM
riIDRE05Ja4xwkU3v4fDQ+UYtk5jdWIHUV6N/Hrenyorh/Fsg93huUB41ssPc6hA
ZNzsPAwKdNErc3KUUfdqSxWj4/FGjCtThpK4asmC5dZfePvoMqTnNjUdy/jEOnyf
Lcwd9Y4tUaju3WNQFHdpkACMoTm68LskbNueQ7/oO5uwC+TxBOsNguOVD3stfKri
DC+dwpbFJYN1P5nz2BNSog/iEG19Oufe1vk7oj9cIUjxgK+7ju9gqLZvLKg54KeT
6/9TWpG2gszG7geelaDi29B5/qAkcBkc/8z3l0HaE80VYq3VVief0h6VfA4cZY2C
vTv2ev53oAlg4CPYzqiUh6h/nz7mfu3OMH/UZms6AeeNqiePZosLLsAn3+XGIbcE
xCwoh60OS9TdIegoBFlivH1Fe1Q7bk+DCCNYGzPz1dUyIrtf64+MFWNXGo3mUJkc
3c3/laTTU61tC+N7XCDBfkIY30oxcBKf7DXMhGQ4WkRkFFI68Jd85M3rGDrdJut7
4K+w5ViqiingQB9KTi/OvAYobXwQjoyhRv1wMdMf7Nd6hC2bh+gyvBvROEEmrm/w
gPBjIJVS/UjY2OYrFsWEPHiUMNcdOssIJoylxGxqLMrbN2HNeidZUhyGF2wrdi5t
f/yb7nO528ZWYOHhtGCxjgxn5cf1SqC5Z2CwGFWEH+2kkHKCKDSExgknkYGu/aBx
EDzELQMjALg/qGnW22/6W8dOMAA868cxvWikC29n18yvb6VzLTDwIgF7WgSRKaU/
rsX7rZPvi1LJAlpz5OuFEVyx7m1BzfrtOWw7y8F2QepN1jEJyRTBlf/MOVyOBFT/
E9T/zryxcg9UOt1dw2IZ/3QDVsME/mjYrChtktmNzqkx3L/VOqNE9yZlaxAD0lmQ
RuATF3+1oBUG+lzhmc4uMTrt2abua2yffvHUwGlEdgM2l+12kIo6J9wrEkAqeQSO
ht/5cK3M2eIoG7tMdXFLDnRSDy2njccI3+fbPze7y3y4d+5KIAEy0882XBMDsbZG
VgZJdfef07ibTpN9UeUJtg5YLYkF5rlGedo6dqNnfzDmbzipF2pxrG6uXY53QVQK
+KTeh1NGGAZ9xPDCHfqF0qDQ+RGwe9lb4GG6DGFjTh4gzSovalqqLQNytt8ngQMl
c+X0Rw3RnEAJVAa0vqWqIaWV5yng4s5cUudQwafFm5X9C47AwcshSvRdudmxpWOD
nvqahQ4Iy9zu3z0fmKZV4ERe+rIVs5smY67Fa4T88cPuIvmC6ft3Ie1XW3oSMsT6
1RSIOt5bkn7rOwuFAyZZF37TUBKQDWz63ADOu5AGtkgKI7008GH461NN4KFDD7va
rmBfoGed7b914g65HuUOrS8Nh89Psq2vZJJAs1hNwr4AMJAUmJwiK6olzh6MAqZD
gRUfLAkWTb+k3PXOBWvtvw8+e8JCEFAy7LKFp1969xLv7T2y+BqiB4N2vXrOievq
cGdW93L+QeJvhBs91reA6QQtx+8H/SiZX2h92Jg8zn08yaLVWPFu4KYQv9uYHnzm
Y/C0Y5o9ekitHKUarO3pODK0Zfx3ueKqOUa2gO84rzLlw/sgjLHA+RDFzXDoBFD0
blW4PVG8ILO2F9ZeQYBNx/072P9Yo9/VFsOxcgdB0rCZr+R3sbKVOpwMRbTgD5SA
5TVCIsGTvncR9wiD7+uDrF3jRn8VWNjhFKlW2Vg6LyseBlrkNqbuNZSI+ggpu22W
ymDnpOOTIOGJfzKciEKntu6IdJGNzISntbpmWmNgrl7Epm7Z7ZH0S3V7jlFUH9Mj
sL2Go1+TxDh+g9v3Frh7BuU+4AJa/dtuuf80VEwCHdIU5p4oX0DuOyPX+q0um7w4
DKJ3fItgzSWXLF870OJDE9mtQYCQNhmvO/+2pS4fkJxCwk3nlFOhv++0o+gBf2Ew
VZulsUIW6CWoYeaYhqPV19ROJxrS57cUgOKBAIdavbC0O+hxwOSMXZ8sgdX9LpTT
5NrKgsP7HSllDlG5liyRqV8qPFlXFlgy+GlR/VU2R9JYT4Q2yHeebS5MjYgFosdw
aQJqk99D6TF/lGytQGz54fOftyn4lyrXrWQZPyD+JX3DrsYaKahcnga9OfrI563b
PSptX/jqW5Kurc5YE+swd7aHTiLgK+xYiz8JpxxChlEn5gm+OYy3M1+tNfl4StYd
nCGqbUj4QQ50fhouFOgxKOJ9AisdnJpUwAe8bqv6XeQe6G921+Mz2bL8zJhbEARf
a1xe5mUvklhwml8xN+ozk++Emk7Gr2/ytFJbrx+EUBbRrlmsWqPFCHAOiX1NpmVL
v6b1l0uthgLs+tzYlRW8H+ydQYLH7tZFku81RskCLcwQOJjW4KIYO/498ryeHN6c
3sp6Oz7yrY+AiT2jGec99PzO9rGzBAMhbTlK80dHxPJAXg/UkbD5jHjBPsD2G/zk
A5HTfWljeQlBTxrw2Rr5bElJg3D/9+iRemtvhgoApo/Ku14+LzcSstfmuNdqaG1M
eNVP+1/hsaZVi5t70apfWMJkJKowLJ4m0csA74SJ8FPZooJ3l+TI9cQRD+zOtCP8
QT7sftlm1EK/LyEmT6o/5hmtGx6L0a9PCAgVfOA2oFj12ZiygSb09gDtSznHVRG3
CZZsZECGCCnmmpWYibWd0FBb0r7pB/6zEDZcFah7+q5jki4ujrIj7XdrQPrWI6SV
3tZ6WaDi9IsQH9Rt5QzF4k9kh93Ys5+j4DT/7soQPERwuB4FOGNx/TSQ7U1GK1aI
v9M6+isIC0UzikB30hXQTcue/0lW0fFMrC6DrkNKulSQZN1T3nOnaoYlfxUl7uos
6v8aAzhq67r4ydUoR4Z2WDkISxzknbm2o8vZJkznF2R5ZG0ryrkOmo9omIbd3dYG
lDnc0jZBIVQmmvqXh7NVmnDBun6/Y/phHUdq/svAKL4RzSmLXdo9F9W+0+qQWYpj
k01zdsHPAXMlbiky855/TNevbruXqdRYnT6LSS6Cs8LBnHwc8RjVvNIlc9QZD2mo
JtyV6YXmtZ7OJQG9dtaY0QQdnHG8uONFQ7qKuqaEHIxMmDp7Sk3GOcEMp5rrUezy
7yR14CBDj77sv3FoO3lSqKQmFGtiKWbW0VtyEErWAhW1wwuWzUgJT5YILHPEhqoB
aa4EfqNjChytfNIh1GmrH6UMMR+dpLCY+vcy+L4BzRccjdDeEVkdlNhyZwFp+qXI
o6K7W0BFnGpSYJ5KwYUuBHhhDPUrjniwTnWJQPMXyBlt1pGNTw8ltjzS/b1yoxAH
vLf0geiWGJ/PitLCxQm8aRCCbvH7HW8EeWbvjtSh5gE/0ZXIC9Ya6tWyjLnhL/wB
rXRNH0jkQh8f8tv9Cu17FwSgDPVNBNeuh1UeIn46UoxLhrUDUuSadgbb3dMNKFz3
bLTq99Pl4TNJednotzYvS62qV5RtC16+ds0as6LFYw1XGBU3Trm9fCsFS4bL3Yb/
4XixI9wz6+8gUsstsZfWV/69ETVPTeqAjqB76HYIpIpFI9CvgAHYPgh9/y2INE0/
NpqHAKWaQYgt1UN6D1Cv+teF7TSlorUQD5ONMVGi5qmeE/8DGlIn49jl6plGJVds
VO9Dp6/RV9Q1a7Pav7pZG78grFwRb67XTQr9FHe+NWiNiic3xC4mMKsPsifssDAV
3b3rZ4cWJy8W52AdiYGLuoOhQZiJZ3IUectDKj2nqXYRi2hyUSAVyvmqjelQrQ+K
t4dQyqFDl1Yvk7C2BIndQJjUou7Uyfnmv/9ZQ/iEoJVeEyBNZncp3nEWRD/sCqLM
DaGIjM10ZQ3enyjTTzhsIzArdyNSfx1JanYRbCs4CvHVkaF1pbN/pq/Im1vLMabo
z4obMroWbF59S7DJNEH4RfdYS18fImsa7RzfhCQs5phGpET3RAorQE9Yi6nhicDV
UI6EVjoTwNQ5wBPglqMEI6FohF/GfFiBqdOLFZyElocDhH5SDKm+XG0bz+bdV70A
7HlGdSLBgbUWXBNiu90PJ4iZxEySx47ESx1Uaen49NUEE33cwc/+Ob3WTIZ8T9xD
/GJk+OMhrYqnJ5Ik6rqpRMwi6zYCrlSnoeRYqghvHK5WjVUElgCtBLL/PxwDD/wP
rcSxaaUyF7ksdFZDCJYKXDh4AmhLnEi+yy6qOsH60VlNaV+vVvcyqT3tvUPuI3tu
rc0xoZn0KQSgivfMU3dYCg0E3VTvFzmD2I2rGir1fU/njOeIOVzaFOs2TpLmZbn4
VpR0GTj8RgGti/55YDUR77xBupFJm6Ndkeom7JQRdWo9R8LiEjx3irviJp+cKzCL
3ychc/sJy43uzAF5/Xa834VCdUdqsoYq9GxNhfaClxQ7OwP4Cz0PeJIPQd33NeA7
qjlxB8NmUbdnyrZafaOt3Zaq3UIdxbQE0X8IG+xPdTJYDwa01rSSFPnERYcFquSl
J/1u4AZfkWfaUiqAu5JOSqc8o1Auht/LJgr0NKmV3y75v/aRaFLBNCEoZTgp4p+2
uHAy8YIYTqw4q4gnic7hZvkY8VKAEpkU6AejkdgvO2LPIcWVZddFBxm/PA3O+ALw
x9PUrbLX1FLHBVBQamAaix7qBoX5j/0F/Ye+zzf4qq115F8v0GRzpzwmck0I8OSf
fXLHHXZ8R0vaUDxoorqeAELdk/3LvCfYxR8GNQ3gPyDWb1FTVXPOyZ1FwNETma4O
d+lb9NyiH03ASMBSKp7veyRuJ98CePfKt1AzVzkS5hza86tvmYQeLtF7+TTTQ751
gWhq6uoFMEoO/uhbEZqpoERn0rMTmbGCEGKqB8DQuxcf3hnyhXK39/GZjf5vznJs
3ylhXcni2BqLDZFQy3q75MKrcD695VEAgWaQL7Vzu+NI+Mu5Gr1qjEyl3QywkmT2
peKDIrqXvguwbxGlGvBs/0GgD7lwHfcP0tfpxM/ZygZNT9n4sslk2VVtIUM2B3S7
QO6BZFDQ4G2Fydbhu1VjJRNsQMt5tYtpBBEN1f+DjHwnhVTEGdYUXKA0CCwHeF8u
0bJ/eJyHZFRwRfLAwPNSrvnXFeLeHZi32bgAXKSyHWQ7c0A/Kdj2y4piE82Rtgij
bz0vXkzVDE5znPTkfn+WhkbpVcoQybkzH4W41OhdtXMgafQ5nkU0GXM+WqY/O+iH
psJo720opIeqUYD+jFodtINOND1Pmnn2ZYVX3FA4Syi1KIiFfgPAudvnMK0kVCYC
qT77b6ssPs6YghQAw90f5/tsvcqziKeZeUbaYU3dpHvA/fAsarSLFoyRraETr7WO
adgqcbKMzGNMo+SMaajqcA5JXTjgstNAzXePIFBRCSLX11DCVysiL9sGIJ7kB0HS
QxSt8fsqH/OAJ14hz9jir+Zoc8FUUdJ5ocZOy0z3XP7KcMRbIfiwg3jO/w+IeD3c
FOp7Ayh+QHQHsbm0JdzUBiy/b5OMzMXSUNpRp5r4+PuTUIaT+NlkDUyRMXStWu18
BBN3D4PtJSHbqrc+KQhBrJwZYKc1/IVZ9FA3t5eUPKCCZso/mGVrVpWyTSXwaKhW
tdp0CeWBC/Kac0LfC4/+vxR2dVLSTzs53fWPV6BWNfKhDUThYgsiUFs/0XTD21wo
zG7pVwxzc6qElRWB45o3cZCSOu7Ap8sH0VrgTzykViy+K69O9CbWvAj3B3kGG0wO
qtZX9K3pN+7iBg6dvjLNTts0GXajGLYtc1J72gYsEX5K3Yoso84xxwr19d9WaINe
LU/qJrYGs/d0jGorniHWq3dftxq6VKjNvJk2Mg1Ds+p5d1DSKO9PK4cXUYZLzAgP
/TWNtB4ye4SyIXxesRqtd0xG3ec9df79OhXDuNHWH4VjUuRRmel4d2266QJb4icx
kFuEhhBqx1wWmIeceXpAZyqnL/aLovrereyt9ddv2VtA08473wp6ab/AjhjLHmtW
horVJYM2ZOXiSwAPITOBlvErmclZdanEPvJrKEfqfiih5dOpqpWv/XWE997N/xE+
vBtk7UuvW1dil95LjG2gB8ia1LMtzOb0ZY15zwlU18pGyhGlL+v7sTeBehJoOx1U
i3K1XYXrTeO43VuhKBeTmZj3RS8b4s7IPiFFh7fgBxFVf1YneiDUt1AzOFs7vz3M
3Qm10WnU5B7h7I88T0FqaNp4NIXJ3L/jSJS+O0B/iceIzmiL4FvmjNgENSP6cK2a
JWNJqFYsFuwkcRo1BB4DaQ4HNDdfFu3DthsMrWP/aJRnv/mlHiqqXjMtGVeJ7DUO
VIddpHLF4+/Z4Os6kCnb9VUBGScW0Hs9KTPYjViY6tBYRRFXo7K5MuVIXxyjSaek
4uB1oPN2YNftFLmtRCqoLNEfEqK0Tolxd8JSgncpR0+1cybyFxaW1G2wnBbp9rkE
bVu043AEulKmUlgbigzYUO81kEmPPQmUJDC440tMrMtg+ptfFXRVdtn0DnrsWMDk
4z0XXmVUAX93Hw0Mc1jQ2WHa3rFkhIM765t0M29/eWQoGU6f21DJ8e35DMVb8Txd
Q8N0H09mobyLl29EBo7XdWPv1Oc4iO4q5K7uYqyKKbsmA8CXlnivRaadosbr/GvH
KG++iP/TFNpDJhhcNUgq2U/HyEHAyd0bJ2V2StrLUjCzm6mVR9u0gDKrHwXdyhsa
qH5hPLod6B3fum9i5vm+IekxbXNXTX24/GBzTS0KDzndQ4DvuIJlTqmZ4YrtBBEg
w/7zGq+Ostwt/naBwn2aeXRNpUKrdYLCI4pB66RuhAFWJ1Hj23bW8TPFKGbfjvdq
eotjJFUcsvGckYZoF1uYeskRYmatGvulmk5lJgKeUGkSWZZPFPJN3O8XlX0Alq73
aCv8j/MzudJ2Muvph0PzkpwUUQWNzkEwatdiAjIfmdySUIFwD18++4sSIReYUDRw
XSmLU1gPUNoA+b+yYzKiqd8tiNxAr9dmu29+mgvgHtIIqIiAkqsDSgNx1UYXxnZg
YarOp5QY2KjUfNAgmiZCDt7tCa7QaklPY333c74FnSVBr59SGLd4IHrHmyFMkF2D
20Zuo5PGdW2kpmHGEuiGuJAV9+Oex1tOsPuzmTVPoqKA5lokJHfTEbfRUCKlrE8Z
vXaIt1BDn2yR2URmiUMyABx7dqZlKt97NQQLXEalbLSmjnSrZ1C/CZq93ko5pnFC
8iNMIUnUrli6jYojA6M9p70JHd7WW/n+VSTz3M/fZy2zmtSwiONewBM69g9lvHrY
BEXvYQUCLQ+c2G9GNU4GIJTYk5kpyW+wzrRZsC3gUUzT1TVtbiTuE3U+nFaMmz6z
qnzIsxYOmkWzbXVLYNNYZBjolnYZM8TkY7ma75a2Fpd6oXSywkR6uPZWxBwdlNfv
Q1GDlEC8NXj5iaX06VoiFEXTxPL/yatVVcxEu+c3NkDxvJtFjFmfk6hH+FFF9sn0
+760UZHw8m4z06l2+YpS8Cu3fCB8UecwkkdhWYxKZRuqZxQg9FR4Ma4y91h6hNzH
bNQe+1i9275OKkYKEZMrhF2bnmUwBX51Yg1tWnerohyPsDBfHBwfvKY9cSXMUOT4
0LWhCv1eRVYnOmftEhR3PGyL/nTXuWZIVUwTiYXIrIRp0L3d3CPHU9+eCHf5iCB0
IDhrSI8lGO2+xqn0Of8T85J9HkPOrrn7hYgWUfANpz+o6vD/glAlqt4j1copSL/c
1/pxhMleYYXBxentkaMidASxYeZW2MdXoqiKc8AG68qDIk6xmCb/jIyuRfza3m7r
CEGsrNy2qY2QoWqmMJbqK+yYcKtzMmfBeSI8McentD6ZqrMxzjYMSmMZK+0tAeuP
8070HM5ph82SIhjoAma1W6Zb7ZeXj7if+yr54tclVENjFlauHc61jZ3xgECE/x0J
6vLT91kS0o1GGEgkU1hFi1uxK0DXwBjsW99AES77tR55Y05K39SvEg33KKvD0lRO
h9Y7DDuRhKa/CUBF2VHIsOPaC8uimSERjvDsZ28kdKa42+fIvWDw5udCiDCnS+Dx
sLUlkQWrCUaoRhxytl+ccPpXtusTEehFg6uPq2R1dlGe9rV75hAfjKK0qQpOkclJ
3WItQYVtjlrQ82pLx3zyZAMulcuYSO0mpVHCTC4fbJ69dhjf0Tge6pGb5/rF8KyO
TP8MIHAf7mCL3lkgWFQYe75ICh2z+cMmYfexj/OtxOhtl3yTahFCOCZpkBxcJThK
/K/TvtVNwByF21AqDULqSPAleb22jveXLcd+DZrmOE/uQodVkv97cSNT5CfqNYIp
QZgV0ULV01LFBLoeScn1TP4w1vhcLPRf5fkkt5q1nwbznM6yeVqGC9aVgD9JdGYq
+x5IDjdmsERfs308gPv320MWlxMQGjGduJ1Ju35dbtZ2hbOrHnzIBsz1mDQi/OgV
heYxPyeWEExYmJEpAV3pHfh+oaebVFTlTFKZZy4R/rA+7tLnqEFJ/yxZH2B9NmOp
aHTNeS8+E+oN+oOo0ULYFlk9XYVc8t/NSNIRqlIYnCdhs8bwYCt3jPNyROFeBi+z
JxTdgp4cQbcB4BsNONIcSRzRcsBL+TH30M2hCSxk7Ak1rxCJjMc+7reJJwyBTiPN
NhjOWkHF0Zofx18XDMYz4FYBkaFH+M30Z2dUdSjhvsDz8B1s4+lw8J1ncgzSVGGH
H6GOES2HrF2x7l1NuMD+0uk+CeMcNialTHHu5GEVTr/q/W2g26M4EVdIFeckpkYL
lmOV5eYEFfAcWx/nr7/obyX6+Mgm71zuiWSLpz6ahWZNDYiwwc78tK0c1UqTHhwg
JNkMwvLdRCJPK69JS6ollifli1hXTJZ2O5xK63SsMCeOqW/bauSyLL12+6LJgSrk
NNqiiE4rrOn5gbZB5C79SGQT8RjlKA63evuz/f49+V3g+/vaDhgARTRImxLDLBY7
xnQYAibfuJm7+8dC1sil2Xx5bVbsUzTpQs0VGMh16jgw0k3WiBa/EKBuj9ctThU3
KP7DSHbDpB9xPZ/eHgsPdIaceLDfL1pkQibHLq+A+6eTwGWWnWWeMNsPC0eadDCQ
ddEdjKoK+n2kJIvMKcoBDsbEY02tcTTP6kzFLosCJyn+/np/oDOajBgnPx4clnsg
tZZtU1Lwg+klbaNo8ZWvgYmUmu8RF5UHVd9DuwihvNYoL/iNyzozbiWCP3LgEahz
YKYxD8qbV6ZXaIWT4njiuWa/3f0rLuUgF5Zk41k+fq9sLZY7jOdvTAZUxfKAZHzF
vXOO7DW8mlzdG5eA4cJN81Z5zlVo5gvN7LkJ6x1Mb+0A5fZdCI3aQI4YzTLbhnba
HHAZtYy3MbNnhxtacKhmELZfPNNsChIFPQbw2sBydOUqurvT8zGVYpnLNnJxbA3F
alVtLxIMY4UFlOdOx5dj5SkAolOwGS/Hg1D5BKUrlymYlNEnwz22E74Qg9+8HScN
P93GgMau+zioQ2XauKVhAM5Abs9jecEdZaGX4mXWp8i0OMGf3kVb+B2ip/KRRGQM
5X4wfcoNHsm6p/r9Snew6/N3EhnUjVSTlZ66mac329y9Tl9W51WUkCXkzw9Ablxd
yh6/lUmwgUGn9EnsQZ7+OxkQ208+cLkeR5ikzX4aOK8FtLVAi+jKS9J/e1hxMsBm
1nQEwiiIy4kAZ6xpiOGuyjnTMWL8sw3tPNqdA2P9ZkglcaIQydzypxZvJpqgx8eG
/+hR139V9uRC7vAxTXXILe3f9zhAWXRiX185QbnONRS3fT4+03JNuTATJ03AoN52
DxuK66YPOgGNIf6M0kiL7H3z6i95KlhmlXzOXXtmWUxOrzQHkhAaZ/kgaFmBsmFw
JCBTn63W4Sxo5DEnQolNH5W6xTq9c6J9Qd8F0kTMP4WNmykYMS3PUYgN31ilhing
Rf0WLgLCV0pJNZa5CZmNEB+pB7Xt0JODJSdaA8GJ3ij4IwPST3Zs9W0CRnHqosiR
U9LPOo+Ny5Q65cJTgHd+02UKFGpxhDhonEaqeBLEXqaVC2BUeLvLB4w9fmmbzcRG
aI5pLod5GuqyNJ0C0PAycfX8SVvSFMCkPuq05KPpJ//RhGlaTEEWlJGxFl6yOJ/c
GAdzfdRKwbpILBW9fLUxO6IGllMtQSD10L0/n++L9WAphjL9DkmAYi/jAYIIn1nK
MXjAUy/29oUz1VCP9jedR13VMmmX89EMVkupTqiBykooHkIncBivOtGxQYS/IbIw
RmRgL4Zq1OeDcd9A5aiKt4WhOHyPQY7nBgROqv21aL6rS4V8Z9eGEh1hmN5IUh8R
BYHjnsRegJcYXsE4DdE33nnC6I4CT6BQnnhwS/uVEbeaYLGeL2vXxoDHHcUIHJao
jBe0lnYVbSTHJVZwLP/3y1NAyDivtfzdk3H//Z4/vazL9k80sk4PvtfDbZLY8eKE
Nm9sTIPUheQ4mfJLD2ik4YTpeyACk9GbLoIk61w7h+6CQ9SLdrF4B4OOiTKpcbBP
MFVSVfjo9IKS0c/nO6+DX97TXP5VG046BS3Em7LMwfly2IDRMuvH28V12byGuBGu
OA6NLHyBLaXVQbCM/OCI4zs0qNrRg7PtdJoIB3kfc2m3fPuYVYkfyaiVobzkOkhV
VFdqmguDC+lML8KZ2jAplGs3QYRpVd2wHMLoSznJZ5b/br1AUbObuT6iDL2chZE5
9Pgb6xj4yT6K9ncnNbw4HocnwBcSfPY2g0w0/kTrJoba40h/hjFbcN/vI3GYWHzv
llwdVH9NC4FvJ3Op1dxEwjVZjhvR/0lNOZx+M6DWkLdLUiVLUo/mREqPVCNrKoYW
t2Hh3YDYtYPFdimQD5xGifnqS0sGtnJlAPgakzomRzkDAWdgpEz9o3uVQXSI50k8
K4ooYsXOwsjosNl4iIsVt0sCjJ9BKxfjaCvMESN51DEZ2pKL/aP6y00GqBCxxacH
5aSctX6zbQqojR2cn7sWf0fgT+zrfXnS+9XFqmJPvjuDYBkmkiDzMWk62sPbalEZ
GgHBlYWxTqo7TUCXofbO7LHLW+TOx0DL/W74LPLmvjPDtjLvOoHuPjigk96ND+E/
POrP4IdlZpNBW+oq/Cr0yDbE1bITXr/TPwZkYJKTJPCY91NzEFhsyZBsawfWADSc
ECH8Mv4CYiuyrNdZaoeRdn+EpKAN++OdwkUpoXZ4xd79ooEkBle814lJQOAeMiYj
Pjh9okcVFWmlVlkbKJQNhEfNg93GVSZ5j6laSuh4Hsod5J1iD0MoN2eQwgRAc4B1
NWDubMRA7LsTeHMYWKW0s6w6m9JxBeMgq9flrFM6uqSYPqjMHHlxqsLoJlUHF7YZ
EhA+mas0liEMcg3rUpnvo1gggCIgGa4z/KcVge0wM4GR3H2ge8lE1X8jD/l6LZJ9
UNNQcnwgnpHe0ASinJtz8gb/lWbhRY4uyYDsSYLh1ju/daGkVjE+F4Ujevm12Qg/
mvHnwkxRnSDz5I8a39oFCE7wpevAX3TO725n4W3gfHwLI+XCN4GhX1tJ8YyXu1rl
uen9y+MRNWpErR3Wt1bdHSi+lr0rwnSF6wHNeGlkZGRdN2tzwqRyP8Bfi16qj1mu
xjdhS/Q5UqbxrQrqBFDy/C9fUaKjWb9pNW/3je0vMK8ojkVIvq1PyVgvJoZXhAFN
+oSoPZvW93KBTnX2QSwmk17Y+tjtxUinEJJs68xE4FpTEwoKlEmNMvi3d22dxuXr
PYAjrbOCNcrR8b61IC+ckndtsqWZDQ1nv2F3fl6Fh1zzdAP7V66LYZDjVmkPPEXJ
ZdSX+pxCIyPiMxHTwk5+keKboiXvdeS2fO5MhSWrEqcfBnmf5Ll1f/lwJ64L4c5M
baCspRHztj5NHFbHd8mda2QRgnKYgecQ2ry/dcres+zPndUsBYqzOk7p7vyYo1dK
NxnSuJPcAeqc1SdO+3X2qbG7/hiYyBzncFo88lyV4Ab6yfxooTE8wRB6lEt4quMl
wQa2Ll9LzgVwfK7RCrRCYu9nH7vOVP3w+5XIkuGBug49ALScPGINdzOfUz/f+/PX
yvdDag4MWul0YYW89lMjMwihka+8vnap88Jvh4/O5NVzfKBzRHTAb1Na3IH2BgDd
qAsPf9p5XydBMTlKqMwUj5Sm1dH0zR2zmbGooGjf7dxlEk0OZyu8w7pKxiK5zpmc
DLWRwetVh4Dt26aNJiFDOOkAdzUAM3KBAqCSbo2Qedh0irRe031BcHP54yqlMx5P
2tb3QC6U4QtqU1gRtt6sm4/PlP7Mz+OdVE96sUMTMXfittBlMYAqlW/aLg22ZhNw
PkOm3myAZncoGV2M7VYkGEoqr7zsR7k3NxPXh/VB5vorZsJgNYKlPuI1mv6sejI7
2Qu9FMzaY4eXAV8LybZJEebk6j9KWjXk5ozm/7j7vZUXc8Bg6gfSh4WzTu5V2kA2
6Y9kMPoO4YNj1ZH2S+j0LseUycfRb2gtn2SajL4uYzmz5kHzgfCHF67hlMspabdy
kSkLOunugGtCtUL36Q8tRbQfudUF98tRL/rs0AeU9D7UhZ/052JJlWa0dnM7S9mH
56w5kkkVQGS8mm1N5tootMAYxkT8Vc7kPfc8rtcfw5tcsZNB/y/0dgWfXWjcAIJa
F13uhDk+TBg1iNsW2f0qGtgfewSv9Yj1RB/skUUpLeV335wRPpc737vPysO+XXvB
jD+twvYstsOQtQ9gXRps7JDLEKyn/hK2lmjqVq1xUFbAflt0uAnFj3W2xAbgydp4
6CO2psaZrjN9X1WLi70qwVK1nJ4cB8Xx7jYJ1MqFJm3pbZfEj7bDA0yvWVPYSo15
Cj5F5XuN1/vDpFtlr964wSn6Ui74SnkcbBn/2cE/lgI+e5sZ/vDzakg3xc3Ubz8V
1vXqaVOhrJc8LDfRuBZygjmEDMNxwRymebq9ls7UwEWfXFU1WI85V+hpxBMa1bET
e/T14fhgoj1e68wxN0teOwKl56ONfe6TJPDEyuUcWPPZ2logCGXuL5561BTsUA4e
C03Ip8l2in4E/712IJlvRRj38EmyPJ7y6lDLANe4iR5z08uFqujXmIxKCwdYoUHe
YFnaUu55CqrMtTuYijSzaDBjpCNS2KaYXD/564+kyhL3AgnV0b5qJ3xo4PP/ybqs
qAU4kh7skTpo/+7yzaP6BkgwMBoKVLpBMd8pogccS1hbwG84AxXnTALtnKsdfHsP
NSkkmx3nGKcbEzo7BQSFEPmckHLfS00XNyaoHKkz30pZg/z7zTIV5rQdbisJEobG
tvXoQ15bVuNROJtUP6JkRQYQeq0tSPi3QUCsKiPuExENGVTqUx6BqqvD9C4aBBua
cP2jDfVd8LdNHjTuPSIpTkZC4Mm/thSwE7julyFlGS5OHEZt09CBRfD43hzkosMr
trhuX4oJj41uWhniT3oM5caSKcrrrTF9ScxUSVUhNF5mMisHZyhTPyevXGiC4a4o
6wOm2xeszpNPGXBSCntoeDZZSY1ChCt8pLu5zBOW2yC2L+itYjzxX+d7OvLXqhXC
gTACSwtPHzMpfFdnLvZ5ryHbcjCYkPhHNknDNGZVo9oXBa6ChWS1XXg+XN4Rxwyc
Md6mP8HCk7Q7DU1DNMMGnCgLUgHG+ATNCXNzrMAW9Oz4DyZJKaHtuJc3eC6kgwt/
p4hFSe+Wa2msPGKU8LpBqp6Bp+OusPNKEUIdzjU2EVupvvDpn7swYH/hnZ8zp47V
2g58Fqne3HV0eJCe06ia3YuaK8lv9KNJiCWAJ1NBVFayWZeZKmVIBLsGKLCk1uxO
t37XORZq6CB2IM+hsTv5mu9aVY6WaK77xvb1qMH+fmTGLF1GgRZhcG7UUFTr9pSh
exrjjQ8PCdrfX7uwkXv+Mpwjr9ajFxjPfRZzsJNF3CkVnTfeJ95GovAJlBYh64JF
vh+urITCG2TnJ6LIVD8srikvFMHyMLeNKCMykJqA+TsK7d+LkH7QSPuUjKmISATz
7Tk2bZzitKxmpUkJP2pao5JF3HaxdYAMUxEX0c2yhYwEA1Lnc+yPT4Fs8AFFwDHl
sjG76QWsxfwC/hNWyXkNh50xq1HV/mPgApzTTio47icxMUsvfKvz7oxR8HW6aGeE
TYGT3wZootFvFS6jCXU9fxwvZ+BaxrVUhkbZQ1DoEYcMX9ObRHj+TKVtDDGiwAqP
FvvmNq8qCb+iSv7RqYT04YdTsZcBB8QEbVn/UzK8VMTYVEmxN8Ln19p/DWfYRUqh
Owcd9W43lwbicfiLtptRSME3NlSgJClzyISg+CFlFHDxpBzzkI86nF1IpdBQX21Q
FGJCe9PuBLU+ZdKbWb2otQssKFF4Xz0oUYRvpQg4NozztjFtB7feW0GsaSB7Qn02
l1en2p7vAipOa17QLN120ILrLOj6yvSQ6WmFobAGgZIKdOdDksp38apZPokKW2dB
RlSBTY256jebNKvvwx+gyRgE77Yk/gsfj6lN4IXsBiAQk2C+7UdYVzhhkqccno7f
5GunSQUUTv5DfXwGhIsaY/P8vO4Zx67m2XDCtoXhmkST4zCzkoyL11FiyldiPjDq
QrqN7eRwHcpc9MirVOMUpllC45+AY4a/geiR8j4XrRyLwMNPFPAWMivHoqkRGNZ1
EQmouYQ84GN2jqU4E3JM+TxsxhekuvG3fN39lY5LHLNmMD/uYSdcqBe61S2cBpN/
GClQipYuR/lGrp9rLovJhIZzpCe1qbhuCknraEPxsJHwLuKVP9aukpqsxwJNtahK
YQjTg4DFN4LCBEADnbadD5nUODh3rVTHd85gVPBRUUrZD9rtorrIDTnPCZrLnFf6
ID/D7W/jYgQZajGqvDSNYRChRpgVUC6oZmzieNIj51aszGMer6gvbeyrjlZkbdl/
qYVTJR5ofFo9X+SIudKIBOUk9gSolekAA5fNq22QHtFUL3IJWy8PU8lZ/Gq0+KXD
KbByKGkhER9Pg8oIsoLlJ+YElzHxT1fgT7nGZR2Oah3/S9IevlYI6DTZwccWUGvt
jTVDMHauUjBe1QNcbMoqRyZun6wtV8FVSBWq3ln1zDYGcOO1vp6nJsiOzhTmdFaF
PAH+pREt/UwiBZ/kQLLg8iVQJITJJPsUiZ5Dtbr/8euKZ+EpMDwBgpgTfM8ULaDF
wvGY6+Js7ayBOVKFveGecY+8oSSqJF2e8QKrCS8M905Al30K162m4Q+026rOk46W
bE233LVSHxjBeekFh2vYjOUuP6MHYWFEyo4QXFPmwsyEC/YPAgDJvr4T/A2Xpsto
0f5bfZDnAMG/oyf0lJXf75SbCBkmXKTQZWF22kvzuwaIDf5Rs/Tc/kULY+C9c47n
6n3nOWt8gb6INz++AZfohjsyleamP58/JFACWSwihZMwRlbNkLnwA5XRRTeBU8ck
Qqz0Nl38Fua0ANxCQGzk2Oy4KfLR3EwmmvQm52+MIzEOYQTZeHtmCFGUfHALl5dU
Tola2M+j6Ru9n8WEL96s0rXHepvpWFH4e+S2YYyl1Mq0nUYS3R1lLxMEntLyHVYU
mp0wr+g1xgu26R4uRcRR2on6Gfzsrmf8qGqal83eRS1oRxD6cXXu2H7DOW4yknLq
nZaYZNllAdrM0kAbwdVl/jOZyPweIDMjuMnw9U4mccoUaBdhi6194rehx3EHSVOL
3no057m8iZS9O1OLsF+ECy1vjfcNUzdoQwSbJCeFRmrq3Sq6tQpYNkwZ1zYrejEn
Ae8nkF63HQvIt+Q2cmAl5B9VBX5DFNpsPEQJKgnhAS3V9oCMCqtMrd+iUZIub8/r
90CwPOYO/NKbaEaw7UjCmxXfhZdyzKgtkNydu00QaPVL2capXMWIB2JXf6Fez6Bd
b6OXCoH/M5TkBLM0nPXDyo4FAIUrFaLkJkfotDNyCR7FT6o55ba8RE6DZUaMCjdG
7Nnz8PswTRmlG+3jSUETp/xAsX96WumjaFOy9k3+MlgGTiO7sEKHHQswdrT5ZRHQ
3lDrMq8mH2LO/5kwPU3mRbu2WPb296jGTvlEEuOzqsP5E36OFTZYHTArOsJ1tkCh
F95vLuOVg+GhakGwWQYpu5LVTymVzmwF7xu/90jD9guleSGOlp8SdRRvJcB5xru7
HfHffRB+UWLfUxt+uKa4SXE8QweBbTee5zD55aNXL1idnIQsIdm5lzDJ59ynZAlg
HucIJlOip5VUwZ8nOz/iIEkz6Oabg16Lc30EzgQDIg5G47Pt48m7uV1ZRMo+FGI4
dBZIoVUBtjEXBWMhdqnarL6g0rOm5esqValw4AkIX9ReCF2dBgvTTA8lFkVPbKcL
tAXXdccK5kMtWDqYI9+ftxwT21ToqWwgyUBPSOtlh3GwRHt4hmhh59wbpgVFbhJS
zV+bHoZNpwGiJkIXKYsQSTEgM0uahUbLWC9yqKGJrJjJiliSBp5QMLb8aw4s4JHb
01BC9o8N3KxswzVFEdixrDTBeSsrTqB66t7OSbIKN5Esr8swuyJvIZUVmlOqazcG
AcYYOR8jHcCKTtS7ad/u0SSrsVsJlD5wSbBExKZXBu++EneWwjwbQ+wBYJCqSntc
nydjFvigLLBz+/Urr57tYC2XKfH4ldZ2fxiba4iivokOvkbS3opIeAXVbKxelGl2
AinZ8w89gFaMTdubpD4Kyv/pNXIojfLNWCjsBqwzjgrnxWqEN/agQH9Z/1GOjqcG
432UJ04DR0csItzt5iahU+T3zIdzJVuySIg8C7sq5SUGnjeIFAMaHcoD8whwp2QR
it9DS/4l9+pTykIj/Jeagb/0O0IIlhVDRQ+ym/Oo4+SpZhdn+TaflWOWuc3BezXY
rAh+0rt0hIGslyEgfs6yL85wBeD4bUoKhOhw1bPqJvcbwjDyVoLO/bTYzfBgmb54
4jYZitUSD49ndR1Len5M8UKhP0B1PEyE4mm2GLIy8+MtnO0ewDRVmL2XHexG7e2n
Yn4XE1HMvMDWmZJvD2d17ocuEny1aDBTvDdhHvGF4c7TNh2xOBjw1xbusTqJKoIM
sSG4pPB5uHoYMxzTjSAklthUX/C1zg0tsqc/3Lz55TQ5CUT6Gi0LsH+dBJ47hfs6
c3MSbeYnawkMHIOZSXt53wHAPF2yDQvkpKb18IViz7wANXWwSj4Nk4KEBiXVJqHw
n75A36ecQwELqyZuei3PCn8NwOA9oGCm9kIgrOFKC7rmBtdNGqohaI/gW9zM6s5d
hXHD/9iY8scaAqVmN0Bv6rJoy2HPqTgFHTm5DttqhC60eyPjPV3eX8ENOCLv1PUP
Ef6aZ2cRgRvvIXp0ZzKqO3LLE29zBR9Tx/SN0iMCNJGoRd02M28/J/qS74KWymES
GuwEtUxS2P1SAeRgxkCxknL+DWvExvZkMaF9hhVVvDztJFGUHpjNkjkpy7iQqzX6
tWfcAVx2dQg0UUZ2pDC6XaQidXQdIG2/ygr9CSTRHskUNLMuUITTJFpsIgr0q7e1
pMbSM7rVn/JzkJt2sFCECLZWZJKskiymGhGmv6QE7Fz99iG5Doejak5/O1BD6BMC
c4BY/t7NcoBvbd6n5bbtGLugdR9eT4o07uGzl/sL1NWOysYfCgunSVs7SPlS8VJZ
E0TTGmPF6BQn2Voky7YUbs3FPD7KCxtA9Fo27dyKE+VtwLoDXPJ7lqzKTnY3zgoH
MtughhqVwFEsbfTRGx3HOv181pcP/R9WmgamzWme2iOBAD+9CmQBUjcsPZ6QvJX6
Xvq7P2Jnnh9saT5ri1xjQQI9IKlbkS/PX0jNOkhb34A1UXpIrfB9ySTLW3s6urVs
g0VcfPhPR4JrmV3Q8FdIbp53hmNbe23U9ZIqZGzCg+RXDSm+G4lKRYwM0bVFX1wd
HssrkgUSTLhx1+zTXz8J+nh6DEm7iNDigF7/plAB7QADDIcZAoFGcQu0NEsB7WTB
npj+ZsT45dZVS+dHBKUaVDUnlD9GfbePQaYJLThW3G5iwUEoSI/xQeNWNfeQn2om
gEYZQWqG0G2COPvvzwwUr6126xDMQNmmlxysO1b8zL51AlG9jmA4BZKaZfuk7j0y
IXixTa4BJqsbWr3/PKNus1pRd3M2z8kjOKX54lHU9FbAudFfrHUms+hhh780XfOF
eL4+BUoJA6qriqH0PHi2O+FizSpg4lUDMQJDjKVf88hhdnkK8V9UCeAwhzgfbnsN
D0hlx0ep4VbIVHw8ELA7XeU7ChaQzHlIIDYnwJV/bTEvJJoIaIdZLuAzgelzqq8a
3KanycuXaVtliD70VwKu2vLjLxhBhfntyYQjBZhIxxFJppL4fxJLIxaI8eo7v1mH
rga7nYULnbSrzgNO1pcWFFf3efjdD7Xt4qM8rXkpUbgTW8ALvv68Uy8gvH0PqKO8
IwxyxOse4eDgRo+eYt317zL1jAlOnq9aye98+TEKqhthDuLqEdkiVJtYdhcBpPGM
UZrxlTHqn05GePNthOuNR0ZUDzvc9W4LNVTV3EUPD4Qw0ZF77Z+fBCCxhmFqBq1i
Xs3fjNteoq0uUv2C+dhKz5AVRuo46sHQF8gGk2kLT2u4VH5QZu87emhYTIOw0MPe
wRC/qn58Xkzb90m+Ab/mNsQ/sQrAqt3We+zdSIfICXo1JYv59bIy2ddRtPXiPLnk
XWPepntaUCrTj4IMNpa7POQCl8d90IEFG9xRSTBSPU66OJh1X1E0AxiV/uomKIjS
lG3nGEnf3zGBe0W3zbIsS0lhH+6M4SyQUNCJsTM903ZNzcO5Nma+gMq61tIIhUhQ
Fg/vqFFMidXn6mmNPa/sLDZXJf4XQbOTVuoEMhe81pyCsV0Ng42kacH0D4fomKvF
/F+J9b7vdUGOzFFcmBBStbA1PhDug9ywDBBth0VGhAX8L040D2HfmAluyK2ALEsT
cW5J9GnR4rjry66LYYWx1HS7GX/tQzdGYa+3tNgi4ewwjZAysyNO++SVrrWQMhpX
x00v+/dgHTr8wLXejlOFvt6vOBI4PhpAf6U/gck5YRrocY1EtphOxw3kL5Xo/I20
yJGXBV9OcW25uXvHVRX9VSjJUxe4boRpZ+8cMgogRq9VN2K24O1BZVtVTrF1ws4h
e4mRADqSAaGlA9o4wzyYLGfWSfbH476yABEQV1j5LCxWdy2M5ObGfshkwHf56y4r
UCh+0bNQt4NYbYVisTeXOorZKgSvWwDkY888Oq0BEIcQTlciM3HnI45+xcw8cTrv
60kI3yzOohhm9EAcvdJQCDMuia8HxtEuyRcFXejs9eYU0npjFk64Zte6cu9WpjRx
xD07Rnu63ARu+HuMyDpCr4Bd7sWALtlglWeeCMsZp8QgmQzmpJXDUVTVU1sV6N92
kodVKL4g7k0B2rqJt44745YL/bwDaTw7SX0HI6YcWfpfjJ7Y75Xf31+m4iQeHHuL
CMuYNvdGAmyfCvV1ActavlLp680ueJ8Uk+9HZiuK1dRjtbtyNmhLf7SoiWPuWDl2
QnlrLyxRNzN4JIW/FxU/7Af3l5my5QRrLgFgbfVx/VpUvEz/CtyeGv9oJ440BpQ2
U6RaqyXRIZpEFi4NcQ9GQIpm3XsezAxUepTzc7PhAL/x6ABOWd+qcYrK1Lu6WhUW
oIK4+6KyPGB9wSJNkonQs4PEhuNuAQTYwFX8WtnheEFxFOZxMdMVjXvB5qbs2I9F
ofpQF/sJ+j2RDBPI7GdgLE3pvdCvPQ2nZ3PLw716UeS65PkGAPyn2GpWtz7TPOVa
XIzsZJUmHJyh60OpvF/1C+QvoBpW4KTqx4IbiQw4o+jwsLrRk/GT+hl1ynJP9/eK
rT9/KSvawqhkm3nhRKreZ0wRAq1DD5UIGwHM8tNUDokXB7EZwovsCuCw3LEVai5W
jO+LmeOxAASGxB7Jc4KxQCg6MQGEjytf0QnORpnCDje3esvFumYA1CV/ZP9y47H7
N6IUYOe8oE8Azku54WVLZ/cOPFEtJubtPQ90rv1mBQED6ZF44p5oxcRaecsL3FKn
TkG32Muh1/R7AGEwKGmNgm5NDJmc3qOLdI+vW+Kn9Rb8uGxISV+WWrihKa2euEWo
goJok1LN1/Yu2s6dJiYtw2rX6Z34PmBt56KihFqpiL+ST7R08lQ7Sg/mWwsya+Gx
YKf0qVWzNszsS0CoHsbBJ8n7APnXwdxYJMGCyJwMzUuzgFdh/XLna6LcuokjkdTA
xK/QsB8Yg8eioxypUEEVZWm48STmYSsOhRVcgZkoL8cQRmul/M55MmTwJ0lXydve
///o0bXKFZbNd3Z2d/njZqjl9egjlRqCR9bHHifrD9OhgpzKR1mbjVLmZVG7snvx
vneVNPuU2UvFA2p7ilYPK8DTSIT9yBP2/sGwX/rHL9qxO5SNROp2cXo3+qI0SzUP
wmViXGFyYnb9VE8QZKAZXzWHUGse8tL8Ip3+GZ3iQyZfeZ517XcepmwchR495/7D
qmZH4v1wy4Q2y0xwyiAd91ZoM9eGVnF6VFG4KzBlIxxzTkas1iZgt68o5q0Bsp8p
1m7E0Kd7wUrFfWe2Ck96alO6QTDaI2jaoqlMxEjwjR7zLS3SM7T9+vLR6RndFi8j
yJ6IWsx0OyBvHaEhB/TkcKB2O3FiqwWTpDAJHjReqxI5x2Unvjqgv/218OzBSnMD
vSNqZsgHauYQ8nGVnvN7PEYjoQEDO/8/eJN/J+83JUBqVMy1oigUfIt7iLFS9Bm0
grRRvmb380rnM5QbWnqn6QLv5gy+uAJyuBqtEMyt3+0nmetKWnM2WKQ7IViae2tp
eh0ulb0sYm+ERGfZ8SciGp8QsIvYPpsHr4KUAp5TykscyCZZXhm052o4ANDGxx7s
pUnIrCQ1nhOxqO40EDmw9AdaXCrpvyi0VTsZdjZjc3mYdWIcetV8NArQ/C5SalbD
ouig9OD3HoCtR42m1d0ALQovH48JkZssSjC/1zbz5P1Q+TCkXeWrox+NJ98tmEDM
QmBmZMAHD+s0waa99ruMz1zNiihb0hT1X2ruIqPWriX9IOc4qualRZvqxRBioWOT
P0rAMz8OusmgEFxVpGKR6K5YBH3DyW6NXLtZn3+T4Jlt6HsW9NaKEE8MbGaW8Gzv
3/CyusZdVfY2f9B624M9RFHjjkqBd7sJ5XYm9b/XMC71XIPn0IEJkjgp/w9XHnTs
+AtKx7Yoi4cqjNG0HVRUuWwcLut/iDMk3ppsueuJDmewa56V7Urme8QufX8etnhA
14iYqPB0MOW4PYJCnfw1ulOr5UdOb1EJf30nhktTevfMkrZOISUA3Yw7SLuR+IsC
6CpkhQccdG4L7NSyUvIFhWP3oaOJvnsosJ/nR/Dt4jNs0Ef+lusB20PErvzqc3dZ
KdfNTufp4z1qRdVYAS5UrwSCXKSFF/ouwwSwkmQjcOU+cr/7iC/qO1dH49pOP7UP
7dzrtqZVInCkWHkXB8ai8/WA7YIvhr1Yb4BFkJbmI+dvXaL7UsgOrjO7WpJlQmlt
6IVC34g1xzfoYuoKemcg+Hr6+tuIKEbqtRGLStIS6y+sqv8WkpayTM6qVRRmmbDJ
s7FdyjTBzfDP7kseTfGeutnskNVXLUGagsNmG9OA+WlIUL2OzEWdiQcJusm4Z+ma
mn47pPIUNeVSiIf/X792jM620naDrOjFO6kAh5S5uefqYYhEgVM02QwNrvOAHmj5
xZFoJlBWlx/s73UP6/wb3R+cxV2zpyfa/es0v5yHkA3vB8ct0LOnUNfmh00Tlpuh
UeBbXdOURVlG6kFtksJEZmYFE/r6d/0gVIaGZMYiZwc3XEYeD8sgIcLsIXUbBICd
kkC9wlcWlHpi1ykIljsV3QkLeZ+nXsirviWXZy1dpSzRpu17z/gSJm5Npf9Wwo+g
B5LGBVyn2fmwnNoR51rP4P1U0dQl7S7248L/5ZmmY7Ta9+fbB2Dtp9OF+kzVAj62
mAivAeo4QDafSWenyCCB8xz2ed2un6bRJO/7JKjdNxssIvmHPxuTmpnbWYunR2+x
8H/4p92HOAa1o7Srg9UJc6kAqlsptfP3qE00IbcybIqPJZrKAHnVMDuwrkLsZFXF
7x89jUPDbx7UAo3eirYHeiVGwf9oC6ktnawBDdPATonuuCIuwYM8QDvcD1205uAj
EX2/0KDRJ4QlTmPQoxTt2s8E6zE3J7mDCpmwtNDT1IG+NHDC1AEQHeFsaUoVsLhv
MYxZruxbwM0LLQPS25mvxxZ10eoudsFlUoLvHZKAjPPmjOWgFvVcj6MpunpMtWOM
ywM5GiF4Osy6i0mZZzwoPHdNqYAf/+uXb+8cHn9uhuQ/KUnKKtGRlGB2kiAjqCXY
g6sy3Z+6e9M5wvXM7AcB4iSSMZjzzz90WLNSv8o7a8BeLvdhaNaL/aI/V5luMyHo
lcAF3/fz8X09Ac3pX1lB3Q2ojtnsR0UJvt0TGDA6EDykMUR/rXxI1lVzsWw3Rrdp
UqPvB/IaogYJGPlxi02JSsnWO04efMgQ8t30polFiKjrVMGPg2sEEmoDgnvKe9do
2oe+wnsYkbxvBSKUfsSJY5rmpo18UlaSqDN1OXMD7tATmy34x8hd8ZTc+Nykxymv
JSmSTn5Gb4cwCwCjuB3MOJpez+IwlKY5lzeY+1h244aJXtz9pMCDlulry2XEbDgN
NlQpZbSw9lZ86o0gXGE0JMkSO5EMQCo3IA+JWDb/UHjtFM4zUt0pQLjH0KnWzLuJ
njoALnz6mdkR2NI+TgzPRC7Zk5Nj8tQ61FFLM6UdRtdpuI3MJPoVVKTVi5AigheD
a9uhT26OBDdvd/326Nv9qxDIFk6rttfFdk35jgIg3QIFBcokVjKNvvEWjUnTRbwG
f8UwslcoxsXrDZQhq1I9PHB73xrCnvFPMzqLzQaHGAlJ/TfV/xe7SAmgRijaWjCn
62DAhHuVy7+fi1AM0w4nQ4EwSVRN/5FM1I9NkRZs8IXdzPU9/hlq7oqJ9Z6yvJLk
i5utdhIms7BUR36S6oNWB9+H0B2QDjcsNMZ5/Sj4BgZX345vAVGlVZ8mB1aJLJRM
355+wpLhvqD/xqBaVeeh+rGEursi7YRAMjOT/dr1/FDu6jaMLNK6oXI+6qcmPF/X
te0ajaBnvRPmI0F05Fi27NO15e3B+Y1c1jgtrQ2TMHjqleEhC/MTZoX9O6KaU0Ws
+ZnkhKTXeoAxywy+n0GwPBtCSbbwyFZ8Nhh4MY4lKyYkimxDWz8th0mbHGkMJ2UQ
m9XnxuO9LHA7DGsfY9n1GAdfr7SQMtSoiA9NZ6roEyyA1lws29lvDuGSDz7RljWs
y2UlR7gXZqqdOwWBePkvHcP7WC5w3m77sHzblBmoGSvE+b+zriooAYxNqwxHnpkr
lEvdA1wvA1MaGSVyTFqH7Vm4TMqJnXlEmLk0du/X7obqzojkAQZVNTolbSZNLntr
YztC7sAaC4PXt5tYrO/x8f12p+z6EwypdGXn4u6YMka3SFQyvpzI4HFASk+uj57W
F1NOpped7HxAjHMg/oLjERnXFiuzSyM0oyTz9SaMYu7lpz4BIbDZaYR6zEB8HB0L
YFa6qLg9VDirnDaBCCy40yTWj4bQuZofwtgyrIp83eEPMNhhy7OP2RITUCsZBxgm
WB6zHOyQav3ogqVPz2nj5yCAB/LJgzRpRMUD9qm+roBdxRY84JBcBPy7BZzRhr4X
J+xM4b4Ms4eXmwPPiBmuAX4I5y8HRSy0LObWK3El4zoRpGOdB/yHuEaRUiU7NRah
NDkq2+QU6c5ehFFPNB7W7bvgbJ2Wuwe8d4Y0IhpERu5IKGfwUaCUXVwzdqSLQ8jT
u6oq8p26lPw5WEBLwN6gnYcJgYYaN0oHZbC5YH0zMeG3UsrBWPIK9LxbKv/P8Xec
5lryedoHYvuDBOOxC967xiAyT869DutnIfJjUEroC0mxp/4Gui6759DZ167462yg
L18+FHHW5QUh7H9TlWgHKWVRUEPGkXp3TkA5ekTkR6VGtV1Q6U1+ClYzKOjXmHi3
TZhSrlrsrHBfA5lqaNxeCZiLFXadZqiQ9LYDDBo/PMOg4k1iO8j2NdxLyNeY5kGM
KEwGZhYvHCtSlESUmshT+Z0fy4AB2IYnpSWRORvL/F6hZCKy74R2W/js3t0lC8hd
MwqETpBY7wRZM9Xup5vADaud/cerIIRv+EnKlTOkxgtn8XDq6zNrnUQvH2cjnp1y
2GRpNvnKGwqBrdt6X9B8MJq2BT/DlLzk45mLIzyepfOhUkcSdbpFyrnQRR3iUlwa
AGHra9ebtu6dESp0kP7H3orYipMp8Ync1nUBGudG2qBH3gJRBwA5V51hQgIC8HAd
QezMrvkJL9/yxnGb2O/eivq5ct8Xg8+mCGCpzoRm0JzN+MlI1xotaSTwoUeNuXA2
ZLg2+qb3r3RpcThzaABOFF1nScXlmy84HeFduE5LZlUGSRrqDGLPmFOE3NvCmYEe
q7rpSc4gzPau9+JEG2I+SeHUvLnpUv33D3JlGJGKn1uk0hEqHcdIZe4j6cu2b6bV
s57N8o97MdyBwDy+USVMchQGwHqha177gJMdZQ3op/0q5suyvqG8nPGNBUtvQvtI
bGMBZ1/z80motL8lBNLwJlSqN4RnQiuCcWBD/TU33XA9bQkEASDYgzY2PfUAxMRM
i8of+9uOIVdJukMcSsSnmQZDRpAdehSjUUjXSgZGqXiDXPFIhAB6TrXjReUHdLDp
/VOERAK8WzlRSdIkyLAf4uR5sUe6s8GMlstXEJdfPoK1is+vbKEf0hQ3maIfNYBU
OwrXjQTyDnT0hjBH2J/hxdjzj4OPGogmmFt9gNwL134XwkyZiofpntd/lmqFLUme
a8HhCs0uS3+IC7vrtKR+YshedZfmegEjRGB7cv0qGL1ZNqAtwSxwk+tP1/gMR+pU
oj9+y7Px5q1Cc+Il3Zi06q5GI7L8TnRDyXhEM8SYwDSDfUQ2gE1BxvdmEeM6Uexp
gzEO2IvlUQnaFQ4RMwGhgV8g46buAdFCAhuVy+MI2Xr8ioTGgTH/Pb+wbl1kptp2
tFrtC36nRx9u+UlOnxQY9fpQHjc1BrCo+kWQTnhwrBvudlbVwrqZZD6ihyLEWTKf
+UKjS6MdDeQZc8ND0yufSs+O61OGoW6swxzUut+5xy+zgKa0UHxCk5V65Q+O4gGG
eD6CEnS+7l+0WIsfH75iWaHp0W4c9zDjBmMlYku+Ip35zb6/MxC/fDHWN8m2EzLb
rFSWizdMWuaWacJg0YTQIGaNtOIjnUtOgIC9HVuGJH0rz4BaeJQNej3UNtmy+rff
TKi9HKFXbwCfyjL+bfrDY72kSwB01sIW1sH1LUHDp3aoHZtJpySLUhyu6t7olZnF
Qd75F70LVscMhIlG8bmb2rh+Q9SlKW/rSh3ln78oGnPHuCikwCEBdA/gRqysp6wV
GLbn0tcezZaLhh/JwiUj0QwJf/Tla/5RMBmW3szeIYHRaMAki+NmTvvnJ972TwE9
cCLtBi7FygPKVqm0jFy9OPnRo/QU5L8PEjbh/lpFxHxZWdPGfqaNl4E+sFH+++mw
6vgIQrYktjloPoTDKxWNHYp1xBwqw0wyVVDbwnHuLppxCpAVrt1+hKisdT6XtayI
L3Vt1w27PUWfIDreYAAU/74b7z+771d1oOVZY5d6DKRhyoADFvq9kOY7L+WsZ3BG
MvpwRZ9yuj+OFqoskFItSAdIbG5WQfQywPPyrX0ceNn01n/gfUCMZ7Xzp4Tsygv/
WJx71Zlc9IgwzSR0T0H1O3Lf79k3BXyBbyK8ncv5pTPB0prpqPX4qxPZ73TGal/U
4VWG8osRCXAfakVJ1ZkuPRTYOoEs57sd0ukdX6yNAklHngH9r3gHd2n09HltcSFu
5tgyYvEPQsxT13Jik8NXecU7u7l2c/lVQOEIn7rBsSnldPC2pkj8njglqcoKZjtp
QUUQpnhhMIfQ8i1bB/FuRbdwToQGDJXsPPeIOITKbkN9kjz6PfE3jpgDjP0jsQ0S
qa+Z6Uh68o6QsqkkpaCMoYSZIRac+69yNAbkLYyHyBjpSDesbnXjxhONHP1G8Dlf
bJBQ41KAO4NdZmnJtzoCesGeW0nY1d/SABvUcevKNoIQexBOkPMEV1szFbfH1otc
q5TMj9bLm4up1jWZ4Sn2QghcDKmiChuexZ+7fN/BnfVSlDPLRQdByrVbq5ygQPwC
auuKBvQRvKdhuso30opHEJ27cZzZgpr3UuhB/5bkTV0l//Xx2jQVGJ1F7B7oVKTj
NeTtdy9I6PZOKRvyOJSWwRb6JxOr/jW2oOUiHFSHbagcCQHbv6MYLdfZuBB2oHGO
7ZtgmY4GdhNhHZRPhKYNU3IN01gZFnW7tNYVAdA0Eaf2kdMh92fyAmA48rNzQ3d1
tY0i3EfDQux5pwpacNLuXqVYqODMo5fzYupvV0cODbGOoLf6NhBi6JPyFIXB5jLb
9mWwA7HH0j1PQFnXD9NfSVe4I6lGCkFvtgenhDaymPhkysloPqf8EOTspDpP9wBf
qut8b/xMsoq4DSukWh1ZjsTxeU9eWjpYmgzuHNQiBJvk9A712ygtm7I97lcXKJxX
DBOvMjOUI60KmMjUrpau25yhkMrUXvOeYJ+xJ7zOd97US7baGG0E9ZqIdvlDDBCj
nu9N52L/xP29zbqBc5q9dSt2MJhh4ZEPqykNEliqdJK2ETAuk/QRGhBkpHhOOg5Q
Sndd2D7qg+1YSPe1EydyZfTK+tTI0sBBUondppc43Q9yeE+9JZib87wAZNys2zBn
tAL71aQTNm7t3RIP19gwzK7uKdipJrpl0fVihjdSwApDKlxbNFgEh5ycy29UzG97
xpm7MiaHVQl7wFrK2SUlCE3+aZ0RWa66YLOKIdfxT4o9YGRMzEkx0eyMYGXOyKe5
R/83yE3KEpAe5qzfXAs6tq203RvkNi3VyIdXPuqRuzq4VNSklffRqTO3l7/N5yI6
/LkqH9TUlFEvZN/bR4V2EXtmAiX72Irf0MxPD+rEPlvBcP7RtZtKTaf5VxlGWmKg
GI5avxY1D0vnd23xXYyOjm9VnfTUUe17jDGd+vUQMT3eA9WheQsv3R6Bbl8DwBmF
urdnRW7/dCp3tkdBO33E3mR6nB73t3LmJGCTBr5LPL4/wDThoPkZgTvJ+9EcuDJv
7LwcBA9NH/INsHhoGdEXoxKti1YzvDmT1cSRgTiD9b/52/fUCdg9FAlPhqxwqnbr
KzmBHy4ZYq7hoWRk6tlmoI2MvWW3HorpqLeroMspX9IyX2ItRTnso1RwXn2R7qHd
09IBNTPhC+8N0f0p4gSUhXnAdyX/EF4y2t3ie7yGunQnqVGhiwXTtl8TmPMF36BB
Hue/bjmRky6MmCWaBUmKO6H/NTSABNCSsjgJontMxuEDjn4o35uUyAd1gvnezJAM
cXviKh/QoaQ4sHOeHHmH710VdnSZ9XhWDQeIHoYCm7GjQ4X5M0sIM4FAPCAj5/Og
HkbRtC1A5AKH9AHrzOlK4bOa4+aT0/V7xgcN6qE2ZAuz+txgSPZH6l/kH32eEwTk
aeH/lFIrsWwc/fgpd1t/lNkX8A6iju/Bgie6SgBEftbOubQqARsnxUAA/22ClJAF
AoEPh9bC73K41PO+rQVpx/vWfINc12K/Y5QJDZtTf6ZH/+saFneXn6rtX/31hFFh
zZbcUEX0cS9VA4fcc52j7q06YYVnLx0f+4mYt1DgmEEzvIVQdk8Gq0FLC7uWtnDv
hxC7FbLa+l4/drRieef71VT60wth3D8Zq8244dhf2LmpB0cnwZHv2G3+nYJt19+4
e8qpM3UFDO9eED8MuaTkjziBQTeBRsjTg5AludZEnIYRNM0CB77VOCjthHOfi1IX
apixFtGWRxkAdr3cMoSZFl+cQ6DWT03NObkLQ1p66HJlvylEpSNrHiKuhyh/pwEx
b03f0YzJxRaZSa91GvgCC+iNEJJBQQlB6rI3f3iBvovZTYeXXW/4+vV0kPojN1HN
VB8We05gvFPu67qgH8laI8iSM99hImNcn/CdzezBhYZnPV7ACw/DmjSZAy0W2oRp
FgY88wx3Sb82EnaOs2Y7/bJQdoggRVDur+qc6Yd2ejnbnNP56fYUHOv+arpEmoMA
afxMW1wNFK8Rcxadm0zIA78JyGy0fYChQwuMSjLcqpsZErUkJd+AzyMVI7DLSQxh
1zVPNw6EQ2e2KM7TFAh2lxdOYFQdSJPZ8nTNCyRi6NIPRtamwhEDnlmSgyOhVy/0
gc+ofSfj+Ml+kintvAK9Ums6B0bYIxDlbvEc6iWWSdJIViuSZP5jXjrpUlb60fSx
3FrxDtctwTVyAaQKuesb3tT1VjV7Z6ZQ0XqdNbIwClpHgjk4kNTDWyOlX3D/q1Yc
7ZyasBpsmeCA68VMl3s6U1lBt6TgRLgElB7vz+fDEaCPWjyD1Ew+CEjzQM23DgKp
OlNNktQcVZLU77ZOEhPRP337SiFmKQq3hghIsHayfNzcncNik64MsPf2KlJBVe5h
izhbedHSBF4eoYVh7z7HvSQhKfR8LXsw9bit5uwkDKnLDO9i6Gu/9l1g+uemUFP/
7lsl38Q+cWw47Vyra63+vsLvHv8zO6g7NXmUs64uacL0qwgqf6WDoXo7li72kVKt
9T9VA3632XzZZRkR/QXQeagjmT9XuqdenwnG88ecyo1gki6CwDYsVw9ijXCl3hvt
L+FQvRdOhlFYqwxY2Aian1FuKhNERKGlaiEDPYa9xsFrA0mJPUskHcMUjRqohrPb
hppifdpG0kePkquz+Eig4peNUmlxJPJbGO6/JSC8oNBo/P0t1nPMtNbKZgV3T5Cd
cIZyySWCGYwNwO3h8HomsB96v7ZmDpqF+mayU5aEu/oXtA3AxkkNFQaaaLF5xobS
eCPiJ7e74awfuxTkoJruqQL094NN7b1QnMKWfZ/1fli5ZSY1rEruTYKVwWmZivnK
vxFzRLGYTMiSAJKoS6qs7ohL6AhyFM5rHE3hrRmuPu2l5fwelOnuXbePTRf3LEJ3
KxZgBMpboc+Febo7G/ifsRs0doaQpQ5iPIJ9T6fjatjbhv+BOJRekkrrVlHBG3Ye
rKM97WWMoaIOtO1IAq/n+evLCZA9kTywvHnTtJUBKrsOa7rz+wghy5xGPRJoLU22
Hdea2JJpnZndmnRMCnqLsgxSexq84PaRaSF9HKRFaesYDXIOWGaCg3PMIu2tzdSS
c/YLaQzgHt8VEwVhBXpE3zOEteJiP02QRbYxwq3OmKCu4xVJB9f5fK7Fy+A+/jHp
OHD9I8jJW6BtXzaBscsOyg9sPKwWhTEjCfbCigqCu02rb43XN3yMbKQ4bdbMalUa
2uQBQ0GgwnnIvCOss1sNA+9LsARG2PMXXOsUEaTK+QLZdxwwChKPJ2rkePzk3wMA
lnxRXiewI3gV2HVVIdeeg2edWPj8Zq10P/1PebPSBVEVBeF28kIBAG+lwEa9C/iu
YN2+n526aBBbR07nb9Jt+FpUdYeWWd6FrgoY5SCqkkeWlbMFF9np2gXnt5LW/XbH
EFHGjadWXA/28xbyliF98oh5TESaPBDPsUi67f7ExIUS8srZhuU8I7l84jzQHi8m
j+sWscNLZ4O3zOoTGejw5SmNlbN3uqCWlHSWW3MVecQweXcWoi4yRVwl5ARGUVjR
AngBddWIEfY554Jx1oQzAj3zaqqfrG8i0pdXt6qeJbs4Tt8T2YvHcCEObf71xo/2
0FB0KHuyieDvJcGtqyJgqc0YcDBRQMhB/zS2XfD1eX7zsqEELRxGgB+wJuVFQHVP
2Nbz4ugVlXWNEAjGwMls7nRnC3iiMCtknasDDbY6i3ZS8bLFry7vGK/BsXXd1I4R
6nKSlyQSK0Mwy0BMQ8jR0PFlCGw2wqyUsSTipS/nhuDQt0MIdZfmZpbNSL86T5cH
uZUbHgEK+69MJe7+eZaBz7o0AuJStzZQewHCPDrL3Av8OhGjPxYFUED5HauVmzfF
uXNdSL6tjUiEWXsoqBsAGM2gpsVbZcalwezYLSxmMNjouICnR2cE1FIoncbIlJpJ
dRjLCvkb0Coxv6f5nhsJrerT44d/x1rJRU4g7dqzYpE4N2LxU93aEaT1VDQ/cH4W
lkGZxJAYg5DGbwgg6efaCzPp4a6oONsgo93aDGDW50tk0kPvHLqpvJfJIQTnv9QR
FrR45qkSDo3GdD+A0QgaLGL6Vsic4m3cNtbIIzpIosaeN/pDeOLfvxMX9vRUWyzW
0x3ERxW53v5yfUX9Px7BmD6ZIgwTNG16fotY15YQy+5BwMlLPHU2fO3pE6ROduoD
hc+jka5BXCNZaWHoxAn2Ky6HjHKy57iRhoa9xTyTmxMsv6OT3GgLEefQYMs7YSrH
suzS3WYPZLaedW0XxIrBgvyPzSmV96z+3PiMayxKNQwQI0J7xfvwEeG0R7ePQru5
A/PMXC/hHLxPBegi2BtrPSbLErpTw4va88hKJDldDfXdH2HiR7ZyZEDFGaveF7nM
vhPvLUccw2lMLTMsGNS0BqfnQ4Q7A3gNHwM5522YCvW7EUoyXwJzTgNaxggQCBwj
Bx+rK1sYgAZELg9rrT0gSk1Tp7JInMgEXZjKwyC9e+mXhec7xIq6kMges859IVIF
Mw+idpxz13ZO492D7ebn5yTLAvFCADmQPDz8Si+8b95NkSNS4btHvSWFJWkkAfrI
Ii3lYYMoNyJdsmP6hYmfWMmNukjHheiMTQ1a+ihdBPWlkB4ADMIadKeL4Sc/xJZ8
ECeCcdhcamTw7cHTaGrEKjEd7Jidf9zhqx+F9GtZvGiQlKknwZaVJKkzv0c9bbhc
qfrPLqT+S7roggZ3pXVEWngN+28jiQ3FFsKMLOuduGH5S1lDVO05HImSsxsb4HJq
xb0ttf8dg3VBVY/sbsFeoiMmpPpLQF5DKYKfPyYBc45+8BROYvNoiqdOQJNmj3ET
9sELA5C1bLhxvXpZ65FtU9d7zbprPYrWJahHXCeEbrtwypc9Zv6D7dsiX+mp3Cp0
8LPV5tUJOVH3WxAa9QrV+/icFqzpkpHGer6tUbMGmxixv+bK5PG7ovLd8E39dfF1
lTfL+QAbgmBNM0GO6f3DEwL0RwMcp25NHgLURkqi+QTSyeju/UNBjvghEoH0RU4U
eNbRj0AXyJQijBkjTI27ymP8A+//JpILyfkw5hb97Dr0Ts95BXpSPU8nbIYIcVCC
KjWUHdJ3kWFzi215HDgteSFcvXuDHj15/zGh1ulThXo2SBGn689GJCpJEc/qHh7M
ppIXztOxgkdBMC16VT6tps7RHU0+Ggv9J7y17hK+wTXMvEANc4KRdKXKCm+pfA+R
vn7sBj7zls//rba3D/C4djovCJSR9oxvaWTB6NAJohxYvJNCdMbgiLaYkHpdLdXb
kIRTfOw+Cef87eOOcKSp4UmhPv93ZvtMdf9u8mfCAHppCS0h9uwBU8Sw33e248d3
kwRzpNWZABK/uXnEa+HrbvvFt5VJhP8DLseMyD6zbrBxmrJINCNQPxVQcp6WI3FF
RMq+m8LrXaSG9rSK4O+6RId8ozzLgwxibtte0/ckuAXrWmED8kOHAK6o4wf8MOC9
k6haRbL5wsZTYfDxRXSdkhuiWjbtUh14kD2mBNl/4/Ky4atjQFZVOP/kaF0QCsdQ
qNlIjqgYhL02M6sLyRPRK3OGTn9wzyc3F8J92VA4vIG9Iv789kuNgG0qAexsfiXl
TuHFtdeww6LqFrzok5SBpp3Kfo75JHHJliuluGSZmqf02aBBxj9nRNflX7Hi9iq1
Gq3uS8B8x37TOPs4nJrKrXyUKCH8Hz0oovwyEilf0mHCF+9Qc7Vv4vFGUYDj3acy
2Bk2wkBMEMw8tOalTSxtprIHjX25d+He5qD1pImtFdncPrdUgnJHCreiRv7dhfar
selhkM9D6Zt+PMspj5wcGpRz66oxnYLq0FCDQ5yfozKnzJX9EvIvn3IQNnBTxfBh
90EJe+EG7cO59bVSC6UQaAyA36+eDTga+wP3N/TuAMZeZ/UpuM6JHWCs4P9GewhW
+VWAMhqhcjBn4csBqofg0w+xoU49XqEf4/Li8yDSSj+vVtM6KAeYqF3uYzq983ng
hhuIBS+8WbR8RhAogQK5L83jo475f5Tk5MZ/bXeJ93Ge0llI19Stpwz1SAW1Ry9r
siDn7OlC8PC0ZCynjg3eEvs7RV/+nRJjBLv9XLDT/aZsX8mgpZVzEtPXKGF/wp9W
T1C43vmSg1hHekvQR2uDH7YA7WuEFH8e8TQYILKNAOxGhZ2AbuJj8XVgknQstRjh
SZ/SiZhn0CaGmuUqFY631mr0JlApniHhPnlwoE3Kfm3f3+LYFK/dbmrE0o2S1H3X
i20NpCvNQgG961KUZiUrmprWntreE78wi83D9sIhrYXy+oKGeqYQqfi5U4IWEoKH
QnWRP+vXsmgIeGbQIaP2u8WgT0RKD5dW4T9Y5a3tH9WBLuPmF4ZhqD+H2P6w4dgp
noFaqVRQoIdmhMh4BA5pqKkLFvMUMBTF2871QfqmmyQ/YhJxo/HQ9Rn53Ccv7ezx
eysRY2czGWd4OPJjlKLTYqnVtQSrGzT8/lgW4buQ0qWthnJ7q07JnCovc1AmGM2+
OtKcOSV67HlVHTsgG72Z1cCk+RDn552FQKsVaYNT4tEpw239fvfwo+vMIdfFIaxI
UPIkQfTIGwjOUIU6N2zUDJWVQ8MZ7UeETd/Ce20XEWJeuQccqDEptBlvlflcN5Ai
X13u7iQiqBRUxzrZDI4EUs2EXnBEl4FUjnLNVUwM4SgWcj6QAPwkgUj1G/CG1NCa
0rblX6K1O1c3rZd2t1XNGnwzIBuKS088mn3BU3pQzuTsOxw6rg5+lATNafcuL/CF
wZbieWbJcrr0a7HYv3r2zq+/9c9RW80gtWAwEIA6BAUJWha9bxnpSP8Qf0REEem4
+aopAj2DsOFE/IFEIXn6bLUjcnZK4bRu184ILxknDfVj+BVFPgosnyQPDh0eFCt8
6BuV1r7fh1EBZd9bJaCbMf5zoqx3Z/RI5cG647bODT9DaGseRI/YP0DrO4ftc6xi
+hlS3cpE7ZUJgKaocB9d2MHbyaDtG0MxT7rol+B2BGpXZLS2E3yo/5W56xxTL4i/
LfDaERTpzcrOUl/tr4yu8n9azGErqO2FUNo75BBeMJYIMy29mVUS5b8foLbwuR3v
nL2BRKLxbhPGsSDiuDxX5bcW0iBj23njCv2C1ySPa7bmsZ3TQdd40JYwx9mbkdKd
qb3SJIgzLGGZB1zsM/bUaUkS2JdIC7FraQiUCdtx5EoCdBq2Brb/UiB7NAwbgtaA
+Cg60G+ZoOgxcOPVa2v8cY1Tv4o3xIREXiiaEqBV1I6VF9q0SFhrRGpijONrzl34
SBqjOubhv6i7zwn+gMCr6mrda3oUBucyadN1zqqE0kYm1frxCRxWXPGsYbArvyh4
it6A32KipKNXDuhswxMFfCSDkj5a6lCHlV1XAaDKwmh6TCtsmKaM3r53VzUaAMgZ
phhKUlcaC541Ehz4VLk+szGym/D6BFo66CtiGlaei7rZH8/tuL79eTW8VFQzHzV0
kSl04fIMGB2To7YBSms8RLRSLi3w7sdrTmRHqDwM9itBmSvjoBRiujfYuOQLwxIh
gmPCXyg6RHBcw7Xkq5nscQRXtTI+1xdXcmyg552p86g89bzcnjGzGSKVjHOW1XoR
wSctnz/LyZ81LQGW8vtAU947sDl2vOZs2bHc/7bwqNLe3Lha2iN5DqlhRRNObw48
zIjmyxjNUYJflh9MFulzLdeE4X9EFlT+iZUoZ/3N/Do/8yW2tGi6I3KjKTJubsME
bNAZxIW+MuH7GKPbEsnz2Sj5w7Diie6rzciitESO/s7AYf0bU46b8yAy35e9Dii1
+sZn9rPfiDt6Y19ZHMWhi/s8VLPaHLrLVz5RZu5wN0UfaP/gMZu9kc3QtPwjjNfG
VhC9w8aCFeoqSzZJ5tpW6/RUJYoPYDDKeYk9tcP2PFVbQD3fxdtqRsdwI8hIElXi
8wGeJ0C+zFz8eT9slTQt4GIX96BwvlfrNBavFCbTaVoagmHx57GtquDixmQTmDQY
yoLUd+DIBlvptwbcly5CTKTXmtoz8DDcaw4tA6Pn9ILZnnm4dvn+tMTMrpKRnnRv
/ZafqD1FVnogbdwh4BwzosbnDN2/htOB3MJY/juU5aTD/HyXK/L5rJUEcRN+ASzE
Hf61KEVwYEvjTrmdbqLmWHiFegqQfjaaq12dmPmflVkbwHhxWhMbz37ObVvWFAQv
QKirVlsPyaSP4q8b3eMk43OwyWCQZK7wFS6lxJ4Vxelq+QUO95OVpl5EG1l79Z9N
ZbFkcwQxT5ShqEFZyiWDCk3fNubX2qhgMvi7TjJJcdRl6Nkh2wwfpIhR/pFc3BhQ
5PQEvMxTCToCxWDNX0GJKMynzWX4MMMh0TPWLx+APMibMcussvrdIv4ABSeFPp9y
JUZQ16BaYtyZQW1WdU7sEjnFBGewrWh4QSesJ9w7ly1Zs4nvYciZpkYzSWnGirrn
doqdfekeaL6KiOvE3+tMrv7S4voWJneOwgaIji0G/eDI4wGEBkTlTARepXIt3Iof
bT/vMq2cp494Imlxi61M0AhNnj2bn7Z9AGOAahp7hHAumbh35etP7CYowHOiwMoM
fumngw3zFkJrD0rupnIn4BtI21wLR/JjjFdqYu3nps0IKFo22/F7Kvs7S//6/ttv
HcdKs2T8nA2yNI46OT8gDE6rRapdur/AxtobotDZAjeTtosnv9Li03cpr8FaY4e2
73Cr23yAqfsv0BU/Go5at6eCEwVt9/5FgQv1OEeMIw2VpxnrQIOotxWXomy/G8Es
FzhZJplAkOzvgvfns4uqcZ3bGUUzICBUP8X/d/lTo1EVCMyKCTKe+z1Igq6+lTX9
AeHV34vOLRX1HNa4AqwNrOGxmrN6uLbqDr7aC+Qq5/wLgcIna9v7rqfZyyNy8nbD
zXBM1xkyMzV82GYY4kLb0SDWqdBmFmDjXDcgdasDpQOspp3QjS9yHMbRvdtK3PBn
pWRuOh7cknpboTcTACP5QLT0YGf0PDth94TUZFVoj+T5DbGee6ZDW7lwV5AICzcI
Hgb5wDkY8BdMiWKxhXBw3kLBOAHQrlVyN+TmMfVWX35dM5KfmjdKqlFfVAaSnVTC
bwucfuJxa18vbCwxlP5DonEo/QV7FugHpbuK+PVr8T8mgptkS20KDHdOIdxFNzkI
d1h91AKDInk/sXouc02hR7qGtLzovd8AZuECDtnSq6de1azHHraFj1vBXmq+D36R
b4Ax0WsmCkO1mL/zgQVJwq6k2kwSzERefpfSY2j1gZh8gqVMb3VudG9ght66kuHq
KBEfLENX5KMSkNDLSWPBgAPENEdkW12a9q3eIGRNFBOb1/h/ylALl9PEqrvBpXCd
zn4MrmhjwMJg3HtO52wk6fI7R/NoWyUouQqz1ByX5kIG/CJEQ+F1/okihnnBfqvY
eT5TlyA+aso3OCt7A/lrGOsSdp4tcSj9WgU8F+0jcrBMnaPJtHq7gADFJyq7Ny8B
8ZciZGpUC+VnSLLmsl6g79+tyU/4j106fMO+hmI79cGQ1WrkJjgKX9r1QMoxppzG
4sz7xpyxf4iFzseu3fixNGPtgAg9MR15b/X/h+T7oQ+Oenw18swB9HaGrruDcue0
b64gUkPD1pJOrt97Y1dAHhZYjShsZ0HVIKt/Ltk9M3ssPVDz0X5RQf9cCrDbRg+q
LgVR1ww9WRuzg8S1SyL8W6yqLiMgdF4t5RnnSGCLTLORM/W3ACA+yXvGioJl69To
niELPc4471EUXzUSUPVkeoyxdAkuaDLbJMWUwPfu2iamr6j6fvxjkro7RYgqlIqc
nC710G6Ee9B5jw/jEsdzmyj7wxv6vfEjH3CflBfv0lXqPXIAgad2viwSyHXboKE8
pzJS9+jGgwhDUr5uyKZpTJkmM6ARw9VQ39ahn/+hZFRPfyCUicfPBDJ4DkYnVuLq
2Hm/k6ECDFlfzlEgT0a8VoOepkuQCS7gjHwTzvWXc5cFMmgFrF0X4hq9jHoHKsUR
c1tSQT7zKmeBXSHAH7jVDtYKhZyVFraJsu9wvmYwBqRg/RBnmj0lep7MVhWVUWlU
XH6omhiLKLoQVjqruGq2W965CUhHoiX2eYDltNPhptsiZrCNo1y1HssxJdSfgS3r
X/0cJIBgj/U6iICjtkWrUzYlZ1eAEe3B9Yc9oHT3XuTaaY9sgCEOx3QVTYT9Q6Xx
veoXNGs6f493gWYpukigA0AhaGOPH43YLX07y19vxGkzUbyNl5GYQBMAoPqctNxH
gXd5R0lY23zqYAlz6dAENzUmJW6JUG+80O+sV4m1yEwYAMQtNBsDm7oZp4HBdFDt
WSSD1BZj0Hyc6d+EVYutaU5OCPaNJrB30Z/QQWhR6LFPaA7uihW7gf6zQNLIDzL2
ENU66TOJLIdRkwAyzax3AK5xuu+VqPMGoKlWrKJXpOPI0C0+e0UArI02QbYFuIpK
EZ3p3QJA/EYzGiix9PG0FySXKJxplJkf62lVjvh3sg0vt0soHhXkZ14nszoY0CwQ
/kNBEQkcumHsm9cgNGDrk5queU3CT8ZIFBWiqvylLyRtfEr7RjscbgveecSwvZwh
AOyG3piuT4Yutm/N/ht5jNYY2Nm/3xPjsweFbIruLeFt8PlqNs4+UMa6zQAFsOia
3sGsMUkRTUmyPXeHrU5/44sRFP7vHCCGz+ps/eRS3iwVkILVP2p6uGVyAhtC6cnN
i3IF0wFDFvWrnU8G+gqGoxGU+fOBFdU/TaZsTD9rMhmNqdVLkg+mZwsfFXbePU5y
csLv/yV9ZNjZriayPVeYTMXsHbgPh6sHvBMM2kOqJImShau1r0mrYnJmzyjyS2Mo
T+uIjyIDKvrcmafgRdTLKUOjm3+5RUVl48LcYc48nqBn/DsiFhD3El5yBCDtEaEo
4DyjHFnDj04IQnO7hgUR5jfiFBYVBRdvX8IGttp6wec0pDJ6aG3c7SL30SXAfcaE
kw8dqtdLJ1AhBQKWmjDSvW7DYGzqJz3c2nfXiH8xkEShkExeQALXEIClN8/aw9XQ
wr84/Vda5TVXIqWOwCU6FpGWL2aV0h6mxylqNeDQGlzgKwF3cO9HxVMZ3PejgJim
LyNpGupQ1YFStE3DJ7pl1gT7mBkhZwKVvY80AEnF5lM5Tur29uXF0vhG3i7nWw9V
keQkNLN31d15LWMIxXmUBRkBqddbM67EnPzEstBpH2O8sqYRib4MgvfwcxdWj3U6
/b+2gqxx9B0LountoETLMtQ9bpZLZbQ23hLkaNsCBsQmtpxg7Gpymae5Jfcm/52y
TDr+xYPRniQbqNfsXTMtjF1F4RiKBy2ipGVdHg5ysiVrcgp3m9B2cn828wCf7A1i
ijCLgRTL0EQ9DI2URzVX2NGJOOxIUzYzPJkLi+4HnuvDUjmQ2GFibbg+xvXTaJxK
hVGBEHPJP9ilDkn1NTBb2+fhH6upXq3TZJagN/5yBJnI33+tt4QNnzkKtTZUKPnB
QcB2OIwpyRJ9Bd1cu9xrVNmdEurAbD8IG+EC2KHsRXuRx8xoYgE18T2+mZ7E+Y9R
ZUn+s2VqeSd0ZMlqWihvJ0IDgmvFYT2BTxXsiYq9bZuYIXYM2gr+fLCtibBZnmmA
ePnW8gtedhb/vLVZhDInMIDv+evCCkSD1fn+mMDW1vDR/w/vdqMDs7vdhYL90h/d
BP++Ixou1uNTezzfGZdDHFF2C9aSwFoUl0yESfLybL3NtRJhmNrPbXdkEu6qUNa0
4R8j/d02zxWAfyyFmuI6ir5ndseNETni74w5igwgfBtzcip0xVYIbh5LZYkQzrsH
m/E9mhjKIlu2FUC1RamU01BlLAxoOeEAfizQK83NAewup2yg1vMl+TsTxT4MMROu
NvSmazYytFZDPRifQMtWOlAcp5mmbjAwqFIc8YoD+lDUiIfvjVtvnx4x3fu+vUt4
Mien8HCnb5wDEzdXTBlgMVAEI7DAWcBb5pGdh9BjEqcIaPbSJTGxZCaGyOHIUyhN
MbI44g6zWgOzXtSYJ6Qt9hyFOEbxnVWqlPEJBAFmFAZpVmz1yKzxxwrPyDS4pnmR
Q+hOmbsb5u0fsPmCxr6Zch+UimegIq+Ch9cBHVb16eA5ZcI1CUhC7o15XC+LhbV2
XhM55Sepdnie727iL3WFDcX4rZOehIE1epVCZ+mA88Yl1Xw2OZH/QZEO9zjArJrT
ga1eXqLUdiAzHTOummxSUMb2BEjEiUfOTDn8tciHuriPE1u1vSTc4dl0wpMMcVF5
i8QIrfnuVv+Q6jUHKUJwwlQFqCNrZXZuyF458/skZ+oLyefTdILQRWd8bqFz5/UT
x/zCuQqpTjN1xGFpKtmn57BdMd3yz4fhpC58Ee7jHfGigHoF8fzqZjoqkxThJeAD
b2JjnrewHYZQ9YD7GI3CsiFXIR/2IPneG4ey6PRnWkSjA2dgcNM6WXW3BQhSiDQA
97UhfkTeO6VAOnSrrXwsWUFxZAA2lAhjfFCxX6IMAqjtZmCWX3vRcsHZoWaNTu7a
v9yJg3rUAKnYxoLWviFV4ontpDgY91H5QXI1mLzOmpLxfgsaMKIw6AViETqvC3MF
7ZHaQSAREo9E5G67LqCUFhuA5bTb++q+T5ECfD1BllUksYSHK2liPeVLY23jTmoZ
5NCfBnFtBmjA0mL/LiK1pHZH5zo1I/HnmSBxY0MVVpJ2Ui6cnWAyL613kZYMvsNx
03bF5trI8i7k0vG97eFtS1x/ORx1eEYjYZh1u4AdIXv4MHBuS8byxprhXEeI18kV
pbUKDWBL7ma0sB0ZObb14PUg/dsGVODmlQc9HS4ww13uDQ7wDDJ/qcSiTaZpLMvc
Rchc5B5xC/UN3vi/bBlWIPo1ssHKJ9DA4jyF4zryVM4PLyymbYpZ0gtE9UulXws6
l/tYA4u6aFY4o48cqiP8zIA/NyDKRHBcRuqNhgDE5mJmE2P4/Ycy/aWGYRHULQsx
FSWml+DsLxwpYl9gQratoTl8H94fazQaHtx7CC71KC7QNPlpIqUrYrhRYZIn2Pb1
Fh0kGqFCIKeMT3cMx1MvJVckRCid+9iWkAVpLdRHiSRXexn7lODF3z/W9CaUEg8N
k47JQsyE14wJVpCiHVLallRTcWd3sX9Bgpdjmfzu0sPc4B96LQboWikNykTgULCg
e5IppHKErhjMWV3Yzx9AskCwYgLI0DfIgbj5SqhWB89mLeX8Wwm2zwDhLiERPqDw
I2QZ3bjHiU+PTrCq4XEcS2sZ0j6r1KGhQwSzI83+FUF3hCFN9UCOoHxn9ElZCYk5
jh6VkL4Su6idhlQLcA2h7NNyNvB9Yz0PayPQVFmlYK6Cjwb2W8UnMBqYhs4QAISx
FKDXWTtg3ZlViL+A7o6X67+q6qtz0kW3OfdWqq/FqAAqEfldpkHuStSVmlYBxetW
osN0qUdxygRClh5EOJlg2mzEexztuvUHF70/T5nqbrDOG7g7s8TEmj9YURqVIuV1
/41hLJpVas0TgX+SnHtwS8A/mu7KxjxpYaTs9UpXBZJTwTAV6T3dXq3sH6sjxc83
jmKyfYHTvLGlX4NNA0VPg6WTTP6ubNKQ36VU0y1p2YjehafaGy+2xE+Po1RNwU2f
uFLBGYmoi79pGbMNWXUHEuQywjAg1L04sGKmU9V3sEYOUL9/MI+msX77VJ26PiIc
rtIfXcRXrpTTFU2Xlisf24roFl/xUoXRIO84R5yg5ZnmXTfkxIY30kz/rNQsW7TV
ZhQkhojDyFpCjdxZg3cGFWn8NWnVHW/7MEyUwscicVHo8IuJbxkdFTPXM18TCHS3
ucqBUt5016mADTlLZ90FwHnjwUjYns/lYVCh7cEo4pDTPukF3YNdNOUX/5AgX+2N
8t0OVgiZ5JjhGa9swfpSLXRKiwjAD0i/nPwc6uYGojp/GizX3ohnFynAuBYs7IwL
AA6FSlMQYwFn4x8tQWrtueaqgfqrd7lbbMBcTzqrecfe+gMFSsXTOWdJouuee+1p
+FJtHW1eAS7sy23A6GOSViZBrYM6p/vg4YxizA2+C+jMQP+AO/s2iV5IHHom7k+T
ZgexS9cIJC/STAmWpHkt5c8nKyaasKus2FsD4U0n0CkiuZgDhv6zGl8yxtEznP2c
eBvaJTfhTC2+7y7J1hD4nZqSD4Gi3FT+0/MHDNly8Xb+blteOzp0MD+27g+828RX
uIxCyJpKnN8m6A/bVzR8ax/gSsDUpVZ6fTeQo9Hxi0mb0yDE/YANDY1Ip2FBfMdD
dba+jcNzDt5MZn9Mfoj50EWDyxItJpZfwktXHkIQFJJAZjpkN1JoTrWb0xCWvjDz
MBOB+h5o+ZuXIscwUr8ZB0A80VILvMi69i9NR93eCUgsrUE114DgQYr8RTgROk6/
zl5+Onz/JcjC40m63O1NqmaiRMHvSMFMBYl7KBtOyGmUF5o0dDyIY1LjpZ5Qxb8O
Dsp8kZfxHWkd1yBgNWbxesot72Rdc835bIgoWPINz2how8SEbop9rhMlY3U6k+xe
2v4mFtNQJmJrHhBoHKhtfGN3UN54G1Xbw47LcatMktuDGNwl6cW5AsmoHKTXm28f
Ycc/Isn/X6ZpEjRKf90rlLVVQzZRSgBdlsufOwgR01A6V9zgqWmyjdNds8Ha6p0k
RzJm0mWTZpdr5PtsqSjsDDPFWQ4zbVTaSj6IFRzxvTvUiE432oPG0cZXGyA1pfXa
OSBYUMzlzQQ9TiNVxVuEkRU3wuvg6wktZWqyjw08yClA5gTohS5zCe3e20a+YjAS
unZqVW7qq4HYQ3+urB3xBpoFHmNEh8QskBmfkbQqL1+P1G2RcCcTyRrhcJ1Jvn4d
CEJE9g1tkjQaagJduCj9CUL6XY26QzEqylGBDLdj81W6zSndNGC3w/nBDR3kbnon
eI4UiBLB/nRP7uOu1uZfn8t6eiF31dwSd6nXlGHrxUYCwbuX3jzdEgv2I3DvKwRd
AgwsbZam4XSiBs2XvbGAQ9AviZ165pZCmsDUEa6PsdlwVmcTZi1uF23XPWLQH1bA
DXmg+D6+w9j4dVrf7AVLdw/aKpfTKLdtbZDtccQhGXAyJTumA5dJZ/i6QZbocXif
7Rmk6vu0WwnNwQr6RxMEwfxBNtGyj2z8otYHvItARvwviMSP7jcHNrmzC/eUC9nU
nnIjmg6HcPdda13X57Voc3zbYUPnjpAtXHvi7xW53HrH2HEIuNN/CZrvJJeBs/e7
p+0BvGyodXOywVcdHn4TmuBMKXUmTrhXMdGpKI4Y9APu9XOhQydNsHULkelNqkN0
Vbl5f1/Q3WTylwYW05kDw4acb5AcN6Jr1Nqx5e8a2La1xfOkBZPIPbk/VHMaZejV
e6BoubKWtiIviP4briAiTvaCsic8MmuqPUUwdKyGEH6hwDXrFd8Zuhh2s6yQkiy9
JQ90H0vuoX3zTACDZboDDgY9Vw07ms/bemetDmBwGB1GooAFjHLak8YSqh60AnZd
bhHgjc3aLaqP9s/EjovZtKUKGzCy69dl4v/l8lD/SJxjJF1WPmLydBdQzwQI8yxQ
Sr23H3910JcpOrBLRmE8vMavi4j5S5dr94Z8hi9uPvljqVz4MSMl6S7T7cSfVQOO
Z+B9haZHSMuFnLDjfAgwsUpmVrP5UnW/g1TF9WSODdsPVQXmxvd+w7snhz+0MN8X
0u+r1lGZILMAEvzO2PWoQeq7fJmEP9SZaUy4LFkMto0XMhjCuvQ5KvBqPcEVAHJq
nrimBApj70gkhVq14Ec2Xgn2C9yAnzoYAIv9CYsaIijwKmZKoSCTe/2pZMmikJpD
3nqA/sGYBZ2Bn7pALkL6WCeaO7Iukdu+PilQGaIn+8lKMwVJKte+M/WeE2IiiLyf
K8RReu5WhZyJ30A9qJj46tfjvVtCULRtA9jWyn6z1ZabdsGcq9Qms9itTpV3PnfH
D244I9t1Bod2PILp32JAUYjWfqjgeRpDo/KSvS41s9ekmlG0M/Je6Cg/fF/Wv6zU
Q6k6/I//FVNsDsWG8uTypQhzmoOZT8oL6zIjjc1hKpgTVaraCmwGGSw+U0mtvxzB
vSTLBmripKJ2CQO91qObUP0vnC7l92eloloJrlEiugIifa5nsVKoA2mTMI4kUMsa
l8JrA8hiyZdBks78gqChcu8+nCLwWjoSGrkOVD2Tj8ju/AlCxbgy0WV8wPZtY975
P7AgmTCC4kGBTVOdGxH8svNMn8DkNMADV9bbaR/a6/g/sZlHfIS6zrXkj7z5ea1f
gErBUfZ47XUPgRteoaYqMWJo7NPq/KqLJRVIN/60Ede7YACWNGDL6qPA9vrGH635
X5UNdvCbcQ/DP4JGNzw4FxNTrLWknoNb7xcfamv3w1dzrhTVBx+Ay2ws6pfD2HQH
Sfqnu/teMBFFqF6ItkWKiWpychzGWGRx2XS0+tSF+wp0sE64qUyffYAs5DhwibQS
9uJHOCn1WyQpKM6My2C9r7YJqhZBk2h83RFNyboSJHkNAuzvgrxdCFRQuDjXz78c
Bef6LjcYz+iOVTRwcsmbb/37iFt+zUPMFvnxEW/MrBoxAaz9sodUXywxZ73BYifa
uAzNnaDeNESMcBCJ9f1iEWbfpXN7wRFa0KDZKunI+ougEi9gc0OPx5bKYEPK8yUC
4UGOeUlkLEC2fwecEL+4LUr+kU9ZfXs+K2tUhu3cER00In7sTG2ewEiWBq4NmRWM
+qVmZOWUppiQAno3kh0Imw2jZQMeHL2WCkLIye492KUxKRRR9kBn3nHztKUY/Yuo
lG+ioZevribpgruviZteOmNeRUody+L5uXMHqXSplrA4CnC1U5546VP0ERU1mvOq
yldGAA7IfufPHzA0blcCYbzttvv4G7Z87cI8f68K3YRJZjpBdETztifyGy/mY/Vn
gV2KXX4PRkQEnSeq6XqU7h4URR0FyR4oQ/tgFIRc/AUmLUTEgPn5UeYOcg23/uDj
wOrJqeU0LDB34YaDDCRv4OhgA9lOrM9Zja4q/GcPFzjM/gIUP6xRdPFgL37pBZm0
jT08EPSoRh00M68XtLdkzjTl+6VMXAe1WZN3nlQwM7GJBeJbocfrS5PGj5XjTxc9
CI8xhV8AOFREEpPkGgKJ3x3lH3GI1Byi7QD3ypW4WEmcscmOg8Zkjp/yW2NppGj/
cn3zBFI7FGcumq1zLUaEm0rm6VsWWQ0mdpNx+xZSJHPGHOxg3cG2sGKfuJXhdDnH
65nHppAufADWoHCj7TG7bdjimmMW+vY4Kt58ga/yr3LmaIGgEg6wHTea5/xAvcLh
g6cf5NHosFQFMuLOP21T4Cq3Qoa/jJvachVb5kcV9JkACsoHgaweb7wqwenpPSbu
JINcS2TaeX2xUNptjV0hXen39CGFih7mYSbqj7OBezbD+IWM5SxIlGCEjNfeAmc/
OAG4B2nbGLcT2FPnDC+M/5oexQYV6DLQgNOAEq3IG5EDy9blWYFTMOGVH+ktyKpf
8m8s/0YhjYXZy8Mj/5H9/VURWOc4DR5fu3MuRMLVL3yWb7jqonO34Sa+pZ166cbF
zr1juaHaSfSwR+F8OshQA55nc/BbwdvLmxuII4yPEkR22R1Ny1On1UjRnoKEf9kQ
2IZHp9M6VTSUnPpwiagKzRp2SiuEQhUpd+FsyrKdFBeTv7xq45rpDAeZBtoCQGyf
2c1GJxzfLZs6EGJfUgg6F5xRhnMcRLW//wHIuCa+u18eD9P8MqH3XGuZg4/5y5a0
U2rxKSFfp9Pi9vYrwHCU0e3OHPuvQBOt5792qM1v4I1VoXOVuEM0ZjH1jfz3/sJW
ptyyyPWHAqqsrQ9r5RxrMq40xWxcnxqGsmk/vAXC5XL7DJA0DK47pLg/TwM+NMn4
mSwIEx3IsNhZ/XZN4oenbaMU1NG3zhkGwjOVIwHqVR4/L4tAd3fJfe/+JmhaLLUE
SAAO9glqJ0ZIaxpz1ksHCNv2zdXMeWbTM9wC6ICLJGs5Klp/aQA1X+97SNlVxkuF
/GM3Y0ZyYP39MDLgSpCSnY40XQ7oweHS/O7sw8PLR1n6pqrGZwhAb1vsJwvPWfwt
ly3yezU51JfL/5chDzSt2V4uOyCn/zCcytdOCvY748EMdcimxfFX/AZAeo2nYYnW
+ztfbdcJpRZ1HIcmTOm5zYkXL4NZ6kD40rt8UcLKblUjgKHe5/rvzAhtdQ+04Y0X
8hGbixd59AstuUKfSybcOFdOXrft1B4XO6RA8axb5g4qPH5JiMR3QG7yNIR22jyH
5PWoFlP0CO5+fHbgiOEzrUsmepwXIVQnMbpltWFmakCZjoGtuBmb3neGVdmlcDQf
Ml75btiV2C5EAHxGaHwJmFvMfbbemrtkLwwlJaQ3WCp71z+4K8xcbsCX269Me9av
6QgiGlNAypY2GVv6sCBkEa/DkKFjqLqweu6Cy1kjvjP/9QoN61EgFNHnty5rfHpd
cvPB77CtjAoi+h6GCHkMkbPBvy/JkJFSWz8ReVSkmB6BWg0h/wo5xlGxmhi58wgB
/WS0cDCLKvB/37I+uVa1uPNTErzvT+glIx2XTnJ3XCxu/sRoL8tJhTFc6Sal+375
h69ChOIXONX8cFemUvYjP5AqJkl+d7FnEFKU2iWRxkv9kDdLePAyTJd21Oe12DOf
aFbjzUCJruyRfUJbju4x41ckFUgihTmACw5LYGjOOSAJZVW5VdgpWfwdcXXye1CO
loQpLiKlMFSKDNTgKGlISFDy/0Ge0ysDnk1blCypAm9pzL1z16XF/gTVnt+41b0w
i1u269ZNvtwJmr18bmxEG5jUlDqOHi0O11WTj47OGDPUVdgShqwUELGyU6Ryyl4Y
fAtgKocyWaTlTrOyGW/ocPq4wketrMvQhKRgSYcKMlDpzbv9pfzLH9DcYRyteh2T
hMSp3Tlg+PlFCennLmt9ISItXHvHuP4c7zrBIfe+tL9RTLbEUm+AZFaUiJm6NnBQ
j3RZa/2aGmxWVzSyiKZLU4JULGEXcoafNIxTMkKjjYOT+wKl88C2aVeo1KhRMDVx
NVsOR+B8mWV96cFiwirdhKhJSxf2rxVQBW+a+/c32jf0VaF7r8uEsmt/Srd86wSK
+9V7GE/tTJxOzwxHhSsgz8wmTo2voAKoAEwQwV8RLD7uFvcZK5poZ4IY1wbYiIgu
XbDCopEbCgSnDds6T2seqL5JlLduO0bNwBACxz/H5XG1NmgtRk0KEYZvHIaUz0fj
Nj9DcSYDFTHnm+TxXEC3glGh8iN5z471t5h790Z1J6kuj0ueI1oPX8+J9Cxo7YXl
1xY8MqWW4AvKepp6UAm5DH12sVVlEUxKCphwwUUhjwXMSnVz1gzZ0KVuZqjM5RSV
YJoYhm7AahaU4wFJA7zdvA51OhZWzrOEEUBOOddK1Cssjj+eD62VscmuxdImmOsp
IzU61pBWVS125EORm1fXT5EXSlXGrq6O4nIU2mp1jsCbjPqyy60OpK/46o24jqoM
m5YF20DMBahED8Gkrh/w98IRZocvv5Gt/b0XAaepMffs7+GMgztlTrqQ/hC3ONSr
5yQNOxtcYIjHuWWEcCrqWDNxQgHvJ0ya7gDi/Bp+cpV6RKWS/AiiJRTlji6xwI3d
mz8w8QEcy+aFv+Syc3/yvftWGltJo3vW/FHuktAWYcYhkUqRjLlf9nQIsFRv4iby
RpEscbDeK0IJTVki1UWgkMmDstN3/oJYWWvwBzYbQManyQXrT5GaTsv5ARptICp6
lbcAb3LWDnZU39WtBOxa7HtjoI2CaI+33pP8sLx7+qYs3/Deu5eOknOCN6Op8Qgp
O836CQqbHw/qlNAkvHNOSgL7GE4g+fdFUahcR4PukBbJG6e161gCJUqyChYMM0Ap
exfxTxuwc/3iIDK9xfIEQYvrRA8wTiDf6SLWdQIERjNeayHIgdrCO5UrmMoHdv+E
9Or3v+oxxjk3lIVK3jxmMS3D8Y3bC4UW4NtqxHxXGdBxvvr3CkKal8J1LaVzpbUh
KHvVWedVrasMtZZAqceepkz4fbEIdmQap7hBrT59jC2QflJWFlNSgt8lZ8DOof1i
PTT71JbSKvZngpUAxFtZEHomrox0n/xnmTF7SjyqkpWMncz8I7jIBIsC7E07u+hK
2IqSfhkG1u/Qq83Nr8PKMT2u4uhVBO1HvAR6Wwn4M/59f+0Bvcq1qJCa2UO/veL5
osWOm7eFbR4IxPUev6eCyalvK1/R7F/8oxzhl8ghFxEYPliyUv8A8OxrDaMkX6Xw
WLNnnoqt5PCniX9e8EE/4GP3bmUqo8pj6GOGBA2k2w6bjna+9tsZcYJfDRgJZyBS
xpjgKHBQRdWNsqA2Arts/xml6GZB0+bqapQYf92OxQ6EKfFnjzrAXCUmurDZASML
2IC+lOAspDDFczdLDkbbaziLdtw/gImuCPdre18M/hT0+htdVTTNCSkdaaRkHL7O
u8EwYROSKh3qq1PHj6l72XYR/sodtZRGsTtK5Ew2lOrqw9wRhwgd87JenTbikyAU
chInSExeNiCJe2fgLV0ufnkseH5hpjIHtPcl5bOJaWEB3TGYS5HC2Tf+e1c4nR0Q
0tlm8hPs8QXXxZeVAOQYMpdxWRz/G7VBxxyrRvcfDtn9iHahHjuaaKqMfzOCXHMN
CrSwPNwqICb63n3Nlv5VHyQA6oCoG4R+XWPkSVMOnIYOxypueJyBgWb2ATrNSQSg
FuJIiwxqO68qPJWX8lDygiMk0TCGvCj/XwvtuX1q2xUbMBCK+T0ZxMjE9GAW9ns1
v3xM3QKFhQ6Jdp6glYoeip9JRL+HPzVFnmpZefCvmZFbEu6iQHAa/rq84IFZB3oe
rsdOBD03Bq3bmm6LCfe5W0ohiXRY9/xxl4FKwkRq2jvKXoVrowizCdEpsWnWSMEg
RuZjBoqhPNXNebUpbW/3YQX9f8fPCAu2a9tVE7zoIWdaNiwMT4GP9Uy7vWB3kx8I
OFKZQwRT4CCNrcT8R7Y7Nho0Q5UsS2BYVH5CdD5xivDotpuTpi9/n6rngES/Ira3
3f+RP5JIGwN4op9Z6JAlv8dYxjyp9XMrcGMPGnvTBtJc0+XRbTlDTSWqqa/zdRZp
P8BuaJQRB7Sne/3fzvtZINUIIdieOsDKHsg3KcpQQk6wD6nL0LAxNN39nO2RPWw+
Uv0IUah3gLbHeFE4xkLezaCi8MYGRmDmHe0m5Aj4NrvaTeGd8O/RBuhAto+hnu2h
0JLSlrDGDWAR61p0Min5Gi4/glT0HtTmmy4ynzwwuPJ+0m4nYBo94+k3PrmvaorX
Nosq5Dc39GNYxVudg984JThq86vNLa7+gn9nJGM8LHJwKwYjULmvmSFKzA7z6gOY
kQTLDH7eBQhdJ72idcmSXaFbWZ7J3gIKJAJDeiKwx4PBhWDydA5TJJF57hFyEwLM
RCUp5uft7GnFzrxbdSmt1cm7ENEulfJk5OFgsuorqlvM89UkBk5DYPT0pXGmB/uD
9MBob0IiwKJxk1ZEaM4DEQuI7J8e0JmrE1eAMcyNQslnZ2SRX2R42Uc3xs0qdKv+
N+TfVtS+cGdEH/lHlgD/sNm30mBD2s3UIph2XSway1poJ7jqiQb2AcYAXWUN0Fjj
WMv/SOtGFSS3Hbucuu6+IzAsMIl8ynAhTtezOweOvYVxnGFXIT3hFdwatIzFU2cY
y0s+9KI9lHZ6O4UmkxIVRFsCoiBHTPsTN04sp8KJ0eMC+62lWLM5zle/+8hIhk3a
iwek5G/BCCNUop4RQxyzWCgXzKaf7qZy/KhT5lLIwaQyWCFvs0mBNE5KpkckLj+t
8Owo/nbs9mHWUDITdpLMjeIb8V/q4WkHhto8oBT1koOBvTQDBwJ9J/0Inna9y9nz
VlT0pckZ0AWvK2LnCSJ+DJX9syAdZ3dkqnalA3XfP0aUMDBrgAt0ZRumkwc6uErQ
yX8JcYhm0Z4CV2lPx9KSr5s0aMPPI30hx3nu3nYLFQZ7yoh1LsB8lvLu9me/OaY+
OpfxKlxZUSWeg2HVVHRZcho9wc85LpqYo3ASh/7Yd/q68joCe5iobRseROjLsVs5
pKm8cmI/jGfMldmIMzBFm0f2pPS0zvj/nOosLJqUQpTC1q+lCzWWV7tESV772mmh
gQ53pBGemFXOGU8nKrW93H0g4KXfYgCQ74gz/a9RFY1XTFhFOOHwlmLSqQmP4Wig
V9TkpZcv0UTf0ukN4AYvTHMNYkampQWT6Q6/5zwTLRNenT0/rhQVzA0SNzXjyT7k
k/YbYkE3PBuElhWBN6l3Q2wa+m1Fn1nMxcqWbWlEE3fcCLpQMRhti4OsNim8cMPC
CHhYiQirCqvgl0ie+r+sEUiQQnf/S8jvtuf15tECxSA0PLOtqXvx6aZpbADLh18s
aZPn0uBgZc6OtLi3l3iKI25kRPgp6kKjJ2XmY6KJNSEudryy6Ukz0wK48sVYzGhH
e78VLjLymkUlMZ2a9/fFoAYON6GXljhl2oMoBKh265sxe/Mo7PjnSQty3o5bl064
13Pd9V9oFoUjJLrdU9DjBElELrOeQIgiHkdS8gNJQbAsabhu5KaDwyebIND7HWyv
vZm76eNzIlQv9w2TGs8bizj9UFDrZrD6gk0KgJ73JGiIIFT93QSgGJGOMmyElVCH
wOFj3mLT8fIsVSTMDTU/NEjctQi5fpdr6UHp1GsWKg4lthwmuO492lH37g3nGBug
3Y//Pu1VRjSAD2raJCFNqnEEnkG0pt77ypZ+71KkKIhHDIWtXDuc2gwUN6E21mgM
sA0pZtNec96MnonrrLGsvj0RPaFSIY89e2ws5/HlXS3NWeGuVcusA1CL7W+vn4Y/
AbOfl5roktjtajf2Xgoy4hDl5iHj7O/WebQhfoo3SQR/GGOsWlmP5NB10semnPUw
UpQ1lwaEQFcwWgep1j6Li2MoEhwxbGZPK7GAPcsNT14QGIL6AF0ZH3YFqj+mHnpq
nHn0FU193RqD11qv3oGq4I1BN5z8Y0wIsSEOWlHQ08O/FQyR2qlffS0W+HXtasH4
QlxTjMGbkx1YOQvDbC7kKFPYEqbUbGgvGYcsJcYmUM+Qf4/lYs5i+z77mUpBHokU
nMWG8N3WuANqtCjXwxQPRQ/3hrFRBKf2HQTO+vI5u1urgGCJBFv7HjaoPVqlqQeI
iOVO6moxG2vuQNJ3OtTG4nzuLNDJFtZdb/nQ4aNrRNQ01KSvzfxpw5XPUuV18T9h
jKR8F2X7zD2ksd98i+4lonUcGoEVfFbHqAmogbfgwFAx8QM9AYf1LW0lAT7XcSrY
4wBnGp+V5OjS/Dp704emsllbwR7VhfpEwZLlb2b9iCPPk93E7U9pHI9EIGIXpRNS
81OSudwv8UQDqzma4kzJ81L1jYBSZ1OEC8MXhnXF6PlE3G4XU3iO1VFbAzLAO4eX
M8GPzUkfCLa1Yb7xrOymMd8a88Vw8j8o6URhNpdpyyLutR7JbMK+tiiehxaIf9lp
MZz71S91MOK7/WIgvCxoNq5yYxz1YRgTM6Z97GaelUYFyvPCKVzMLy0SIiiUfkk7
YB7m+Zypcb0v+6eIJxAb4KlsToPMRWY/oLjNPSBKBqdCknZ/UnfRFyka4IqPlzhS
EHvNheVBfXkDDbM0WbFj3JyNgZBv6McewqbqUyg+8+4/swDLGPyD9y/L7tMqEl59
oyzflHSZs8HK1vJ92u92oDyltaMdhI7sdSBdeoqVbONFcgs3ACzIpUmPhlJB1Kl7
q5IpBxK4bZhd8BXQawPx9ToZvYpcQLydcL0eJmMeTE1JzWNwofwN0yasnwsxEaGn
4YTj25MEfsv77gw+I9hcwfs/66b5ZmjWeBCWAn5ztZMlg/xn5YzzthHTBrF3ER8j
ITrOtMVnwdYEaKa7xirjdzkzuZ7fXHNu+TXraYHR+SMwVb1wWnD4RU7TSQgeZDil
qk3MEkDO+4w2abrZ+5dnrfxjEn7UnO06H6BQchPtNXrVWciuDOmtj79Lq+eM3u+A
9HOQYaediRlx8ivE17q3h85txKLHUX/OBIstUfknWEn5sfUmJ4J94yTcXnn3zmzo
RpD/pTdigvz5aGSmUWeIXlkEpPsqwybpaGXsYHY0xnpncwumzIjjcooGXgTDdvSK
ZvTy4a/fr3bG10Il+u2sJzaDq1IX0xOTQQfvGqXxpBsQPx4Rb9TZ4XDap4In3UgT
8j5gldMSZBI8cPmXtDFWSpliISmf+yPWLZKMufI3mAGcfHgQK6FIgO4RweZEJszi
+5yK/Vrx+0UWLSRa5IlNbm/kalUpt28yYzIMNf8Pb6reXXYXgxEFJ6cPYWya/kYp
LquusUT/qlainKt+ZUCNJPy1aW1DqiDDGrOgbA9l0tslpaLYvk2jrGDktQGQoRRV
k078cg8EkXP2HZ+rgwplq9/C+6nvB3Fgk/B2RQzoYjFsUgLt3DQ9MYhivihHDY+G
/snf1uE+cdTaPcEbNDfq34C4gYFEQLcZlLoqtY6hKUrZf73GHO305saDyVUnprYZ
keyzlNlQh1kpvvD0fN62Xn5Rt8AgXdLsHxQzzBjKLAYF1XCHdEblyGn0RTkItvSl
ms/CHViLF/6UKqTIBt0KhyMDRcoS9H8CKZyBQwAunRsCtGqqspf22EBr4ExYCD7K
yjoa0TP8oCLJo8hIy9+16Zs4kRNq+DRVaQSMAb2Lnz8/1d3b0pBcPcZ2Z7JYf4jf
ULDsPmBKDybWLqfWI2icjhHJKhfTfmt+d0DmA5Mq1M8YRNl+/S4xgFCEeHgh33ng
JXfLl+J6ZPDBVweYny+up5WhLjGvpnIjpDoytBZZ4wcbALlnMs2aNbBqJtNpQDLq
aV1KHhJ6hS4Y2tF2fBCnlTkeezqN2MMg6TX0Qln6Jx6ouieU+qXCTX5pcZ39tDkl
ZTMEgyi84u++IqoxTtHHYxOrCIK7Dtit9ZcM0T6QR0ZXIkgJXQJj8dYcTevvWXtq
9gziJJ6laNJ3UEbAcKdzXCviJoLwY4WwR5vvJvGcbWG3w2N8sQigZDsgCGO98bGK
aayAbiDhCoVJNKDYsrTljihTiz9/O0u34KNbywhuxTQNJ61QC4kROWM/zVjIq3j8
Ixv6CQbbzgYEiy4CT1MNnAZyJ2T5kBv6BfhWT+moJCEGgWzpMhIYLdBEQjfeIWLu
hp6FZ19RGfgnTwghHKaxJlpbMGqRdbApx3FpvVwg0W2YkyMluJ5qDl+/7CN3ozU2
CdGFteffVV9/ZwiQEfobXB7LxEgnNTJJlqrBrfD7FsLl5wkMzIi7zLiwnI/h0hGH
2dyepKSTQc631fe+8ICwB8Y5VDT7GQunogHSep5HDHa0+h5SC2pYv4VoYjy61i+p
uv4g+/4iRzEJZhgP8j1nNaekiCLP4AWYl0qhdmEY8AtIGE/mQIxzD4K/cTs8Przi
SeQ7EQo4SN6XLKbSin4z4gluoeoRaNUKg6AgxeYpDEiQ47AlUy5aBkDiNzkbt6tR
DHzPcvz2mHcROp70651dGR9Ty+c8ugWO1ZcHDu1tHEAllwNy2gApZsKxVQj2ZgzU
+WTfcqnPwpSvWodtwghOcXjPmjUyBfQLszJZalPfQpWxLMl+I3vIAczgjyrAiEwJ
3ZEhxkT1gSuAi40gnW5OIl3xn2J1dLINgI5rng3s8vTs4kSVooAZcT1Up65fbqu2
2pRMpH/PIKY0CKhwd6YGhDtakykD54cfETOFHc58Fqe/bxrN16ceK+Mqtb7DZkqk
OXOz29fIyAeAy0b9TbFdH5SetPvpTotj5dG5VGU3Qc7WZHlRP9ynE9YQseWg6kfz
SqhUNWcxJpOAKjjsz+a2ZvNvWHIefimSP6oDffXwgtVNhcOyabO1qlDqNh2H3BAE
KJXhYb8V9ql1Wrlm/WLoLSoYHBZ+NWLG/6ci264lprDnkl791T90bH3q+UIgSyhL
I4dZhQUC8VhsVqcBIxntXn7SAa6LLkWS1Z2B9oFY7IWBMhfe+gQfnvoX4aPBHpfN
0+UR410iRD8K3y+QE3ghG7Q1ZmZ0xRpvgdTDkyVJe4s23hRfiLBxLBCmamWJ7ipg
dcJmK+FM73jiz3D6aBKlYbeb6JoaDucA+UE3Bfpq2a8UEkgEbmKnWXZ38nsvt2Dc
vkDn6jnK9CurIMdqMXaoX+0OnVn9fJvSyaIe0tb6mGBJSO2/cVwXNQqKzoH4F9dy
xI12t4sW2JO5j1TQpQfhcqdgdyChfSPGIOeZjitzchYcDoo7mmkkcJsxGuvKN08p
VEQR0h9DjCRakU04mDYPPjJz3JiAAFfx/bbKOU8MiYbs9COL5Pyv98TowLPIL+a+
+4WKrHTLxqPVxnVSLWMUkNPXLJSAy5MRwi4uzFKlXeLD8C47NLpQ1seBDj3lvgSZ
zZiBjoVxMH5YuUIe+PIxPO9WG2WKVfkfxqcwOIfTB0bruIg5flnzLfxKeVRkaZG0
c8rOkl+lkst5VyALqDKynSFs0mNTbE3sfpoRGhWlQtGPExn9Wl2G74j9DApLLTAZ
sMeBOg9sX0Fpu55jODQQRElaQsrOh7LYjKdBGELsb7gpTv2xE7x9/2fgGoz2aANL
3v7kwg7ETAYaCDaBepLP1c8Tjp8pC3yar4PUOPOMSwR499WOwEVsOeQyWpv43oeg
7U6fE+H1kTfhAiVjbVwjKvct5m3c3/b7m70WSRSTAnLEpx+L/PCYx+b/BtGySrQJ
7OE7b6AOOTcDpVpuf3vzsq2U7N0EZEA8VCxeYPiBM6VsZU/vW74wOtSUu746ZCsz
HyEiGPcxk33juhCUENuHMuj9jhkj4Jm+hMrA6kKmfJKARLFAXxIBuAriIURoGwfs
XQCxJ5WE/om/C/CeV7dE1v2fZGTAC2iL0xnQ8bl10WQk3LOLzNLgAGYwe3pzheqV
S67h0hRswLlgMhbA2xTUE/GxBkJTbbAVGrrSOuBQzKD75tulIQD3B7SZT1LstVmf
ZcXXltiY6N/DCTErUmhYask39W6OdOsyIc090Sp2UEmZ5L2J9iMy8fIub6UT+X1G
wf4Sg+Jb8HH2On2xF4qNmolxcWsACJxzlpakHb8vSl38e3r+K1luRVT5D76W86w6
4/50yASczZMPiwKeZxz4D7pBVPrqracxHLqjL8F54cdsu2hh1OE8vqHHmaOGP3XB
tD0Y3nHyTn89lbEUiC2OaFUdsD7iJIFuiXu+tDZiUQSXxpV/5dw/52go80nb64zt
aIKpHhHT8MIs5HkZCRUdKxrVM2ZWu+FVXULWbeVp4Dv+OdX4AiHwAjoBcDcW9jMX
7HVVqVbq6YivEDHoNdSUGFHSZD9xvtfmNwS8eT0DApUzfNEpJqnkwrwhBYFAS+3X
gl4Noi5FQrH44c9fi/kg8N+FNzXAeuqTuccSXZNF0pW8Nc7zWQClvYPTODIwfRw4
18Q6KLR6XDdAWQRK7pGFkyzLnLrWZmBMpCbBmpfjIMYdklD/2fh8/GpbfzDc/gCT
hPfeZOeusYkt0R4J6uTW6QfQYF+H+DI8wtWnaZRC+8TguAkC0rEnOxpsWYPiJcTE
fRmKg68cTn0qrvWS9sLUYsQjW03lg3q92Klb8OhYT8mnSrHoJQYyGyX7v/11dR3l
SxaXPMjB73Y1QL59eDBtBtB/WzG5wj9NRXYg9b6DPYFiLKXuD9KXPnh78sUJcS+R
7TR/RUz9r+5AAT7B9Tg31hgE4T5uPz60f8yCPbSQw0CECq5XXGj/Tu+fu97PrZCm
13JzioC29oa1o+1WdyEJemr18Oba2PpDzldvfHNGfvylrdRlUO7xM7BEWmvw2aAN
JY1uQjIJ0JFhCAwVD2xtjjwrrAxSTYE3nd3jgQ6K+bEpQjhEDTxBdQ/LTRb5QoI5
UxVuIdXhMbK30MoNBFrgEicLjvg0cnqCWQXvQnW3tvWmjJ+CV19kc5DJp1HTnqLG
gNCglfH1aBAYUapgeVmSCmNu9yDzBtbh+H1BP42N8MIRY/qgmi41yjfjRM0bLrOW
KVpxU8W9Bpi8QH1CGMCNFH8pzSw6y0G8ErU2/Qf4r+obg0iQ5ExTkHdftF6JmY2x
hg/XPOK1DeTQO6GLrSIiIRVl/4CbbfOsR/IzpDniEyBWwf2WHZ5xrysBcPp4Zf5Y
s7TDfL14D8SM4geXIyTJY7YDhKF1Q6f0TY8oyR2H3Xqh4I7L5Y9CgFoUD8Zfhzi4
9FL6fjpzVDa8N33uLVbrJ6ht5b9MMjZPOoriN89rjPkDiUrbk0TKHsxu2P+7Fgs0
AZBRqJvr5GkXxsxFZCyT3XfpHy2SzZwlA2z5VF/oJoa84t2090/v6ec9aIgSm7gM
kblOvZDqIP30TOa8OfdU5aCg0IdQnOvqeizUQwdHutw8siD1daymIWvOf7zWfY4V
PT+xF6XvWfBfyHtrdwvJc2XHxP1b9ViPbgGodxvogVrTDVOkYuw26+ne6VfVYUnH
YL68jrMB9JJsekuG8a/Cz2X6iEu4PADkuY14vMSkd+O1ukMZkz04KQ6XDe+srzL9
K5jgM7WT63ht8xsTYKfsiBXVbK+XUiNQ/vPYE0ZSpO15hkKBnonR6boJ2TkxwiWz
NKJYPQ406L8FOeSs0u7k4Mx66z1xvz+lNSSvH/+JvO+Sck7cbwa4ciAtLSIHTdMx
FxyRix9/STSArZqMMgOQbGLhDRIxRDCJvPGUZRbVEBardQS6Od0KE+P9TSpX3f97
E02KKXTLjd6IA1DwJ/a/auyW18AH8Pza69hkN+ETjssOY2u1pY0/6eMVnq6eGJ+L
p7fDrmK2wm+H3cZcKPskH5uWF82mJ9ERZuGy47NY6yTAiFBvBu3zrkKfPBY+1DY9
O40DHlz2CeMZWv4j4KrefxpHLZwDlk4IxQJjRCdpm54OO9BKU2H9agMRll/YoCfp
iUt4ECkwtA1Gbe4OwltMd3uq4sPn+j5K+RH3CW8lH5d7MxtStntaShSWobm6GjnA
wkVWpxksrX3hFS1fy5mhu9WC48+sQFXctLtvdUg1oF26Q9MG8/3dS5kmVPdaL07i
U7b0auSqFHeJ5pswpKRwkJ9px15fVgHvSFuGDHMLSYM2UhthG0zggSOzLzahsdj3
CJDLIqYmDfw0EOOr3WfAzvfl6laJq34F/pGYTB2mhwdQKtlJODdf4o3Ni06OtLdz
BgZLAiFrN8nFxHajxUd8zwYByb5218KA8OR8Ph5rGCnVkkW6GIGT6ccRjB1Lj2xq
GklUSmL4EiQKhgk0xB0nFgfDmaUZD6GHqgpFupogL4BLKQFnbJcf/aKtr88aI6cb
ZGGkOHwypYhGZRkn7kKVjOJemS3tAbzgv25s1NlaV0bUpFIY/x/ZFrDVIL73AMmd
1MIBW6V3z06oZGcpT74SAkEJqYUNBZcLzx+JCAAHvabovBRgzaGw7yxtnfLrIJEC
1KiMfk9VINRBU2SxsnR5pf0wrI+pgZ4/lz4W4Xy6e+E36J+bO43ZgD5vwIlJhvBn
RvWaLjpYflCXK/osE3DMSTF9XoEyCiRrUE7DgpyJFZsmwY4iORZNIjNqusknnAYW
g/7esO7va8ue59xBpl7gu61eeFm7muYXR8hGHkNlBx3LewrVHb76ms/6Sxp30VM8
e/lO3zNUZBqAFx80fMeiBMUSPAs77QPkrwIFSN7WBgIlMJyWa27bUxoR7pz68Dxv
Q6o7Cde8/wNqrKqTl7igvf2CJcsH1m8xtIqmz5kSuDSeWCDnG6U7sbwxUczGJdRu
5d15oqe36dugPRF01aYSvvgB2YVmJQnOKzAteozYC4z24CJKYTHzLGDXcUP0uVQR
o39Zw2oxG0xn+0ll/tLaqpOZPvzf+WjruwQ2Vy8VZegIGQXl1rZgGufXqoS1e+CE
WAspxeCpoBp3w2mpOtHBfOAQgoA3Dlz7zfSuRjtwZCGby1QSU5TA8dqEdk7UCmgc
MY8hQrOncvZkClRW5Lj/Y5I3hkLpg8JItyHlRcROPnYysvRYJhj9U8aY4+8YeWEk
fMIx7Ic6m+v8lWGu+EqD9gmdgBD+bY9TO9WPSc84R/wZCM8Nsobd7dHzZQNyimB2
vrbfcrILcV2qxXLmLdtuI09PUF/BhidDGSj7xM3fbkbut3ok2ssQc1eyc/U8wqUb
+8aqG4LNQfCX4dtL2i4vJfs0Y17aHQ20yGQQfitMistprsKSh0WfnBxgX6WiHVPR
ptmBiHdr+tJVqD0qQPxrijrBInyTkBIEF4/IF2HPj7GZ53a784TcACZdJ1CmBUml
Qrg9ARq05pFWDBUAHJiIXBgOWgx3LTcqi3t04P+nfSHpBHED6LbB4OTtG5lz7V5c
ypEBG++lq9iraFXPyDueteTP2XDBR7FNpTe5Hkkomik2yKQ/wNJt5ZMF6+AbeSAg
wWzuOsYxEE96ZBWbKbkxcQpAxfkIBLqQWtNehjsw090KBZBr27azw76rCB9BMxe7
cc6O8IK8CBgAuE0bv8pvRT0qP9A34NSbq4DkRTuUGYxaREJXk3eQOdXGEadLPPyJ
KmgDSxnQxZHeLilVOAWuEWtH6f0El7Rx0VL5hB9v+W8wf2EjysS35i+3f8JydSpG
v0HDi3qZwiYUe9MKLj7N2iDPHeEeNTwWvmMjmHOCEEzVXSq8J+n6J1C6OhgQmWOa
FVrZhj+oLmhtOJYB6/fYUJcvdlb6ImCkj0zmK7CBNquWwgiqRSYDgjqx6M2K/i/2
B5FrcSrXbQlvZlDFe4fo+tu1+8j+866vkSgmFj86KIyn+CTjcZsXVIrG5KWrqMHw
uijcuEcpWnpWyT+ax9aay4+lLMvvDR9dl5eQxzO+AUH4C20dZuzZTYbzRogAVrxq
p5pOub5HKwk+jZSPAv3kjNTLkhv8eNi9kpeu6f49fViTTHGVVXL3pbzqHPqmgQ7I
pYJijCHwEYfoNbE0VlDfOmBQGbssmZ2WB61DR8e9DwUDP7MCe9ceLD49Fl7L7+rf
5C4f0Zuvx2lDuYAqH6NKI1mRyxo61nuOtbjXp9zk0mNzKW3T409aoxMndRZEMG/O
spK89WDiO9IML7GV+YD9asz1b+4jTFGHp6I5ba+eWPOgZM4r8iUFsXmj1m93AQOV
c/9r0Oup3XgltUgM5IjEDbYArwI8qwdXJN5NAlIA2f+5AD+qAzfXGVQk3HxTf8pc
93D+VGtO9e0dMZz8H9XRW9eJw6zvLlHtQW/k0axpiIkRMg1N367fQB0ymUW1TrSR
P1bIFpSIN5hlNLzZB9yNpJAb4dDLPYw2iUcejLyT+1SI3NXAk9aZjbuRS3vUToqn
+5md6Kj6Wb+0HR1NBkhyb090r6JnHyM2h+/6iBHrMP6HV9EErh0rtnqGTLOpI2wG
eu+9qrb86olcIElqfsQ73QZTDzAKhpMWUfROs8RFzL+hf35i5XcHbraXKxOW/vyC
cAPP43jFOTuRlo2gkeTJLJufhRXXVVQQ2o0ZL2BZGMmnWkjV6xfxzyNfhlN3Gv3i
xwBjBqYCo1BC3d901OfWYdjQcaELZtIOF5fQoj8PEKHM2Tr1whX1WXhACMS0QzeC
DwLkiPpmbU90BVmA6q8ae9LeUvDpbUi7kL81tqxow16SkXoCYc5ms3YIBpWPljEW
IJM4goSahy0rBffIEeDz238Bl3aAF/Ts7QAhqnEynH/uI7M2CcSIuNN2M/6FPyKJ
sAOY/DV0qgfjEKkyd0OTG0Yjs4gqV99dkHlmHk+9r5322m5lLJlPzZ61s53fwLHy
VMzjNwd8YV3L6W9dfEoVAEykEOy0fTMsRrJt63kKUiKx2HEAwhL8f01SEwLnYDDm
FyCWA6XcWC9kqG6iGni7J17C67nm5dpCyE/7G7COYuMEdwTxB/x0LM2Mr/yAaE3q
jugFtZKuXXnCEwd+iTDEDDyCtuUCVktxdEy/j3GoC6qvoEY76HEio8+vK3igfsJt
zol3MWjT5BXwxhmJF3QKvCnCA0YFYZLyixpR6jFmzdzwMzaz0HtMWCJ6V/CNSeMj
3pEOmjvo9ZaU93o6SrQqICI7QrwFXHIlHpdB3cjBOgAAb+bZ0iN4NAFrjSgryE/z
d7F6VnNFce11eqm0EJpWzcxRId5B5LLRQoXe+V1/dk7Rn+TpymRRFeJAiV664q0Y
Qf386oMF/FFCziQIH2KMiVoGWCgHNYYkiztAp2RLlMKbP4pdR8vJIGoChOirp2tr
cRNYmo0Uj6Um+SewrSp1AxijDq4i6HeHTgDm4FkgLzhuumXR10OAbG/QkuICvbdb
zh/3FDtVmWFk1MvrId06ZMMk3SIigFBFKCzPDOskaav6syZ0ycn1xxiCI52TbhHX
1H3N5BtMhJ4alHNDT4u2LnsncXehHUgz8MgrD3kxVIbPpLRMrvvsNOc2d+W2gpQW
7BAw89b8S4szTcqA16pDVxIrkniddiGppqzyhdJC+GsD4G7TYnPDw9tJX/JV5KxP
1LFpk0wG7fSiVM+Pz9fKXqTvfwWjAMl3rRhX7Ggj4oQL9/x3a3pzr6kpyFF1klVB
5GnHRHlIV7agwuBPm+ozYdxwkOnhBw35kXuea3L8d39cjSNgCY9bZEMhid5niCUI
EwM13QSyZcSWyWdm98Ln9yZ6INzf1kRK5Olwo48lJg/Q7BqLBsjL9aeRjcDC8o7f
ddAgJutxR56MxQkYVlSRPeGzGpKs8Mg7elW2gvPNuucL/+8/vL5NL8nKkUf04Pin
yhOFBuskYJokJp113+pq+uMxObUmflSl978uRl+JTtVOZP8GzN9Qf37yLtAOLEWh
mGoIAw4CTmIIR1ZAeaRuBD91eR9QaWhftnU39W+/gHrV3xDqbjCKfnB9nONkFvdi
VSXxvE7xASgR2ZTr24HEdznBkhDLWqiNf+HuTiWVTUXieO9ShDvlyWkEO5aiRUSP
VN9WDCRhzuEae/a/H53fhaCPGiEtz9IeFzMNY3YiigpwsB/MXngsU/mc7PIHHyTX
P7ZCMTuDhcwNH+8EjQ1sUKZiOJftWV4tJ/1V1UKOnK9dyNL1Fga1PSMhOsi/nR8q
qhQqSCvbuwUyyDVuJApN2wayz+sa6tUYU9399VfcgTqLM8qGW52n56mMsl6L9PVT
9x7n1bCQMFdTFxYAlUQEYtRRVdTPUE9nHiL/calm61d3bk5BnAnab3pfC5DdJOUa
g1nq5p1sTfHgr1yfI1VuwieE7BlCCmREQ+nMCR9rNWw=
//pragma protect end_data_block
//pragma protect digest_block
0S/G09IHx3P2mRXwH0qonk7vNd0=
//pragma protect end_digest_block
//pragma protect end_protected
