// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
oqVAgfHjuFo0re+mAsn8miHRmZj++oVDGUyexTpL5VU+cWxHcwd2Ub1VETtmzVZl
0eKDLTUp5P0a2n7nC7t4/Rrto20Xyr4RYzYhCgPw8ttKtWj4az9X4ByaeVerxgo0
mLDIPHOvGhHDlcaIgq50Ub/4WsSSHpvZczjYIiBTvRWpQpVRf4+ygg==
//pragma protect end_key_block
//pragma protect digest_block
nRbIJqHQeY3/oYOzNS6Azh0c+HE=
//pragma protect end_digest_block
//pragma protect data_block
Vch1dbw+U/2vUUaHP4yU6Lf9V3S6HkY/nbDUMYXzsvMIC8QdbBawLcdR7visuzbe
uX3+UH4Gn5B/zEw2Vmvv4uql7fndHVbbXIw4D2Kd0pJKTKWxWQgJre0lufXRkGoJ
kQw6Lb3ateGtN41kWKFVjHc3b69dyyJ7r8YYPY4cZ7w75qhbH97H4o36Izbs9LY8
OkOWubGyfdr3KpTZgiKvEFu2IJa/xuM/447jBEy5b1SA1BW67NUirsPE4hJ7uTRd
BBs02AqOqVJ9R15Buo8r7HHvGA3Yk0pswYVTaaRjNXNfYfRVUffV0LvkFiGGvtRL
DMV114OJZKEUpYDmt200nvbtRaMzerivHb5M9Lq6d2ZqR0TST+KZhQ7J26bG6+as
s32CI9d9UfDkqYMLR7iQceHIQTmu277Zt6f2d/QUdakLXgNsGQ5ZllgYu7pKUNtF
GkNZ9859/nmrJ6PiqRQC456EzDiWN60SJu8l/2oPvDsHKwWnIjKRbT5QsEGC9afV
sDZGVb9PQLEg3gbujL9fHeGo2wzKj5ADpOkFiua7gEcIBSVbYgJj4fq2VJTndTyi
njdTltP3UsVLC/vsVEt+Y7qOwNgpUaTHZ3lAowiSZ8jcTcYIwNb5+vNPcemD7InF
hY88tB6idjBCWujoy0y3T9jF6ptHnDEr4qyoPUgH5p2A0cnDxCbfDHL8eTqZIQ4k
heC1bK0frI4GaZJeP1taUPDDcL4/HMGKEDUxgxgL1kNOB2NonPS2RyBgy5fac4yb
JQn1wON38UrPASFGFxZcpJl8Oi79yzKmSYh+5zASdtoxxdrL6Yxd58TSThBest5p
ufiYkkw4mLguupZOp655fqWxnvm5dACRBqwCSKUlLoRqRMTmK5hOA6Rlc90dGUrO
YxMFF74iPaSU/99Hz4uWjiOMR0uefdkrF3WpsUIZsaoMb99g0//VUY/QMiK8Te9C
rYNDTDeSs3O/iAEvFIwy0ZleSCqfPH0CNjx4Q9d49l8Ly7Nud7vwPoo9YuKCam9f
4Wsb50zEPm/Uh4ftnHFl57wijjtx2hxvd82lP3VqglMhvgm7NMICWy/PWVRTteqC
4cUWu93sUMwhi2KtS79/Kc5/MCJp5Rkv9s2o2mZV8AFzA3f+U/6ZCWlnzZvZ+fZd
iCVbbmJQ/olPY2EO5bSyX+GKGOCVUNwD9oiDJbqx/zfsGEbAJmdE/gUDGXSylfc3
d+SEV+eWoWMiKI59pOoPE5xhXuoGFFVWd9Akn784vYKhS4eIzH1Tfgf/aNM8atHJ
yOXfFQrR1vPkIEVUEHqkXjeVvPfgAMTHUqT+c6UTXfCkeVkTD2VoxZPasXD1DOFi
F8SwiDBJbBe2skZE+EBW4eMHqLs8D2zkYR4nrP+ihbjRsrdxkogQQOgF6IjHZct0
cXu/H3VhvXhnQylX/3NUnPMAm4r5gQk6yuCdgJHAPkVLooR9GFXA7Y7EWjqxKOZ9
I02cpvY1tuLoM6SL7uukoy3o7EiPzCmcyuPHguhAbVU/WEg/o6WKLKlLCm2dZQkp
qwiQsc7Pimqp7GfsvNMHVvkdEMVxIVnvNQQ6VpotaHCpVirFX78vG3RjLrbb+F4r
PmRb6nNte3Seg2TKir3MArGhJN9JW/i9MLeENPP5VT/iVMcyUYpXxwvF33zs94ub
RPPk2vk6SnukdkIFlwwlBchJ3g6Ypu8XF5RBCLb8iKLhog1ftxQDnU1xnjifW7H0
MBZMRyG0JK6CeR2Drh0nru7qUKfPQSbe6GOHmKAnlMMzCb31A44C1v7M64BbBYfh
0ojlAoaqz2oJj5gNo76w0M9cZsk3SXJJW1IagikIEQrziTZALDjwCzpMwxzJd0hF
h1MbsyJMhjSVVn8GZ43ksajLuOYFOxhwnEY3+6Ry6XLyliF7Dp5Hm+bLCADXlPG1
jSDjokEfhbhxFkmvCbYfMWG8C66jMDDXe7BFkX0j3ZDnaooRL+Ue+HZfiz28X8Jg
IT3kJXUD4frUKR2WYTzVShaSX0cHIkRdgqFfRq3fkSsoWODDj1mWyaB4qEhYDHKx
anXLUcSss+Ffa0iRYd1GmthRV9Um9mE+OF3wdEHW1KYeX+YLYuhwZZk5ChMNKFOr
7Rbj6fIwq+csreKzVwBqmcbP+LmG49H6OEzNW/yBqLm8q6GQXdeJ+tMazOWXUHpB
8mwSuwgesdx/1jyGl+JBGq4XbsleL7HGpOOlE/cEqMF1nm0KWhnfBx7dH1qqbvCl
tLt+O2MMHNyoQlQdioUD7kfs8Qivfsphn42+2AwvZRNl1J+6WJM0rR6jUNkXvF8g
EmewCksuCiYQsMZAV5r3QTj/Egnmpzu0rltdGV+RyT+fUw6DHeqpaOxcKQHkx9hW
uXdnY8pthEWts42xaxLmYyKfnEMmjwY0lRWLccuwA7bLSK3pXgZrmOC5pLfvYlpC
FOI+pp7dQ+s+9idLRHirmYfXuLZiDNo719kX+HBuh9AS5PN0RY1qkg4lts7z67sF
KKg+8ovQhgwIxxDJ8qUNv1rAxA1sHVTm/33DpO+iSBVDKqjdZNZ2f6mqYbseNzHi
lQU8xeSV39+OO2ddI+DeKaX94R0ZtqSD3xSnnTGCtujFykVVQzlJdlLKyW9jbegw
CIBg5PVar9YsNdyK0zrYYeIUC8qYBVwpCDm7g08iRtP4IDIIqxM5oKQOShHlU+s1
PEbEdZF11Mk0XwTYUDIe1gtDi4yYM35fewIBz/kYzj5MofFGUcb2oiV8tOF8+uuc
fvibsuNYehg0ZbRWDe0PsekMULqcsSZjEgzQ0/JwxD4djvvsGadP5T9ZVb5Mug6D
vIQoYojYNBMrL19EHplUwmM1iPT8IbXkycougSWghbiu+hGG1OsFQgdrexeFuVwB
ofDLzn3umpDca31nEfKoEPC6D0s5W7lVnVAfS5w2maRu0nOUOj5r8DX1UY3xTCIM
1f7BBAmtyAV5MNhSA335gkHjI0teZNLf4uQMknWppf8UVn5I5KRZw9zg+DuRQdHN
+g8yiLtpq040Euuk5TpIyMS0H0Acloidm9jxPIabzbV9VvTXl04jH4W53rVOtlAx
RQHvJmSLCDlWdcIGUjyzj/RXm2nXkImAHCWk3EpjQgN6hbSusSS6xz//D6waRQeA
Z4yWrJtiQRsQQW6xUqD/iQwURve8lCt0oHfzidRb50VUjhUx06j1FQ8TdkCCUzwi
0zekvTFeEDLHSM6EnlOAYvNgn84c92FhdCiSukbUbBHs2YpzA7GBQXHAdfjXMtO2
ys+yeCi/AgqXu6ckvI7FuW/io3qUUtKhw8wPgz6vfhYZSDArN2Ou6wp1GCcBWGir
eZBxDr+33TQ7B0v20UuAmwlR4y+bdWurPWte3FubNeSN8E89QclbMT6T/toONqa6
y/8qnMEP5uJDBjwR9vwQNrDzZbfaNtMb/j6ZAfFwNU3OFXgrInwP2O2LtUIfEEtF
75EjCiYUJOVKafl1y7UXNCd7gG/+al7tGdaYSkhHOLyO0Z0pd9kOTnxhdO8QhJQg
leeLX4E99z/nbI96VP6r1kuAPS/2qh1sXr6dJ3w/PxPZylGyEXTZAtJ0kLHb5lsq
30Gd13VrXhMgeGuvVAoZdzv6cIUD2AdXqciVjVxNmMCJHIKS1GxWzQkprUGstraW
nWvIRxoyhFYMcTItb9Nr19vJntgzEfG76n3VPT2TxnpV+98+/IIQTkejaCpa6v5F
Mf2yPSY5+nAztQxe6rwP2uMBnwY0DcdzERr/gWUaBonaLrv1JuBco0HtwUqlqwfH
K7IqKOTrxZ1FQJlMIoHq+fTNJSY36iZ9ygHl9XmhmSFauXPVIOBnXBIbSRmAIpN5
PyHKzFo69FkJiBajSE6qnf96hnLM33S1lZdlcb7uqsxdos6xdC4xm4sAzmIEgZff
tnatapZtExZBaPlzwJ+F7/YR322ShlFSO/VO9zK6d5p3DHA/pQGyWL98QE5V6Zlo
LNcuB4QqoN6d5S4IH/sziBvOQzYXfJEJtJ9TXDIa4IXN3SM0s3Sq0lxwaF79X2B0
RbVA4EY8UIoOvV0Sf6wk48CT9ZuPrBFO8wlsIvtcXy9jyK3VnqTcHrRQcbTd7kd5
yaVMqS/EAT31DtkmQJvL7emxLasHMSDPpa+RKd1OOTk2RKTQhIZ+o038SypSRk2s
Tncf7Bc9DrzgPIVMOYGFaTXFXbpx6x5TZz5KOx0+nNX1zobuFHzJQTHaMwGcUyzT
c3VN20MW4/SiEp/z10UtKi3mc/NAgz9sWsp6SSI63Ua0qk2HNTUtiF1C5170Ao8V
713yVjHgQGYlEFCXywYhQHgSOBZLX+KTIMqZWR2ph7CRmyewMXzuPSRfUsM4uFEE
U5Nnqwx+MKS2Hkby7QboYrqIepzKdh4L56Jh3+oD803ye2yhheScuX+d0ymBK67G
5S9BZJ+L1+stiWFsbiHygi+YJlPGNjULg6z5+L4/COYb+WOF1keGy+NKpv+fC8Tx
wuUlLr5+w6JyqzaqcqKkK2xB21A9wR7P6rzwkqYmRscSv+wQz17aA5zR2izyNrVF
o+Ya5cX/9TuohUYOVMlyBlGIfugYMWiArsTU2yuam04TqSOacQtEm8HN8KR6heHn
WukbqMpg3A5ZHZFAYm7UuenrPHfaaMubwvucG6wFiZRf9uTxRBew1HKQUq6unVgp
aRpsEh3ukatvltbaWmTrs7HXDhSk2Z0aoBdmn6oImH/6acsjebJvXA/lIVuGEL+h
iPpaMWpOKMZldt3tcZLBECtLLBeCDmppTb7UaU7RUT5Lh8ZZmv0mFqBtXCuZOx3U
QxJc/7jMk43X6mwXcC/dtiuj3md9pja/xZBkLwKBefSC018geWCf0i5ZCSY2vshc
ctVvCYDFB5JQ+ouv29uocJEJ76Fc4zQ2aW9zT+lZc2bZQhmELyjfQiyvMxZja+cV
GQIsxEvqszkDdTuHn+gZZq77IUkarA803ZwiVyhP8joGrOhyy8HHpuuBpOLTQ1IT
+QwD42ydFgp00nYxCFyh25XLZYGRtivS7e7PrtwlcqBZxShPXQmjkrgEgaYFadNt
LPTI527MDLcyDBM6OiiSYs8hKhpFkw0PF1G06DqzZBgdmbT10m5u9MYtwLCTuKVV
/VyjUJEHmH4CzdWQllSRVjaKmzJAQc3LM6XKjKDKw54XiE8IF/+Kl/zmLBlvXxee
FsHmRBRGMJF21/LHVKPV5MkPMFCYZmH0kLcrBVuVWmwUUk9CFKb6PK97xjGRL/96
cfrXO9OTzBKyDnVVpoW4r2BX7EXETg2uv+oQJW0+22LYCp3VyYU5HVLWoZ7RxJVx
oC7TBZeKQrHPr43AeGtxpfLtbyfBoNs4YjzBaW+5uYd/oF5jMxTh2v3odMp+2mtN
nZGpF5fqOyngYOBrlEZj1Drb4APY2ej4h8M/ZXQposVxxZFOMx44kg+G5fTP9Usa
2bOFVF99TvFETbF/7n4aESjg696KV8BNTfpnqtT2iZhd5PySy+E1Z8FdFOeuztdg
Peu2PehhYSJSZcQhUrTEmHPHoGp9ZwGTL3d15YzO6QnpGHDHgJPDHLR7xYFXJjJT
uln7DzvJRKfivuwfGXzlGxptz9gtqoVU2xHuqQ+FbJud39vZNZvSIXe+og9ZyJ+n
gCKi34quB7ZeqgZwCdZybc70NNUKy6eHVzZJft2QlKtaesLCOzQIDlwjcZO9pZdG
z+5Qkx1tfMprojH/Bl4I+2cOPleP2DVGnkHYRGtMbQPP8zMzhuOZedAluTyUtBQL
Wr/OBNM/m9J6Bkc59Gp1Q4eq/2cdLzlubHF/ID8nFtTvvSFpKapcxw4QFoZY6Swo
zT3hN6f/YeDwgd9aYwneKw5TG0EO+eS+AHOsvSRw7W9UdBNbXJQfkgbYGrMw66Y0
B9WRLxnsWbsFGHQYRnZJ06iV4LeubicVkzc5UdEfLVY3u4Iz9N6OSiVtH/0IXHTq
rCHRBBRYCh/zpdDzcZwx70nHEu6DS9rNtWi5DJ0jkS9JHqeLEO3YsfX4ghhqqV6i
vqf/C/Tq4KFoIeWR4BeRPZoSi6I0pwoe8C5lf1qSMuZsk7Ujv64h776c43dcXjx6
xDFI3WSURkx+16g4ASr3U4v3x/fxImMLTYoXTlMDVshubNd+rlU8MwqE84YhEZeP
Tv41apyQs3WzchaylmqYkNl54Q0dVPh5KV1KRU+MKzxFk+ow4742WblRp9PfHMJb
EEAt/QoJ4wZLXlYxjf5VqSn2qMQduQ+V5RweMkWnKlleQKcNIDYUKo1qBrjacGpX
XFisSlqqPwFonwZdeeKOdVoZe99rXUJVE0sWc5x2E6fJp4d0U3gwfptJn+VJN8WR
GNzDnMeqzQbp8c94ZhxNWl33yFG9xwg2jSDbPi+Sv6eHH/6DlgboWgD8po2iPEgX
x12XiE0X9BwFov2bN1zFG4kB7lIA0ZatfG4GJGlAVM0xhfkd2APArB6ymazoeJ9l
CVDnPH3LwxjvD0AHWPzFEqOnH495IJD+fyvLu2sv5Sjm1P2969A4mlUpOK/+cNa1
L3m0kKs3eKnHAOXaq3ZaOGAAwpbj8rI7g5RlQArDoYtTkEY1tCfNnsBGoi+6oWjS
AukjU3sFsTKi4n86QHFk9bYFkLHAFaPgMdLX6VieMJZtKuIaqq6X+qdU9Ax6j09e
HMPPgWg0iMo5N6z+4DkZqI7ufe0bUrzpdQIzuoD1Doos5WN2D6oqTaxwTGwmtoiZ
p3o4zUI3m/5RHeomL3WRdj8OXApn763yf++rTrKxrU9oJe4HsIdacnosfrrRYsUm
a8NNSdeuIPwzpbmPNVdTg0iLJejoh883eCjD4OTo1k2fPXXQeE/kfSqxcxZAnT4J
fT9iR8GUQ52ZHvvlA1qQYWpNw2/LzMXQpMZJJOFjAA5ufYSOC3oz0Mw2Pd2J0U7J
YrS5IcCpvn2afh0ym3cwCxee8YUJgWGE3Oy8RLgVTtMjB7oA4RDDIFJF4A0a8R9r
Qtx0AtJBlz0eNepOV76m9NmdfdjlNZerihetHkm4DNB9H1haNJ41RHa0EwV6BTj4
M1P1LWmsXdLPHX+SNP8NntmheIzQDfPY3R/D6AOV97a0NmXoso4lpPE0yhAv/JqK
hNiaxIlPfNI5IdtQ/FW7gIkdwae8VAsE1dxNs3Glw1UunOiu8qHRXrOYlCv3AzLo
oZSd4itdqTA19OQRxnu9+Gx7XBzbJl5JHpGtVyFQC1fydEDbEBrHvs8sjAAFePsN
qKvpKGi4qyb98moiInoQ2fa6uNnp7Eb4RnCXiCPcrCPbxknYlPPtestc80nebtBv
xkwuVDYzKNBsznkAbJzOGKuwdy4q3bZs6idOH/LWS1+iwUOsir4E7bcEJBKfELDq
9lAnKNGqhFSfF0lunOmIEVlozkqzEFxn+vz0b6VHNmAMo10T0t6UFAvPdMCl6+6R
RQ/c8IRqvBOeApMA8sWIIQFrSU+zRqw3DmEHvA5QCI3a2FmE8QUYm+GkSlZLT+Ox
RbggavznESr4WWLSLiwG1ECqLy59gFUYc/O00ZRA2+x3U2buXSzTh4fA4/uEheiM
RWSaR2+URc0yVPTWhD3qZujvPVoG08Z2Y9kMjLBpDMs8WThozQT43CSeLDHr7G43
DbtqBPVSRS7nvckesha+T4De0/tQz2n48ZR9I5U/yWAZ0ZNEhryVByfz4YO4xKJD
FJ3YkFLX4YWKp1g0q53zumVAwzJUrCIsS8Zt9lnz8NE0rUQQvhpBXVzHn24DBCik
kBpvsHJi3TYmL/Rqwi6kl1IsjlyCDpBWK/zYHI6QoYXm7Oy2OY1EpWEpD+7juc+z
31w5xMeGYzBuLjwiasd/Mpqoex3ZQuof4saoRMtBjOi5RFzzZbS1n00yJkVtJKF6
yKxAS/Q5jHwKJTIXcIYDl6KF1anElqZeG9Muc6+B52SSLKJSg2hnPXXrEpN42xJJ
pCJerhFY4IW2gbAl+JezVdSHV3fEbyEnIXCseBSd1Ovecp9hG0FLOpVBc/hEX4Qu
pXZd59hFzRLt9+H/uSnLlA2owl2eHSrg7MJjEvbKB471KagZ7rQQI5/Zn1ypO1Me
se/Znw0Xfm5xx3Z8wPydXmCXNqFFBcBohrXaWwDyA9E+CfQ1zsqan5WVjuVTiOGX
lzAVW/GfEZZcMMoMaROcVrEV5IS/g5qoP4+/bkJE0ONO9KNdVyyNbqWWV6C6pNX3
sRnfPlqEl3rXDJ7BtrcN0gzppdWkc8HMVS9I0TjBo3BVPIsC+2zDMhrx3ZxHi+Cw
dfmn2Zttl2b4x7hhhSLdgZ4CJHmFrjK2aLlGUnkg4wj+t8+uPrWlOrxjO488I6nx
XAzOm7vb/waX9aL+dQmGCJyY5MsCEdPOE3cJJFIeoEE/f5oB4NG6Q43YMg/rR+iP
mChjq3Q7Mqux0Ni01kkfRADl2LVBb9a9ZtBjtWa+0YFTXR9iwNrHgTa2woooMv91
2UgagxHJ3EqyJP0JvARO7jSL7TjDFMhUgm/9aukIzd8/LfvIxNVkKfej182LZyqq
vBbHe0wYrkXHMZnTWBh/ijJXhR6o7KuXhkkLCf2FOc+sWxxf2TlE8sG9vnL2dyLQ
sJuEKoqU/BY+D1DvUHHYmkxXawXzVtin+JK6I4gj7O0kB1bK7A/l1WCtXFrOzvKV
J3V2/mDiXdWvaYadauaHekgG6j/fWuqlNPDgffrAZp5IwHqrVN5ztgxQT+JIRxYl
oU17bs2D7TYuoxH1R54stJezkhxD5EU32KUQs5nRJVsXy4Jfg3MTPzEzSdYEx+JI
ClBYSMglWJWNSZpnzJ+lx3MQEBRhFHeuRtg6wMm5YpS0odK5HR+Hd5wyYRZA6YTH
bbg13Kg28g0WTonzNLIqm4jekpFlUOKXdgq+Eoa1wKkn3YmWqAjGO+7xyCs9uill
71ptpOg4S0ZlakjCICsPOpGppMNvhGIY1KtkEDGHmdrtTSkzAfttI0aY5/AsSSUC
65/zjmhKC4Zb+i/cqH4jBvXY+zYWOT39ZS86jzoO4N37N5VXxGxKOANwDHuq/fGw
xIdKoXMzVICQpR3fP4C12jQuSyrekttsQc2XZQkHf9yRvWKPxS0kq9P4z7hBFZZf
ImORQtZyFRITbpGtW9z4mEpaIvWuPuBes2ggsP6/60+pdAoJDR85GHCCro6Myb6c
CDC9gws5YXBpc/vsu8KGO3VdOh+GImSRpzBtz9PDR9rJqPcqxsU83QC+1RLQL5Qj
L00jk5EmlocO7RMl3qFlSy5OXywNVJYSAlk1jk8JrjcvrA3UQRAcdAxmVqB3OfAX
NvARB3C/ihD/IMIxOGTub7xeGWW9LKyXuu/T4NbV5vqgsXtXdoKEdljgOEoxRKKk
y4eDHgHGHASQmvQlFylDpM6j0FoGIMqNI4KD4YNHhEt0iFro1a/9T4bqs3W+GEim
zW03uqvjbyMFMcbMbL2lPHAyuen4eBSy+T6jRM42dsieQbDAO2KSTbPLvbVfQQIi
My5vIquLi/L4nxpIOpy29Ua91GLM6GsjhORgC4lDn9o4yRumoi1sFWcMouN1ejdc
vRYsEUr68r64wTEcpOjsn35kwkkNX3g2KutqWtOJ/LFv03hSxSeBz6g1azSZ5YOG
qXzPCMlRwhx5/YT/EN0DgAS7fvICvBpgwVLYMQJ+t1R4kDYG9vtm+72xJyd6voDM
cYXYWsfVLTA8+U4JsoPlZnno3icHg8Z/qx7Wiin5KyWvxNrH0ztRzLY19k1QZLQI
xw+qMBz2nkk87Y+ofUFh9o3ECAio9zVGj3NrkcwsISZjE16E1PzLLtl18yzOzYA/
BG6b4cFczES5djIhB4Jz5sWafPaB6/iBOPzVzvl3OLU26zlBl4/HW2Izsp0TNYIC
hX7WE5Cyr9fSpc/CTvRdFsJ3s8snHO4jUIOu995+1BOF+e68LLXC6WozBhnzbGg6
v0kCZfS1MKNeP63Y9TnuedW3EYaz6ZaxynkivRWyy/eBoZIPwuc2Z3OhGf+NWzga
aI+d2GNx4UvC8WJrkkRWcUgvPm0e+CldMUxGfIcKjQHPZ3o019/XC9GWPcmrVRXa
nRLYaNPraHZWJqvUI0goPkGrZOnBxs2dUcGu3bCIzqiwtUSzQwW0c+I8vCwy8AZB
n9q0GVKowKrpTWDEi+R8F+DPXoLHB/rJtP1YCZMvQ11wHtIt3qq5uLqaKZeQqg1W
I6xi4AL/6+ktpL4XExb5ypbvktFPT7rYS+miKl/RFCkdIMhc0XvcAFIFz3MtHtLc
qjMfc4wgGcHcpvn4s2Xm8bqADoeVsJGw8gVHuwjUTpM+jBZR3oc4oEooC9jYwUEM
7dYABjLOa8W7BJ6hB1z/ctrdVwCd3j6/eYE9RpzeTzp2kbGUuui7J0+dYZP58TWB
tKxEYxyYjhWfZzohmHOuBpUelx03qMTca1R1AZjaXBlZq3/YgYVe+GoaFyyUxWAT
cVFjWGI7q/xm9PxPcc34dUZIIDhxLznaw67WWHP8jwivC0tILdJ2eIqfzUmL8nAy
Dgd7+m5tKchMYQrcOipSzAcG7OMsTA4XTzoBEQlPPG3jCncTFT4l+aaDzCb+iSoV
pN25BVyn9YyrW/5sNJxCB+jPHXO/okdJ9SFgNQwdjmGaaMmycSg4Opxf1ZYdzOK/
WwIzGgrbCve4qj/iYfldoQK17AP3eNFz0gQG8YaQggvqF/CB+k5yUQ4SlBAKiTmj
W0vbrd0tMMlmUJUEH+dvkNRAAP7Rz+ACEUM0Myl5zC3szw/6bAGzHsEskkC82g1p
oXiowchFX7VkNHRgPoPydRuHPXVTJE1pYavdv2rshFe8YIxI2ajPtLtC9ikN28c5
jzik0InN2oAHvP41kHAvRgyabi1qfHoGA4yxtvhs5usAIIUVMwKFRay4fXppk5ZD
8hFyJaeKxlmslQ4kZVKRRkTfd6NJKfafxvOry4kbsz4vtB0mNgXjNifrdG1gv26w
BC92gKMirLXxM+fdShFUmCtk+70kTUN8mNudqzzNpSnoL0qOVF7gLSvbZp16R+II
JITvQlyyWVoXBtTRrK1+Ri+CUXkrcPgmfB93oq9z5VuNZGL4ABC+Qsqg7nBLW1K+
rF5yMEJc+TSSB90nl+VZcDioRi3PM8ibrds5SAuAApk0Iyp6O6Wkgny+ipWlFLhb
rAjsnEZCvn5E6GpgJaQEZtLO/ZUdhK/JGHy422CeNA6FnQ3R5PEo+Q5bDPrgfWkj
q10k6J6CXsR9jjzDYtaF8vIFYRd6pIMgi2wIQL/KHIMPHLVDtGfD9ChX1SEOoVWV
AfUWd7nszhkw6aRY3ZhQLpQyoVGLM4wqW/Z3NkYaBYFPreAZ8VAisYukgoNe+nBt
OlSeyVHjXMceMwCn/kf7kW5+GYIdid81q1a6zNBvoL2Rvm7iA9t3AIJuX53vQOFG
vBDddgnNN3Yg9M6zihAFwWPsjoWLr8LoI19mOBXq2eXj2f8uBA/QMhxCckakGD79
G4jGVv6fy/i/0tF379YYd0LrYnp95rnbVcsTToTcyl4d1XbReE+8Y9ZOjUZLN7A9
ezj4ol86lhkVBEnkyldCM0tgdXirYrucH6lVB2GBJeqfiVKY1jysyrr7Uu6LbnEb
xhttAO7gWjRibnxgEbVtvl2MQsQKSiA7Tv2JAhcacuafYIyhucO7+8Ts59gpufd4
vwDmpNkw6MwDq1KjPfL6nsm1RndKRZG3f7CBo3oF7NgCPYxGbudWdMCu2dSSTrgh
67xfc+Ek5L0H4Q8UdvpI6p0mZraLMFW4aBkEm+Kgjy/zmVVAfd6m2d2D8p7a2K4f
U5vjvrsyiTt5CORKShfQ5YJNls0PDQBTz/Y2l/paJftuFeQa/+0Px6r3QeF919xb
BLeofYQzJRnL8l6xweQWyResp0RjPX7bnjog3YoEiiPRgF/GGUlkLLwA/CZRxOgz
2b2Wq79N5cNN62Ceno8FGpgPiTjbB1mOQJzUcY1Qg4BLKRWqifcW8fFllVVTkZvs
rbutzlUjyv0VrOSZQXeBDtQk641DPRBDI5weZAJ60kaKjtWVN5dTJ1dDm5y6fzUf
o5tfywUcr95FaMWuX4iBr9GJXWQ3dFfYxTfY7Bw5VZMrGoUcbEYs0pCbbTDiF5cc
lmScWK5sgNx44XReA4IDjr+BzbQPaCmgkTRfibcxeNNM4ZiaSI3tZYZPNNmn/nU6
R0n8Hw4LYKB8NGwdubdQvRAqaiJaWW7Ed7OZ0VZ9sLUU/QPkupj74jo/uBAtgwb2
/lU38/CDvLU08Lq03sCQBNoOjHddww2MvvNZEWR8KGCAYiGL9GVXa16gENMNomNp
HpJGlW2kdmoXH4H/Oku+4Jo47uZ9K9JgfG/1K0CY1+Q55c9neTJoE20JYIDdz1eG
XsSqgVb6ETS0K9qdMxNGFuJKHXRVPliswiNF4KkyC+kZFOPvldwbTBjGI1OlwS7i
vwjv+l8czA+m/jRjdf5DoPxnFbqRqwH6wvxqGTh4PcWu2Sae10SQYxaYPoE6nUzC
HMiCux2qrxhyLSW5FMxFJ2s5BRrWfVIXZNXd8+HoJatZwTJVzjreZxWG2TXs4d+5
6FDAsToF5yiC0K76U/ot9jnc97/S0ToH14Pe9cQUTlDPNDrbvOvtUrttQmzBwZaf
NZbrvv6bjAahGQ2rcpa4oddARpzU2PdFg8c0lOmVwzFziTP8Fv7qNJ4cPgECFgf9
km8st3tttUUnstdCytrnBpFhcK6oPn13MtFKducK2dOnoS0QJ+VfYLoVIH/Akoy6
P6lP1yskCTzVsjwuNITqo1X7d/FgfPDpyPcQdpBI4t8fGH+Scyn+r+qVugcKBi2u
wpnKsm6d4b+LHBVefuuptqLH1iKH1RrLZ8oQbni46vcY/BzjKWSeFEyhH3DX8pcF
TqkwPKSa21hjDY0u2BHDfB2UzaUySFWHGbjKAFBYevk5Ig8pK9By1XdO4EblLPfb
sHs7eSeDPmM+GVRZ9AkY1IWRhwSrS4r0YCvlThaNwRcUaT0SJf8Wb2boFGKa3NBY
xErFfdypdBQm9EcQgNZa4sgFv5p38ydBrPYIyGih8UV0jQYpdAfFkSJAJk/mH6wL
s8Udh7NjuyG8ZuJ7SdICksz2j1Wr3jzcaI4/0q6FLIau81YEua/Bh23Z5I2/SOwv
8v/MKD1vFARxKfz0ffdTZ11p6JR2+bsDH3hF9Gro0sn3ciPKPaRcPIANocfYYzGC
qQlV8HllsqjqlbYzapxflmnSwO1xW2V7l+ZgO+mn1nbFiElw6vtqn7BQht3Qu+Hf
PSrwMO7rIR15NEpJznv+Dgyk4TzkvVunkcuzdShPZ5sD8uksuugRKiS7eFn+ILcH
YAADJzcACHe7W/+t8x7CdaPIzqHLXHTQV7jGw+IimjNwvJeop496u/pdtY/k2PB5
GcDt+ELSsfmGFxIpcQg7D8qDawDp1FIw42s1SJgicqaAZ74sBqotmqMP3ortmcyf
6mv/Fs7XJIZ6Vh2mtD8Es3sJs9D6EpcAHuT6qr/5qwECqUfw23bX2Xnc0RGJ29Xy
qIX0V6CSkE8vqBJAhrI01hVjouJwLGLfW71SRGzHZ+L1j+KgBuslJGWjVp8WJH5j
Wmy8670QACToWwuf+GMVakj+051KuuKxQNOakADxhVYBSlohiS/2jfS/XZOHKwas
3njjHtr7W37j1HBY2qkjNhA3u0Tukq9dOEh5pzOySh6ZCfY9lH0n6rI2sC+SCcnT
wumDkoKDHZdZ5QClDlvjxN1vS4f1ktcADiU3KWyNKh6l4SMiE6IBsRslAqQmbnob
jCzN+SUm1Fe/QDqs3qWlvaar+EZVfH2/zwdzjjqZsj27PXZq+/TEufVl7qRtmxzJ
24uC5pnfPeGWudp74x3gVcbkmJfpod2x7tK38+qoS0tC6KEdSWSVCmFyW8JFpHNb
XtA4UFy5Y+aqQrPhrIctMrUraOrJKHL0/lg3n85yJEJbnliJOYrvhRbhqtvXKz9P
XKOu2W7aT4lJV3D68FEP8oGY4q/bArROQsCcioW3g2riklTQHh6VBcAVmJY//4Ft
56LUMTYW9v01KaQRGEbykZHWHqciX6uxEqQJCbRH/OTpVRPUqjOtGKhzsbXM5sSA
J8ijffVcq61SmzDz7CdhpdiRkKdor3fuKDe5kxyjqLMRV0PtgI8kDw7xxxB28hkO
Qt9UmUpd2ug0GRJIzpr0pR38Y/uM5W6covq7Xt/6SwjW1otozf0KcR0YGzd0oFpV
NWytpuh3d1+XBUUVZZnKRo0fctjNxSkLKg/MCJz1T3oVVMlRbKv8bNrq2K5LTunq
SEMatM4uTxM5AxqAUAKwz+mJ4GZa/H+U+DCeDeGFv6HoI6eL2E4gHIUTxInPjzxO
vwQB9PMc9CYoWTnINrJqBREtkFTEs3K+5OzQnwPTX2A83K1s1L5oyuYeYmAdOma+
FlGq7SxR3drpDto0n+9YfeaiIo7H5i1x0A6WmA4HDLMGvp4YCn2ZIynxa1FfTgp/
1mxCXWYrdw9eVev7WUJHuW3mngvlvUPCyrXHO7LIkQQ/WJzrQeCzu8h8jSA4ssrU
b39+ICBzGimzrUTRbkhdTsRgGOFJ+r67N1sU05pjMo+t1f3JtYh5d56akjnl7FDz
YuBOHCTVIV9n7aBnPVKhwZKA2dSYaXDS4I308hahLrWN2wfYfD1sf+6Tn54ot46R
l0/R9NK7E2rpMv+HN89nb20sfXCtNtpLgI8GG3BxK9KxTpacegORgZ8UjQs+u5Rx
UEEURgOnnhny84Hoi0whH47W1VJd5Mbe1Tei3QZn2OzP/gG0PdV5gzjegPm8TAxb
HRAjNEi/MFvJVR4Yj5HqMzXHAiVQFr0zOPoH6BM5vQRRVe43uhZ5HAKvduTgnpx3
lo2ePv0OGskcL5hHXiFGOSl/yNdsGmwoYsZrXe4nZH11kqxcQ4Q65RnHiGS+Ekjm
X+J0wexkG65yk/U6rBCdXe5vAH5b3rfDmiUdr00geDOy8nkK2jLhjrlQdXhA1eZo
6Yj8em4Ewe2GNGXzOFmju25Ocus86UKEUk/bjfv9feNdf3XE6jRZ9IiufSjpxD9p
u9Cw9NMFU3BWUZjgu8lsBNl/6sjPonw6MEENvcP4bTsDIHrc7IoUT34jhpYYVtOk
K2im2oKWBctKyh0lLs4H3niqx7wHbgQjxanummIP73GXh/Fq9YRH9OFbgxkW2pnf
ZlW9+0H+nXlK/JrEqnoc0UOMtl1/RBDgWSWGNmmfbMuD4U9fBAAMuVjqFEv3AIfT
twCKNvvnbv/7Kj+l79bOfLJo66V7jC/0XbEp1nSu+q53KHsyk9QCEpMbL2s6SNf7
vt4mNF7z4tqp2bMIG0H+FsxVnLTSQSjUiwx5u9tdRtWsjMRD+fmWNs5EMBHfRIu1
iJk9/yyNDDINV7WPJd9FsDswxzNyvWH7BZtRZ27L3x1qR8x2IDk9CxOAWfwd8iaN
AkvpNHX/cxnZi6/9aVtlMByTANZf4ef6CqoGUMnDbCenr3jCzeBCLlFrGfwseC/E
DFoXtADwSkrcAADxztYQf4voARihJ3kyD3OHQG/cAKtkXdnOVCLQsdU95l8S1UGx
42bs58gZKO8kJCfhBi381Xx1LRfJPlGxNIc6+xFf+l1N+WKIU3BlT6nWOMJLiFp5
aAVLfNwTiTMf9HCPjd5OqbtcvDWhB2ffuXAtjqVM0wIoJvQQE9xPOMpblzxQgojU
wvtXa9flqhxz2aAtgvfs6Z0jt7NucvxT+JHKlatXyBAK9smJP3xhVYMrx9ns0RVO
6M2386t6DKeT7892oQjEWNaCbEJ+BK6bgDTFu9biFQbd1dKfDLcvZW/eHxW6oJP2
tuc/cvn39RoE/6ooQ41kYT8PGqEqhmn26qK2u8jS5TBJARW36fpqKjKkMjg/tnGv
kSlRYX3f9OeZjnMYLlrUH4nEoX1qKEUFbTIvTuhJexhShwFGwDNJxhV71UaggiF2
z87sorF8k7A7hUWhQj7QRpgMr9I879hxB8LaHU1pK3BsEslmKi4UXHc/hd4ys8kQ
B1KutOcEGeX0l5nIL7pwl9mBXbEbZm0zCoQp5ohfTzZAoD+jJyPtDCJTcvebDLNh
FQhWZAgXuqzRq/eGRJVKuIRPau3bsNhI3+QmiAntQCmxlHJyHAn8qnKKtdQXfK1R
rT66Sm11RWQdva6dbgBIDWnB0IoQIT+MRvA0QoXPwNCMjQviHI+jq6vlA0D+I0H3
rHzx0XpMUeRvIou7K53v0+9Q12S/L7ockEWf/s7uyBmnuwiy/L+44FJ/kKjCwFi5
4lAMRDpaPDer578BNvW+FhV9wjWfTkQ7RZd5Nek/++gbePsQ/ql0ciYARXMDvzib
BLrFT+gy3FntagYeWBqs2RadGwteC4lsSMYDvP+3qf0VTI3XIqb9uvJMHSCIzgX3
RU0N6P9DLBkL99yoWM5hh1nHm8Alnu37gUZN49ZfOiy7C7Op+6hqLseegiA33qfD
OUg/J2F2FxsU84cgOf3Jv3EOG12tYWbSlEuo6ob/5Jog35jxakgIiQk1I0Sh5UZn
5CtHD18+Hw/JlzmIwo5yOgp9P3yioNPIIEph9gVJXLtKfwm7tagdhupTZCpcG4ai
f+az4dN43XH6mjANhMSKMzMWAE0+iWVBoLv4l3TESJdKK400C4rNAqExfMgWkGEL
m5LXeY5BwyCaKMU+e4CTB2JJuBOM5cSDPAUD8wkeFzth10/wk3Jvkeol8hOl7DM4
Kc02mHJ56HnjZU0/i+zD8omb7IAxHW5JwANJp5y35oHI9gIgaGgAtk/sT5y2yPK9
qc8aIrmdQX01Zm1Uyouo43QVCEY5fYEmVy4H+N2aAI6ivEwc6JeBN6a+cl55zKBj
EaNf7WVWqIkEaJ5GHxMRbQfsOIi2pITdx/6s1rGEMe3w+fA5wec78mfz0olxjOU+
7RIWh6RaXIN7Snx++BQLLOx1AeL1jtfOgUjjodEuayrr/XLl/0KQ1xXKex0OiAaE
SbTGCO/x2S+nvmOM/RE9yT+NsEsAeS6aWlTyX+QMXk0V2i5kYF39U8ToEJ5gBkPm
fo8eCYjY0S2a/uKvqdRBZdlB5YQgiBecVp0sUFbamV7k7la5Pd7g6zVMyjZ2zjRx
k8srTH3hrtG50BVVN+HJMoUMEqk0wkNMzdNClMF9Cep4+0U9mpF8XOGbnI7Ulkqi
/4XuRyUgK3puyNrUgm0dBol302In+LofiD0vgQO07JXadCFRxbF5RHn9gAHrDgrq
nLglIR4ny5KkQMeS+znQrInh2sBaJBysrbQQWH+Psi57wYw+5tcrV9RrpO4Fvzww
67v7qxruMFT2+5AQDTUSuliXjbE2jxkOB1HBj+K0hDKT8XLA8tFkCZzo7heCdHK9
2CCAK6WOaC22jyqr7zcWfWZT6Bahx1KKLX7AtnzqU7Ea3vr5kggMcc75lARb1uKZ
zY72aVQ3i87QANr146fAON1MhMRiQxDjBslNVpLovp/3qTugmPsVkxO5P6D0rxsT
GPfUgSyiiStH41St0mn03K3ElmGG4vDgNQ7VwdkEYzsJ3ce6KzDqx3U96aGWBn4l
MLtoVxX84P9gb77l6futHhB7Blv/vcNDl4lkXzszUGlBPGtmBnIUlMy1jWRpcMb4
jtfzic3ggMqclUuRFLwIqzpqMG1MvsMwsL9rr1kTIm213ZGjYvL4tHJ+lzeiIC60
BSfeTDOJLdakTT6d1Ibo1SrgrAXqP1i5q7WhczTsurXrJJ3xoDbbzjYPgXZe2nEd
HYAdu6pxboNXMaDQtxNHMi+NFi4ihh9vnUrXMR7ltjc7HEnDCGdmmogsdAoueAp1
mwLkwXzOBSxGNN0qW7C9dl+5xcOGiuVEUL+sYQcPSBU3PhzTBAgW9U20yFbFcdo7
JO9DU33fVYAgofREuhTijcRWuSAQekq8mRuipFr4sU8Wm9x/yhA1MoGsIwNyz5tQ
KohWtO7zXNdJzrCxe7wAXxjG1BFmhmHEPPLOzDFpJ/sN9njZVbu4YakHkiHbC+fL
X4BWMJDfiKyuPPS/LZPWH5fBFQXX4EEAhiW1dU4lCxy5p3vGdDipjFRALdBD8IGC
KIA/TVqNFIl2gF35tbbW917/lcELN1dSOPH8l/KbHXwrHRFtcd1IlwEY7j95VQoe
mSqwmqR1nZ/qHO5LltlAjbjB7b8IfAshFOAAOcKTZFfoUT3+TynTn7hxvYxabN0n
OqFSMJet2Q9WXrKPm+8TYKq5EJu6WMX1P0oK1QNzTbFqyN82LXBA3Ka3sc6S69Be
MqFDtsh2RX8vVtYIAeFuBCNgXkkC8GHQW2gQDpStmYXUKJkWxtGxGUYI/2gAamO3
Wu8ERaOccgnqmnS1WwQNGssYwUmMAzC5KENHEdw+GsrfbDTf+aw5p8zVMB0vkQoW
8rytqDWa+UJzZEkv3V3qScrWvAkvje2Dn1CsoLhikU430JteVmT5jOGzgAwrXMTS
aCyqfwhx7Kvgz+PFYs9As0vv4D6Sll4ppih6LcNzUENwF8yKruQafh/MosBCtoJB
X7rl5I/DbQXRJfTnDQyUdgF4GowinQ2l6FX0BHA84IY2bRXQusvoviLQ0P+tCGaK
e67F8Nmc6JxA+XNEqEaYESKJQqADvnN99gOUZgSTZD42+phkPJPvz/4jVye942OO
KLSwBx79kL1F0F8dAh8ZTVqsrsQKzVWSBvXoZtMjpnU2bprEN181RCUHsR6Hiw7n
9hE3DZXN07IksNPdoSHA8O3P96zGPRDQaS0AzupgUoY/p2KF64MAJru2abcAD5DP
gVloknPEAGmtun+MRjHKbG7I9bce8Km/yjQjsoRf0W6FZe5qwIi7tEk2dJyEs0NB
DaBNIh2F5/Ot9tRQoWwTxfOTZxSS/iC/ozvyh5aOwYNfSCSgYmzy2BjcUUAU4A/B
wOu2bquoFrK6dqUFP9ZmbH4PYoAH3Z6LwcpI7fSCip/xl8hwzt9qfztoEfZKzie8
3xRaLgbdsFX9eAWKx/FQyJqHJiCL9P18Wvi8noVX2yh1pelJSNrxHlYwHQ5nxSqu
eBRympVQ04ie9yo6HpuQ4nIdLjASF4znonNc9m8ZqaguMd3jWFh6W8zvZcmGCxSA
ebhPBCR2wkHEGcTX6N+CzpWquppvqfQITvyscdyUzdYBiZJv13v5AbVDqf6NtbFX
HVM3ItCLxFV7EH8uyL72d0yenI/srZ/dOy9LfKA4salzsycUvlFV/mDHRhrBsi5g
nWOc1OjiDlC5voE8v0vd7liIuT7JJ/+PKf7kR+3T4YWb/qJnSiHwRE50qhmzsKLk
+1R+T38C4ksnOXx8aw0DHHkqvjoc57dO7Tmy0UC6VBu4cPDZ/XEStrkZldQS5ZWF
WbkqfNGPY2k4YN6/CerWHYZ0+qeJTlk+nPmP5LkXotLjJDqutmydGSO7IA8fz1au
8YKyLKE6KDuGAdIYnXAih9IO/8R9pcDPURi8N7SM/MbwQyvDqThtTRt+ttZpo/Qh
6subok7DHKk+j12sNMLcPnXp07sT7wHrxYC8Hv/A87r3tWTCU8wOSxsY0EnVVleG
kh6VzTS66rXTuIDYPxTl695Sx93EGuIE9gqqvck6f/Pi6DHQl2wx+GUTlMFwBif+
7/LJvpHrFmTVlEjgCOlnLcLoQLAJYj6+MUm1Umem9CgK5hfjsVQiZVJO+7pmCQ4b
8Vd9kj30Dku7RKlMjFr4Qkpy5C8PQCs0YYDRfk5hrzpUxQDgd78OH68M9woELnop
pBWRO/IBhI4/CuDQu9IKfVLZN7PM6gu6yQKlHxYPgL+GQeW2QS7Rto1Ix3RozbMr
+wFf4uCwc1UU5tgnhGH44EHo5njlU4664DilEEBhCJBI+NPokNYjjdld0b61uINt
yx3VCwBMpkZUywUewIGsYg0WichJ/xvv3knWpRexpN8NR9WN3ynj6b+4GxXzbJTl
b18resAcmiiV6bCJTmCaf8kfVW8yClbjE3N998IaGGLbal0LvqMjR3nah3G/wsP4
r6+NYIy3KRzaYWCzcoau9MZrUE0ud2bhHqAlouI7zzEBJTiK2vIz/Rk3yLoUo+jL
tceD1zsPV51Q021P2rWdmNmc1NM1Rhbh4WHwZi4teXr8Fv+XgqmbhrEQ+oEOmWeu
90VFxudy6WWRmVTUYuHb4f91L0CROb+ksH51QpIioaZEiZfKW78KuScyKMgF290e
J33fMspXsAT68y3AvnCF5uIIAVsNbW5TsTXRFH5PVrKqm0sfqLR40TIxM+xbP8KY
hAK/tAAyDrVSPJN+wFV3hg7PZx+H7KthuGClMEEqEMjXkSDIdqTN8oXWt+kinNkA
OIk80oPupnsbi+vWp5HmE4Q/AfHNFmjr+YOLYAwdTkhlYSsYRK+VnDRYdXJ5kMBU
q4s2UYTpNdG1lf3f+HshKechDJe767aCCG8MkF/INHye62dh6fUmCT+O1+/S4dJ4
hWJ8vX0ktdQyfjW8gW3u4HGKuuohW9se1hhsy9w2ZQQVYcusp8U+IZKF3SDIeXb+
rGAtOFCFzpwoumgRGRZw/T2vY4n6dD4oxMI2UWeBEZGvJTrBoIXra2Xjfz6Qt9zf
ipRztW+zMU7Z0/DZG020oluX0HEBCppEG48QDnfF9zEkZJbQ9TXy8bd1Qfpbm01U
RTi8M2nZvhTaaUAOyBNGk7BIRlBlc/qxYUQHc4pllNkRJtC2pcWE9sqsXqqsz6h4
tuqLQQPoyePDe8u8Sq2kVFx9D3iFIjHVU3wT2dLgg7aUtlLjIPbJ/hgdvxira45D
aXrkZt39Y3KKiEYoz4gZW3h1wYlXupFPajNJiXZdWKRp4mw2Hp5/JXSNImO1vDUi
tT2F4osGfkH2ItnuQxBD4Eq1eFLKf8figlgarxGytGM3hcFgcU+YMiBcwydZZmwO
EtdoAdExr/8BMK3MsFOGKorZhhtjyZWK0vaX49y+AQsDG9xIPFxhEENel9YfzhTy
SmGdJlh6sX3N7z5d8EPqNKp9jwYvYNYYU0MeR8z72kqgoyWYv5P2kHRx7TApwYeT
jEWPlROYPBk6tCIeuZK1JQy978tomwCue8wydU9gvapSpFRUz/sazGJZV2ba5Z0m
Kmff5UEoFJ1PoMXssPFRX6R7S1Y2zM9q093VpWCVlASYdpHUTInI854wlQoKKm72
2kFK/Mzzs2HTLomxnTYBn+VDf68t1yaUh808bHqw8v9isoNOTNuOCF4KNIKglC/1
QXK0oCgcZw8vqNRtn0v4c8c8fvF6JRH6gSYUOAmN10z25cLAgVfN6LHtS7yOsELB
0xqQn67Q/6nHc95ZrNd8AJxOs6B6Qtvxw8/zH+8JGvPufmaGTHXHYfMqV/mnMbGx
tDmdX8f17Lxp9XOoJC2onRniT5KBLRllVleUq4V+qHv6hWz4rH5FCpjacO5x2v/e
p6miq+cgygVEBN1Q2cl4D19Q2PoQopM8BNMieErzOFrdryl70Awfq8ORVg34Fe7O
77jrqTDgSRTHw7cXkHo/7L2WrH0E1XRGtQJr2a5kO79Nlh/NK2kbzC0sDeLSJ/rS
Q8ajxoYONLDwDAHXCFFeLx4G6MpwZeusMLs6R207lBcsG8yRd5umOVEhE0PrsMFD
h9RuzDFhw45X/XShJe+IRiZuTBxqqDK8BUEXhYPhRTIXLTd3HYodf5tZd2AMbyQu
HYbgIeAkToYpmR3qNRt+BU5F41pAIV/zxkWV0iwF1yi5YkARiTSJnnEq/2Ix4NV/
+2y8MBgzFDfiTDVCCKmYdRXlQ9slgFZxX+V7lVJl4scbOSLS6c4W6e4fevRdZq2D
w+H0csg0kIoq4TYLKul+4DcphhYxIicTBQm1owhFlk/kvLJDQdN8wiUhCdT6/iwE
w9WaFQvs9fq/Fr1ycYoYmBaVFoVNJlTIWYrdvRzbonDjTd0x5yDPVd9TuEq8NOg7
65uvLKk+wUb6S2fgRmzEgF70gdBxTihJhBg23xOR83WCNE3a+tqo6BlSBAuoMRc6
o/8YcY1SOSISR1MJdTXUQav2g7Xx6BO6/MJpgISEpw1W6saM84r6R0O5x2ucw7Pg
2laCQ9ogcvaJkgOZAbRsy4y09KRA0iTygPht9ard6PNC9L5zodP+nxAAN2mYZMGV
2zwhxkvqz3gfZQvkaTtfvq2M8p3nrgvZxNRk6A9Iug6lI1WiIv7Rd+UtiwULrr67
U340aDZ9jSj/2qagMJNyQbHUw9wD3MakvRtxZ4uGm4QrQUoEnuOBa76iJfGD7wI3
uny8pigtBGVmUR7epvp+1gyAFGENNkGsk9LseqvAo0I2CNxKIO7zBJE6yPbeaIS7
28s5uXcXyvINOw75GINKGIGS+UIijh3K289X/lXWXa/Kubt6z3eIRTg6nZmtj+tZ
uXnaGj3djCdLhtlifWykZjinba/QyIwyKys5IAJXh+1GwT5BKQrVZAEwqMGVdROC
adcHiPuQ+XaF3pDOZsW8K2h97B9VdyxpgZIRbnv049vCvwYU2/wXKDcbY4ULNdsC
DOTMDhXCUQEEwkjbNC9ecj4AXZ5a/llF0+ChUAIRw/IdlW7NmmZW99sb1iUl33EH
efBlMC1Dl0bxPuxQDKA06vWWZ/fOor+/KjkfP+Urn+6ag1EWWH3wZ13ONT1RlotE
aqqIvbiz7SdJdynp8WsKclNA4SJ4/0xaPS7GCDnNn+PeH34Jj7XAiflExQN2co3J
ooVM3Y0PPJzmIyDy07zlgzgaOI/7A+lh0+93Ke2dOGcgLOtqSaEMVhr95EX0F1Ei
jMvP9oZueRiiCjZ/qEchFGNRCsT33cuWDTaVBxxwmw/922SmKCQelOWUbzwXnMyX
Kh0tf/IFd6MixhqGWyaXDZAnLpOJfT7nz4YfIKD4ToCE6Z1BJu1E2rQqeSdvL/uc
DMlevYVhxE781bl5KD5z4U1ZJW0Whd7X8OZ9Z+iWcuPVvUwxZ56DjUgfMj6HUak6
xblsBRvYTDtfNi0lRVqq6lrn1sJboqxH7/+zwvtAXW9sPhU2WEldXfVUF6Pd0HFh
XrLdGYlb2trnfCpCFkmRlx6xOX8IvKcJ2jQChu5tBM+dhA9X3Cvg1sm8fFZdAEH5
Wq9bCdMqjO42g2RPdEok3CkmgEJsTzfVf++QTirQ92CJQvbCFkJqXBXlJ501eOva
5kV6mi1GIMfGUZ3OXBi+OnqE/S4XNqu/A4q/7B6Kd/ffR92A8O+0aRVpMctlk1P8
0RdMLkJDG08sicNDQJhjm3ZT5Fp7j54DWe3delH2KT3ynaI8YOaL4Fup4rPcQdf4
rQ8Z1Ov8vOXdL32kLLvYmBai2/KPMDpaxvgJjf6uBySawc6L7KvclonEzfGd80io
kJA6pAiGApDItdJrPPG25u+ak6N5rekXkRyxkGhrBmyqF7jfnxbVW9zN+W/ZprCZ
X2/IyB4EQTsx3tzf2/Ss89w3Q/LS1CwKbrOoRDKIrPeKmJZsGpZK8oHRiryI5oMd
1ShhOiLnx1llBGOr89oX5ozwoBwDmwhWllKiK36SXQYkQeahOrZrw+GVWWYUzUFm
NUeABkFBZZZUQS7/PskATtVQHXKZBFT8+GLZDEh14WqOhSFEmundBjZAVpBwc01n
m4Y5IemnbvLG7l/UoSfcwJ+2vq9z7qIm36qjX3eT+ktLQf8mzddeYXRQarN3OaMS
b2imvoD4pJTHSd07XZvI1d6u5fT9wnIBAN0qXRi1aEMwieIkDd7stHTkLMmMLHpl
LRQWbDrtAo0jJkpwHYqMbL1woMxgs+IQ4b+MDS5+12gUjIs3UheKrPMARPqjyOrc
yYaAq7aJxSIxzq50xG7ykakIjfOyi1qeXmTA9bbRQXLb0UZzS995UZXLc2ubChLB
Xd93G6avyRGA9Oe9wzLhWku7MWja4biCbF7+6LkMevgDku5KDcVgMY2O8afQf/rO
Ohz3n2R2IH0TUxP3rA3kpEhewIisdi1ZEe2wSjHMh/rFrVDgdChO0dKPACgv8H6q
v9ieVksNv3dOceiwEqUKcMedwbO1FgipU7j6IhkCPlA/7l9E5UO2G8Pjf7qqsfCb
M9g4I25XIsVFmr7nHPEch7hWqejWZKT6hn0dekLucT/XBl+PWMocxIWc5d/k2XyZ
gEGB2cEyGga9IN6pehNAIaMOm8HBJE0gnRpODUN0uaviiTfLqkwcmPcM4Wu/Bw+X
gMYW2Y8QHls8qSoIoUFAcTHpanMoHL4r4XdhUkjalL6wYIl+5YZBuIE1CA8Jz1XA
A6jqjvGf9fzWUTjVUzm3ftx6UPjzDESw1IIT2dsX51hFbipbnGKNQV2msdyndWJs
1PfA/2qMp/IOuyWc2wzi3peGdYm2/7Rhg6RtMeJUoCGSJvjXzQKup9hDQDBRvE2Q
2zGdCNjQg+7ZVzSkNGvN4rcN+eYCLmyAx3W9FfljRBc7Oqg18KOBE1htP4Hy0GuL
Cty4ek36A08yHoKJ+YRQePj+pFIw21g+Aisq/leyxzjEZ6yatJ4bjh0eR3g67wAj
gSphx8/33QHQl0jXVzWWpsRfqwMB38VKsrTpY/bKxW/zvmTgXCsmh12qyS/IkRhp
Y/KaPywFnZUE5RqirSbdjM4jeUkGYWZ9FehETrKU41HwCW3GN1HLY4D1P+MmD8c0
7+/FwRI292VY/duvakRhenBia9WsFaSCIW7yYTCyl02M2+VGGFmcj/T2OGdhNX0H
r+DyQJA+J29/l6Hji17Mu3CPETP94MOuccVP6NLL7tO2EDDCOdtZUUQQs2YnT2T7
9INfXEYGIJiEZoe97JVA8qWkVadl1pb5aqy2YdNIdj1wDwfOoEqA78CNL/uMKh5t
kboi33tPeymfAfVJyadx07r/y5zEoO8oCUtIuCjwofR7hyH4t/TWQQL9lY7XIXt/
bOHAzZOGYE+TdpN9KPd03fgJOd48fojaYXjqSgtafTjxDXhePow0d4vz6GVz9Wr2
txTvu8AuWT63n1VA6/clkNgCyJ+4eU6CTpgShT3W50WUCafHHaEpfAqAyuSCiipX
uUZj0hiR1rKC93Yvrvf/sVbMVGcjlVsJFk8LUWArplYOsFxG+CLs/GBGJ4yS09wg
wnbJydNeJgGJO8N5/TD54b8WaXkSrhAgXtz3ZGXztwtc6rAKQx7oJpVeno5fWTty
AnqCjJ7oZUIk9qt1OrJVBCaq3Tz6Evj5ZudpBDOx2NO6uImr5yoVXmDKSX/MOt6C
vbEsm0P2tlg+U6enNJqRwu/WrqfxJEJir0O10KZlXzw9DrZb1r/WpMvLxe44yS4A
gwqjObkj2zpvC5V/HAiMRo+cgq9EuO7XTqIFe1OKA8jkalWex52OT8BvALeYivDm
su/fDu6xvMdpUgCxiDg3zKc32noGGTpaNQtnbi1BiOtPBEfFpKoGIvxcgLW/ybjN
75GU5zXxQ30UIn1vk8wt5Cwlr0BJ9AGhaJd9yG49R1sT37TbeoexjGEQSiYOB1OM
4Ny5yeiI17OdkbCbg0OcqOHEB4wwQ/E6g20F4bEiu5r6wGj6wAJ78XuQOEWhcKw7
o7G1/rqgOdpqykxyyHeDGe3729sO9nmoS+p37HjmNzZ4PZG6eGtEW9NP/VK6zyO8
889IOp0aaH4QOE8txxzLwN34McHS29Rda9xNeVjwE8fyPh0bx3pL15nP3jwe4jmK
n6X/P8U4JGL1QH2NNvTBurUv9hLyoKOvWSiRSRm7Yxc7jz/FIVyLt20Yai8IZS4K
xYRw3edYm21Mpu3miAFkCkKuafEvMR4xq3zdAMuLBVWEkm8+86ZmXhnOwhG9lODG
Y/XDLri4N/twZgpLGDHCabIIdmUjzypR0U8ARUyiDR5PJgZsTserqk+SFvMYQ/8J
nzmzqveu7qg1GuKxzDe58mBwNKSfTZIPP9HSjzDUyDwvs9l6gLxU7iSL5p/SWLpb
lfRoCzoOp7fuSnzc/h3loD+pTISkXxE+GC6iQXbkpcEWPwjjuHF2RRT8MYZJ2q8R
D0uOLj1TnbdtI/9cnzW75gmODKzYalB+NXvH9PX/+RZp3GRVjBIPC/JI1nyb0ZXE
FYa5VE3zfdAHQ3TICuwKub2ogcVmeAXGy2+btUVkzV9xpnVwC2luaWIw6T3cBAUA
aum5veggD9jVGJvDlVf++gJLkFe+itDZZ3HikHjIkoKP6a258+K2OVpowpFpluss
X0m8MvJN8e6BYff5YQc3N/7QlUOCcrwecvyG+OD0YLRPY3KY9jgmZvBXkhq0u9Wo
et0LhUXzo0VUMknNwZtv1rCXgOAiD9pYTpoJ86eezFCe3L2Ad0dwQDh0YORIsrqi
BdangIjOcjkHQ+IoBlF8TSK8F22kc0140QWqvz4rZZi8jBTcSK2+Zu0y7XHP1NAE
3p3gk+gKQMlOJUoLDhKwPPmfSg5rT+3DFBi+3F7daH5+WiyUNmJN2a/Lq7/cmAiG
4EwwbEQJJeZWom5YVPMBKSochicQLPttu54XxB3bCXv3Ix7Oqjs0vhZJhinFcagQ
s6JeINZVEP6BceifoUKu0eFMUbv84V14LUqu3f+O4K/qrUJgzWc3Hp8HF3LZXNlb
z036/mgceqMFJD4Dgat00qoczQLcfF09HB2IU6aqMbrSOsEcBJFYX7HV02dmcbTJ
K1tVdf9nEQ2yDw/t3H5sovFbNq+u2Ll3u9c2gXxbRNe38CBKQN2uaaKxWLayJ2SD
gYlvo0S+2JFMBYfH3nXUy6ehXD7VI51Lgm50OlZ1hZqzjHafhqj3HwBzcJ7Bdw+T
pEgbZ70KvYPTquwhiFzwnrBdLwhPZEZ8axaHvf8w9ZOe+mx/IPwR5M27AwmUgwzj
YsO4lo/+d+cJbKNYwN0FwQxWFpdtXTvqP/WraNzUey0w8gQTbjKMZhldJTa7YHV5
2FFCVseaSWK1J9dxyObCNBUBt/yPhrU9TBtN2e6kJ4AB9Fk76eYye8SA1DL8mgfo
Dv8nV1nsZMjOsfAQWa483WkfgwjD4EbZ2OYkC0URq83eQuL4bWRTS/tRTiABhdKU
2br7eQ2T2z9mu12cOajQGgNIn9SXYzL/6F1ZjdspK9DHrhgtwm6Xgvc/r2Onz5Ys
lWumtq0kLjVlhEcEeSZYvHIrXH0am56vWzjYZYi0d3YKcaEDCKVrAm56I5ww2oru
wZUn2P4dS6cC74BpUK6tDfvE4gk+LAkeBu9jG5NclI9D96sLBzGR5RdLqiVDjIgi
FZKQWtHsT/PtNCKR7J2w4CxLvd0XDuuo8Cz30xYjl+PqfIVUPSkxhP8v1Kx3SX3I
fEA0mshzN+opt5vLoCD8sbOVmrHV86a4RilLJbXYA/tn0u+5BnqOU1fphnEjW00u
zsz73XVB9F6af12i7W3I7PuEX3e7L6DGDljErh2RLoBkPBmYiRC0KlJZZ8C+B/or
htEFRe9dxxjsdPxWFYlf62BWg/2R0Ue0WP7wJSc66vwWVv2CucPCBBP8rg/E6S31
guZVZ9v7rtmne8u64n63WQOkIt306TRdNO9/QfrhY+0EhmA+KmIY6HVIelA3Y1Ai
ubbBUDlOsQprRs5WRJdiXxFDISoC16guqL1sMAQ3ztCuDRVwlfKnrWBNr5Va5kYi
wJJlKXwIY65KUJwskYs2C0y1JCnAO1jiFEMkExNAbBNc0qTQt8/g3gy6M1IU9KFc
aP/tbWkewxSKchestZblxBq7Do9tQOcoEwH76Yqrurm42D5XGMquSFi/4fzgtFC6
olzyn0VbXXx+65ZwhDy5Y046efDSyM+LYTOexJqIdBwWV6yT2cIq9FqsfScf+SdE
d7kN4z1O+YdtP5qfMAsxtsEb08Hog/i/ujrcbzkwflgsK+pC0+aerimq4Yz+YHDO
/lwDpbchfzgy2d/u2BGiLKL8bMqkPIvXUhvcbBJtPwDYd/1oauRnRT1QDycf4l0p
SrU+OVIPxtt+3ZP5td/b0ZH/2LoL+pCeBWvYmozy7m9lEuFZcOgrAFN10Ndydbcn
ObLB3kBxHIhOuuQ5jOSCoUHOEAZMqdyvP71dPBrym6T3myRHuCiBzPlIWrtweNKp
LKo9S8/antNd1p0cRdX9VXTQ08+5Yl+cKhmGXWnxAYlMxgIczay9FCE8tNlZOgQm
4h6Q9i4TWyUlIicrfTOl5DIqQ2NpiSKz96lfJppdk9etFzR6AV9D7uUSuPZjbd4F
BhnPlQ180emqIbJVdG5s1EcNCfYdMFmytzrVcbJp4jQH0r8w0ueAMQkxixefT+Iv
lGY0rJFxUyrCoz8JAJpwqRHYgypAGKtiNze86Yf7R4BC4c7GP7wv4WVaDODetzRp
/KKIMRLo5FKwtvdFHQ6H5MpeqsNaxZHOxwspEOtx7qpSrh48DU+7DbuUdc2yhPsd
M0ZQSrsu/IWsulVt0ULxHUjD4EOw+ZaVz4Imd1B1XaShjby6DBa7L8s5tqtDLiYl
K+6zPtdVJ+Hx8WQ7NrvFLzY3W0hE8W2cL06wdrMgnCHEFcrEcNYn9e7B3SODwBS2
VFr9dfRS0MFBlygvLLiY2dM2CYUtaFEloWi4gtMO3vRDJpvGxmvsvEWqOqqGgQ5T
Cnp8w+vcO7Fm2uiJkXscC3j1J4FlsJ6wA2iPoe3GkZG+AYMqsPwcRsMWjkiGtfIu
uDa/Xrcc666eXTl6K97cxZqdthHPQYsC1H2Dz2DUcgfOxviy/2AzKhO/p6uYMAuI
Yx2+23cd+IgcmAC1iVx6hhRIr1nynl9RQY2JcriHkdqkZCgNOIXMTSzDzplYeHzu
j5l+rAMgoxROJJqQU+ntrgaRf1ls85uwSJUBdru/3OE29M/XXKrjukBB1ThKl57X
kWXxMYOP0HXSHQn8OnDwvtjFZA5zinlwUydho4WKGurvcN96NMWImnW/oXW25Gov
djnP6uEDjauDnivMau8QXckwKxK/XkPmBeIejmQHwFKz98ReNe9cCCVBBVHAK/+v
v0J9HqT51KBzxA9cfyXhOgg8Cg5zq0Nz2lNDyVbHS6QbMzLKqd9B3yRa/O8qAHM6
GKGfjBF8iko2aeqSZ3d5r0W2ABLUvCMi6MUpQWVImW5CGwJMEqXQWL3y1mD5AXTj
jmV0E2hcZ2paTwqQIJ7VjEZUWCnja5o61QXct9D873V+29x9IbBw95KD4uDn/cl+
nMdnZXqSl7D9ZE4iX4Ider2/STJTBXYFCL/ZfYxh5wWKdO2KE6DjwxeKIHqtqVvp
fpYagVCHS50u+2f/dn39f2nJNW4q3xqg+XT7cfMu0kKYEU51Vb1YrR/cSLPzeHjX
oDIEvWijXrJGSk5TOuxVLHRmMQInkDmzVvAJKEVLBhDOtW9ua0ZMwI3melrzaPX1
7hZegfDZyfT/U/Tm3KJX7k9Lo2+OuHb8uppKDNAR139neJYLN/l7PWuFGjFG2zuT
ts4mkuk/1PW/tafvcLYBFno/G0CHn01YYh7E1la8rpgyX5vu36Gs9KcN+VE0qSat
5rEX4WFHssDw7TMaTw7TGeIC02LAmPSbYHJyDhcYVhfBKtWXRC3O5FZVMRsaEETH
ovwrrGv+hioZXAQzfV9uvvW47WPPJaWcQ4g5g8kQgrs1aOVLNhOYhJGg+X/I2pY6
MYLtPnmhaGleicpt+Ojl5Kk3zmNvL0mBC9Nu+Lg70ckxSJQwLS/3Swf2OscNj5h3
3HO80HamUjhfaOddetz8g2C62ancyJSSIk1zOBljlKuP8D34C8wZt9v48k6sxgE5
v9EBomnk9+VQ0iWZxsYwmEXQ/r9ytzI7wM9WUVoVWEHEw4/Go7O1PxRJf9q8uvvT
Zv3vWd6Xo5zo7nbRjEK/G5mEESz0bS4MFr1Vm2YL1g3Fclk6KAM4xY1/XwB2I+WJ
QlmUZnVUgvGfnj/hOYeOmSC+BddZlZy5PjqJzineTGMKX/vnDbFvXi3CuEX5E217
98iKx4wKPb5J61IdkD9UVaBtlFnKEwSIAyVevMmBTDvnWFGgcalpUgM+Tp8bmmPI
+zdbcpwAcbQXwHgcIKPi3x48Z569xsI/gNBC3pXjdCcyRr/+RN2thwJXlCIw4cjg
VD5wRojuzkcQE2nPfBIXyszO/zjwtTU1KyBbqHRn0rJQ9V44Yct8O+R8Ism0oqZ2
m/PEIzJfgVUe70/X4mgAQO9rKfLRGMk2fChN26xU98PTjrwZo37offKl4mN3Br1d
dj/lDm3KVqoC4ZXVndgIHODD5MP1MxMlwKY4MInTJ0r58fpM1X5ref8eZHalYU4Y
sVH0CnSVL6ejOEvNpJMeXEBncHiklRZFRKXADvUlbRnzJS1VvRxHtIE7qcm/RTXv
kBgvAf+xdo3/9La8N3GTk0EEnWX+zCVe8eZT5sEnmGl3cGBt4rFQaPzf+HV9mDMM
E/gVUDVaMjfUr++94yX1CAay4AVYGTUa93SLTbiIN8vZ1Q1ScEau+iTWvyyQVtRJ
HkDEhaaH5kf6ZCKxrdM+Pituf9hyDpliEtEEs4Zwf28Pzm5ghRdH3YRa3Cps5Mii
1CMo2ZueH11g2gIqhfAPy6Yw0iqqG6wYZ6hU2h+CLq9k6xB5Y06rLWFgMathh3Jc
vXSTILg+H91NztskAbN0vnBI8r3/o4DqYBX31D/p308Mr54822lhKPRuLKqZ/X68
AmUcosACxWEg7u7KbhTL0K46xqNMBDS2CryCPOVwEh7KgJvZo3dwlGrPkaWARW7z
K2aEPShZhdxJMqa5GHixIdcjnpMgdgiJk31kKdmHGhxKb2nW4ULQEccl4G6ZR3O3
5omsv1FKGTLWxjYsFDHY+IHlvrQYWahaxAqAoNJMUc57ly97Fu8LaCufWZAeka4x
JHqQb5M/4dDKrK5/M0gRDnMstlChhXg+5D+BCfOfVTAKgWrVw4Ow5D5dv3m2Mopn
V9LPuGr1UQfm3+MzND22g9zWVOCmN1ML+hc6g2l3f3Mv/7hBm7Ml2GnJOYrkR7WT
mReLIcO3muSqzu99bptCAoqmYSdcmrWnyRnwMY76vyQBZDYMckuMA08MZgsEiLOK
8B75kaVYbm49WmLm3NjcYY1h6JHUlVBpqg1dRIEAvXH1/xZxFI5hHjY1oF0+Fk4E
tcu3it8iyMXGE35yHY8KPMLT5rjFOa2tNS3iGYpDnOkRNuoPNJ0Xvk/gAh+8qSlB
yEOofqu6OiiRq14+5qlpRtbdR7Xgutyl9LfUcMizp7TjIbYXCeSVfcj/jXlYEIqO
7sJODT3f8j+iPIOVl2Okld/VRpmDlB+QcvfUq87vo5IAcFZtfHbx1FOo8YL9L8+l
bR24dSYlWwHThmtaVe2Mgbha79BkbwrWdU0kfElS4+ZpXd72MkHxn0Zro4QlIzf6
j7cI6y6ep21K3Y9vg2YVPJWgkbt+PnxX+UyZqIZomf/j+xEsCtnSZ8YBsICYEXw8
cjk8feRgy+3sb0vHlCbmHollAxFclg/dhuMaO6QIH5hV9bWhobPe1ufxNphjajDY
iCjSjW4JVPI7qNK02anRboZN17ywjzqGmegrcTv6p6I4vTopr51ZOlw4BvlIXMpO
1Y0awSnqDE5Jd3KgJrA95+PNa90PkfTvOPCSdVg39Mkm0YkaHyXfmN/DxeuOuuSM
zg63VuIvgKgh8DG/e3Kkd8nmks9RYE8cTY18/IFPplN8tu8rYUHV92XO0ddF5ERG
DnHym5PItFlhK7dDSnzQvNs7U/CrIDkjNrNiCwmReXNCZ3PtqZjTmJiu2Fo4XuYE
qFFLZA+oI+MYMnZYP7c80iEzbG++rq9WdEMIp1zqtN52Gt4asf6WDVzRRW7nEc46
9B/y0/+QxrTruyQvL1Wpumw05JRUDBJ58w7nSS2Y7+LLMpxUsIL2RbEm9dhbaDDD
GOjAGEbuRlsPmkQ+K+ihnzQkIrcxX3r0MkCFEsSp8xvDTrlSx4WcF6Q4/N7nze7a
EzpiChzrsUwdLpYscHKIyJmVv66/7E5j+lov8aY4iHJg4HKtnkwK2kQpPEvlxod8
UBCP1fABa5EEC0wcBmOPkjq2hW6lbZasYJeuv+vZfwyDSxJLOtRnkqnP7SQ4SFI4
ajwDeDgNYNmEkZz/GQLeSvfgOsYumBYhZS/Y9Wb/WUA87oB5b0fHShEubTxnViv+
tU/qN2KyUUXTdpVm5ZtLt7Bj1/T6Lxx8UB52zO67bqh3NN2guEujysF6vgpVlE3s
OYe+//BiVgMVnGTrJbXECNNQLmy5t0sM+oykVJqAm8fT1lNM9pysY0HEQlNxNtoN
L7qsx3vx91byhWZDVkynVVxduylJFsX0WEvt1NO+d0MkSgT2Oa6FjGcQ8RvTSauX
DiGUflvLMJ5eYga0euLDy0uheTrPPlZq31yyidUnqgbZP8SaVPpPMHlAmvqF9yq2
tohQj/95yT930fRHSU8zXIHjzmpvIXbIyN+nqGrn/dI37OKtj3pCIdUiIFEenwaQ
ItGiWyRBRYVW+Aku2uCKN8unap1PIoI7yIxRiZJq1Flm5RcWZTUTA6LGxVpS9PQX
jQ7iwut8nFX2lvAi3qwsxdGlcix4liSfv8pLe439ZrQBQLRkqP6qdqlIF7smsPTS
5FEiT/bXJeq3ehhdc+gcID8FUweKIXEKw95dJYczFUSn8i6HHOwAmk5XRZMkrqc1
Rtycz5rgJMwydPtv3k0gQ49CyA3NflN1hn6+xPRt23+WsQ7nnoWZZg/3RZj1AYLu
LjEFjY/+hyM1sn9Xc97HbhaBNOC9cveu2QPuNTYJ6tKN/Uxi72FyO2zUq9ishixr
4l1wVbJLJ/QpJHE2bGKpTey61nRb+dIgixPaA0eIDNPyh/ydIDMyr+7p+nTpkbA2
3TeNdWm/IDn02Hyp//nb+z9CEwogkHNAg8pJhTZOyxvH9bJtn8xjVjCbxAIMGR4j
bWhSJdFPEvVk8kLUpT0+bc/eK8LJHNUrdmWimuzLu9dnGWculj8o7kw5m6Cq1bkD
7GGd+7TZGrzBNWzgVR45s8ZMNcxaOheFyfWNUkfmHfJc+bE2xzHajKGuSVoBhqmm
PAiEvWZf4nMVfd1MGK2C4IC/U+vCJ8MsNR9FIGVj32iPEXI00GE4eHNK6m237nOq
WLxx2fVMc8UjGBZV4O4O3g/OTql05kouWLogDiq6A43XwJKbm6Khb+cf6PiZW/SS
P+38fwnVExxEKDEj6TrNMJ6P8Xkj1I0D8t5EP+e/pbREJkIqufGA0cLZ8GyKUkhJ
Hs4QfvjRoRJYMiAnYdJVYr0svivv9x9QHhvP+iixdO6hG9lGqEIFq0mOZ0A+DohI
a0cdhJkdWEpx6xRghPZy0QX1VIr71W/EJKBUiTwBPcItFm1zWUdnVQSvLAPA8Ptb
IKSS//rfJ/JAcwTCSlXzxmcj1l2A8b/v1mvs5fvuv5UcvfCZillzJwIrgHtx1CD5
bWY9CYgTl65DyjiwaUq5WqQWmSUrruS2KBw6lE+WVdEsJ1v/0bvk3JwCPwtdeqBt
ibXXcBIpkknDgmW1furd7uwUzfLYHf4pnOVakLx47BK/de/ngt/pYAWdAqiKgrvz
oJH1CPvcUcTuzfk9ulg7xSBGPdMjS/3bgeZFb8PAs/XDTVvHXb+4pWIyKug6Dbms
X92cC+l8yPVlmBhRcK4sCb6dzqhbpIwC5rid4BG7vTr0DdC3ZcUKR9iKJRSjQDSJ
nt7QSjJIOuTpUuKb8xbtf1b97rZtXKOvhNkTHYWU0gWVWkgOrW3dLYgr1vhUppgk
MdgAAE+Foz6eIKwZCJ0epGNbRf64lHvm2cjk1DonvUixWKPupmg3wopzh2F257nL
6G3uCzpBOGHpPiev6Ru0T3eAWXGX4rfS3H4sRqrsz3cibjVv9g+tVdedM+9+ipmo
Hx8yWMGJT6txR9BTWvZ3z9Ubz1+jJ88QhTCLND0EG89SrIIj8H5BaC2r4IZpas+P
mbF7cI7DuZKPGTWB43tLoNOKyDVmYUKjXQi+FqkXdH/oonPeX4M60sODqJoBDIZh
jVFyzAwcYEWCrJhTj+lkmhapnMf5xQifjn6SCdROJdA9v1eY7Tyy8RQDhBreC8MM
QSOSexczx4Z6qiwqvFtrLqBsnN4M0RT5tiTRzQ3tvoB08I6L2EB8VrKy8uYjqqzt
VLKv3clBGzLGdd36e9/Dqk+81jK6hQ5CntXJ/FQEcrXFvfbAvtbe1L9iQj0kRtKZ
1g+lUdrrZ9Ad1s9X9uePCXZSa5CRtM7s9FYTx819675SpkAirgvVIHUilMvgqRxU
BSXawuQBo6jur8wiS8KYgX9Eb2O7Dwf8aB+QZPz9nzGUxW0IoP5/dg6o9U6TCuul
GFnIUeUpvt5BOXEo0zJhcZoDmQWacguIsy8dOPzcJBvZLd7Tu0e8DwJ5y3nNCrZb
+6rcflUsDrtyc+dsgJNI82TsAdvcbhyHm7Yi2SEdynHcpeQSS94xw2t69GVFMh5G
ra5EIAc2x0CksxeqB2bNal9l4qc/pHTznppAua3qk523Cbp/A+8eJeXMfeYR7ET6
ZBqBMxFr7DLRIpBOTEL4PJjtkoWT0x1j47Q5Hz8Y8+R4FDqlgZ+DwZKKcZ2ytMt8
xjnumdWvymKBDS9iFmZMvEyjkflY2CucH5AbvqcblmoQMnHB3yFichN87CJKMPfr
7b+BBFX2S9WYKs0OuX59QUd+v6ggtGGcj+rh7c/0xmWCQqt9YESKYQI3aXE5hRaV
r/8iFNluCkjhrsjt9RZQBsr0HgtgDJXrHNtHRLOe0NQMlySXvEPYZWO2uINPlbf7
yFIPz7tJc3OfP0I9EutxierrJukG86z9viiYUlpQl++fdK4vbWc65h1uFU3+iy9S
0BIzn6AOLXBt0hM34haaceEiG/GFWqb1RMoeh8BN2Vv0Jzv+shKY7bhaSjMpHz3Z
EaGDri27UBcdy6bCViy2Ghlk2DkzE5Wrua9lkrkdszqHh9TR4gt+yxlL82pW6zlw
AQnXkrhxAQGzkof7mQqrGr9SDA4ps2c1KViBTGnuBEjVQjFl3f+Mh1USaSHbszGy
rOoo44pr6NVEJvsvM2SdJqFlEKkn13GOZNhNpElzuox1LW3eta3w74tZ5bPJ/Iz6
/8+7UuTKfLeeB0toKz5fQnqjeVTOBxOd3+eR2Ndvb2RlFd0r0sU/7EkhA/TIS8AQ
w9mCc7TN+2VuQaWpT/o51blwgaWMDq0DM8NR78miLLd/NdpIcGzMK+m6RGNnOgTr
KvPOs9+aU8uTiAMnHCaW3DoWpBfdOg0XbLcIfLxt11s/pmfXTockM0vfBVMAYLFB
NV831hFWgKZdEG1mbKTbx0s9i6/0QUJMfdu17SyREx6h/nrorpkU979nrxUSoXLJ
HtAOw4RlXKg0Ac1DVVxc2SVVRqyV1EzrPli2Y5uueLMsPa33AQltWDLd1RjG+PHJ
xnvFEHta/rLOpD/ZIWRKAGpEtWqsasyA0O/+pGjJn7fg3Kz0kbJLxp8Ce2fIoYD8
2WEdW4SkSy1np6CrkOl2VwikUkpwJ/s0d+uQMGaaozaQ6lol7rBqyzXXAUNeW02D
0pb9+wp4qV7aMzkihpzXXHAKe7cMZKa0qiFHSy/Nr7SwP0dQPBMh8KKdjVy96NLP
qXufy+0Cf86Hdxc+ES617wnYT4u3GbF9dellxW4nhQ2C9jCUd4wv2YGMW13bXfAa
3DFW4bwkwbjHI+k2YgQIs0gdGcgQxs/cVj4N1DE5sRErjr/+eGNZ7Fi4mYIh5WGS
mc4PIeDcrSefg4S2uzF7ze1l2fek6H6hxdfb5GP3rRFZ1ZtHj6rqBamqXVFQMAVI
GWz4JEkBL4RoAa+cZLtPltidE8/GFDyP0gKd+yS/UOMkbLxs1I78Jbd3tabqnWUj
668UsaOpyXwn7txfdh+Foh95Hp36f9qOak1PshTgPQiPXrk+qfjLWmXcfAUtRVkf
kyfd5DyLoXBE1+1nns8TV3AQBqRqp8aOQnao8KY43O4hSrut/jZnPozJNalNz/xt
maWTUiH5x/k8jb+PYFRl6Wl2BpRaGvSvbHb4K3S5wC0P5KSHmEuK8sNrmrJWFV5w
aiQpZCyxqqvJcV+uLq09KgsfXPbq32tcGc7J4w4JotftOeQShLs5dVzUXICHKY5C
Psclxfu25XEccGBtpQ9nyfCcBtziuxn4g1LzpMWFURBQDcVJToA+oKmCsVEQZ1L2
ElIMXFHsivkd/zA9bqVcYq4g2mpYl9x4d1oqpYv6626HCdtM0C70I2p8WiHrFrMW
4hVaOyzhHHukFHlS8qv18ynR02cSv+cPayDmMgY2/muRK1LMJ4lp+W7KtbeC54Mw
3aAg2tRmelIZ2z7ijGTrKcquUNilHz4H9fy0wVAy9Zpt8wkaQ73kTaj/fRPCJpDC
RFxmrTsZhy1jrtEJpepOjUml9H2uNO/MjuAQdekbYM2Gzd6jUQQO8UhgMuLpqygi
NqZ+ZjtipeXa15YNcrTfe6AvOo5X7Yn1eLC/B/LeErDD5jafhgFIvNJDV8uj/+xX
JKKxjCVjEcZLR9eFmfqhzLDIVegkB7ZWptv29Ch0eImfmLS0w6z9X47UQWonTIHg
PE79sSZhzKFKxUSPmh3qOeKNs3FORLM+H6grk0jHNNtbMNFVFCzj1vHX0LdGxRKv
mHKUtWnkqB3K6/B5CNlb2r4HbC5mcu+qfkVxLutFAMtP0O7b/+wB2bNI14Cx8Xht
CLPlUfK3/PemBLh7WWiDXCEU8ssr1g6/4Sq5cvqAg5Fo/Dd4+x66tXWJa7R4PEax
2G3XP5dSXBHrQSgjs1KTm6UquIP+XetonFBusWIsWmxj6z7rDHveddQKxoflStX5
/R8Gja+3LvG5jug6L8IRMAKjqlRzKH/+DYvf7gm13zcTzY2NQxPZYKcplneuF83K
KK+ijXnJWvhqlrqWpU52Ry23ie6JsAsoChfazkurLw9vJ/SFppfnT228sA9JKuXq
0aZ0tAwW/Vfcl5yNXI4R5JhW6neM9a/pFTZ7BGY2Ael+N+5Ruk02E41f7BgdNiDc
qNTgc78WgeH2fBzt7jkdEd7kuWp/fny4OG3ZDKsIK3puDpy08KY88bvh09qKh/Hc
W27c9AvklAxxovbHcgmSMnMK0e+2SglQA3Juw2zRnZdhRm6RhvMInOvNfpt5rIcx
+38IJVmhLbsIHUBZWD5pQxSOEf1BTg3K2CcbflCK0P5zsY5LYqtfauERQ2/CCk6M
CfLwQOC6LXXRlr3iGaiGvkDa9XIRzUAUoIvXJU57/HtBymuY5VKvK16/Qm1RtYAM
AsQb29RKZpjVwWG8uxu6NCuhhvB6TFl+SljBgPOElFZdGtQTd8pBH8RfVuuMiWDb
txQaCu73alQuXCn5yTUKqoK2qnrXSDv5OIrsZFvNqNpJot7jQdWawgdywM2dqHx6
mnOr1I+C1dazRsyoOmpG3PB8RQapiREyBazblgsZ+APtJy25T6pCci/31qcl75c9
KBzTOgN1ed88TpRvMSxdwHHOEv3/3rIdH25uownB1VTAv0n1IsnrSLDNC5ZokMy6
fXKau43Rc+V5ItvkymQX/p4W3ASSZRDLT0d6k73LJahUUaeKGjzKiYfKPK4mcUPn
QJZWC5RLD5ECEB/ba9XOhnHe5mf2pkmFBiXKZE+nLZpxQ7Bl4vpOJBjLqBTbU4tI
81GEf5KkXThKS1ttnq8axHlFkI/bm0brpxOYrLefDPi6l3iIFL8TC1dNAa9j3TwK
uTryCfah4kO+Bd1qmpkRJVzr8dbPqWLEGqlwbJ0w0aog+y9Va7XA+bHj8wEZZ3De
um1ZLc71qCVPa1MusCNUvCdhStOlRAUyhZ3lNuiLUlWXju3UxJLaKwFhV34a11j0
HRFhgNZ4mJzlt8GBH2doX9gek+r5S0kVwGzsOO7FKGgYlSwrg3TEXPD8IwsevdmT
EfnF/V71I22mluUBFh6dcOoOOb1STXcp298SUb8Sc5TfOAMY0AkFPfmUHJqQDvG2
O+vdpD9rMYvB1Au6ZsYCGWYRxNBLErvdro+6wDJ+0Fq7LiJjLahsDvONnKj8S3PB
RxGuR82xVEkq5oCTXK8q6e6wAqtpUaYUD0oABt2YM0yukgJNGUit2FqP4yQSockc
1uacq40jhwCdjxJin9aLqqEVEiSB7W+OpNozg8Njc9qgZvbJHlH3Zyi1C1gAMpE7
/sNNnKqCDsS/G0i8LZRJMsAq3hluhZRVFkkzGX+vIdAoURMqrhGsJ5bIjY+pshyp
aIBeeGJsMYdqTQlnHhrZw8qlKYst7wcU12nUR2fRdijL9NDrHPKFZGaVBFzFTD9r
EHtIIRPclphimAbpDO5K6EWK12OIPYJTycPWtfXZ0smKzuBcxL2JH+gWCcvrPDwI
K8U64XXQKpl1gUkZXzAPTE3qeN+M0lHN0YvrEqwWp6lSvnNMS6XDf1N1LfJYbVm5
VSDAIG+99c2XDE1MASysPd1VyUu0TlKIeLQIpHx61cIAAD6LAVIfBYiB6E3PcbKS
DUWi7F/dfYlKxWUY1Np//ufbr6PIOPjh80N6FvRgOjgCq3ACkxj1OzKUA8xtPa5Y
KzJclgM4tWe35w/HWGTcmD+TSeBoyhTYwDTndRrxeM9cMpBaI+HlpEUMopIGwNo1
A5hDH0WAFaiWaWNaprLDQ2cFuxEYTKgFWZUCXYpa6PdKMTms3jb4nYBTQ+04Fy3A
nPstLqUoOmRc+CErxY1OfxGLTNHYjbhHRKgydKGEU6+UBkXGHZAIYnfI08UhTRyV
t9oF7Wp/ik0iZOdGytuz6P2plw6UpBqeLjhN+4v79CoP0THC6Eivhtcoerc7JHSA
ShZ9EDUscZibS/PfsnEcgs21J1wJUOq2HlMFBZBJdNmNLJeC3NVsKkNbS/dstB2T
N+bE7LA5oWmo0Miz8CE59fvBLRjmcUI5N2MtP/YoJHlzj394E4moHzofoEG5xICW
dTUyT/e1GJQZD6THznIv//MewUoq4XNWEvcnLNk0TEhmSrcAX4vD40xHu3x8AgsI
PzQxsUQ0/RR/+7yDImTtdHvov2mD5CQLZ5DzK8PF93myOTE8jzTnoNRm7oEzvotc
14VV5U+cTU9PxhCgZ+bhN0JM9S5d+1F3PItt/ABSGfwjQmVxhM2HUESgcRwe9QYI
7yMgx5FOReuxnRjqetsC/Otalc+j8buDhL2ZLP9CA8WZnMseP7Io+WCPS1oxKxhG
hlS2EBMpdtpjoJkEUmiUCC1m/XzoEPDXdalBFzoB4VBS1p5SVYmWPJ+eUpJc6R26
ggFbwJ9hUqq0khltFGHLjpeJUZ7te/hWESaifPQqKkZ6Bq/Xh2NnB3XY16jCaNS9
KxtKUIBZzoVdXfopE8qsG70YP9pjtgZ6/6zgKI1kWkTbfoxh8TsxFs1882efapMM
u5ryHXqHeF0hwxts2g7JjZabXXqGbl9GHpe+hWvEOwsXwbzizcuDwO/5XuPps4g2
IFJGgipVYhivJtOW8FJZjdlv7ETg4CUBrzZHwSjv6YExVgECx7xbCdiPG5yjjJuO
7krz85KRtJh/MTXrRNvcMtRNS0hpZPq2vVDVQxIkYswSoQuQdTf05gPaTSvmyMaV
UJpTdnb7Et+krO8luOfE3w1nDWiiLfsNsdCQtjFK1pJB0HqCbpsbv2WiWAO27msd
OvrTyY4JHF9N1v3BkwwX2CCZtpFCUSZ9RvnUeamjAux1Np/iHfMBfsT8XOhTWFYi
eZUp0jCYYnlLFlaZ5hO+gRcyB5UpXmOBLty5DaX8+IUgdYIWTt3VsIPD+u1chyWl
oq0X5k/0scw5aCzdadjofRzJ5WG3ypUTv//chZDKkTHgtYrrP+H5VSVG1d4l4lc9
sm0x4c5dK9mGyz6cgXrrN22ulZxGogGEJsDP/dPoXD8GNgyXYifFEEyECIzdvz0a
4aDbp2Egcp8098wumPGgB2oRGS5Afe8fceMrP5kZcH1nzRWJgQGUZ/moIf+7jSN+
SZHY6GjAhwj9gFlD3avMdpGPDSLhHh5kNSubD7AnS7TQE+9RiU+qTEd+LbGIncae
q43VWMWnasE6DkhSOyS+iuLcNXJ17A4mxbBd8JQgZfIeV6o1VEVLGkUu3r4eCjjN
yqrhVCmgGPWsxrjoVz80z8jOmyIcXhnTdvW5vroSJtbMQ7V7dpM8DRn2Ztqi6nyf
+XUtL2c92oYFQ08Sb/+sJtCcFfuwYspVzD1/oSXZqpAh7GooHUCXUa5z1gyQxn9J
S8h4FNlB/fyWBBMWyGkZogYyI0FC6INSl8jvPdE0yQXkX5JwyEYiI5ec+C56NYgM
xQnaBIgtKj6jnTZZf+1DnHMOUMhdgC4Yok6osrnr339G81p7Q9WuLVRlS5UEqCBl
gT8ZkzsapBeJPsv4/ZPVVbDvKo4shPOQz/zbehbsKaB0d9bwS2vmEY4YqFDAkuHT
b8D+4reE4th6VWJPbSL0pTVjV66m+5l29N+RjUabtSkuZNkQ5sXnvhof18Yu/wzD
JCZymX3uBcDsw21caHFxJoZmDpUXxKaPFlNc94fE5BtiPA7zzxsin4xsB9i3MLUg
tHxRX2fugA7x44XwQjk1XfhnYhKC4gR9cnwHb/eBjIKiBqNj7amyIHb7WZasI994
qP3D9UO53PFM3k4+FOpjGpPkFaJi6BpLkOO1LkIvqs0jtn3qOdy8d14aTUsnvq10
SNsdq8Lm1+gtISvBYP8m6gRToI8xIigyWmueJXizYO8ki/BdY+uZfxtmMagwgsnH
Rr2pQkXKBCkMOHLREEzk9rrBjhJjXwrpmH2qzlLHXxVfgsAyqKFNVBp+npTk0D2t
yR7IRICa+JIY60DJBlvtAkl0Szcn2pengbpGgXGO8Pyewif7sCLq1hWgl9gZuTiA
UR67BAE78JZXfJMOXuhX7wLQqh0veTfVO2xdPhG6gSk2cxLpaHWrbwjoFUckAlhW
SniZZl1PFCIoyWhPxoLylF10s3NqVNt7pSgNTBRhWIzD3B9d4+onHEYt4BIdLOHU
/bzU99ZxAhKiK+H6c0yjKx7rvMwwkyiDqJRVoYzOevEQ8mllx+IWFIR5G+HRFJHS
LQBhSU3suhKuahrWhwH1Ow6AF5/8U/r5xClaEADsba64Z5hLOJ80EKWN5DNAV/mF
TNNYrUDcn42/HEhhsdOYond5glwh3v/g8VCXlrwn9psHeWDCpK433Jm7uKEu/fuL
WT+iR4XrKqfljUhbFCuw5PTj/F6CWcgiC5W2gZoQ3H1KJ78KdcjQl6+BUmsoasLf
/Ukm7mrp3FgTC3atp6u6XDP1EIUqrac9vMOy718QNLynskaMlM3RNjv4KyogvdKR
eryUHVCvHpNBTRgGXcjeQY8YhFavOW0yBdXqkxqrp5Sfrog4R87dB48VI4T++H4w
Dn6wRgK7zCAGK8ASU5acgDEZuRRD5KxBo0BixwTDNdV+nvomts4CP0bBFnMxm85P
StAr8Wra3Aex4iq50obw8AyXyi5osSjUNjlXEaFobvO5pP5bAww9moMREnKvlcph
shrF8D2b1GlmcKLmpITSKZsuzKLm6XwQ8QvyVu2aLtPJHvLE3D6x051tUnS8YdvM
ZglV04r8SarQilrk5vTiBVzbEXOyTvy1KuKCAMSYXtSh4zlKwAPVwXrSb3Z8or4o
XkQ3tBf8fo0eTKsjWWemD2YhVEYPubGX3nBwA/AG4Lybg4cTc7Zng98VxW2m4yaB
6scT+YiWe3GQcbR112j4Vyt8Lsr2iwmXQs+VgKPauTO1bpfbC3YqeYxTRcgwXZvc
0ENKILEOClitMz5wWs8fTXxuL2I8ZxsIGQIX+rHyDPVnoN6vUE2QNPzy0Zor3LsY
z1c1e3Vc1AFB/XSjuIBifhZuEnWL5bC4OQNsw4efPxNEgBSR6Krxcs96FhSlU5L4
RvfeHm2IKBDcrk4fKD/zSaB03Q2XrihX/RmzlWXSZ5kYGj0j+KdmDS/linl7uHY5
ZTS2eXWhXDk7MQD/TkYs59ej4RT2Xyv2DGAh6rvlWJlY1V+EhldUjkr9MACgeqNF
vpPpPhfjf20qAlTdBhQ4KmTf4CwtqyAleIE436b02VThTs9a99pHr1MB/RRBPCMT
d74wPGGg4mxxSbwxrTNZr+9382kVrk7NASo47+DUpgw/OShHHrMgecM6V2LrKLF0
0FPfxURNpk8b/qRR/M3KmNZkKfEJt6qty7jgoFyMFC3oDFh9NGdFCnK+JjnAnb+P
BEk29+jYXuY1yAKhlKBmv50lOukfDOiLTBju+Z2o55fk3loqD7lVHzAJpYMLjtCo
wr7NnFc4jLS0Ychjy+5/jmXwwVOxOvfzld369xJBWe7twk8DtYAX5mE6uqZAhI6C
ptEhOhhERa7df9WyHL2JUvaTa728jWa/hsYoTI0vrDNJ1e1tJimBGs6Ty2QR6FO4
SZKTMyhREKKX9d2RlBWeMjfOpCZHLIrfIPIpN0XjFLvKG0PYjWEe7DbYJ/f/wx6/
3bxV+8e45cFv4g0Q1/zOm9KWLZCuA8qxzQNofBD5TJvPKYSog2KH2R1/gL5IGNG3
pFU5jl0sUvxQuteZHHIdLqZ3p77VSnwaqVg2PWmy7IaAm+siJ72gprKA3z4ryilW
Ke0begfw2iYTwAsZxkartDPU6KLK8yoqGb+v8ta01fvVprXvryykJFY4fPjroR2f
5e/mPusn7q4Fl78hYfhWDFPIXk7cGXB0Xn+35GCb+Bupm5m4NdWXstlow0ndsIzU
kxTq/j1zEDIc/N1NbDHYrP5jLhKN0r9m8k8rEzqLN1tSTXKOG6RVP3NjUMHF7vhL
OzH4hlNmr++aa6C7bt68JFARaQ1R+iKJY3N9ZThqeL7nQ4XvSyKtLEJeXUuSbp2K
r5NHwdSy2vdhR3xbU92ZjXh0qeoTEakD0Gz6qyEd3eN0JggCkg4ijp97L5I2VGih
F9EyT+jtO/ImCLJ5hGnvGo2HVgjA1brafFmV86/QBKfCS41VwLgRQfZGEi3woEaS
FLvsDpo8aShr3b6MqxX45sXB89B1mcTs9u7GY1N1DQr73P9GonHQqizvbNuJmYZW
J1bMZA+wE5zJ8My1004GwSMxq9FKMhXNNU6dLQr1d4jNGL+Rnm5iNG+HWngG0ypC
b0gZSzZ8HN192Yvz87C8I45VJiTJnTE8Vi/Oyh42SQDVkI+JJvxaE5ulWvrNNL/6
BxM6EOSDXHPz4DcDS6WkzQ4EeQLWLy8Rn1HZpbJzS3LzLcCC2OwuyBrHebFQ83F8
OsrZUkJNH/z4+K1thEtNszSAXvAQRiN6P8FT0Ct5C0cDXyvQ699JDlpNsU14Au2a
Cge2+X35BhbaX+raSPdcyMwAy9bi/sC71gT5mZAidemwiOBjdGrwt3qlDImpcHZb
FcBs79E7b9Be9cI/kqonx4c7YP8v4mO8vt2rOq/PWH2yjTOalbGV+++RUrc/s1sZ
RUrJhliwv7ot7fFunnay4EIibLDBbTYoEM/LWVdrmHYxMlL9B/C0VQtfjHv/RfSs
/h/CnbSV6I7zY7lJ/z/yOjbltLygFsVdH9/y7HuRuuSSEk1Lj99Mde1/ety3FqJI
XX42XMH8PIzviljSciXapv2rcKHoa0ILpaL7WjRKPUgPJ7+iPu5pR6CNnDGaXHc6
R5QitSqeuInKd2j0FtXePXMbUwRb95eHJOvEFZn3KAhonQLM9qvQvs0yMF11PdAF
6FBbbcsx1F13vKqbRE4AHXDUHvBzjB9obhebm4fMzxZYq0UexhyrelGuBwpAtoH4
8zQh/EIbn5oQCG5UPDt0CtgVemKlyt3NZq4mFqSbOd0j52D6qn0ypBfWfNgrN+3e
Gi4AuRnQ2Hk2kEqsxDOAkoV6O5RgKJs2XYqucpsy9crfaMxA63xRp+PbQeEI9zu2
gSLBurJqxk2I5MxF3jmBhIyaMqoW3ynzTWtY4yB2ck3fE/Rks/EYYoy4pa83zNF4
6QDPRk/yWIdeRyQxzDjLxTP6vh9v8dwEPv+k9z36muxJ6PCYRloNpu+1Wc1OWab/
ygMe9j5HYuqKzjPrYJt7j4EsJ7+qlxrnkFj/pLafcsFRXduA7Sn+aMKKrmmWIRU5
PITZiK0lxJ1ygi4HmvL2ZZYOw17P+2jq5pDSfVnra5bfTYpI27QVlVPoJ9lB2f9t
NVvuCwqRHIfOVmjfnX8+HK3o1e7M5y/xTG3Saam+xbop+UEuQ1apV5WH0qzfOS8W
vSd8HR7v74BUcifPyvzARPUu+n8pvxEmW5d1yx1KXdYu8inSmEhgkST2pDCbYnUV
GgcLYotuaHAfeN20hC3pVAZPUWZcBOn0IOZv+MQnI2oRyN8rpuIQu2uulyg5/iPe
hukhPvwtAGiEcBfCVP4A3V+ajaifqhATC07OTu0rVPCyRIEE4MRbZlcMnU+dfwjk
wsNS5B41khvijIqfo0LMa7vzk2WX4xqDsZ6mQzbSGhqnsXDWj6KK7XoGJrC+C/ZQ
Vr7Oaphqeqoi+FilfRG28p+DeCg4LGkzlGIs4PYkmtpEoEdFEALwGLUEyGfDHfhN
/SCF/nmCqxxTV2c3cSE+XReg2bN0vzJFlLGOlzGuMB0HU1Q/dv4Ge1KgrRVDU5vH
amHhrrH18s82EU9ACYhs+SKE4ypDj7AE/Xho5AWzTOgOKmQxkB0WljcxdZ8Ybwo6
8ziadVzUk4gcFr/O+4z2ZNDjlkPew0PbrBN6OPucvqeHZFtwpOrvNRjVU/QmwpN9
hOE+VZ55YRHtm8DcQFpqm79SV0S+AhqooMy0M1n3uaLuPjPP1viVPM4TSrhdJkyD
T0Ki4xzUOLjRPQNr6cQJ/UDnA7J7d05GL8NAbnZANACAVKUHPXPm4bb52uw+xGvj
F2+INigBXwYNiKTvasw46eiggJ/lLeqewixknvJKd820hkHJOFNzJeUV4z78MWo9
jOyX3y2JoEYZlo5E3NJI5d7vyOhB621snDtLPdhQkMhJozTPIfINXUALuUlXoIzw
usWLcuwYkl73fn6mnM6ad6npPEs4KKBhPZQbhdrXIqroupauUxHGp9HfBcRtllDi
AvnqOqEx5IMkZqM8hDHvPrJrv7y7N2kGa0hnuPHMFGkxz9M2pfP5BJTYkVazUegF
u8khxrXyJizkMs94l7oATmsCNoKQK8zg3/b8bGVsxuLR2uU9bJjcjJAxJtyBWn0S
pDJZRgy6wyBzMabYhRwPK2iN1pCjuI3a4qLV2pTjAISjInh+A6kNlatSrfN8PBKm
OaiDcwTxVw7Om7fwoJl9+TS4etZrcr2nD2eOjaoEUfHmKEklwcMLIg5GTqXwOipm
fnMDtPfisbVyeZELqH77Pj8Q3WYV/ZRvdPtkkia8+2kRUnDz01R6zqu5QVkWBAiW
q2kGUiYhTA0Tm140NdStlJhuUX25LE2lQq+DztIjxpkbFEk0eU1piGKgdtskoelt
Q4cPFjwEIMIlS4yxM6Ex7DDtA9j4ByJR4jdp82NNAfhtmfBNkUTV7E1Gty/7B8Cv
22vbQoTdhiB2wGFWrdR60x8qPSlVUs4pK7bzQ4yPZIqrzf87EEPxooTl/n1NIemo
d9XilKKAcPyuQ0PeHKNkCV559Bmpja2VEt4RVkON1/H2HABLf5jAAeak8Lnexim9
XGhJ2At3BgxYdPBNEwxyIR6i+WfZHGB4RRZ/k7RIXFzcirO3Fe/JaOeh6jAwynbA
xxt290LfGuJVUatXi55vmWdYUtJb3EFf7FC4lVmldkNjGBD1Ep8/j5WXPXvrsXog
lOiWkSxNyZVSCuBwccrZfoPGGT46C24F2uo8Iv2P8kBpVidbW8rCEYFwc4g3xu76
+bOrSD8OLH+iwL7Z70T4aMN6CL1V2DKxdt/XcZNR0CwObhifRF1AV148SNBTD/bV
en4q80H3f4H5uFd2YdUd7hK2aMdo5vwCtxULvUQxgCue+r76E3yQXi63xYTT10IC
PoqLUOHJOgGr7UERVEKjfGq1/8uXemWsTHO1eZCIZ3tdiuL9NP7ufa6WhJ2AiSzT
IGysIJTw2lfvlNuh9HcZ6WMtVT2+A8tGpXsGTASL09M6Br6InKT8g+yhvBEwC5dG
twAaTq6RFPE86hUcgn+UZNwCF7V6Kz4Ks5x8zCtH+NnHmSvBzGMiJ1cuhpcYzv5N
0Ht6I8YLC1qjL04gFA20n90+3K5EeScNyIatp49iI4TYIzFwW3RWaQnXaghOsJ0R
sD1BSo/wuVkso5iRaPMNuESlKdAxv7dvDRI9p6mc0W5ykRe25H+IXaI9pj08NqU5
YU594Cdf6+doKKKP9R24ShKMKGHC4fnAvKRUS7OZKf0CClLh23xl707+f29BccJ7
CMAZRIlTkgpyKCuNDZiKqcUF8Q5G9A1Dk2Td9pU3AhXUZh5R6xx9d2aAviG3YNIG
TBFv3xkj4QAbvzg4MpqrTgn4ag/JU5HX7Xzq8VgZpwRPJyx2H4mPjh9rqs0AUSLQ
GroYAxdOJEl73ScTr5Bj/wCfcHz+YTPFiMhzQNvwbaCkAUOJOVIO/9OHdnneh7Fq
AHPh5EATBasfRnYmfu3+/6IqOdFCnGDU11LXo0N00tyMTg99zgNxIvEAbk4c42ZW
Vhn8B66MO7TBQGy6ke5kEpdXJt0ZlOUuRLY1F5DUFW9y7UJsHJB/ULQ52Zn9Ab+w
Ug7Xlr4kkWgRkxUm2TFYDkkIx3+0vCM3iAArMSt6FRVB+bO4mK/jn9eve9Br6FXp
3JdNnE/A0P+AJe3k6o+tdrpHtVNizGNX9cVnRFuubYju91UqxvNdnXeJleSySoq3
XCBRdT0YlbV/d//07VOzYgRZah8qsKyZZaDbSoo7oi7zGwKmKu8hdlgbrAA63+FC
bcL2iJsfZJs4M20v7Vw/HbD1OqPLV/og3ZC+hwWLu7N1SM/yzmJv6lNjRN3vZyv6
hLDewxM8tl9B8+USr5hQwZq6ZQHE+M6FAN4FPqnbePSdwVwVLpEixdkIUZVI+zeI
FLTtpbzRLAfNnR6U7yirmnp45q1EDuID2nNHRemzs7ApRZJY4NfNuY07FCvRArzD
Xp8hIIR0r9r7nIcRD4MyGsQRxNJJzhAcomWHAuusLI0++8FYUcZgfO+n8o4DXa1r
JhtDx+KUnQkTmsPxpHhOZF4DnQ1mqTg3+xCefaK/BoQM8EMBugPP9ikP3q+nN1Xu
90Om1NeuWpUsbxs4bsfckbtNQvPjdGHUBoHEr3STs/c6bA1cYuiH8kZtJIvgOUKB
BNjEpQazVnHgCplUOli2jSQCrxAg/cgELdLc6+Wh3zNJyeqKvtt4rmYJEcNdb+8r
tC9OChzUfnnEn+bOnEKjhZVUwQkZVeIt33mStoghOYtqELYhEsLrRNGQcspA7O7u
hnIwkx60N/EUVYJdr2Hnda2SKIgarYxbeTOL7u3TZY51QIbtB0B9QAykA6lrcwAS
oSeTYu6rHwVPbiZfHRk11HtZ4rcDBQAcWg7rTdQhqayre2NE+YKUuNklInrweUu+
8vel41FTgqmNnpk4Rt8ijj82fzG0Dknl3T4Rv6aXBazdY9SC7WVgjYYcwXCHovyj
OFWYhPWqdylAcR4dOhAAWkfC40S0Dca4K7Cabnto4BA/gZlZ2bNpeFQzBYinO3lq
8s1G2t73OeLwHYbMiqUBHdCYj/ql3HImAHAG5kDkaNl237D0dkiA+ZbwmcW7DSq4
M7eQqixSwUuscrvJfN4tb4LsRTPXnKTLaMCfb+/z9/o7MIXpxQIeKZwwS0FJmPkf
AgpbaRufkKjYFp1sjBIgZKiTDAHjOzA3MlfwRX+m+2v4kHZBJ0j0poeZf5a0OOKK
DzfVYuHbVZ9P3HF7ZM0I7wuXrE605gZdEDTscQ6B6FE2bDwiDj58fs8ROx+1Hew8
8P43RB941DGhrvLjKsqEqbE59kFIfbfNMOg85TltVL4OSPkoIn81jDJ7mioIVqJa
932/WD/dqyBtFyGgQB/ZICN/Ix/IDm60XdklivBBKu968fOQXel7HjA81fPhK1uF
sgfm1xaeCGRfxTkwxmhy73BntoXJTNTwXe9N2woxU8auLAndwkwK/CEqTrcacrpZ
AU8M2bq50iOgztf5wxlDmQuof0AcbVemaFXhiizdhE+1BdQNdf0YHcvQvMDMI8Ig
a6T7zaZ+KRHuM2YPLZwcZfmmpPnV/hUrA7BUKYIET7GCwENksnFZU/cxYf/BlCG7
/2U7zR9urOCFtMgS0buidCgo3KpbsmyTy6ibxGbzumxCtmOR3jev7wLLYCiyqvZY
hqDgBVRCZeKMk5kcDS3wzuzWSa8IML4So5XXWKv9ZiqMGaNcwwE7I2Gr7H5xVVEG
sXDVs4jsZB3QmdVChZNAfzYFgLIgCSi1OmyvBXRZnpXoY6DslZ/Iz5Od758c9vHL
Y4yk8M9645beQzNKCghfuItpRAm3eZ96dUamcl+DuCyF9vf+3bXr1RMBZPTLTqGh
85ixeDApv1E3q1y2Ud6sssdLzB8QsDQR1+mWgnN5QIGMsUc7ySZV1s3s7Xtmaspi
aphpRnTLwq+Ct3IbISuvLqfnNdR5vWS6ZMADiIJSr/iGx83BaLiS14Xf0L/pFxKP
djOzEptnKvaEANv7lEO/lg9Li30cbAHHpPa3TJLSZRgL4yzay1Prkz/yqFQ4X4XM
XWvFoMEqpGw9540JJh6R182r+lTUf6rN/Mu0SJAqdh8BYJJ2aApK/AGF/RBuPWib
7c0GZvYW0ic3esCpEKaYstQpU8/gSyoCGq8eC+CX+QjsnAwcezwl9qX55z3JDWxJ
3e4SbpxFitipPeIcpB/TMALI5fF/j8rwN3AF4tnSTjuipMBOO0wU7ggPvQGM90p/
A3LdhRUvyL1zEf1vpdqcbY4qQiGRBroFHlFGjwXDB7JZZqzzPGtgxg3UlIQQLwyO
X/Xoa2zXjqkHJlLuf/R2Sw0C2RM4EBM2LOb8GZPQKDcXC/3QgbOY0b4uoBnNpNPF
liV8E7n/oo6CC/673cqAhIctNYoAXJ38CYxFcG2ZDS3s6YiYbwITdFteuVicMDJf
DiWZZMtme5XVkXO3eWcnRy4WQy9J8IQ2HQ0bEHqq/T50IdMb+PkeVQ1NZUOilIVP
NLI8BEVoAsrFIrPeokz/bSCMUGtHzs73aTgEHeBVp7Kal4fhxoAmteaxHrUv/A50
8rux6XLVfOnOkcUy5ZmldpSQvJDcLStXMEZx/o2K7D9ULLdCWyGzji/VsXUKe7aF
+d1sjGDWPUoCVt/kdGUYxorDNQra+GP34eGnPNKHmiMIuF8AKgdKazeU0/NBE6NJ
FJH0Eb//x20RmrDbD76ozR/vIayqUjvQRG2Ko+KMpO8izgScCXiQJDmg4r6BL2ZT
7CpsAhkGCmzEKD2yas5BHIuHCVtY/atFwXxtoArT2x9Y4ktM/ul5QoWfYVOPJo3S
hAsh/M1hRtHoTzR/EJYHQ8gEErx2JAgAJa50rX07WOrheqBJq24rsus93BJfMGGj
mSZInvieY4yMQsskQBCH6bfYlscRvoOnCr5tju+3/W6qNkCDTzbsi6ZMbNQqlGk/
qkggc8sjDh/HJjXrvGY/n4jglpI/fYw6BGJh3ayk8yu+XKnld9O9wCHCMGMg9huv
fS3blZtSqbxH5+VAds1MwNqRPr9fOOaUQRqK3WIZLNUFJFaxfks2mhqGXB9/Ztei
3yIXPoudyQXEbenbSzsT87bFWif+5CQyyqPzCVAc34fOHsR27KJTejsWB0kdDI/2
tZXMG9QFJ0hZ+hw9VNZSDwtdyeUL6vmDJh+CrNBfv7wvA6yg8APbBhcJTv3MB46S
u5VSDzCiDSIwoNo0T4LZSHp1DJwF/Og/SPCfRYexIT0p0q6ws/J2slBee+a+x2Fe
J96DeJONvhXvQKw/PVT2ACgnUqnH8kB99kya6uqNdZmNyQOj4i/PC6SUFMt9w3pU
HwIxZzzAO6JvvM/mWkZ4yUVho1hp4+0MjgHVzPEOiCRMqve0J2AnOd3PVZ7xVW++
lxeil/uwA46ChUXUg/G5GKgMSDhBFySsI5ZDDedgsk/3Ri+4bdMznleF/NSkxn37
MOs2y0Toy8WEK8M88E1e2vd0O8bmLiXQkxTypbLX1HSgIzBjDDRff9IJ3VS0onJb
d/lIrvXBdRzMog8x/W4oFkiUtxR6z/TUzrxJPzDzxDq9QK2/CsokxNRT97TekY1/
UhcnxluFcgCkOw1Wb8v33w9S4raPQHOSpkD9WmA2g9aYwrQz5EOuvi0DGwGKnI1x
V9g5QfcLHmAvZ600DMz3kA5GmbtwpLK7HEBahunuQROgXxsNXP7f9+k+NFysGdTH
sGj8obQXJTIX+tidTKS8rWc+dQSTorLSrIbZK5MAmIfEz+9bhkyk/4iccfBkhKER
ejfhAuMuTE01VsUeZXilhUkCdgpAeCeydqXeEtNz5yEUEt6vMITRtoSp1DjGSiq/
fdV9eZ/5fEipzYo4DOQm6+yKMyyd9sfF8r+RwskZeubPOFHOCC1EDKsFQKf19oBN
YF6MeFndcBK5bSV5dWN/IXPOdtVVYmFmdKjPvQeDToJPzmIpT71oq8O7fj3T0SYz
iwbRnkkIOUCJPNZvu21sIguNGAsrW1akbaoVQsIyEXLcJrQm11UeO4YYT5tqTjmY
UVQmDBBObkDapZbXShV3Yeho5TGUwF28n1azlgTEOKX9Ptu+cWQ6MFibeYWZJRYC
WCFSjCoUyta26N2tVbLq997ciCjR8crelSQIf3pMCNg9np5E55BveSO35qZHDFmf
5znBPbcoB0J7AzHJxGXOBvzPCyPxDrN+9mIbpFDpzsv6q6Vof2e0WUytgT1kj8v9
UsvQtYsFqpQOPoYlJadvf5i+Dn6qAgXGgD2tEAx5p2wBTHV73e2LPAZnP4bMCvgd
bZzr+Ia0khItgsYtaLVVmrEp0tNTrlpdcinv7/wq9JMgeKTw9SDFA/aVJ2XhR2lJ
vG0cgYw/+o4+Mv9OdOOgNbGFR1A7pC92NfwreCJJb10sskSwiWZRj0aE3m9kni+G
MGOhVl9JwDiLeDSeZm3Upue/lFsLTaXlNTAtPGviV40aLNgiZ3iuhQe4IKljAlCE
Wtxq/I85JMipCm22Zachjtz8UsVknhFvvDJ5/5/FhG2gX1eyky7R3NhjzTB8RPPv
caklMGkXIKsGGainBiiW6uKfcH3n9shcLx2TmXxzmAfB9aOOA0qiYa7L0EMDPltX
269mDjPRim4I6ljw6OI54yflWNWd55mkYi/uh8+b3c8ORTHdOocMQV4kO/iBtEnq
jEx4KkIzTb1R57b6Z8o0ZVjx68KsXcUzGmkVkKRc/pTWJviRiUrhgHE37mFiY/it
oEvwfHuxImqYuZzqUwdfR3Vajj//ls+jr7w8oBuTTrArBw0yP+KdKrqsrfb+oOWf
q4bNMlwZSCHwWpYzQXysXs3ohqAiozsg3NC08xnMOoMNgRGQxDArbSbxuIhRS5gW
BYVDFcjzbsguYKAxGoiS0WdVZdowqqjGrQqRbfJyl8iVBAKZqFFt5Zzc/gnu1YVM
5EFIM+dZ2OsgSKkgQMLVbk5xda1t0zKGxj/hg5Bj88nyvJWOWW+rgueIZyBDC3Mp
8P3Dguom7vO+yFcR3tOvVs2+asd0k6ce2A5UdYHNcH8A2LfOgeH7/+Nl987IDjlz
Iumjp1oLNncSPQeQm8p6xjZa6uEOLiMnUln2JenZE0z4RsPU1JxtUZFJ5t1eaDTp
ogi+xxz2yZs+i/TgwRH1J6s9S1CmartZcWSuVRRX46Vusue5rVguDZQXc9WQNRZ0
7+QwSVL9J2hf/UE3TUMhOIe4HYsUIlSDrjp0AKc7L/ZtevG/TQ9R4VaPNoLkNK09
WJbWBKXhtY0Y+iK9QXfxhZUEK12uWATjv3pqBc0BWfzfCqnLFueRZE8qzQ2/QSx+
1BbIG6PvskVYQOPtv8rrDTWGm7f6XxEEgK4z6FpkUx4s113fEkkdhsTeosWxNkTT
WZHGIhCzTMBLm/0LFbaiNtqKXctAGdFiiBcIXefQSC7oUzP4G3PU7BfBVMYSpFH8
z8XiZbJ4gbF+gD+a/XeDoZXXOJ0mbshFhgSN3x4dpgzDDNlvlH5/3DZh3kYDhRSw
f61shLf401vSr6iXelMWEzgMNA7Fo2C3gs/SvXtjZ7jjl5YpuabD0WwQ2QM/SmVr
94J/2YTviveAjFn/w1JBozzorJwiKC+a5DPYxVFKr5NBIWeauoF5ltIzVC247LaE
j59wH9zhR2mQ1HsOpRJCovm7hQc3ErgW/SGO+nvwtoM56l3JDv1yVdR42qBd8yKC
14/aohynAJ7JZhj38zQPEvZ6IgNHnqOOydJLtRvmqNQN6sjspBQDKRHSQ7uqPqDK
50A8lId4sgjddAkst0BGjdaGKVa9JhQdK8cRwsZp3Z4+86rpbv7sawyAfUvJeWvf
YwbQz+5VqFVLWdSUfe05CKbUliyEDyOOukk57zXNcbJIYv3MXVRcPbWcQa/PeudB
Yj8yXiwB0cQhxcTa1gkOUIJgps2Ux4By5E726VAqemd61bCIUlpLmFE/nikLpvA6
xgwKIai9+m38sKG/wgFv2MW5I8aFDTGz181jc+ttkHOcsj7T3izKde8l64Q59Fn3
k21qO/k9ffuF60RteFkdJdNU1POhnjAx/r1DjfgOvhIexDp0VP1gdb24gCwdu5xU
zpAh0JlRqiTGYc5x8VuubKM5tm/Nc6H0kjVSGGgAhjTzz5L4okBl2fhtvdvW4EQ2
Vv/m7LFvhqcZPtQ/xsqyKzwJxo8wcNY9zRky6clUOq4L4gtdFnoOyT1siGlWyV+u
bguaf8G54BUDLQhiyEvg3mxnJRT9/fN7fA5MnEuqEZ/B/tCSSBUahnHgErdAQlRL
K2LSOaXzHMBa1dDFmvTfDUvH2hnxzQ893hSTvW28HFpJDoGfvdK9vepK2QJ6yLrX
qhuussk3TM5bw5HCDT01psiA17Gq3LdwEbqpXgoiVrSMKWqMQ5apEI5niAj/j+PW
JoiVc6wzNbaB3rSPNDGzJwVwrVhGGnhb+FtwSw4jJ5utjp+mzicEXEp+aZHZwccR
KtocknWXLeoQsOYBszG/Pl9Jfks1e03vmXvYyIK90Vf1qeq9D3efa52BMLiLSlCS
Elv8U3qe80/Zi7Y8m1KaOdubrVoqs03AoSyZ/sAymKCsGGCAwvloICbFnjP6eOlQ
knlLhn8CQa7Vk6/dmBERpTVbW519vqZsQHxpa/PW83oD8oSjjkaQLGcEfWyh9Iyn
eb7cxMS/p4RpH6ztQB3hCHeXNM64+2ZWYWc20R2WKuy37TGt/pQMZeufodjfvDsh
CLBkBumJuOLXER8QsCKSxgE5TawR7N2J6y+/WYMmXa5cE4JrK4m7vbph+HTwciX1
PMixOXBuQM0yiSvvPNzKoUv4vF14D78zT8KdzL0UwmWIX1wyi08wy2dVzzXKY+8s
N1rLV8vm00ulMKDDZKvmn/Hb7aruXieKwlTRcBm0hqXTzgkLt5+96TIY3jHvZZVN
fqz/ZB4J/05ONCvozSBgn2QsBKkZhbxws7nJgmYCr2C4FbjySd/K5wGgCWxU5Rqd
FzcTB0Gky0lHjXtJxVfRoewgEY5TDgIbCNxDIE0XNIIvk67dFrEX6ORNxMqv3TRO
DGmSff4g2SO7Yr4Rfp/LKBojuEjzMgZroYPSgtIUDw6ifTtCbzs8egNOYWgZVkJh
70ajfyHmn0pGXy1dIYXl+1HXq+NMu4My0fEqr0F6SkbdC+TgbrJdvCv69vVkQb2e
T+0u2/T3Hq8d7J38wKH0u3IhWqTURPfUPIplZHfCtN4XFPORTfEJH8T6zUO2sfCp
IEJoekQKqCW+In2FJzrf6shldKeExZnnJFXQdzYy+ypkUztf4VFBc0DAFBSlefd0
DIcmySF8PZJ1W28vm8cQaknr3xANmw3jQYbJJFWscRGu4IfITyKBbsWBnNtVC+tO
XwqDH3nKgOR4ObM6t0O+kbFYHAI9+D/wGWVy5LUVAs3eaHn84oSwVR1x4PRHWlBY
jTPfWHwbmSLZnPiZzSqHtUVVFpHOX5/THUY7L/9rNGjqugTZ7YcYxtAdG8+zTXFz
c6iL8SpR5jsJCRFF2zEzFjAX3a6WD2Uz6rs0DIIEC/8pnbZljdw3VOBZ23erQ7yH
nU8yE29w+rF0tDwlZg6PasAWHTD7dinDLmNl+XkW63+l+/wOll6MB2v7pfghKifE
nVzatD0ro2YBEtYeT3N4biTnfQzywF4vkxn2Up9ypGgqi/i3srKrhbb2jeCWEbei
2PyqNx9cK/dYI1lbClCj2FbK7raMMbBHjtIfiFonjOd0LBqtvkq8zyrcC37KePoF
pEjq8LBNEDrYh/vDvV/3ejubcR5haMM7l4aRNRnQr/HOspFfX/DUUE1VLKnhd5T2
xrZPHufCBDOGOMjxqKABdS01leXnQupiNBP7nwTPpyAt1Ed1/pWaUB0Tg36npARN
oyc+QBVfe+Ix2Kk+kM+/i/4srQV31UW+V2wp47SzkrVpbjEqrnbT8/GBclhvV8cP
H59VdXN3fyZ6j5veerzQqUcKSd9tXst+ANlHNVDPt1PLD3OycTD/G/vAGFhacZDX
LezEVf+8WwEbGVUuefGJsxnv0UBAmwFwxNboGZewOsBJ6GzoStrWoU8PqOkbGFAo
eCg5Fp5EimXEIQFMd8BRytszA+jDZ1tfbK/xMkrcT0Nt1V/hcJaJpkxMPGuY5m2v
qIj8UwIdlBreOr/QPoAi0Xj3uxL93862Y17GOogbTeHRohU8FymXdTzQyDmQbstu
YqmpvVw9KPrWk+XSqBGDh/N6P/xYQJ9+xO8AWUA2KHIiz+BdO+7BLUDOCqGrHejx
btHCVP4uxFlLvVN3pP/bbyEf0Uf3KXtIjyHzwxIVAxQC59XzTKbgtLCNNiBhOwA+
fM/guf8Bi8ElH9nsd7bfSuvTEhfXhKK4cOkl+Url/DICM7YNxYyImbLpHip6tgeW
a1Sb8AYspRSotpukNt+j5OKjZqA0hpWzYNF5yFEF7rpgkfKaLkbm+JIHLxl0+kdo
zWuk3OaRNVdE0F2YLZAPDzPI21oZbhbB22Syrjq11xSzGGmvDjI59jROgK6A3md5
GvM0e2JjELEUoadBw1p0VI6x7iSxdw7lmwgoZyYnlwj/HXceyCTRSmXwU2DoxHPF
ctPTDkfnuTffGT6ilvywBc+PO81OQ++NMBOpGdBcCTgBRKsjB3vztIcNEIUL6A98
426g0abP4d/AinrRBXamV2+SjnF0qVD4JuCfIOMVM4xBPru1RWP2J0IiT6zUP/dP
Iq+K5jXr0Etx5QO5ToVOFmhKNjVfDHt0Q8vC0EjiCzz3rdBiuD+rd/K1Ar+79Fmd
cLa14DzZyi/yKZ7lS7EGkYCjQkYV+1BdVPaZeRDYXgQiPPrvbNkkgcZhMiGkZKwZ
Zt6JnHS5F7Au4DAccBtQF4WELHEObgPAN9jcfXrEqF7yvq1HikfhNMhw8zwHtfnc
yWc4cyV+IUW22XSt2of1sAXVcgzp6UKnTNRnk5p20tpXHAe7I949A1Q1F0iNl4bf
tK0yUDVfqXMJLfoxlgMn1POEZCrh9P0I6TV389MBjx0jZ+AKi071m0C5vI/B/2jA
AkwZEHlKbziNtyzK5VJC04lWx5WFmmTbkO+LOwu/LmlUit+0RSCdPqunyEwOcYap
2FieZm8cYfF9UO/jXio6ikUIfRvm6s22chn4py+/a0dEvep8marN/Ly7ryW1Wotx
1nFiefowxOufPOtZt0ZxzKeXEABEG+AMrBz20/nJE7cmqQxNEHtZ/ylnxVCJmgaZ
VfWChIh9BhRwaNrDHbs0rqQG8ggAbUb+O1ERCH27Iok9cqbFq/sgPpevU2jxfu04
kcLqVPr6nHgu+d2084paYSVHNd6YzTcaA+CK+r0SOHXinrw0UQ0NeVxTWI+sJsUX
dJ4vqXgfHoxZt6hZzxAsQMj6gIHe70kyEwyzVAInk7PywLncMph5vwFhkt1PTBYy
TcNOKAScCoFICEgXfzM/gOgcAp91GlMp9iNrSGKokOPc5VmADmN8HJxRFpIy7GfD
c5xmSm/kldq7i0nLJH8XIow09fPGwHm0T/DvK/sGUcDUjgCq1Px9FmsHoMWxBzZC
VLKrvTTHB1VY6wwnS9MhYrooi+/13xATUJH5fgdp9QV6M5HE5BpwfcHKGTnhShA4
jZrv0cxDlYgecmrT76IykjY1RBJxZvnAYUDTwENwtvEyJl+0uRdEsTue/RmvSZgd
YF0HRtrzBNq3PSrgrq/o0jJd6/YEpJv1F7ZTmyajWzni8eKremFyw5C5D9vPNZMC
I5QYHvDxNYXhXlYs8jmwDbHw1tqHiALBPwu65eenssX30wbAOMn9jRbW6n39glIc
kySl7Rb1y69NqPFRv/DTC3R7/UBeE6mrdNFLJJx8eCDq0Nks0bgZqkn8sgimsddm
sUXWjnyn1/MtrhMqKnUkox9cntNcjVC0srP0c8I2axlZIyydbxw7MlmPrzfqHk8o
Ii4nWtkpsv2FMJKHNYhQyrPy3C0onCG2BSKuC/kS1MKCRB1o8xNZ4XlhVOBlju/Q
Js65gaFewY1cAfeLUlEuTzm5lAbn4YWZ40koTuXO2unkkethT1s6DpgdxMLqWMbZ
nAYQ5V7WyC/H+4EDXZbQnLEsE7mbpkA4aary2FKLG6OWnb9feH02UnfjcmYRqQeK
NjzM2/UM0iYWDrgI8zKoGNuqpiEysllIDcj2CdTOuAGtZwVYa8AuA4otqAOYDOKr
QNPPMILXD8FwgFyRO1pa1F+ofFPwp6hK43j+trG486zqsq8B/eeJPh78FVwHuaaa
QuRgaWphxMWerlguOIicAUGwbC+tMBAvqoB4/al4AAQAwTV5dDj9D/yxANJqSC8Z
i8XmzaXaum/L6gpDgSKCsozUdJC8roikhm4gEt8mz4jf7nKY/TVTqCuC7UGZy4bd
0BOuMVE5ZBD+WR/yLSA6XKUua6rjlB6p/3HBAD0Rj9G8XEIb9DyWG3PiKXKr4Wfi
67nvcSjaFu8NPWY1Yh9eo6BkrPTovdmgZXZqExA7zQqQsej3g/mpj3EjCB6MYyaR
TBruPus/YBlfm0VECA8l2SNx176eZNYoECtsBm5+08Pjh6N24SYpR8Y56Mnm52xg
Wth/hvri7in9O6gXd/FBZcqSdiWYxeZWsqt8G1Xs9WosHV1ra/pynIcQrYP1jqIR
bYsUazqd8jx/vjSH8mA0kNZ/1ZuzZfl9x6iWs3GDuGWqfV6ZwBwSaJGwFGtdSVjn
N1H35Pc+3dnAsfnVYZ/ieNOzlOYFiRfSEoXz4GZTT47n1gv8cRIOYkFTi4kkpDqf
qGdIjxzB5WDxMgFhYljLKtBCHQV3s1fZ3UskjQ70W5qez8Mi9s9nU+XSWIMqUt06
t0kDvfI98Xbmuyyq55jciX4OSPbWSI7dJCeYlkVoPfPMn9igl7B2890FvDtmwSM2
w/kQXUhmmb3wk3oKq5SM8bvQPjbgj8MEW/aPlBNYONbat9u8EjoT7+r+Lf6DejEo
bo+ExFl57KqlnZJmzvKrPI3ksT/++83+s1X9ic8WbSkyaWfpjK2pxtnA9D2cLVYA
dMFrBErpgV9w0SrVfBPiCPfFH34IeRUUMOqOM/Bqq8JNsOFVFfDXEFkz6aqE+XLB
f0IcNd1kB26WmYGYDniO10hRelI2W24GmkmxJpR8MWojWWufca1Bg/Y7X0q4Fyz6
kOKMXqNsMqs7IXvTZam2AYQVy6FOyTsw51aSskLQqEoCNvVWHSiC8nVrNvgcKFrh
FgCxE8nbdga2GJ2z3TQCLf/FQVUkj7UBjJ7a7n4daxCDc9SiDBErdYLyoUSMDjF3
CGN36SS3jhPE8JkbkseElLUl+oOpSf54sBqSBQtSjue62m2s21Oha46xFf9vG4fD
im7uE0alxINcixDzbea6mlPfHqx5i0O6NLoUtZ++cpzBUXrN6RhArCHHrhTYZpwt
bY+xVpTZdXNuWqRX3ojRyRvxha0oMHTnn5JWCk1SQemA1lTMeYk3BOmkf36j2guU
g68R74a84S84jVCJ0Ikjq8oy6ioiy8t1y26NXB0Egg897cIYs8VyKMYhTzf14kJF
/cGJS6p4zR5hr1pjFXhfg8aV1ZvchNIiFRm5w6TpgGwaEMXAdSkrxQnj7VYsYIRj
sFfXGveuruSUrJy79dyNpi78Wg0mRXHHJckFL9qvr3qm1jmuGgFa+VMhQ6COaML9
tWGKK7XdeyOijj4FhIKbogy/7pdMn1pPEyqm9DAeQMZOx+ogta29cHBXhWyrNIQs
ajB4Nh3W9diL38xKCPnrYjX+y68iyOMibY2Z79e+xrIaaVBNnmLOgZqCfPfCgHZP
UrM413wiqjAFxVelaV3AnzEB2NMy/1npX+19fcpzApUM1pcHqP4YgimiJ9R//T0W
iZP/XS4lZwz5WsEDOgDi62CrCheQeCOsAmw0i79emW08W31eEnB4DJmVgb2tifCS
22HbcywUIzDuJE9OQ7PswN0uAHlhP4v3kjqqEk/LyoWckALJd9+gQSfAT7ceX1m9
EoJE/o+YXphVtRXAZcepIilWXLhvQfgpxW4orbD0Qy17h+0UTb4wPGroMrFnmLSC
tzp4t5HhA1cX2fgFgOnrcKyln9Sb689TYWawYJWDeaHgSDyEKfB0nVSezu5GKrB2
2HgJVljAVs+yoxlpS9KOkq2mO2VCTRTYlXgphi5UZ0ZhmLhx5iOGC25AUZmQbAuI
1wtGc+kHo/cYOzl5GWK4QyT1Mb4g0Ie9lKRo8NdoOayHOOJMFGVZRngv0z9QiDDE
dT+8gC7+lq1sO43Avcrq9YF5H4/yO8p/SA6NQpGGtMlZDCM4laT3r8iLHXfnKIdL
DbNbieNDVWqNJCs5Vdj8E6YJdTOG3Ye0RWzjy5JkU0SHBQSPFen6y7p4eCTWzqdW
zHpsUWmVaISRMrS1TAaRIkwfBXQLwWtIITezxoJHfJT3JPyOW84XInNQT9GtddkG
DLSnZLNSc3fpdrNt8gP0JmBvCVQDRgw7hfL+SVbIvWh8hZvyGvmMyC/YYQV24Xl6
PQF+Ji/M9cz6WGErnAMo4vkx89GMfNP5I7q8B3M8hSRazLMrBYUdrCFSxvMmMTK0
Mj9q2399rXxw3s8eTwRmA4u0cNTKQZNY2tFCAOoL6HS4yshlOOQh0NF8k4s3J+dG
I5ulxHD6ZBpf8hGWe8dTKady0CxwrLtci9OZmpY70NJBFLs+1LLH1wRwRfGHmYT+
0vZ+WRuYZhjbahJFc+C49q2EGAGSZZyfmq/yj3Om86BDot8+rQHW5FAcBQAbc3vb
8f8Ry53iaMnlIIyBJvtax3WasZHMOpyId/uqjLPs5yqKEgD50zlGLGWxC7cN9YsE
vM1wdfHdASm5Icd6kLEeV7oWorPbXAtQ7Do0a6sBa8Z9pHJEaefUlIcnlk/ghWFI
ivgHy5oZx5HPh4tVEVxgNYhP1Fvt5i5buXZpn7HpHqQsBd8LaEX7Dro3qHWelzkp
Sj5zH1fw+eVw+y1PI+z2le0YxDrQYUIk1pszv0zQIm8+d2bUXHVEO/2yDLrphYQM
MUaYWmg8N5Us0Y8a2UGCqMYOpTznO/ByrLtelP9ffvQouEsY7Jk7c22dZ8PKLhJC
5nfOvys8ZpckPWaiH7RAtaWMkJH+6Wj7ZUHZQWoHsmC/xKvQsBvcXyYTp54As4dX
H8klmWrN9/87ClmeY3cOvVF0iio295IlFv+YZqx0BaSkr3+INwcoq9GJefoVtOX2
hIiepw6SPl2+AM8VSmsDChSnQqCfBzL2MVLL/upW4JPHhBdHKoW2jawQbbKTto1x
bwKjpMoZOJsq/HtG5+/ZFOWN0PVNYlghGQwYlkFCmqeKug3HsjTA9j21NGh3lj5e
eJXtazcleDJzjgcjNArWQ5KOXv3D+E1vJuvX3Ez8jBJSklqeDqD3IcMZB431gbfp
PHQ+Hs6ezsrWE+fdUBy6591N7rQhB8ODJwPEPknv3MWGQDwEnP6/xaGw0zqO06r2
2DxrjYdBAeio+5nvtJEdsRlXnaM4/yWNO6kp4mVVDT661LSYjT7Xu/dn50Zcn0bQ
xYWsJ0IJDLjJL1IQ4vakXm74RI5md0UpVaQ9TZsBqqY9UWQ8YubeHJwFTmm7zHUu
LgmxxCG/ufLG/P2JyLdRvnpoE4mQ5NrQU4S6SOZcDteMk2sqOsznjKvRx11S5sEn
DER4jU+rHuoRxKWTwxU8ZMv/kujqPCGXE2MUxtaL689KFsxHHB31kAzlaGINkn1C
WGBTcmC9PQnjOXOLdebLdSn7vwDWkuQ3jbk3VD+dm4p4Tg0l397ZSzQpzvi9/iTr
SB5CmUBxqr8GrrZvCD63VvgrNtvbKXTBDCBC4nFZZTt5T/DM9rzd6JrQjPD31v8y
jrCP9Tz6QP9IxHVnnAneJ/o/5mF8GQJv5CJU42ASXZ8bD3Kl9FEzUsnvp1pzYcGE
V1xSWS5xJIP7+LoBcXr7+J6wlIou7F8rSftgMYND6Q0lRpECooUHaGSxAHv+PZnf
DMFmXSTgBQHGmKfQG/juLjt1bOuO9LTrIyJZhLH3w0LLY8E4zrYeSksbd0Q8LV4H
Y0WIE2vTQHLJdBeuMtyyiwNDYFombmeTUubB9ovl5iIU1w098PYe9NuKSBxvDpBk
Q2uUkQEFyAHrseBNoGOTLNOSt9/CjhXq3RvtQHIyT7b6PEcM3lY5yr0Y+Lvtxo4B
RPXwpMARfE/zyGHL8efPwD2W3MiJsU0onAme8IC58y1CFqBmu9avBpT7mhw14uAG
PzMnXFHxkHhVPdEE/ZmWuKiKn36/q3rqV6HPo/WBPpdejM4fy+lbOcsx/MrzbzGe
PeAjTQ+lUZCygX0PIz05CEZ0TZFYqdqGWDbUMtJMtx53rq1omJrn1MreKHgPBimd
OJaAhwXEt3KTV0dMEnLsyHEvFl3CNchqqUJAAVVSqUEltAYSygTSDo7IBPOJc1tg
QfRcwgG365vjc2HBO+FFDjord0v9mI1YaM5sNGzBddNZENkOE+XVzA+rgWFofuh2
XVotZFX72/W8h7Sbb01RXjGprriFh1DEqrQTDlRfwKsiG2yQZK9++PiPyTZ/xQw6
EpBOjmmBKelvl+KhhNVSrzgDvAjfPYiku8p23l0FmXhqtImhP5awyXMYs19fxoGW
qO5bnim4dTQAnM8Hl3O29OnZcbCFO7n0gxSdDWzviIcr+/yDEXpwKBjQ3O9T9+Hg
GEjmDd3Zt9KelyOJ0PcHJk3eJSjW/6mDU9jlJFbfjs0PH6h4w+5e9LT8LZpNQ4/r
VRt9j3LRh3s7UWi4VQf8v3EP98i2KddcXiJTQjihtmWjOEI6KH5wipyTZkI2Rd2Z
eDIjM8mADN5HoTVdnX1GQf7KJ50TCMuTNbU5SpVz4dTDfJiJ+H4XTXg73hP3UXxw
hCw0HYEJdoAgw8Z64cIrzTfTWZVCwpt02xaKLR4Dm5H6S/95tvfwjifUlsxqrHIT
SeQmYZGluWI1WtWnQCPJK/4rWO46FlNVVZbAipfzKM6yxg6x1WgVx9zsSh30Frd9
2jt3DAI/kTpH3S13rtb37Vys1/hDX2WqJuiI7LS1KB0J+ChXbf/6R2KOohLr9ONG
TxCPeCepvf0RxqiR4BhH6WwZc6BXiwxH8zkoRkm6Pt2vqqmLUNupUOCE54bo9vev
BaMBelEL2w+qEnx3sqYcoNLl8m63+jdO8/VDikxvQnnC9H+N1PZ4EN5DlLCJStf7
C09gzxDJVqUQUM02Tk7W+IUaA766wZTsSiWWpxBFWP6Xh6eQY90CSGQ0+9qPBoG/
+nwjWskc8K8KhXx9xiST3sKoDdog7ybnNBlGOnm2Mkds1cMAnilo6HvD8LJtIGVe
TQRcQmIm9PTY5wbZtdWB1gfHOUmU7AB5VxlMy3oxUAztdmyepZ9DmcTklTDtDdRr
mK0JCMQjWsMtwU/T304dkOnDrgQdnsaXAu+OYLiOK2SCOEKOHlwnWSBGd6cJG8bR
K0Z0Y0DWGcrAMFO5xZk0amn+eLxFZl7L0DvvgDI2/UqFeO1tb0QEIKiLcylz939q
fO1wMjJmIqaomHKwEwC9kWCQoimzZGj0g5NonMykTU/NI1kkhXuqxnZakDQdxKwz
xTCzAMSiuVcruQDOPUdELo6EitkU3LqZox+/7YGqm5e4OFG7DBOv+t7Ap1xiwiJm
TzfciFKoigpV2yxdu1+M/LVppnApzfzWnQBupxf055B9f7gygpK0+Pd9YNOYd1kW
Njkqn7eVNncKqUxoepDAjRR86jh70FnABGlBe2GNdQL3woSGGhjKrEs7rEwqmr6b
oORuRO9jH4ei2wA2SHOoXJ8k+HSoXJRvbi9E35h7FUA6zAYy0wEHE0Zn4CDhVIsX
9iDXt/gIJGyjzvvVg8wCPlwQ5cP8PQCb/afLDK4Wc86FKN5YFR1nRHLrngX9Bbj0
YsVLiVttWpkyLVexTQnQoGqy0G+kr8A3N0PTqvO1jd58NGtQX5lC1n4/3+TFSAAJ
uSeMxI50W5GyAC3DuFbvM9N+9sMy6drs4pN/JUnUQZ68UN7mDy5YT/yXz323BPNZ
iBWZMuYY1Kz/5JmqNPKOwYsw8fh5BrJhJ8fHPuealx5X8fcpaLF7ps3HL9h1jPWx
ABknd+ClV9KnjGrKUAbfMYESAPBn69Ta01AI9/W8QLWaz2dILKYg20Ec/UFyIVbw
A+RwTFybBXlLXMHcmOTPCOHpsvccIy3UzQ0hPi3PUnHHsRHxm9LE00u9F6NtRuNu
wg3KJEDPUzp3N3e8MwcI5EHvxCUvd8UUezMVoOvs0MFR9LISuQEZLGUt/YrYyu2Z
HBltaSbYZd1mmLZwurkOwjDaSZIm9ppgBErYiPy7K8QgXnZOdWGnLnE7vq8rwsDe
UyxCp+y4yhYKZdUsWW14Im/HXamUHdbssaK0c5vBezZfUuQKNs2+usQinNuvKuHG
OgBA7hpRkzY+g3CbtMcGtPuLSCAzyfn/hc5gNsCeQPY5pbFyjyFxFOF/AKFsYfNZ
INix46JJpP2c9snnOxNUiqdew3pJu/tK3Ohgb0wT5DXkZhObIS3SRQNaP4glp+pv
J6BA2AVqOHE0YFL2SSpHTAtB3nC+rg4OV4lgZeEb4aKybhTxKN3D/Oa8Zd4vHONN
Z+FEbF/VEdop8/JUci3nPcYY8KJKoDch479zdEwhrNo1ZXFiYn3DMorBBvlcC03L
gsGmhxgBa22v32It5VuoHVYe4UcsXE+rTsgf41lRjKfiv0riawE0inADiz3snYbw
dJDYQoHZp4KDZipXxJJU1hLcctxPGu6iRAH5ARrrE+ZlEGueFXkBsSLuI8tlTBJt
NMZKcTdO1McV/PTC49zhELPlqENQgcJgkSM4juSKbeMGRd3wUJVkQBt8espbV/um
aqA4xCmz61OYfjUKvLjdaDKPcZImTEPwjDdYsjuH1HxRntnR2Ry/S8uon41+Kjxv
+JX9HY/3zwDzsR+ijtRitVVWQu7AK5b7oOtcXHun6r1YBIt30vqeLXc9geVRJOZK
ljsEf/2zvcoY1dLKJyAY0fSiYP3sg1g7j2Cc0X3/1a7SUsuNJ4RreesuNAXw8453
7DThMeeJtjFYApECRhArcqp7ye5UX/fyC74hkodYZzcMMsrL1aE+MgXQHj4VxMXM
zx3S00a76xoT+7vTqPp8b+eIZ7gUfaJu3oyys0zdXi/7OmGyEACCnEYMjO655yYU
oaghAqVNFu3fc/Gr3YN1kOwp76RmBVXb6osQ/mPw+P/S3C6Q0qeN9k26d78ZQiPy
MiXYoHL5A10YHlhneT93wV0FU+w2/itptsjDJqW2cIko2Li/0ZeB40pt4ACK/1Bu
CRzdsEOvMJ2nteUNyRHr+04XhzuqTQViTK+Prhgh24KCBqbPdQeT9baDg3DjWKf6
Qsp+Os2UQ7HLxCCkZwlFLPhdx9t9cUPbhcNl31okVSCixtRn2ZDzWSLiCyJLKDah
FVCv97+LaIewHWuBBvgG4FGLtbDOYTpAdbBKg7IvH6KcM581e3LvoffTlhLGupz/
o9a3GohhntFhIFddRtRkqrAPXn3lfXeRHd6HijNsYNT0o6zcMUc9EEiSrwCyNZjf
LdHtgFlrz1bQ+E7hHrIgQj8iCejvwUUs2F0BnJyRAPv/3mNEKHSYmdM/tHW4T8VS
/175VARuAq2est9nQLOvEVbseKc+ZROoQwfFxi/IvHm6sTq/zNfDEp0PLJMmvFv+
tCRuPanbP81R1nnlq5gU7A9OwU3+IwAeGHn4UelqgoxC3qu4+wIooxGBu9MqxvBe
2aY+nyndZOLJge7VpReBIGVW0vtj2ZOrbc4GZqywacOyNJlXkft+5WNKwfWDlDBI
qUNBTbr+q7Vc9m2+J6SsSo3LAqVj81w1W2oz0rN3S/xvvdRmXYGMu8/oLSoevgi0
i6GriLRkX2gY9MvLaGduJAhzoW9CE/SxW9at5h4ktbC6QYskikFE9P2wL1338HBN
W3jP4bqvdlQtxJHHP9u+H+mKyEuddiCXiPjypzmO8ooLuz6mbyS6fkFjH+Pjofug
Tx01Kj4ZcxM0rd2fLew5ZBZYk/hqhCOiofZSklcTwRLdP/+zUH9FJvmAqQ5kZwXS
LsXo1qUavCM3wp9ru3kZxVO/54CqGqxbhWV/zfuMwQlreXEV+Nu0kGIVMSreLV3X
XBJWdh+NvFuWQ8XnNLG6tw6sNT9ae7gxWp2LT8arOdOVXqXFJTyh6gb+M6vIztYs
30R15vd/h37guJb3DUiswKNWGFLIkyrR6YPB9FgdI0IxOyaF0/OPY/wA28nbxbl1
/J7xybYUcu+UuLbu8pRj2mC7xZ3PBXE6oK8iqnFUHQ3boN+t/NN/DDL86tQ/1SYe
ffTfsy2Tntcs74PC5UfLDz7dZrmcb2FhPVNYzHEIKmsv09xjltwbcnWLgXoEt1ra
sUy20zZ/BaLiW4x4MEuSFBUTzhIuCvDJyoEv7L3faKXbtgDlOWtZaXe3kRI3s9Xf
+SYRpnNx9i0HJSv0Ud5lP818k+zD1Nyb4/HETiQZztVHVt6ZZxj6cvB/1kXXCd2u
SK+d4O6VpSkxhUN4kO+ogiM7+Gnk6CVzcikJ3H3DDjEAIlxDDZm+pJaPKkzoDBvB
Usi2Lyo6Pw5zpDQOAz7bmYBzq+XezJBQqfN5WditWMQu3eohny3T9igDpBWXjSc4
5LR2XflEEyZvwMXRGRmPQi6juiVJqfOeJjRJ0UJic3gshhd11kRornLNyViDmUm2
dDXs5501BHZX+XKY5HWpLGzlMtrucy2t29NlewqovSBkPVoO7ExKOt+NBD2Parcz
nvrsiiA6h5Gwp2yndA5zWN4X0kL4CAXQgub/edQp3wkBcT8CR9wVQagBzUielOzn
oxVX9Uy1e8CVkN0myAnlFnZYaXA31lwyvWWAvy/XJUy5FNZGMRpnV5V2xxw8kazI
hE7gH3RrvJ+8PYYXpKMIlSlOYdmvhWancFfWMXaAnvgAWq7NqJ7OtSbRdkoRParh
Y3zav9I2JBNDnqb/U8Kb1Yjw984vNGe457N5xBRNsNZgzAOodQh2+loiIiAo/uCO
ZsqWFH7zgc+x8yM4e6aEFKszbFOD4bdJ1Haqrj68P0i50UZohgB0NJXoUHYPH92V
RLD2Ljbx7tYwvcli/XmYHAecboSyweeRmoP9O7mqXOIR8yEoBZ+Wb7OldU/xsskZ
n3ScP9PB23CfStZxFrde2H4T3EVehI5IQope/Ymlfciq4RIHgY2/s0ir/ciQT1xm
dvQ3jDrImHAEXV4pUYaoDUPnsYsCWnhAiL8/moJw7VWn3KGuWtR2YeRCHJJArdJc
vABHbu9DEmV0PFSa5qwwaPhUo3q926Eyr4C7pQ/3wdjhzkv88MW+l4+IBigm0lg5
5qsqHOsEyWYZVQS24jVxnRibZI6AIGb2VVrPrAexj9dUvuLvB4UJNPUCe0AEpEAI
CRsS6JtfsBunSyTw1lMU38blO/nePxnS4yuB7Moo8ZR/IVRebVbm+oRZjLsUw7AH
MZm/GBxVH/rUAWS1lGNgpQHIiNKmyWEiieed79Mkkb0fyJiamUGHDS4i6KPmhO4I
596LYUJrPSnpm5rLmkpOZ4GmAE5VQtEk1i0aGOeu75do/sZWNegJm1Pap8cuoT+i
/gs8130yP8o7M9P9mdtTgFIs8LqItG+TFkkEd0nyO0umY1AOq0Abmp8kH6NMtW0x
AM9dhey8djaUfnBltfg5hqcs6FkMwEr//IHnKNo0ts3NpPASFnDCW0LcBvzsGxau
Ha19AJuB2g59iRxSHq0Kyg4wRkPLsAUQBjD19BUwwcKOOS66jL/grHRz5tPtuurz
x4Z1G4KefdEIl+5eW/wZBLzDnk4gNjUTEU0+jzCYv2U//M9T4HoNXNm/WeAzcRiT
wYMIN4lF/V++FgzIRXgVb/PggNXwENwiVyoOKLJJKlmGy6IycpnB5ksbZsRR9iDK
v/p32v3gTjH3RMExuIDCfqyQHqYftcYIrG4mGehTGZavBOYrtj8ne8YfBXcA3s+B
2OQKOvG8wmQ4s6iZaSAOrLN1gMrsxaxXDAAVL/7X16t8E/bnsIPlNn/uVZqXTG2s
tEWDepszHP8kdvE5gTG5qBP0b4pPQ07ZSVWmMDoWXNtuRWiKjIIyxIf5TVoAPAua
xeY71/lBwotVd7md1nY1+/kD9iX8NpdpLwJRWS+znctV2oAHy8vioc9SMYt/Plhi
ikWS/xJHpdhFhWrihtYClY4CFavD3+B5SEi7aq3Mh38Z7TVXG93yEdGVhGx2ORN8
LzQAbWc0/8t4hDcZHecZf4LlGXZhI91ROtE9HsxAM4vnfVfaoG00HDPZ/7lMvYTs
evrtLF7hXEd9hB8OQyxt0SaIkvYtKu+qUHnKEhwZ9Ji6kZgN1JUQW7aCZvMmfrbh
FBdCUYZNgMmuSFIGQVoCSAE5VpD+Q8qrdzM6cFqmU9F6OKwbqxIibUJMLzlRjs9j
KG05Ua66oKDVW/W3kiBN4agjO3uBo3LLs1+V2+GtdoPfeseJTV647I5WjzFH3sE+
XmXGp3R4By+yJvHIpmm1Z20p0qdglepTHbOaNfFmUJojo733YiRNQlp8jonlBngw
q3Q4ytm+mpIg3kjrZvpjhw9tEpi8qchuj/795UBjUCGE8B877jWxMeR1/6jrxB9J
pYG7Ddc3od2jvdAGGoNw8nJmbAoYteOgyZNVBk4K7d0dey4+DzV4cZBsad0zt+fV
p2mDtCYIGSbmtm4G6g/NejzN2EZVb7fj9qWZkVboS73QWnpoHbZYpoUFAT34WcMI
StkyTYzi4l/AU9j1GJzxL8r7DBpR90b0GkYLdVh/Wah1NxNxQwhANZu4haeAWGrl
FBY+NH2yQzyQ1LfV2jhH59x8j6cz1aiI5Bbhm4XPLk2d00PXdQFE7iScqSLEnZpI
MGpwzHSnVO2MsPR//hC17TYObwLNrR6BomTt0iyVy7A9pdKDH0VFvpAWRD5fQcm7
fjf8MkI8GwBPmJrP8K2HP53MTUgnAvoPcu+E4vFpR2LStJKY1trff7iPfGnpeEh1
6m+2gr92t4KFQM9PltyFv/T1jBQ7L19FPVIhGnKt4jxqsI49R4x6W1t3VEAsmOGU
B5ss9UXz1ysDREkzrfSonQMV7ou1Fqwvc8qcoUTFnHxHi3OOdTXwAvMvR69dVKQd
1SNOd++6IaCCKtJO6YCSGUBMkVtth0qnpH61hDdUz0Pas9Mut2IOMECCApi9GYNn
fHUMIQDTIxyDqIMNAXkVmTNDHoY1jkFfNU8tSmCDq/m8gBOtI13fTVIP/cuNR9n4
hGHfTBFZ8UoQtIt+RB3MKnhkxnWKE90HmzRxOoRiS/B1Gvp0aUQl/fW6DSywyzOH
7HHQVnbt+rGWA3Jlx6STDmF3xKcUJ6qtrqBOXREsgcvX4lfoo5uD3S9wtETjJE3K
P8pQmJFG7E4DlnrNED8LKLKlq4GqlYC8+rO6/39PvkSP2RyFAiGB+V6Jb60ddo/c
5vjTjovNjcu7Sove7D3dzpLrii/5IQt3vtcmfSpALsggUOiDx3ZgvQBnz9EI/lE6
0rbbbGnFHowPQnUKU3wSIaNerz9vg7NNQN4N6rP8JluZeSni51j7T+4nbrxEGY+N
SZPu/VqwnciUP9kGBRyol3/87SqyREaPAFm15GO8o5R4wu7bPv2ZgmQr5/Obzgtk
2BW0x+IsuI6CQ8n5/Eu2xQF91/dqxCuWxlx7sfF6/KFY/hPmtvIdDRke9assYfUO
oTLWNfGNSSvl38B36Sbh6QgSVqksQRl7vpCBUsvSStS2SCAC2HEbAhkYu1cTn6zK
otstZ8yZRjgbzKrC2JWtnS2UvijfDSqUebxF1lYIf7JamGR/nBHId25DTREpe9Je
pL65Y/6WXr/swpv6VlbIKoGoJ6KKR5mYXciQie8U/tfrRXS8CgH0/QkuCmTnDPck
qWOz8v47MH2FC8jjC48wizMpJ71HhHY2x8+YrU2n1HGCllog5X4ndrzu/NR0nOw7
wGZ25ZjNejo4AWHfhDeSD5ijAjiwKo5nK4ufOLgM65skYm8w85CWhd9tikp+q72E
tsr+WpoGOC8rx943Ga5b0D9B7bAm6mDEm4044asWm5xFAuG8CudydVUTUgiJYCAS
JaCe9U99nCL9V+QZaQoznbSMUhRG7KebdA+a6q6qiN8yZb/zQs7/R/VSE3Pt0OmA
h1Ag//gge1QEx7+c3h3771zmnn5Yn9SFmw9VweYv6pDNqTy8zranTlsbh+PGhQ5h
mcyXR7+dpNrgVT9krIpOu/dGV0+rtUiOFRczas4pqNvdnMpIIBnA0LgIDa0DqSWj
PahHKqV4T5lY+u9P0jytssUXJlUk7PwAxWdJjH+RAnoawd2G7QzUHXMaGTvse44S
o+KPSjpW1x5CrPDGuwCSOyYRIDaNU4i7qv53zG4/YJwo3NoI8BvfL2rBI1g9xFLJ
qtuP4ZCANVA+Jp1oufTvhkwFf13aDANL9B1m0CNspKLXtZn6iHCI0NjWotVG7v1M
AZxO+o1dE7mxMxl1/vgdEBLpWAXCLJyzj+rc9xDpFFtQEE5XgH9yT/3hDsejvbk0
DVeU+mYMWLjvNQgdPvKwC4qCr+T6G+AfflmOwzewQ2QQSG8ltVsYVAJOm/gC3TW7
3jmnN8oBq6q9NjyJOW5vhytV9MnvEG5Zj3g4eD/iZ+1+oScb6j322V7xJTGadmW0
Rccruxo8QWv8xE7HONVx8DNSa03UF0g439tWSgzc7vn0E6uMd79V6LSThWwkqTky
a9+CwPqLbGUgFRxSFjNJlY4mkcwLUhlFuLLfU5Aua/DmOiNQKqDsYu9JtlNspRhF
vIAn9wPkCTXz6TJPuB55c2yO4rrarg4lNU/g+hLu9JpcKmi6fIVsmifBxtA2+Z8n
vw33m9i2Y3OqU79n9D8JpzIzr0MBjeZh/l6pe2XFRnDn2KAfkLOMpL11u2XQGvQ1
y1X9azwqelCo49gxrbWKTJnd0jUU31j7dyfrxUa+lNgVtPyWWQeuVXqXXmS4mm02
MOAXAfrZJWZqV+zk6gAzMRYZXZkfUKpBkMshqZ2zBV1zS9dNNovOOrRU5d6kmmtD
j2O1kLo+df1ttE9elSnYm1Ah6ubIp+qPGE6Boi5kR2uM2CKp5dAN2149nI5fRCfX
qgNof5roG8QLYRWqrnQbGF71MA5pAHng9/jkBdL2kR/uR0T6+BkJpFIHmrM4Fey9
jck4y2GhrdchmOSpxn3Q5EyIJlf9mgtzXUTifJTkARGisX8mhyMZ5hSQ6alPDtWr
W66EhDhg4aCrIcIUgbk/LwMnwsFFAYodHB+KETibRwofb3WKVG6M0FU518sCXKW5
MI9Nt3CS/3Gn/vY91fsEGS64j3+X5abxcBZr/esy2lBNvq4bUmw/KhuxU8eDYnLy
e5QFXWKqLdQuIsuBMmLAMIg5uoC018GfQJKdar0zzh9vDK7gT6kDBhtClJUfXEVG
7JXMYjziVN3OXu3GpBocKDXYErXmRROky89E8cP+CD41VOOEOdbvt6miSP+nJzQr
VPMsVfHsphSSUNG9KjsITLaOMGrqV5GDoyCmzqOFkWUjb1JPLDwtQdVOD5HstO0l
HgtN5m4ARLp9+qqxYlDs6qInUQuT9p+nFMG+RBvEdcGNWjfUUVqwKQkz7YbSvI5O
cZpHIZ6QRNMnVz2BSdFVkyhj0FDY7Uq7U6ZiNX4TsY9FiWkzAuDS0TJS+MSIb7Mo
Bu2UZ+Y+wahWctobnV0svA82ZUaDzvEuq6+yjhTXVRNoCv+41SSCtUHr9lW7um5d
3Hq6+C1N47IqhLSHYk/2HAaW4hlm/aRecEJ2BCFHmglDwOT4Gq/eJtouNdla/q4P
zZK1Eicu1L0vhAy16V2mG6O0ZIEvL6SyKbzDUfzn/27u62APkHbejMACphstAuyy
7mY4DyBeDb03lWe5NE9l2K1IkIYj0PdEDXdrmWkTJXFmtfANq1vx09S16Q4Nx7dH
MNxg/VrlALGNmSkyhYC60ShbaujNbi2yThQPuinJgQ9DW379hsLcrXmnl5Tj5IDd
lVu2dxk8fo7e+ylKkOTiBR+MufqDLkpYtvmWkVrl0srUihG9RS3t2lxuOLL8csKJ
6qStp+kxOWVqoP+KuXGrnfk0cla8/L2kTR/jS+Tn10ju/aHDyhcz4sOOOk+3vkjD
e/DbAEXhUVxRsYoO5S+s1vXy4tXKvmSNJT++yDRIaaXQsRCFkUAc343YlVSnDb9m
O26uVIagmP23CxpgfsevmT4r7ql9pVyW6aeBu0Zi9eywwLywXEyRa2LcwKlBvveD
IxpOoRl9CsFynxaEEtGS8NYRMH+ugTeFLWycYx5uyx6Mtu8fpZaR/AxNLDjGQ+wJ
4g8Q9SZZuASuttoKQw6SevzGf9koL/RVN9Eu4KahNFwTk+ds9eTw5u+Y3wZJcG7u
dlIKGyzGtNCK25HqTzWJLQZ/cPI3rm9/uAfWNEevd2HCZR6GBqhlzDyjaxrszliz
dWXyLv8GliavWiN1+Rojt9LMBEzPX9OZ3Qnrzlx/3OFTLJFfKuy23NHrPTdhGFjx
6CtXITph0TVdBRa6GULTaXNXLz/h7taRhv4aKWIPDvdYL8cyW15jdvoYlk2xeYUg
PAVYatqLar8nn86X4LZL/ggCGbnewY1Kg5sKhcKxVsu3oOrdSAXw6CN0AtaSgfzc
uhUfhBlQ+UZWyPCsxfvbsIpw+aOhZOrUjFe6voIyZbxy34rQeWg4jZcQx29UjvGP
u1/bHoih0BOgzKWW6ekr/MpRK8eGuRfBM/KP0vPmpQ4zbQF00ZMbZHsCyVflhzN0
TSrJv2DP2hnpMVwwfqc2F9jygjp1qqL1SuF+99U2KT7cou8aZ9RvKjioQppeFjAj
dhDjCy3vnzPgxKrBMzqjb7DdaOUcBaIAM8NIKElldgABg2PAPlG7d78YKGuQckfc
9xpovcsFNFm1W//X6MjwpE7BcyPd6aIgT9t6Hfuedz3CsWiV+iI+yKUfGGyqbrCE
o+CssMm1MBGAILhh5/X9Lgim1KZ1eDfKJ4ptYKC2dMI1NY6PA/GHaGk8egkYyYPM
L9U6FGu6WSg/cHNtcaOfqrZYNK6QsQc238Z4jwj2XVVcx3gXdqwlNfvlkkeGwaJQ
hCUsWaQtC4g+rR9H36JV5QlYsugFXgXBotwc+lRYqxNfazPvSXk7dROFF1cyhZJp
gFzM/AsImQzJLd+zT4a6Zt2OBDBLi2WNr0KWvAyHsbcZVFCBALF7eaZnLEJdT2Ul
ObNoFrbMYZN5b20M5ALHXTmJLR3589faJY9pCgGnocYjnRE5gW8iJV3hBuvUWmUO
ld7rfAbMN1gJm/QgqOoZjFfrD3E0fSJ/5U2iETaFALEY8PUBMRuvXYDsuW3Qd/Yb
rc2/0Mebs77+p4BcVUjqYuNeZJ9JTLD/+9Xf2S0BT6f0tbj1VgZU5UgLi2M8xdpN
MICGmk77JfK2dEJ6XAa+QMv7W0J5elJlGIiCVKISBiMEzsmPVxvEvpRpTgkBIYlH
+GVHhsqHmolSgoZZcM1WaugXbN4aCsKDHi/MSB6MiBY97GYe5xycm6OS11MgYYrU
fZwT9Ybh+VWiqzJAPgTZ5MnArF8Fa78H5H2GXGFgDZHMG0QGJ4LdEaI8u8sJTnvG
mTH4uNi7Qz2fub23zxTCAsuw/8I53JsBB+1S4Kkwo8cXIjddROBmwGFTOJmSepTA
5Z3oyK/URJsUrdkyiecKw1kiZ1BqNhYVYozZMxn9g8GwBZk9UONmyt+0qHekv4qM
OWCfVHvukSw2KhUx+K23mwN57B5N9oSgCxF4g+8NY4GHoCFVPyBsA0dWrWOuSFHb
8q/x0vIjJGpf3Qz2RbxdhVl5Gn3kloVPBaFDOAMx4L/VRxRaNGeFtYOmRY15mVEl
TYLPVWTL+rTszZTg4+Pgkyr6NKDV4bWPEYaB6AeGgdyLhkig/V7hiBk8NZZbAA/P
+bh90FeIB8cV5Wc7mifnag==
//pragma protect end_data_block
//pragma protect digest_block
h+YRgsAWm+W4JTTgRNO1LssSXqI=
//pragma protect end_digest_block
//pragma protect end_protected
