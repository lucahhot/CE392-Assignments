// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
u5yLmCIFob5n6SKNMFMWvfByJg6tBIjHX7mZquPe6Bz4wdwabZG71VI663MSov8CNlKeI4S0q0AS
IZUmmCBXwd6wPe5nnmEgcTTNMbHoO/A257uia9dsWY5p687mWEwy2lGYnifmt7wbHXoR7wW5zjmb
6Yu+vtFQB9FhVUt+faXVzofvl5P+nqZza/AyFldJn4M5emlYoRQDWqBSdtdZdWk2i8MRI0Dhdbgw
KZGOGlrTs3RZ9Of5jM4VzmZCqmjeZv553mpvx7uN/uob1BuhE7nAYafJChwqIEkiUiK9bFw4HLxC
OLPpBaodvH2BxxUUqYbtAxV7nLK6P56mu1v9hw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9472)
gyKmPgeA9tXzztbBFthYawD6IhdNUqWLALOOGtyFh5PYDDiPJggcUqcG5v/isY5cVzLsNzQNxAxy
ZLg1SzAXJZsqsadw/zKgBzlcm8MXGtkNpf1cu8cJPoUMU2b3yFSBqCAb1lY+0XgLTCnyKjLFbNRB
911H8mFqLdA8TnXIj3pTxjCbTA2MEr6N5tGwBZQMNeztPG3C/xML9staxsrJI+Dt+MlyxkFs4Ow4
dMymvhmPOTDFDZlSR3krlp5K50Rc0Cv2EMJe2YxC3bOlgZiG9n0cwnRzPfDURPuOoXJ7HH+WRKIp
rhYS7yConXMkf6vi+Srnn1E+9tPLi9ChF+FV6NeB8g4AphZfVf31iw48LmrJXBlaSgg6Ll1epnrr
MSlf+WwfSiw/fDmbqKvGwmxdkQcYiSKYreMG4v7/PTT23J+Fzn1nWr1/rmRu2eX5GVLU81B/Yzw3
kNqnfcOlAeC38pObkydqw7LFr3utIijVF/q5WSTXW7lwdA5XhSR/NxlP6QPpNhuBq7xngb1zUGT6
RpxcQP1euS02qhZLJU6tuHu6REHOMZU6qWhBJYKQhbdt5GDFBMFe8XNMGDmQb7O3aIjp1k5BcAbR
OoMzE9eIxikjKBGygQlalGkGv6cpPQhBI0e8W+Pu4MQXUgqlAmGu9rdqUX9UxiFTc5fJ7jiaxCp7
FPzHrkfG4tBEPIgoSO4pj2JkEESAkFxtK7uHzaq2Kkbvp3hHU1iJLsISvwn4mu1IMq2cvNCVQfde
RhXKSJo9tqANKwPB7BeR/FmQ7l/eM1sme2MP7fd/6RvnUshvo+CO/7lo6GMU4b6r6rXT/coW+uLs
V2tGbSSpTNM/AI6WXX0CVOZzRNxx92RDqKkAalCAm9EbYwbw7Q/plMevZnHRSgvnByI6iDSD3zY1
Bf4nk6zWprY4Xel2fh0vAPdKWcydRBCN4ob26yxB23n5UyUwF1oeZdZEHgK87miRpHN7Hz6xO1xV
Rx0u7SzkcKXn6qplNG+spuYkElMHcuij1vMvKtQYzHI6ma7IkckDUpqW9FFEllsyP8nUbXH3mNbG
rMhQId8FZ3tMG9Sns82OnoJlSVJwLksoqHcW3dr/ujid1yyX7eeKdoRFINGl/evZ4X6vbGxN2H6L
bTVaJoyaCWxCrL2BGpCfkThI8Lne7v1HwiOpSw5rTnHEOdeS/SfsjYueQoMWDZFTGPrcENSjtVhq
GKgNJK1UqbQk+uE1W5YSPsUkSOT7m7W64biLF6xnGxLWGLe7AjP4p795ttlDji9eKNiM63ndN/i/
PSKOPZwEbaD3yZ97FcI5GdukmfajCB4luLu+Z7mxc3LzviwM6gQKlOuWcHbIAEqLLhc15kg2eDnv
IWPOe6JcvZEqGS3WzKQo9kcmfPptxSjyRuSKqXM3WtYTbkbb/zMkWZLwDMJA4lbX8bT0G1TzeqqF
/0HyVrEIO2GnEGFPABAZp5ldyYxsu4J0AK3EPrLL7blaqqcCrc29kWa2RSUUARBF11Grj+KYTaWD
sTBpyQpxKJfyBgpszqFuTuJMB1lsKBXUd4+3ZNImp+sMYBZ8YqJLKqMDRgpQ0H0pn6vWyN7AyxfD
bHFxQxB2a/E204Nc/SAKF8yyxxVFeS/X1/q69r8NCjBxEh2JiXOlOkO3nbsb0/xrwySNu81e917F
mBivvmfuWm2IPbatV874Mh6Q8HL3nbZkOUx4X6H1XSbldLD6RY38UGgAS1q/j+ApCA0/u5UUwWIM
IgnnswTAqBM0Sl4SPqLIILwi47l8uXewN92639fxckCVx+ZyLZEmKwutquSx023ba9eu023UONYz
d+Nwy6ysvcxx5ydUPPk/ESaQxwTgtYCQSvQppnBOMtZ9BSzKnqwPXSqVgl8I0CpI2X9eWmmWI6Dw
s90Srd9syjBAYFgKbcq3YToKFl5VGt91/kCK+A46x0K7986BErDB1rZ7+gwMvs4+JgqnGVuR/Rx4
mv+JlD/bXkcnuo+KHwN/ikuqqP0afqk8hpIWPsBM6dbZx8O090q+ubiNJJBA/aCMMx8Y7p/HtGKM
RB3wBAF3eP211CsApyKvvHArM4iXJrzKQLBqR000UdU1L1JfAwXj/luPV2v75QqfRvrmABXbImif
fpXUMPP1EYmfbK/VHQb64dX3bdtInvxvGnMwG7H/QX6wxM15yR7x5T7qHi/pvmTKwy6E25PSrvO7
kXChMmZsLUyhrmJS5iUrW1pveqjq5PzuP1oVpoJW2Wmbcf7lzJ08Wz1kKsDbvt0FahtTjyRusWA4
nrXWgI6NSMCBcrUIxOwQQwGjotgxlzCbaAOE7Fa90hxZGjfiiNODPKOCmaf7bwr1AWdrUWkBY2lm
WpTYuqWwpBdeJsX4eQAl9BZceF7V1yaMvYSN9sPEKht9NJVgDFNrAKkkvIcTq6cE7K2kiWp77mMi
tb2y5zgWzN8X+lpBptmCc6c2OyBbyU49qJMRlaQJNSVpPKshEQ/rePmcdzuCFcLHubVCDqulWBkX
L8GWRmT/poH0McLtc3hVWlvfQligXAB8TpiNBxtTfhBrCDVGbukii+40wcDBACQb0teIs1QrK6p/
A1Q6D/z+L5JKJbEyCtd1QHuQBp7/1xk2NTFx1cISn1wznVnujTDcTGZq2l/z6SLHs1Rm/d+PXzIK
mXobDZJgyqCHb428KHsqCFiofmYOQKI+4JC7OlppRg1XUlWVBqxhb1umQJBHPzVRfX8o7bRqwO00
c1TCgVtmyOLfou1ioau7xKqvy9MoLhkQ0G7r1NYKov6lyFqAvmN1Bo0XtBXJnH0rUJ4fMffERQHJ
LmYXtm9W1dYbmIoKrN2yVL2B0UlNrGalqHvrIn08nYDJ2stB4Vs9rcLpgnfJOaVATug495BKpkTa
UZrrXpeM/l1tW9s9qI1rdoPkIgB/rvZRT59UNBYsWUooLnrbWzrCEzwHQHTwwMMPncN9+zzNDaRo
w+mMii92VgV2eian6nGYKg2aHB/XSGN+Em+qKz7uK1GiGgoY9KZgmnpcoTt7lfLehJ1xZ0uc56Hp
NL/pl/mO3OhEMVAIPj52Ciy69iwH5FUXvuO0yD3n8L4Pdx3lD3AyEVuuPbxAjL+AmUBlzYbwWyCt
DxL8v7BDLnN9pwSht03pwGprQXKDZXgRIWApzF+wuFNehzmYlJCmJ7TG1+4fBSZW+VGSB/DHlQYi
RlcOo8YNQkf8tRrDZzNsMx//ZX9XH6Fq/R7BpfeFesmL0nZB52W+ScvQrfrql7MBbqrTf5pxuKuv
Jr2UYqeCM3yLToqYRhwaWaUv11oZMD+/ldEcwreh/Q4DVsinBIcBJtwlbLlRvSa534WNalwBZJFp
Q5+mleXoECOo0fjZTkHY3zWx2zUxVlpDPcGgr4KL8rR1xF/g0iPZhCYFKIU1IFv8aWGcnzSi/cjN
R4fHaWS51Kr5hwJyWq3yejbAwZWqKBiAeS7TZb9fp41if8P9VuTF1QNieK3HIPDQKyOwggNRf/Zg
CBlobLEg1s7aq/3a665lAphwLnLqzLJTFKi1+a8PKFc1c3TRLjAjyTwPzQvDggoCTNh9Mk4/ZBsY
jei3JcQDQlp8pKdBngJwFAU62myvVBeA3A5mEbTMiPDwVZn3PYzed8Of/9ai6y/uqB1Osniyk7oE
ealtInuxgZfa6rjxrdVly/iqWIgFPEd6CU7IPhAy6lp8aACP/HQV66s6XWKKAYZH/b0vfqsmBcwo
RISngH6z0DkCC5UIqhq+LvMUBdAdTtg/MbnfnT6wabCFJc4jybkByxx9xM2TzTeP8IE5u+iwRIw4
QGkU1Vrti8+WFgSj3usSjUlDOSRunDYcK+ve2uDJHG+pDyD9L5cfSm9HlUOlZSseFALRh/xqxe0/
GlmJeuamr1MM3gUmC+14UpcpR4NGuzMgpW4O/0EAEwlPedzSsdNlpZrEwWPlX4qTGDXdMpC5jBlO
Ow9NJp5KSdhHa6QYHxLskmMVmkgR4KZBR7eDvXHXpgUa1+Tnyuod62uaNFXHjim+Glr9BalYq1nX
UWLHMPFwJ2nFLmBzMEkDWII5jX5tp/SrNjY+JgrqIv8AJa1ZZc0f2Pg5IRR+QIsUbQyd/LASxoQZ
1lXpcR084atnsxa3ulLyosrUC1mCLuUMDQK5iAZo4CJlhCLEC0t+/82eIzdT5dck2RnP0EGtw3xi
580LA5n5gL22NAG2Bhwj/6cCztu5MVJObihAVHlI0domGGYf+XsjEBQ0faQVufkjmZZ4rFSXQMB5
i6za6BzbuOLNH600tKM2JehGAifgC3gF7wsOFC4IYVY7wIxCltaxDEXlN/428RlRCYGvS+9a+r5s
zZbeDjQxYONRlEeJpb47VWWpBoy3+Fpex57b7vDeQITvuum9aO3gQKX50OnugyMMs7Fd5hxfSldb
6D5nwQkTJaJxYystImEAsOcN+xYCI5asfhWM+XEjizDzdX2aO2gcaffB7xTEorbe2xwMj+/6YZjb
pR3qGIiQkABIKOzguf84KmnRN5/CLh4flAfNvllFg0rOy0i5OnbT72e/DWJS/Tx/V4zFmUwbh2iG
uFZXs+o4Y4lw4EcGToTD99+AIsDqFDDhH8KCZvWKS3dH3YqGIx0R5Eg+oBgYOw8DXNJNGwUrQaLU
oXVRZqIPO+XCRVgDdtbruqJKsV9WYjwHn0CqakXksou7HKW02A5qpB5XwkyrsUS/wTQHK4CSci2P
L3w5ZH5ay2PFHurlaEcOU+UBwxPRMzGpKa1gcSnn+yemG45+6JnUoJTXR7TJXZh+dFW+FjytEDAJ
oxG+kmHpIl4ttiL4TeSwDQIUCbhMLlH1HlEfk3jTpv+bjCQ6LmSVzO62rgQxx9Y3jSF3Y+xdXjn5
zbtUXN4UKjJRok330Rpx6qhk4//b9+xqO2krxBdEmUJsgnvIaOLSictaMIssGMB8nQMOXmk5H+BY
H4eS8eo2Abb7LiRMaSCcKsc0UJzhHkAv47vrkEZnt8GYLQB6SzwADdP8098I92K2QdpVyqSjHnp+
fpdpK+hfSJtp3iMfati/aZySZ9cNCJ/6nPbUO0HwRKfKsRyzau+twmC0didAFUJHSvfV8srE/jB7
XZkstg9te2m9Dx7cQTgduwbHKmipKMaGZIqJwqv8g6bq2Y7EmPW0b5VJhRCwrzqV6Q9F3hv2Bhir
wb8hS7Q8mMXBuAjPEwSdxRiV4x5lI1FP0U64FQyO+UbdInBPENRI9iPJ3Oeq+Fdjpft3LT/kzXy1
BZ6g7Tma2VWlXndyrSfRAfhL8UWhpkxPmUai+pgEBDso2Xg8eTen9nsf9XaFcpHiDpRAnbGK24+o
22daoM+19W/18njQeVqPDEPLGeVeS1wGrUdXl4NZVQFe4PI/hMNy1pEmI5kKvibJFO1fXwTeX7PP
cLofjkKYjOJcdp/jYR1pNxalDzobPT4x9T9g7313BQezlqlVORVejmR04bbubp0fEWG+CVGWpkdS
taMRlypczWwCzKaTDjC6LK2o3SNFNaZyKQ+gLSHL0W3vG4mubw3zFyElgRFgjG9q5QJoi3xazZvt
QUylIaNz4I1EbfZg5Y8xodEPC9Uc+xC6Y1+JiN9oe+KoMnUdr+UhRAMfNn3d1OJx44PpnpLCq188
fZfRnHXaUPxvNsddZCCt7DMjxIfrgvUyl4bQu8P1XZa0rOqX8CHSnnA4Xc4L53AeQJCLwm0ZJhB5
TQYG9E8CtfganFQMOwCBC9t2RbHaXV8xiubcL8pbxrwtUtXyNuiLpPALoxXe3q4lNH5H6sxuNcUK
inlhuCJwMvZUzA/eprpXfAlsagX1buhK+2SwY2gH4TcB7lnB2tBz130qrQdCuZOpKUfNBtNZ4ktY
vCQEl+pmH1ECJWLngGEbDEPVCNgzb+7wqD3vlgrCgLKIq9Mya/RA7ZYWykSk86ynu/QEyp6o6HJm
fdnCc11CedmvjZYFr9iUBPSw3JTM7spYBKXgVz/Zvbh6RNcjPl/7YxKqSC3I7mBWO+h9N5jdUy6m
pZUYx4Njhxbwax6RKLpsp8x9kDxK5vQHEBWcOnYWQ3kAw2oRmJZKOJHK3wEjUz2ktVK44dAzgRrt
r4hSSUzs04dqIYahQesz95mMukWoUDvieDEiKCvCjYyYt+YX2Vrd5CeB9VG26Zc+/JhSpfsgG0+2
kT5XzAejxBsq4T5StH9AX7oHpHZxGyB43vOLikMGmDZYnWs9WW7FmsKXe0dgX/MIkElOSUo3KKGW
Gj6iONedy8jBYTAaxWn/VbeGkNgesWrsUkDSeA3CFd0W4nLoT5XONhgGhj+I/SeY9PSgOjES+qok
5EnoqGg+JwZI6MI9e1gcs2DE7dQqDfKVKrx6SrAGSsxFdI9zF24lVGrPLstH3DkF/l/BI9j186TF
JFhRfERWt9vAG7AG4LwaiRZYiPIxvfbK507jVPw+hIrFPhVHT/UwVZlE2oiX6JCMdNPsgHDKCtmC
wIOQZh548JKggDmycKJaH498IND0IeOXjuLaXTfC9goSm4kDSzI5zxQbpLZMoWLyAEyovACTOdKy
yPMiD5iKUD83UDHHaSNRjWnwE6JhVC+jqJKU1VLNbHAgR70J9tlg8mhS4lgcXJPsLbRnnJuvjG2r
tM4xBLA6dcCVA3naDu0LuWY7/9LhpUiDfjQDejkMibIVtCBqGNKRymgrS1OA8oBaQkFK/AboHzOZ
Xo6GbTPNLiGD95q8KMu4kt21qBBU70xCo/njTSK5cdsTHWQ6I97T2QnNz5/uJbXNiqLTpyZ5hEHo
xYj8HWcpNfF5AnJmb0pWq9pgbCl6N0jXmv/+hckJ9MgEyfqMUOvoCGYysFhCaiR8AK68fe/9fHVU
k3ju1DhItUEexoRkHWRyom2Jed1kGS2La5LkuNYo4UIiUM2jYCsDxAzQWMoSn6ph7CV4R0fIiRjU
r7rt8jEKHBL/0emUoV+tSGPoCPQp/KM+CZkTHHsWeOENdoSy3Htos7LGGlUJz3Tf6J9Ra8XI+8ij
t6CXGTZUnbc9fZA1IjvbykYwZ0M6xF9Txq4RzJRsOt0A8CfNT7vUS+ZhBqGDF1f/SAxEU3RQpMtS
EGTnjZqVN1GGzpsqI1VOv8VvBfNtbf9pZTUU1FE8iWRkeXgdsNSVCmPK7UvKjTaFYEM5pkcq6qMq
84UAQPsIY3RJq/Z9zrUHBEYER0sq8zzgvBiAJdPISnJgqGck/T1xaurrP/4z+Il8r8AKl7QK9oYa
WCG/j9zU7M8zKp9myObWrUIAFirIaoBCk44a5ArU95Y34OEg1HEve31VgTilAlLOQfXSCOMXT4sX
yG+/6LK0+WYdFP9N2mVu2hQfuDyLK+qEzIWvupiXqLIj93eu2se87fKFsdqGjSoIoyzeP//GH/aV
ezn5xwr4onLgnhWlzfut4LMKZexqp3ns+PP8E/psT8+eLfZDmRHqINWTMTFILh38DLf7dmMmEZs4
P4onQhyGs4DOLy2Y7JNR9CbyY2BS4XFRGZHJR70edYScJnCTKNQvlPh52Pxy4lhIRO6nn83Vs+hn
WUN7R9MB0NKwPW0B9Mdco3sx5yL/pPBlxoK3KZL1+IDvtomXq3W/2k+YhKon4mbNwezsJK/DVY4s
0o5qjdJMp2eQnb40qlViUwCmJrryyS03nyFSAyqi1UiihPol59nRATfG9WIO3dLOCzMXcq/FjENw
aCmf6PYkFPvVPAdA6uKrWN061+yrvFcv3d7ejvUe2izZ7PcQPtRRWzbwnI4VNxjK8LwlEw6hPQTz
OcgpSydz0NXNarY5lfftV6r6nQSmZF7t0iD4G0onxulURFLBByoZF8e/R3HaqDZtw0oKsO5CEJz9
iGI7kKEXO78hHRc95FQdlE7LeMVfgagPt9zO2jzU2C6i/BKR4yz+QUFsVw5DQNvyYT2z6mOkkL5A
sQSnBlCHpTWhTvj1+qfr+tg3CIfVdgvRnrQH/aUE0YUSEChaxAwOjBIr6+KOIgVRfn1dci87oJfK
6FuQDJGIF+Hfe72tUxySpGufGQ7ytlsZf1tSYfCZHyGarv60le+05ekef3eM+Z7B7VVURY4KxlTB
emzmgukf51NBTSpx5/RY3OyegQZl+8d61MD1d7jy6o6ioccrBnQAZckQZ46isPsFp3Jw+fLJROHe
KmM1mhFwKX1PkykDfKn7O1T4qpGZfm/1MjEO7Kv8Gns/Gqoc5iXo5BIMgIGzMCUuf1mpVW/FekNA
s6fzERhEKGyVXs6uiVHL7NA5InWvyDO3LRv7RS2KFA4BKKbfCB+DG1Ia2RunOa9sVNHWoqB5fYt8
mZNBxPossmEU2MxWbRI7ELWQhDv0o7bucJNgrEOkgbz42lak8ldMQs9RoP5QIi2IUubbTFR8nOq+
3K8Lb3sqcqdNkD7tyrVJnuzY1MqTudOfTCJDxTG0mBeRWK9qGC4MX842SNvQM3FqsXiKEXrWV2Zc
3IV95X9b8pkmNSf5RLcFvjF4/izzIvTJYTbRxxR06jxIRRvXnAlE5jN7F1y0yTE03aB3SNCkYt3G
Ldvd2qAriUC00K7T82ZzDx0i+iVAxblbF7DJS6aZujy829icgSATbjRmxhZ7wzCOJdvC+MNqd3SO
lp4yDoffjG7gVQPNEz237nt3BJIyEZtFgla4egTOF5KOZTDNTwvmALENgr6VAgQvY72iAYKZoB3b
mUmwrutF1FYmWdQ9r10Cf71wYv/4B1AyOyLvsEyCY9PhtD3J2a5fOSJexxihRoncOwBq2sdjSmFs
gOYrVTU2SKyMaSwpjlawK0UsvannZi/eVI5//sdVE/7zU2qmR5gIUYxxAoA9trA3o2FOa7KcdPW/
dc/N1lkWJ0NtfhS4sWBd+kCIN0qNfWPQENEMjx4J2BjZYmyb2AK6+qr7OGeYrn6QbgkCc1kZ6yfl
vzXFMkup5lz3hkCR/R0C6zfQUGY07tisFqL/9kq7vEDSJb4k6b4QEz/iUE01zvyHmSoPcXitsXhU
xRQINqguFofC9nfCwhSCUsirOSa/hZuOafhk71qSt6D7EES/hYA8yD5X9bo9hpRBUY0Ewz1CJ47k
8tkH/fNXT3Z1uTqq+ekjKMi9k1IDO/0ZvY7kFzPknngsfRUhxh69xvJg7RssSKl2ABY20NsEX3TW
aEqmccK0LF4qsD585JwZTGjVumipvRaVF6ATo4fr4oRyMtqDLZyv7nzUAE3b3arW6B6+SdGGJRDU
Mp0hC7HM/7IU1KZKr8oGInbOCZrKpp6gTP0SjAf1EHKiWale+wwDEJeJv8kZOipEafvPl5iBWiYV
qnVroToG7gJm34CvE5cdfZSUEQcXNfMyQVNGD8EM3HBLqRFlLf7DG+1eMu7vk8S6RI015Ffidhw/
M4M05u+PyxSQ6VrzjOoAbR5/rQ2KNRUIRAMKMMx/IjA0diEUJBr2ZaUJminKPGe/GV80G6ULZlTg
QgTgNOaJdyDYJvRNZqrZu5WZePEKR277zRQyAIMp1EzFuIxw4spC5O8GilpHaJF6TVTY/i9argQY
YYjHSwvPZkwV8NmZ5yjoIkaE0JtFa36Dm2sPc5U2H+XCQe2QvhBTse2gpCtICHBiTRm3tVMzo/4M
G/gbWYNxbne8C+t1J9zGxtKhutwiT4SKx9mygufg06nFJvgrAToGAf7bYh6TPJSGMHUKz0t+OYFQ
BENoCflxA5qfv7dvGEc77OWs2Lz+r1wHtWQ05C1UMrRyjJl1eNw+8/bfIDbIzr0lwDrjv2fPVEsH
tkVwGXS+n4VycuaoZNEJrhn4mcx1D54BHnSJ8T5tnu1yOpZBdThqSyyWr8T1eF8so1XjmgDOLUrp
tvlHYBuQXRWUxkdW1PMwrRmn7HvUiv0SYPKBRhyumX+tSknLzNoT9Klzg/RZz4/wDH44A70jwKYf
MTBZL+6n+boy3vfyIugpjDXzBro61ge5ipF00haT7zNf2La49hJI2Os3XNpfzxX1UW0F5TQqyh2p
R8PezTIIJ/bUW1ZHdidCCqchw+BKZFoCPHKfSRKfN+QkbGFut2rSfe42hgdKSVSgplebiwpMxgau
2/8KGKMCrmcMTwGwwZ0oUJk6j14KVFOzn93uB0l9ZhrU+RDHBsjBo4DYh78wj0FsgDLMYY6FyG8g
qDdqeUFQWCgx81mrpzInIjtulf2L/KDrkXH7QEUsJ0GSaH1Bb6NvRAuxGGygU2wnlwfpkpBr3pNz
BNFdlZp3rJJGA5cIfSFhak4sNgB3gKn3rGs9bzuiSNsIIIXZ9ETmfJ0DKHQRV2nN+q869T1+DQtu
SsbAlyaOSim7muQAVRzmmX3zp7SMIU+kBAfmMXSIPO1WwAPlxBlbFwEWVcd0s+jY40FT0XYLZbPi
+aJhCCn5yAWTUS/OglyjzMjp/TPEs0Ccnv84gmCSDpz+cFmeZxg6XObNwEMPBhMWg8NkJHtSCaAh
ZBkBn+3sQ+o5NtDjFk1hPVhfoQze+1wu7AN5orlOwwG7fZ3PWxTrxh/BaZLcR1R0iMClsGHQHK++
lpEKla/VPWNTweUy88Rz3K14Q17sHpRK6Tqo3CyIL/RvRyvRiK5oek+1eU/6MI51sDU6XWitl5YT
U/I7aLi5Q5g/pl0/NoSY1rlsHOPKE+gv9RZ+5nzWVP52R8HRGfbMj7i9qbOXrcbjuIYy02dCwfCR
GmbGqcT2l2DCff5Yt6DoY83SHv8OokTsoqeqJ0P7f7kIxPdCFaZw8b97yNt4Eo8SrP9ZuNRIXDrp
9pqRNUoHD9bosBoAsRJnRWWBTtbMTR9CLrld10F5ahhb3lz0RihWbKBjjDtcdXS9s7oYwH3ALyeB
4tx+Jh5gj5U5A2bX3iTNaCO3MkiySatJ4B78UAzZ7nndi6gL0H2EDLGTfZxkYSeBXxRTjMzHk6H1
sf/ol4ZdytJObbNlBY6+HIQkdkuAcgqTgOuMQx9Wwc0MGtGekViKExAhQ0Sntjv14qvc0k6UnVWL
fdhQiLVVqql6L6PiEDWgvtXd0RPaV549opjPP6x9DUgVM0UvVcahsn2HQ1aAtnCIPLHDMXsSI5wP
pCyxqFPF2HQofoWlRR3hmOH+adMWgq8unLqUNgbSPWdwjyHrNcvDgSohpq7Qn1IGTpduBRWgWHAU
e2IEBrQsYJltBXaN4I6uQELyWUCyKovoSA5V61YQ9+9lxQE4RoVaDWiqDf4LloF0yZpwUCayai3W
cSKUNlS9Dt/PSYOTel0gtlBIYRj3Lk5Aq+SNTlJC8p7n6Om7ziJCKhiWw2Pc3m4dR5fJRY9BAeRR
Lwh9yHg8bMfHhm8tV4vRZjciaRSL7Da1rvwozgj7djf867NRBEjpPmrOasO+wROqYrx+h5nJC/0b
EqK1siMmIbpsISGGSn7WCeVe3+8mDEcwx/xc1SWN+McewUyfGHMi4PjZTmt2nJI9NaLpu1iwQtvr
auUQ4GXSqrq2LyA6axt9vn64rxEEvuCrpmwr9rzi4DnctbKp0HOjywOud5hUOAlVLxfsqhFzKoMR
AwhPicLkcw2wwx0E632Ycre6XWNnPPuv+JG/041ElExcEtYYL8UVUff7VWC8hdK7o3kDz1fIwjZD
J6vPBOL1CCy2ZPecGtPeurCfstkIix7/fUimmIYxSKG45ONbthWLNdXzSg6+5TFlyvahKJ2FQrtj
IliCHvWGrEpSxdg+GxXy+/JYeWV11Ch6UxoGHTBx7LFpIBSVo9HcogD+CSeGlGoWP1RLDCZstkSk
GaVQf2L8elDm2+Hv4Ab5coQeHVksJWLVROlHfkXNf0nib6Wz4V1gj8U05gm25l9ix5SariwsoNmg
fwN0xLJThc+vEByNvSim5uylpn7Qw7CB3A9ZosQnRayYRs3quRyVEd+YKcvCDALRcR1UuFpz4Vjf
StCcm0CngTfUfbT7OjHqYior58hbSH1B80PYTpXq05mY8UeZ9xpXqyz1zfInmZq133C929bYMC/Y
fLBoqDW4Q9TQJ59c/7JHRL7cAPglxV2izI2nIvIMJxBhjSCw7xg35APFfiSW6b0lYUPnP8Iey6Ze
Ubu1hpYtMnqi7BwXDxi3/PeB3FMXhttpVKU2pBh6YHebLhwHAB0pV9+BnQGz+os9JzgEOB/o8ybN
ySN+W1vGY/0GYLeGI/1gn5b3HtV0YSuIHRNONfcROQDtygBAU92REbLqwiRw2HBvieZsKfek/3vC
fJqdcPYz1ixBbo+H0EGtf5UV3DQXuoSK3lpu/TVRBymsKBxZkY/0TG1u0Vwez6sDbJsPj17F3Ft7
Si83MnTOzdaXRkZWBLPAO6cqSSDBCybOQigcCMFNVfoLxZeWHL+d7/FyhU2h+iWHOheVekZpfAfX
hYob81dD1Ow+2ETLI6hy4ixwFp7EUFOXDdgiH6ABWozg7v0gyE+0OZNBYUH5A94XYAdRVeeKrUL3
jZloQkgKTE3xVWIMi/CqAwAmLN7j9zrUiGiJrwhBhYDkg6C6a84tDFgbSdd/MYAfXQcTp4ZsUiuB
ZYHwJmtZe8h3u08tguWvDJgGftALe3m4H5KNYjvjbGIhcJUp4yaomLo22GQ2nOwslVuEhSX/JUgi
72WeVI7BTfBOmnV/9PTWfraO2cHxd5VgmVUo0B/Gq22uDkkyegi6V5xyRz8OAqCf/46athMU0HRc
XEZ3RI12YefHPA==
`pragma protect end_protected
