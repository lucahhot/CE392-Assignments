// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
XXF/dEdobqB5PPg1d8jTk7YGQSMyT11IGV2oDuCCxPMoQBFUx9+I3IsFhee6aT1aXQE5g8EHL/3b
Y1NF3XSiXkCi4sghfm+bsefi7HfnAPyXjyA/p//MsoaJfZPLOTWutFRnu2IslMdInEsaV5IJ1SJ8
FRx+au0nQRhiMHDbY890tqRxXo9NXc+az+iB46LfOcT82IYaNkrnjFhWBsBuqY3IqsqIUfV7gWBZ
848B7b+eDPGOCDVqewoXTMs9QhA9MX7XJe1s6F5tl5/558pI+8DU6xe5eN4F+mtaTCYNLH6+fc3r
Eiq+qYrb3a3XPU5Bo5Mq3GuWHzrcQKC9AYa/Og==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 16288)
/+xvs8V6bMV12B5LTk4qvoqO6goM9sJ0EFxochv5eRTsdRL45RKOqeHL2EEXMHYAQPSLk0q/Xbrg
gpw652BjNOKqybY8cHwHG3mtDDelPF78RmUFut1kGgWVstkoNeGEm5mh1UjevKWj2t4bhT+qDc5R
mpiq2VNxIpZwKjfbNqrGvMeK4aoSwzEY/csEeU41oxIcB/PfiND9y9oWxAIfZm87uTPnK3YEpPqh
LyWT+c8qa+evXXtjUeom1iyfX1aC9shAqUewVX/Ci6eN/0d9R0C3VousZIT1OWLWV5k6+BSc1QLd
wOBFBrWJ/QQCkWsmhSbDHwKvBXAOBGrexSf3mD+fahmB6Dhl2PIRk+/MX28jOS0Svr/QLESwrW5J
7KxK1lEU8UcuvvkH3WtPXgmnZpOCcbLCrf2nkeMteeo8Kii3geg42P+C2jc2QP2x/OkpfRoV2JX0
ik8mQRtWY+6CyUsRhIL6Zb8rt1dkvfxFQakwO5uKQb4jlAJrxL+Av5gK2C2zM7aqAd8xp0Nvd9qS
bQpS/P27Q8AkoHgH1JoqQ4YMbXNyKRYQ4hHe5p4IPjco3g9FHKeIPaClqIbMgRBa3ZSVJMa79rua
UhSenJuYNkhq6h5QzVyxJtefn57PDw3VRBMoZ7RuxtAxPG13y5dIAbs6ZWVTPjCYT15whTAzyJhf
jUcJ81QZewSpT3C1yinTHDWjO32CzFClvxYq0Lp5Q0PFLqw5yd8UVxZwoUcrsXpa/nqyOyTsIuU7
9Xih5QDkstuuuCXKM4B7eUbNDNOlA5LKVtr0PglR2W5uXS2JAqSC3lFyR2ucMSFcc7tND7H8H8Y6
Gmh3kyxxAyKL81uOiZ5WgmpzZfGSJucnKzc/Idgf8FXknlbusV8Z2Epc1ig6ZZ5PdpEB6Tn2ueDu
oEej28tBUMET4fxs/R2VPld2vKT6IE5vy8UhrnhfW7Tow8ujLiGKrVl0eJkqw3oHd/FCuDTFusFC
GLxKfRLC8++Wj2H7yLJFlGMiyNOGHJ9VbQ4BIPyeCWA1jSKNQUfM6zuRau0uNjDq6ZgNNrZej0fD
Q8tX1zGzDcrquWNzN+lYuBmhV5qV5hNJIwRxH2ExyR89QLehxZMXeKyngUU+3Tli5j1oG49+h/DJ
rXiFiiyqF9PKUiT77VJ5SNGRp+nejdodDE1rNQs/EaQ8QyUT3RuAKj/1S4eZQxo2oD/C57tfQ91D
D21BAbodh9P+B5kF7zpHqZfk6GV+cBB5MK8+x/5K5fDZkQgLoM7pqFhxZafB4phxSN3Ns21HKvR7
srC9HAJQvKEinLsiuWEkYSnH0uZrn6riZ36WRAPEVXPGfef+5SpxtJfmKMKpHMnM4luKUNQXb31j
oyqY4/1zoa75hOVXhZaSTqgjSiKV4nPNJ0SxhnZCHLjS4/IPY2bRihIoWeoTNLljJVyxr48MRg6N
jfbKVHru5mhCOxvgfcWAgCkVAV+ESQ9ZVyVlFBbbt3x492QUyh5srFTIQSuPvvwElLImzo2pqBSV
ozLNrZYnsyx0J+HPzYG6GhlYvVMMvzaunRLf6o6oVn2YFVd+rDGi8Q/92roPL6iqSpBSgrPwlJl+
ZmfB+5uDoYyd9Y6GnWn1ut6dx3GhrZjA9VASWt/SnNrR/3G3fRySpYvyOpj66FFxLOnPgQicsmQ0
WDaW68DJ8mVSMJEff16q3puuxvQYWUbwLvk8ESyf8gUZNl5jO7+n8Pekk79H+DwzX7pXk0ePWj5P
6RqmD7O3dosnu5Gt+CkFHS7AkwNfoHht0Q0yCyqpSyNVf/994NqoAGD4yxi+hVYMRPjUKvgCWt14
nx1NCYoGMaFRvDROVwRHcHhyF8ohy8C2BaLxHlxd6F1SEnYPKqRa6j+8SUO/n1xKpuT7EC+leZ0N
DfUeRBq3JQd+5y6ccl/qsi5errlGV5aU93EwHQpg/8Q9cO5Q/dJrsZx26TzCEeDlFtMN/k79F/Z7
nUEDhbk5diF2aKTlNub9xR3koAH8dmY7XvyZ1/ZpmEQVbn+iqm52tXm8nf/hjJ0C6sb7AcC+Z8rX
6MymqsPCbEa5twBh/EM1M4sTyrG+TIEKuEEQ4DAtrJ5z+XGuxf4VvY8QAkdRz4RezYcwA8jmQBGr
bn3etiC0Fp+bcFap/5lMiMF0OjvSUe12cH7T5R4K4QCInW+mlWkIFam4t1e7LTmnQtb0SKeih4J7
QWGneq7QWD9QfMsCUm8bOExEKdDl7ez8vnnRLR7U75LzGIa41+KBLCvzw9YyvoJ+n7PcilaxW4wE
c7FcFTKLAJufvICT8Y67buuG8Uw7JuOYs8Q812w21uvwSx2+P5Q58oNPcmwgPZEs7GP7E9Z4afCi
mIMEYREssIwKF6RtPAe/LkxF/bDGJ27hfkosrh5AOJ+F4UoCsKp3CBW55tXAxpdM7Btyl8BoikPD
2eI9L5KecBzzrh18h7dLmA7XR89Kn+WqdttHGKt9PYS+AoIE/eF/MBOzEZbQrhX0HBAcSz1WKmiR
dunjYhAv1j/ZxgSmo28GnaHfcU29/CbsGkcX18jO53X5R7bWH7r2r8ZRmPXz8u0ykOQdC8M5oBS9
arjUT1Gwyg9ektAqhB9WUNMgZPZL3B6KYVV4/fPus/C7NDLPtoUaRAQxOMktzEL3yhGVZkVYvbYN
uiiakeQ979m3GKw3rO8V+tCniQNKx4HJV5Awc8Cr0ZFD97BDzIPAMd4IR7mBkG3MYG1webJeRn1Q
c6gLoBYQh3lhuWNHq8UsDYav8/Xmkd+1IHAN2Qrz5Bm77q41C9hqQQN9xVwqHpClC7HFe0cOiSfw
Yy4oGhjdcEV4EEQcpMrJi8jdgV67QCCHHZd4QGkE+Z1i2cz7XsylZvo90QSFwNZ8ZrZ5gdVD9Qvi
1F28T/qyDXHZwhBHIry81p7kGa162+uss3HHXiz5jbM8lgAlaUcqWRfkuvxrAjbX01nGtKmFI+uO
Ho20GEWhQNq4fV7WPMlz7xAth4C68J6QErN+JPH/XyI2Lk244QMp6BfRcn8RF0J7FOxTiOwfxgIk
9itBTliAJRkUTJgpkjB0ryLU9X2Ze9667wojT4PC53Zta113m2ld6/sAMDNUu869214KQDprIu0b
FNlWHEegZxGrVI5idiSSycOltb13sse/1BJwCtW2T3a9ZzZL4N0XjN/oKaDjB4LiQC8IQj39mu+D
85zQK6Q0BW5jhJYXiXlHZVFIL5UIthL7L9gc6Z78ZqSSS9PpLGvfTI+ltilbDYVKZ/XU9Ttxmb22
hYYxahaFKAm5om4uz/hS3bY2T+1s6L04kfyubzJjqEDxBq4+oj3LDpDyRdk4y0ccNRwB7ATXwQzY
ZebTIRKKdmHvIQk7JEM6AjUmdRiksZ8FkNN040nTt52Upc9SW2GR+Ayb4V0yEEd3yFQE+se2CaGq
0Cgex1yvu54lblz+L/J0zLxaHs+xkIAxSHmbqjrKbP5J9pnK09J7kFQ20QcR5xReh1g9ZjEANLL/
Uh2mp4GmBlxSip7XtKy1fMm+y/G8CNflOvU09bqw4Nf9cH8lwoRIEUeHM9I3nIjcm41I1sEhlnce
DVU4XjKOtcejhXQvrXAUVyqZGIKV5UxxE6f+56XZ30DQyLj8hxJ4G4BV6K8h9ixas0pFj7oYVGsh
HKOSPx3wSUJGcbwXWCh8R2FjYs7hzKwUMijcW06Rum0GyuumxMmMxqQ0b8a3ikpKOVf8KPyO8kQf
9bq56e4FPTAUzLAiD3q0luQ1zEeEDsNmTKY2jtVSzzwc1z0aKsoGhLq2FW8U0+Z/xu0szbYLWPid
4iSnov+emGg4GFA05wWLiDCAnG5zTsz05RHh/jXLl/03zG3bPd5adL32l0FHLpXeOGpfgetFqymU
jNv0j/Pl5eRSZxOABD257xOI9JkP5qsvM8xRw5peQAjiWM7lyyc81uMSprwtp+X9ceEMeKx0K3ME
eXXzbZCOORAZW7BN+uNOwsVrKQ3TmlIs8Z7FbXzSIBpR1QMcxH2UN/KKXjXsK4VOFVE/nR3bLtwA
/BPP0DtR+4HQUi2QiI+86lCjbH5c94vBqSDuNYaJk7Kf5m46QP7AsXcD4aUQLLZDWdBRLWR8OweO
so19emr5T4kxoo7jUK1GweUbFAllMIKNgy8Llkb41lh05LNGxe8LVjAMOp+GVrzRFmnoMNybduAs
DzkNyv9vA0k+S2G66Ydl0M1nULSo9cGBPyEJXs2IylcYNr178HDS10UhPBLy80ByofJnQfBZ1Ndn
T/5Z3X/9sZOux/y1kFgFCHK9L2H5O97zUo3QDhJ4KZ8m6zWCKUbRSQDFdjziE5gEnsoHvWo9TU1S
vB9sXOoKTgjKdEljQA8sj3Jm/DorS7ODsbRe5Ovd94ofxiJTUc0lOeSyXYiqLzDMwoK6uw085xRq
AjCXY3y8HNwyekBxHdJWlEGMgKJZvT75CXYJsq8dutAKDnF0yJ5r2qLHZabme4m1YoNzmR/ftatr
9lt6nZkhff6muZhTapw3RmPUWTu4YUIklTBa0KDuLOpVKHQgoY6rt51cFY6Dky1ss3c+HH3JJTAu
awoensmlZDdRKcTqig7x22zLBfTROh9TySXFtg9omDUVLoBtLCS2qPex+UVqC4FFms/AqntjRoEF
7/l+AX+mcGU092tUN7jWk4td+waVvkWeDndnkBxndXEMnTODQ8dvQJIsC7FdXJU1YqGfS6B5OInw
GnxfJA6AdJ3TjqtLyZCjj5P1O23LCbaP8KAe7Rtc5pmc+dpd/SHktv9pzDvQJ79UgcGOONnJ5jmU
kTqs2YRX78VYOOJbiCFSOgWoubF/KNuPIMrf5I5e8AfE6iTwF5CCwlJzXQzZvoAsCMndlyGCVZ7V
NSHuSv2vqXuhRRY2Mp2UAjAW4VHdvtxv2VmglZubjNBq4oOcUs26VdCTJDNaoLZqm9VfQz/Br+As
Lyv6SRUfk7aSBUyQyqlUm6KCiObtEaAnJkySURlJpXNTGmW30sWr+ddHirKAQmqITRDBhtYOwd8O
mJ5W14Ota/BS2VkJyXkhHvD/rnkV8lmyxo4lYYZubSmKvJIt8ogI9mzaf7zwosmoAodSDmV8iBkf
L4KX6hTkMqFQskXPgvByUWjUSui+FZCMprQr11jH1up101iTjMbVdX5bRE7snnuYEOikiTPiGCDQ
MZfVmwl9ZxqnWDNutjt1hJzaRbAUs39+utVP4lY/yArm3BTi5LhUZUL48hnTK9C7e/QBfLwqqPee
QD+z2CTSU2Bm5iVBW5FQzIkkoWGUblvikZlCtKd+6R+95+WzQ7rrl7A41AdYGIXd4Zc6gVSlLHX7
7YNe1v3J8yk+5ag+/UGZS7da7siSoZyM7C6hc4WZUtuESfRAPmu2q20EyMteoPWt1ECIyJkDYjUK
fyxfkAm/IkO0sXU8xua8jYCdFY0gxRE+BqXBFENJX0JzzDX7nUEvdGwzDLYPuCqUmv8q3MF5uYNd
TaiMBCy7IKUG0dfdz13MK8m4Svc0znDhzCdedyg6Ii+4UcNeFX43Q4ieK+L5s3Yz2t+N2QlZg+nU
GTJoYq31r0dT7Vl9hCHR8bPuNbBgPsy3a3fsmxJ/yTqi3Ravzu2k+ISFFoE+A0OcgSLG4bZ40yMj
IeSLZu1oj3N1okyLKWpei38l6rQE+Y1tv4l8KSZRKyuILF08Ys4Pm1coLwUEvTNCAVyINa+jRtDP
WneWsaD8ZnrpSGTa+WKyYWVk3s3wN/xrOyvby04/2AlK86pQjAn2JAzYakcZXkZsye8H8SF0gIU6
Z3mZnRuN8orlP+yodNzspyYgfWW9T3x3Oyknt4Ufy90Yt1i/AnLz/kBnT5NCryC73Q9ccWB8gZOw
s6x4iD5en5vNPS6L4QnGG2CVj5UyYIDlStA3SHpTmKn/tGJIXsr1/b3hhL6S+YYkJCI8LTY8eKTl
N2oonChL6cy7imafiW1nElUDIhCtq+XTGc4aavfyiXUQL9pbUpsfxUP8E1YDckLYP/0iZyNAwAui
Fbm+lE53ETViGCb4M/c90rlTUqURDVmA7YF4cuL4tsLf+hMx5bQfjFz5QEQRdXF01BGBZyURWxb9
i6Gq1dc6icJF4oC5nrZTAIiQRytvadZrhaPb0O1VIMguQbbKu6Mnw/y9nom9wyXO6DiBCnmXsn/U
Ze+jFxxNFWlAkKhWp+Di7DHAhgdk4TGOeFkcvUZeEZFtfDFVvP7U3dHI8hw5znIcFsVIKNumZmQR
fT6Of2jGQTve2SC+FCty5M01SL90GT/+57nrnHiW7PbntEldf1y2XbwQCufjv6LSlEKbR2GLmWLH
6BpPueQHmymSHjRSc8km2+IFBwIt7NN6hpEE8rdWXrHmGFYZPzrz6rd0V+LUe7V0F7SKOJAWPlyX
3Qy62kLzyhtmuyzEILr4mj+mtiNGShSADLdho38wrQvdPueFe0BTRhtC7leReVBQ2UR81LCdEQ5U
HMIh3b2oSi1Mc3hN32Lyv5egBsOBnaVa4c4L3SCemukGXdrOPdc7i76Tg9k564xyq0K0PYdggs+X
s/eqkvdTaGXcItrpYkGjDMSsSCbmLVn6kMGWmPI6q/4u+pvWvM9p35SGQznWUDwW4caTtA9CjJnC
bS4QhX8v0vmDfnGej3SkjW5yA24OFodecjlc65fQI67eEJMXaC0frSTbH0pac2gXTItzypWpNqQ9
KdLNfXkELl7Da3+XiSdRNT3p4YT1xeLX8dT0VK5GcVbjB32lSKEEPY54Ly7XrbZIQY4G5QJye40E
I0unjuyyLB1WyoGTccZgqYQWrYBLC9lp/RrS8KgmJ5J8ObWnZBGYVGLN7GYUGaDGgEE/f3M94XLO
gRN9mVnBrL/sblbTW3uKnmaBQh2D+tHGp1WBgaC4t/ohEwvlj/eSUwlpS7mWEXP8ThMXP9IR14YH
p3+pag4F0vahx7GrXRXzhq1xWFPIcBpL022dJHvh6aYB1/S0R51ySDETihQeeJaVSAGVIA2/mIt9
x1ftK6DLu8+nDXODM78+EKWfhsGhq89ysfZoxO1w+JzytVB69DbVakj+plbgfuCiOveOAPnIFpT+
AAmcpONrKlu45OY8veM38c3n6JxWOCgN5pH3L0g24lFkZWtCqVIwiCxf4JUad+btbml4td+jC2ou
37ETNcbWvXHbX3pN24l7vh17LfKWnvkkhO1AbOI145O0W6Peyp5J+fa4pEiVwTwcfrr/LVU6I50j
0DAVJNYHxPp5WytnNVXf/uY/kNSYPyjKx25DWJQBzj5Jcw1VaI30JKomhTgPgN39Xk019oqk3v+9
w0OhGPZAyXyNCg0vfRQUJnrqFRhWFgqJ7lJOv0seukaEdXhsJZe/bRpuLxzpx7gk5syW7semcBhq
RY1BkXWyj8VEBe/KGMAwHfT7lvl5yVy9VB/qT227rcHDgzRVYJHno7NPwWWnTfF91VVuhah4s7K9
P1HZ7cCpOnq527y2hYjjMIN5yL98KDLLQ2l+K6GUKtFjNG5/kImkPXyVhCY6GaxgHMvL4Nkaih2/
ABhQ9NgAHkD8CnNTP/RYOek/R9e+gy20njwnKRb66ReArXLsrJSzXJXtjlJ76Re+1X6D5Sa7RkW2
WEM+D+wOVCsU3FuwgM092P04k2wABClNZp13tdRcnxH3/UEF6Oqg0mHCKLZumkYMxf0vhGXWQ2II
ljt0zPEH6zCckg3oOe/bu4Qb2LPEUcaajO0CogP6l+g89q8yOcEO3+r7DdMpl0JA257sauBv8xI4
UUmSUFl2aKXGR6qZUAMsWC3C3w/wEspROYcL+4+o6vYvHpVFBrQU4z9YA3MVatv8GMPSkp8CUH6l
b0rJ548Tmnpb+wruqk9hKfQMDZCxxfa/o2kxpbxEtwULFs0xGEK/n/qumvO/VLfIyANv4WXI4DMH
e8RYrxtIl749qnzY8SJKQJ9qk0QnxSRAMOjP6E2yLypWhAQAPL2aJosbdJEsmSxrCEWlr34Vwblu
IOjAg/kRVfMG2arv0MdiIVYDQvJn8JBs1LRurNktIFRyD3c82+QrGRKPPZyRoXdFRRAcJkCckWCj
GUqn/B6AfzMMSQysFF9vdFnG7Bx2bs+veqCYR3jCsRs61iYtR7NrdzJfgzXYIM7ZNLw8R7DFHJUg
QGt9pE4aDE1+6JJFMWCC3M6aFIMgAmZxzAMpROblOelQ4BmfqaqLRbdzdXfwtm5HhtpeoyhTwkSc
8igvRMFZj/PPGLQ6e1dIlkxE5+O+qL3Vt2B3d48pwjEPds8GX9PQKa2KM8wptj60ClQKHZi3/z5L
8k+1JTONR2VGdM4KoaorN1nQ1njNTtsCyLglNvcthSjChrCuBJEyY8XNQO5VDFLwRtqnCEVh0c+f
O/ia6cFAUq/FlaCgXMFTJ72t6oziIJcDMrCKTq0dt0mbaCsHOUmxD6Hw1fT1sOZyjKsNj+9QWSJ5
1IqhokAGLd20h1CecMO6ySa4NpmExsEvdVCZWQxPPPTJ5zQOXn0jEoncWw7+qAuy4rGUzORU6JgT
Uslzj8W2LENAr0sJeuDRvI7XrX7r2r/LMDHGZ/hqV8xyC4RgumYUYeQK5w4S/2PTHtX3mgo+c/Fq
3tMAiP1McpcqiGD2nvqAisAn0tpvoHkxWtW5J86DF0NKac6ypY4HLUNJqK4QksZwJj2ZiKbJi+96
oAWjOn+pnteOpX9w2E/5Gi0HJWTXDP+Vr8F/wOruWxU0cH7nbPNGaCB8/hjMIoWB+aiwa6emExCr
ypiZ9NLdhl9driWbTCHJnTm3KvsYvEBUM+GBaBt53TzDCbcijJ5cfrO50RAoaDNgDN4ntBx0AB1M
0QiVN8FRFyG3MxhutPQK5jiX60U519OW8VWFrylA97UfPSRI19wtAZ696f3HpS0uG/r65zl3MRiB
pYIrVYcKye5Jtw2218Temd8xFtS2u39qlfILJV3HmyIdWUtZmARDDX1lOnmqmacDnHN1b4MDG5H+
HYmjf7tLzB2/ktfc4H77r6SPE1fHVIfDk5HSVtp3z9z0JYw4xTCD41UEK+/eNOzHPINv/eZW90MI
kc/bf1fRPEgYEcmJIByjk6J9LPf4TWvvH911p+7es4hwmeYXc3VqlDi8nnIL3B9coeTJVyfvg2KH
5zKCZ0GwhudIIQ9kuFTrFrGD/FvQ4L35hkLt9z48J0lwOViHwYKn9wsotg5TWjPTNbG6/5KYrBi9
HEopU+d4o2frkUXaBMm5IVceJfnX6Hibj2Qy8kuUFHkXZqdJkgIGpYnBpgEZYgScD+L4FkMh1okB
AqKO1/XuFBMsdPe3esQdTuiy8Cu62I0QlmpOgBFtpHIengjNDn0gJw/6hULopFLDX6PXOcGtVOMt
dttPXvhi0ws3Rcp3+lJIVkjvQ4XmZOqZdnAttbi1DZmEOP+16wCLenYvDSAE/W0lrX0NdLss4Ky7
ycmIGrDAqaBXAj5NIaGpPJh4FC1U0uT7BHJobQHiQsG+lqU2nqfF44BMymZ7Hu6Z6Q99fpKlNzdU
5Mgm1vYz83KwuVvk8VpK8n+MQvzYFLm1i/kT2DIYafokQfqk0hEQ4eb2b1dA0y870JzhPWH/x+OZ
Iqi3nFo3SXrSNj54GtO09oTTSvtbG877bEZgvVqyVal6VodD+ZwxXktIZEbKHzjCHO+ao6lCGo9N
Gr+qJs0PTRoECSX54dwx5yym9eM0yC2KJzhNzojOmkt0DVKaVceHk4XqbHY3AooTv0bpzbBacUj/
uh4QmCdwAwIciUJmbPAroDRfFGu7LBrrCQbsvyXSJMYijDoPB6ugZgdRBgN7ipKr8sB0lvP2k+sH
61bTrsOIp6zFSxbwdlTTHIbvv40PWDDj/xjpvA/5CxXoThi5y6TEpYtYGFo0OwGVl4HhygCBGzus
ofrYhJeb15aqrprFSHLfhAyenha4Zv9K7oXzCu71X2nrkUQO2XyLPVH8YGlSJJ/g1Ig+spv9JWf9
trwJu8wLsW0JOYwhg3RJVhFmN3AFnPDUAoZH9k7YNxRjK9maCqx044Xah6tUQdzlwzd2SbkNsVgw
5fOnbnD8jx8b+vso2ZujnkQdT4SwFxoHk6o0tYG26+6AxNDEYyDRzVZ40ZeXtjDDVNNONp6gaKFT
XyI8g0o8X4C3FoKpYWD2sXDa8VUznMjrUmiwydr6PEb2tDxs11kpLI3QCavnythsETR9I/iNmr7d
DAUyR/LtXuRoP6MmrcjR0fii1s3jQ86xXJtmd0Qi59nl0EM1WRKeAWbmbIwI2sT9MJGXJ3aRSYL8
oNokZNtWByxvzg40JPtaH7nJnT4bfXKUfqPnHziD6q9XmEq5qrYpdkxAF7kpeXCtmp09Tdu2pI7d
VxenBNPi4d6mN2WjHr3ancrTFDdkKcs3fBtMx2zuUEQy5j9NjUh304MrY4zE8SUX6hZYjEuvoEAw
Mz7hPwjziArqrGL3XKq1EVfNbzycXZH2cPLY5VtE+K+tMSi7j0amrBbmTBzgFTAvV2FP+eRm/Iaf
XCLAPP/cl7I/e+GipHgiIWIfz+lRJbFJtohwCQBQV25Kif36qEunJFKzTBT4VjgzjPcqO9s81nn3
y1VqDC6HJzftcFi+QvWvpDkV/1dvHz62y4atFAk8f0uf1J9sVqBWrECwlbFEUktz6FXaambasRwc
391PjA8sjzr236ZxhaBbIzQiKPAjsIJGP6h7Nn7MvigGpak+YNDLJyBobS82X03RYhBP5hovUOZ2
NjanCe6NdvK2XlGOOQWzFnZC3ZuNwkyP1U/zEpdJbzbXphZbc504aazG5c9ORUo583iHtb73SAgc
Jz+KWsZQXXhMihegGfC1iV8h/jINJNZOCV7KbGCWaliGbltTflNC08Up0a3915efim0hyuhaf7ZQ
ctQH6bYEse+CCblzm8DK9UVD++6gKscAU6xQ8NL176DDZOvQoXc1GHKwsIuudDd/OuhLoyW4bUw2
CfDe4g1Y5bAtBdVDv1uW/dWRXNiAheXGB1UZ52GX8tPxv8pFltewFKDh8lr1mcxdmst01a18v4kG
LP53rn4fzWUl/+OpBUkqo0UBSpJ6BeECtDbShSqZcGgIX30+X68+C2QJymrEPUPO7xqI7oZ2Yn/e
9FSAoMV25m852UmryBt1WScH6ewfK0VyPKi4Zp/pcgYr6sbIVx91FvNqBAdq0AEq0/WgHYkhI4Qy
G/C4k9Zht2vgbKqUu/vDKaK8ZNHQ0/drVywVJfwm13EchwIzEiPNRCe0KjImh3P0cvX6gA2sV5b+
IAffwV2nZAf0UUXXzAKFj7jn9r3NqhV0tOwFkmP9zuDHrMWuW3KKMxWhlqo5ixnaiMx1N0T9ZBSS
/Gy7AfnBXn+I5lT/YfH0watNNvN+hu/P0KYbHUiodBOzvo6r6JXAyBnUnFv+Xx51VyPXT7ZliDka
Jug7hl0aaBk6Af5Br2W3baxO/5I/thp+3W7r4HfeQ1MEjl6zMGepAjPVzJhDt67D4ZiXddg03s0X
zUzMLGfjSFSAm0JCEm4q4fEm4MBG7spjp3K5EtardZqW2rCYPdAbpXgPAdKuUzwBZMq36sZg9rOz
jYT+BliFJjZTxeBjfX4J/z4YJd0SNiqpbN+doEyU4zof7MWTrQPsx047/aPlDIE3E/Q4cAx0lKxP
TF8LZdD1CufZVILCusm08NXVtjmA9IYbcYXos1BMB4+VhMjv4Vb9jsbft3vzWrXbEsR4cGU8or+t
1Q8+IZKqCBqFTP+g1yKwjzW57oicZI8DkutST1FJjNQNpKTKwZhHwNQCbfVEQ6QF9+SG4+Zvid3S
WOcxVD+Ufq33RtB/J/ZXaAvYSqy+SFXuM55DkYpoBXcVVQop8k+Vh7QnucrcYXSel5GWF8gD7aiY
YFfB0JAdMdC90Cnwa+I4i3lZi6+cySZ/L2uWp1wG22G1qKCgGDM2ZeZMYFYShAlHuXTp4qnNpL7u
G+NPSWNpUmpQkIRqxmmigICSIYqPDZ0cdFs6CxWKqLi9CK6H4vmbrefKutH4Y8TegwVQMu7mWimi
SM+NSZYZwVXWByCC+Dgrjw0IRXL2fFUqNDpI6nTJwnvB0CqJJFVVa9px/9pmOT/BTI9bZyyT6Kjy
1CNhTTuukEEhSNnCSL8w8bT9sRJL/WfKpO2zRPEp9Pc4FIM28iW9AgNAJ5vF/OMGcmOAhN6GLr0I
aIKzndgbBcki36CZv6/sQQD4Hgx3BI2O4fVdNCvfqtgt6eS7HnpOVaegvFr0suLwKcMfDVP7VlWB
j8k6Y6B3pH0lVU3XUOf384lio1Rp8f3tCcCNl7XizNSc0Of2yerwa2hwVHkV+XPrUzOqpf2B0P51
dYzevCOnzbqu7ghv9S1mxBKbDhiGknzkF/m4g010o2AaS/IFq3h/FdMknYLr++YhnK0je0pEm7rc
aHTHZqfMdbpsxzdQUiyKaiZUhblmWBaCEPcuizFtBECscnlgmhr0aRQYPWlVh8EEml47vvRAfwK5
tIm9orlML1ibCenB5qjJgmy13apeVpYIIz05/BOvW60oh2oLqNaGbzVwdMqUT3Sgry+oQmDabceA
MCJEYTy1Gz39Kj3SljZNjgazCTOP5/2TBCSf0Ql0RBXr9MTqxEQQfi56rzNN54SqvKCMriHGi7ED
iCGG8QfmVKz5oSa/tSZNYcNbV73PAVo6fwP+xA7gcgT5MV6EUISi7p4pVtag5M5jMUJENCx1p9Kd
erqwo4CYtfM7zLqeD54fTwWPMZ31YuKH+Gov8STtjT8efKk6bYgVrkslPHkN0NTsI/ijfxOiqfPB
G4zQG4gUQg/KIx8UJQLYXyLLPBUDrm6MsMxv/7pvBhdHYcdNmkvhmt4ulH9COoqs426PRSNmkMHx
XqOgvj4LjkrHbraxPNvUjKbtN+SlVfgngv31LtyGCxjWNrtNn9xMXniFe1SdB7ov2JFpsvz/QX7A
7xIw/d6gQf+d95UOr3Mw252UJoIz7KrV3AlQzfyDe5sbUIIBAjS6ernjn9ZRjzRB7pDwYwqmw/fv
Kb+SEkqCm3NCATbBW2cRdTtw4L5jmToANgZNQJRk82G0IuqYz1m5+UcZ6ke2GdQmN/XBRdo1YpB8
wmERny8UCp9ejeDDQR+KMJMq2wjkTS9DmYs5hOYqz1THgiAoVpAf3aEg7sym5//8Ek/hzPGVwp9u
jtSaKYgiFDuXrvu+HWSqlAA4jC4png1mw5G+woAZoezWICm/m4IEpUmnRmUUXs3UEyO7Uy9ZcM1V
8fOmULazojnik9/PAibobjGkNsPAJaQbfHHjJQCf5ddMuo37b1pxR3Ll2FZFhSf2MtaYnU6C9EAC
AeGhY6K94PMXnSj//FZusa8Ns3587aofWrrEJ2tfGat/dGCYQZk41xW/3mkqbCKq3atUNlpz0Wrh
nl3W98DTt3knbJPXzoItK9uEng+Rd9NWHYZWsrXV8NTUzT+UqaJZGaNvSCvDMWxIPn0dW4MfCSqJ
X4oWMsRKgoh3DoUR42+L9267oqTRLmnCAOFPjvcz08CHWPuIbIjnMCBk0wZgUfCq1TimLOVhAXI4
1WnGrvhcihkbki8dj5qv53QPjjd5VOZi9VG7bqGfGYJfboofR1Nz20UsSffN2LOVfutqT+/epObq
p97UXf57SWjaziQQCuoCkouqXCoXKAdaOwJEsKhHkyzZfcHytOx0Hafjug5g9g99FynidW/2/sG9
msmA5dbDOYwbYtu/a94dqXVKYOvjlCHdlqi/pO8KkBNE2fbhLABwzSI39jg+yOLXrLLlxf1i4vdY
KtgYI5FFW0Gvm01cXs9Am6UC7eosn4BpBQJxKQ7b/pxXbT/W403yrJVB4A6XYuqQVZuVoIjcHkgz
MZCNSBIhKUK61SgwWv8y8W/hOnAcpw6hIKEQ4SHETSittGGX+CXpVJXARR/NvWzAGOPfAk+Zoh8P
qhMvdpiXJv49CqfnClNLU5L4DvxoZymII+XgTdWR5bKJxunjN2ygvH/ng/cQg5HYcyGxK4KyWHOI
Pp5VMku7EQ8toHIgU0+RH9I6N1jfssYz5uwxBYj3rRJkX3LNLhNaSZuhWWWNsEoKkCZDfcqnfxSA
jW3mgJCMSoE2wXWvjHnF5MIFuricu7BImot4le7YG/0DaCRyb3s5fc4AqySymYtFLjGjcyqIaSPx
v5kV/AhLB8GGrvwsVW8pfVyjuQB6fEEvPi7LBg33QUQIeQyLyjyIp3lxFTvquY1UcVrwvNHiiOlU
11/SkS3pfnAOwZDOTjMEZPvuYmj3CrEs+taydHh7UBoWy5d0gkNBGbj62wpfduoYCKj4NK5nghQ3
alakZD3ElO9HlLc7t+qJhUVzO1vGxbX0kHIaK5VGeCq/ay8Op7gjJLPYOkz0Y29Lv0iNmJWuiB2s
hLD8557iB7rqmjH7hzpdZPSxZANkQpJaYsakU/b/rFv5RPuLAdJykPe0oJTx3hHpDqVz/dsM32T/
n0HWqdMige0eDY16ziSCp7Bos+ocMaW2GcuRHu8FfH+o/iZVfnpyy+28jlD8lyWeJoH0G3v29LxH
7Z9XNNvn602H1AABfDraCpa1J2Y0V3DWHFEIYYhelDMTWTj8Vl8EPm0dM2TXtzp7v/8PTk73Hzcl
O4B+QEGIUeI38QI5NynQPyc+z+2v/aj/7zS5he24/D+GJeHJldJnvttJ3Eh9v9i2mgK5LbLNxjDh
eurkILVK4jVglaHr2/6GYtq4enn+VvlUXZIWu7mpQCXb4kU79g6suBUt+96p/hRjV9PfL14gf8JI
ID0FVTmR4hgzZ3BircbaI3hCbhakE1dVVagnYwrgZ8pL2sza6AYznePMnVSetiN3JqXciuosF2W9
db02gyKB2WBQMPjYtlK/XquPn3aJtccA6It3Ne2VfrjvM1VKGZDCuK4sY17PcdbsEabLNdCN9doz
IHSrzeaKYM9rhkyqDRSjhcDY4KRHjMMhL9N7179nlSlQ+kMxQ8jIOxg9AtBadcATuxNa+aAc3tDg
KkSARAIIuFBEAZfvHRxdRMRxTnwG1RCr1q9fwBUAeiop4JIm/ESOcMHaIr/+Sl9AisCBPYv3rWDk
PXstj0R636SNOWLYaOrfXw/YHw60fOLnxCobbFjZ2h7CbmX1F3vC7MG/Ly3eVx5VU5mnsw0MvL69
JBUn1SDmYlEeZw/tPlLBOhLDhGVQRSTmsaacIq4bAt86+eKUouFoTVpKEwdoY9DB8cgXmzCDZy3r
VUPeZbMdO6MRTAJL9ZAVF5t3OaneKBhJUiZ1d3gc8IYnBWJVfOZWbvZGcZxUxIHMiE2ixWWFMM8B
xZHYLYPKhfTH9PQQBfFPefNqsrMKM16AnP1thfvMFYn1dYdtrozG05X2PZZwcr+GFW/Tov/6HQB0
CD31hsjrnQ7Krb9Ij0DyhJZsv0X52g1PthCOfT7rnToVvO76cc/T9zI6xUUyJdlxfS8zPEVfiefB
sq6+yifVNMfniIntqO3w8qhOto+bEyxgdPB8uKFO7Vb/mBoFfysPMpGLWL1Agnx9tIn4mwXk1SwV
/SoMMfkxEj191UtHtQJSVzQy+3Dv5OH2lc4D/3AjviKVzC16b+PYhXk4xP0R2OhTSjt+3Y/s/xKh
FYPm9ACCCegVXKnEHKy47oxP5FUtU3ZdTUvo3NGXbL8KrhwagSPVAmU0vwf+UCVyU3nu5Bouq1Ol
NEjrJcIRvjD0uXJudWbW7O3NfLzqMUazAcJsaYtUfiNpBUsA5rWY+hVdQaZSmorhTod4/Hki5ajv
jc8x8OKYub3Rp6ce0CIPRfOItqI7D49G9yD/LOTr5IxB1BhSxg6lxn7faFd8adSQYjquo7d6qlMB
nAXoBQ5ImcyBMMwXnGEytRVf5PIt/GGCTdDaQcQZAdJ9qaJJMbvYutJFxCusMxqA48XrSZ48g662
WM893YyaXaRcd+9vxMtN3Oax053/3U/p8RT65pIMkngYCqGcQk9HtgH2OOJCT6lzmOqh4ed/p0fK
Q1If0o57XKjmWHG1Ej8uLrvDYntm/BhJX10MO8YK77wbxr1S0OksbKI/UUDTjyThvF1oXeox0c0v
fQwzDvQ3h73gwiAOFeyYAE8tmvM0hN+VOLUAVuZ/pK4PCezK+yg3QZSwNb4PxmkY5SG+HDYt7S2p
rsiq44TpANPY3i7xc5gnRCdGVPmtalEU7+wJCHccwRh/0Q0gkFsSUm97OVQEgsXaFzUssXAqfm4X
ITsemN3VleygMhpfqXCosYV6vWGrbSW8P2SdspSuIh4v0Z5ZZGaHumYOI1hKEMA/7QBssq0NGDy6
bRwKmj8SFGXd72RTaBv7phh8VnA2dytqyCxfnna++FID8arK6gueAHL4kCR1XXE+brh7CPARqDs5
+dR0Cuxw98TWi2j8ery2Gsp+FegRc01mC68uI4QafwQI41UP1XQCH/R+0VdUdLVH1autLx6NLVut
bogV9W2M24jj2qwiMlsyNp7ElZdnf7MbDuWcXE2YcLSBIBQLMY3D/9TbRPqE8WYBSeeZizQnvrOI
/TZWaEh3rPXVmgw4pVFZpPXou4oJuzSwjh9ABvhW7fdxzWVSPGYmdVJXKVcisEE4zQlsIgaDZLX4
LZou7O5cC7oZ5pkxq3Nkj31vMr/cyJBCDcMy4aryjUKwm7YwSDWrcLshJVE8kTS3zrgn0ZsGmere
kArE4s5hd5p8jqkrORxsBSELDZdbG2jBHYhGRu7Eb3Ga1dIDmZbOyFuT0jkL+DKHDm15bcwLWL2C
43kUEMymsUc2tDsWeB7e80nj2itPFI0XbBdaj876v60XMWf0jzCteGBhc53uB1j9OtpY1Q0GtNwX
UsXNsWq/2pzBGpQ3BXbTlNS7Z00VgHibXd8IT54cJ7Hg1wS2mrReoNvVsfO8psXLVO/X0lcDMeAS
LVCzfvKfz/GQFD5qYZOkRcMrkZTRMLArUAxOkdMbO7m7B5cbHRPSYWHUQCmtAuv2LTVxloWyeo1d
3E2kvw8FII+WEDQEsYEHkHCcGYXLWEVxavADkh3P5bdRRieu4O7qk5pwv7yV5xnqdRNdWuVyLuT0
TEhkWN5rmDamS26VFlc6HeJHCm4n5ukNyXr/1XBeASLgT//+L0Nzm+um3KQ8k84ni//ifYgp/0tU
+Q9BKhi4iSxv6WESZISOUzW59QWhyhw+rr93ngyfo4teEM34DXN6fok6ZawbvO5NYUl0ymTOgQnr
GxTmNCdMq7BQ6pMnziKmMUvPcfjF6jxmiWrYzR7nfjB45MFtH0+eakAWiC/E8bPtBGrKvkwYxCO4
858W4Hg4/LSd/6a9AKxRBvQbSWLOXFbXMx8mX+u2iNRtg+VvqglmWCNiVxH/dUGDRb1ZCt2bfh2m
rqZ4ZX516T20LQ1N81ASWbJZJkp2HzvHs2pSPYmuBJmIPSWNhzgl1j+SxXpZLXNd1UZ8dRa64JD1
9EH3GeDhwc7MSXAJsRFjBPxwyCgHuCkG+WRWM9eoC39naflpHmuMYHlGwxghw+E7lP9hkHiROBC2
Hx4Ulm8Cg5RrI4tZ5OxfSvwBgvy+AgGzkc4GOfu3rfKSuafig24BKEBenO+WRuwIXs3clxePhyoE
tn2KbSpI0ZoaXcFgENoRHhv31sS5oYy28M7ootvK7D8mmVHb7FO362yd7lEjFBl2m3YG9mj48h80
WHczUw6EWJxTr33oMGDCXXhAa26y3zllUkewwaZggr8CrnOx9hyHqbxJFUGCfwVljCUdgNavplOt
FbEqNvoGXk4AL+ldazEQHfW3N4H576wGHDi82FwXYXhI679nX1DJ3rih2c2b+YP2DgCOH2uQ0LEj
BLWkeCnoeprxsYiwcTRI9CWlKoQmz2ZuZz2U0cEFQmt7zoU7K5wdEahUd68APesb6ZeCIFtWA1vs
GqwGx1/exJiLnckx7ai26uGhS0IbmJ/9gf3Kdmv1m9QtlGvzoqjTnAMkWwSc6MQi7OvNrtkc7SJJ
rY2FWZe2MlxHy1sgAdBcQp+bfnuSjIlm9J681M5F7FQ4TAMzf1wi6iiTYQnaH2pdjFdA2Dm9HvdT
hglFrhN2NzHdpidsrUZZyNTOa08HsJt4kXc275imTW2LmJSePfuiyGXY5rlI0cJu/Z4Omo5sgEH3
7lDQ/X7CCaKbX25seQDE4f5xgxVSlwH1KZHoYnYGJJD4dtkbFcHE55NsFhZjrAzMfk5Cc9A5yljd
StF2qONtVCuA+FkivMZtSQ1cMrLqil32pKVvbetFXh3s3kahpjhdzC7K4d3pae6eR3cud1Bq6oCe
t2eOm/AgfhpAn0fxl++XVjTavy+xr4NJNEScDYYpeoOdQ6ToAaIz/Un+Uj1PCs94LPAKYz2PK0jf
upQ/DvzbwA66kKxzv4Tbg1fEXL9kSBgo+wwuE6/NHlA9UeqsmhphEImKvSCqEDlvQsIt8LkA4HAc
D3VL/4uMxhI6zs6FRbB4+p2GRTGL8rSvDQ85FUgJrYZb7cPZnWTwVgBEPxMYKkB+5StUwMpkHecM
itPf4AV0C0EX2V+d78PWLZWgod7UrCZY9BVX6qMnEqAiIeM2VmqePOk8N0BDY3lG7tl9xz316gOB
IVRrplWUPrYQsdCogsDjCY6lPLSHeusdaZnP3f8TG0ybly72/k/cvkHU5kLXtiR5JF8BptdT3f14
uW6GpcpQeOAx/pS/ir3KCzolzT2EpsHSKkiW5dxX7aGZ+FdOEeikZKevNcVYxjSbQbKqVwVhp8Yu
t5AFGwJQVQc0qvVfoQB11cE9Rgj8Sms2Y1oOrUMK5APV9syRz0Un3GnbTDG4l3LUYywErqmvPHKy
2aeVRqjkl+Y3hPnHi5F+h/JTpmXjB1Kng1zxkc6piSa934m5/v7SJeF5iJZwc4E//n2BShmHzTxN
aaXfrPOazlNSqC9W1vM/sHRb0RpiIu2YOVAHxe4ev9X8K70QZNSaSXRU3MaFIKEa94NJk2v1PvIP
pn9LztrKAuFLYJmQhlTy1e461gthIdYydD5SuIrqgdVooi9Hl3VeyDP07EapRdNheMqrZ3I3djlS
6+pxCdZl0PugVUvK/6jjA7BiIcpWnarbLjkfoh38CpuHUPI/MMwl8m+MaIb28T8b0oUA9Fb4moWZ
2UpcWUKNXBW6ZxxUaRz0o55NVfK4SeYKsntAsPtvw2wD4X6ZbGvfvBtMOV2Km2ctfkvsd6fiqyQk
p3g/CKUhSvJOAoAu2YGfwiVUdPaVsT7dzvJTspeRfLDuf9uhSlO3ODyQo+fZlcGEVDmyUPKLG9OT
RF0jlLWUO4Ndxg7IiwUx3QVEEl8uGN/FP9VKduWSns6D8XCv8C6uHyA9RBb9vHS+P9UXLVL5gXci
QwyrGDVpawUa5ZhDKmUFAh3WHkME7T/ymPlsag5wzLAwEZvyV6mWxhEUci/HAin9m4QOw/A7V93B
mfGUv2XpVmMlUc09BswCdtsWZ3u/q8VmO0sMrIUa1wKZS+Yy9YKYxSxaB7bh0RzuSAn/dtjxVp1s
B6zsKjqeQesmjAtqlQuCqZQGm6tvSfRw9jCaJrIA5YmKIiAbyXAHL9KSF4sZ3rzrhaMxvMpshhC/
Ikxfh1kTSBgvWGuoTeVjhuLkZjLoN8rP0ZG+OyZqrqxALVfFF+RKD0vs/XbDix5YclL7cPnciwm4
mZyGpNnIw3vjtvFTC+/Fg16VWnD91ibIDivKuiPGGCel7eAAAFPunUtupIwxb1Hnfnpwz3SW2a5O
5EWh70TRHa/tdgFsrm65kpJqqxHkX3NaAeM3UwDvAslTDBwtTDx/jrFvRlUecg7g2BJannwcYjaJ
fiygQtjzdDfq/OdacqjyBNX+blP4DgtL5IiqS/B6h5exLbSEA2ereqvzrd5+pHjfhWFOYMu2lrxN
vbTV97m7ytvwBFhhau6YDFP5ckkeoWR3vlJKxqvcuaFNXuSXFiakJUsmkRwQ9jrvnG/d7OElCjIN
WgOh+dA1fm8IQuKFVElkCXCWqtFfH0ik9H79s1d2GakJ0r+UI6FElWWckvxGWkrKN8n5Heb+BvRh
s+Y1AOQGyHQMxR15895bVwuJjgaL4e6WrPYLHoDUd2qnwMRz5UzEl1okabscvgiU/CKVQJuQ8PAz
ZwFFry8azvacfjbbhhOjJ5iEQOlYlbiXG0kDN6QGyDFaB7wBfwM7RZakj75dMbEK4LRIKihljzTS
r/tukIlMn98ySfid4d45XwOzfNJ5+DN1R85iGEFnHtiYy7AfZ2fWnmDl3R/cNrzEPLGzqOLQZaAU
A1XIw7jj8Dq3A6e/xM8W6Pws3Unw6sJ+aTbE+QKSOaHnLgoT9gZnjkB4MYi2T/saXJhCrOViwBMO
6JeaPPn6l77zjbprx5RUjQc69ZFfbakMuXx8qDISlsDZb42Mezr5BAXIkkK2nWcut/GgCsUzNGHa
Z/nI+Eb3QDfycwCzthFRKXgrZIkPsM6jO3hWo7clwvv9Ls6+mgIm3E7lrUmKQ8csFDhIJKmIGO+Y
FvzmQhEQ1pP7lXifxzlv3TpzsPKO/hpPKxXboQiMcDKfRjY3ChiRR1OYx7akcGxco8aIa9EQQXDp
amq1KD7kQ3D3BhlvW0CVJiTQ13FmywNShCYrLVyEHLjoe3REAJBlGHi2ZXzPJUHHZ3ZHla/+IvJd
yNofRENoJ4WwNxoYz/G6gJLq4Gv8+PsFm2+1k9r+21i7D5gjLpNbOtH8BK6cRpV+TuGJ4uk8msb2
hkG82GcfawSPxhVc9dCj+wqjK9RcaETn5rnwD7MtmWxiRwj/mKy3Bfdcy9eWH7to8Vd1xyVnzA5I
YXLB6HuF8C8eHMmxJhVgE2BUbnhGyiYucx93Kfynwye1BUQ7YKDU8cg/p0hhT8KckBtftZv5iY42
Nkc13hp3s3Qn4tm4sNzsx23gX+HO30TOx/sF6L5t5xwr3JYyPO8AXPAdVSJ22JRGhGm2MEaChjVM
WOysSRfU7PhyDc83xuwZZaImriqwpcC88p2Kk+WjNYB2XhCLHS11A0FqBpL351neQ0tJ/VMKBPhY
ePO2cg/smYSNpv8ur3GbYQHy9fpuJGr8BniLPsLel4shhyH5nC5GyY86POQYL3/YFgj74qMz2oJH
+4plXgapULMFuDuqUIhtbVQ1KQWLW6NH4SkNXv2yBXXgniglQeIrcJSMB+bDLdce47GHlU0qnHlg
PSV/bJ9A9iCjNXTHTnURIMXRAOierfjT3mvunYm1uzMGj+cDbCBEvIz8IzDTizrIfqkuEYiXEFFD
eMy+mO8pOjEIKXGoPR2qVApDuvS3HoZ9eiGetHRAgz9qwF7rS3GeZkK2mYdX2otI7/9XuWQIbJN/
huRIdlamkc/NQN8jvPFSdUaPYgwPa2tMV0D7p8sJ9ERRUxo4VquY7vCBklvb2s6lfxT+y5O79Jy8
YvfWgraN+so0qc+L2cpyyjwYEupN0ssyqHmM6l75jRssqQ8+FaQDKjPFqae/DToJY5uRKf4oYE6G
MEKOKtAS+vVSl3ebJjHDRUIg5J/m6JS80TBBmikDu8XieEJ897hXdL0avYG/p+pilhTh/VTxNTf9
tbBZnmMLx5T/zdkYgUHuTgeL0XM+ph0GY668l5PwIbudi157PtOx5hp6/ovESGQAkgleIV5bs8xo
okU3Rcc41doEv76ZuAwyysBNE7s4faT4kaJXWOcREW9k9F/3AvsgFebTFqEbAPi717HocVW7A+sk
Hbbr4hT77483EIHJAFoli+RUQq9icQhDwo3rvXHTMqUGiYO3fSOP/TAAcw==
`pragma protect end_protected
