// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
4hF/nlX9a2x+8UpAZGudOcdJnwsRbkxCBHWGVIdPoIM/fsM/HCnBLlN3HhsurBBq
0pfgzpDlfzqub4xFh2iS6mL3C6J4pVcG2D2aA0OYNr/Ow2xzsuj4Leh69Qhhvd+s
Ynil3Jqy7NMOGwXZ1vWjtUH9tkmI/aSNXhNUoBHTskE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2176 )
`pragma protect data_block
OFX1SoLfH6VGdHPsJhhzIhDgr4ymL2/QXQq2COeM1Q95k+APpcEvsy1FV8cyO/bj
cPRgPM2uLMtqWtfpgOzYk2FNrt2ypdK1K6RaLzFZoewso+ZLge9ztd3J9rdUBxzs
uperjFhz04G/exYxjTiAUnjLzLSoaaO5TSrXIieAPaJLgRb9yyMjw3fhGUKFh9LW
r2Jj0yY3u4JI6Ih61ktRAr9SKPLry/C1mFpCgcelio/9l4BVPi6sjTvP7cKQoXlF
umllHTSenBl8UWe2sBIrwWoW36T39wEYXGfenBUQU4vUCjQQPs8MR7x0lup82IFI
2VLme6nRm/l+NQexg5QnTI0xtZmPukPFA04/ASeN+aYkORWgc7aRwWl+EKyIJii/
Qvj4S8ApTsXAQ4x0JMimSRkaEhKuR2MEejEZbgib49pNVxsDywbTeO/LMURMA9sj
2UExgNVsmBgXkSdZc7gLQRvPL2aLChqaJZpndb+Nv8+nTrqoFffxxzZGdwrrgGrA
w94O5qq1WpcotxgDEgouL4Md0ZRxKXSX52uR0ihcHSkj9ASIbys8wMmt9Erc7ImZ
4e7WGRB2HOR2TNKJB6OF5Qvh481o0VQFHP52sdzfB4rFUMXyKJLw3MzSEutefHc7
d6Y5dEH+6BmVCRbVtWggzLbliB/kfGGN7UB2eSAZlDMxGRdMIHaNNGn8/tBnjA4n
cRm9spn3LrgBTky2FVG5bxfLt7WkPOBwXjNb5vfv1SY+FinO7aW30BBRTXYbfrre
EIttTlb13R9cD80fd8HufvmO7rHFkq8oTdDsKpfrBhZHmd5fWqw/gvUX2T+EtFf1
ywc4Lk6zhKlIHKfifrKxXncXfWlxamXEfIiNfJr8H724aESYe1X3bAPSSjHBLgHE
f4PTH1q3ohPjjYSWfRvsP+yEoDSjDh8Ytkt+C9rpsh0Awf2IAT1O0qCHqPyB1xWd
UA2y3+mR4SK0EEVQggyW0nMMUD6GsusgPL8KpycMixTUZwZ9Uh58vDoNYIUXFhjE
YuPbWP34k7P77TxZ04sfGqT8+WYXLQKdPaJ1JTzaynQ5QeNsH8YKpJesr2VuSzwW
dGvYt1yL2kHjw5D6wHvh/tGfl+/dq7A0oZ1XYnHc9hor4KRpSCoWycRirnfcsP0D
vptxFExpQUl8wcZmBiLFlYU+FbgQzIf0yegGWEzY5euaFbKLVCO/1iPGdLuOLX51
TSOQ5jS48exqt9C16BIcTnJz8Nq2bbwF+7lODMoiykerfeSastaKEcTRn6Th+7bO
PRCNQaQdxOWsZSCpLmPGSY+z9jJFh2gE9JH/kVVYjfDJq18ktWDjT4CHxjv+S9x+
LnGlUjO6+8X/BXXhxsYnjMdgmQSBDteoi3i67iVUyqx+zmeAFKtsFAS8N87bTyAa
UNuqmAnxbIniMY9ti6ULNAIlhjq+9VnyzO/NBAbaRPAuWvqPHxl8DweJHi9c0OLS
wLVOFt+HgB1UjrMbz6UvwFj+n9tbwj1hyD5fmF5W0pkkjAYN3Aiky+1Mi5gCkJbM
Xb+8c070YS3FkKvP0KCYd21hD8JU05UE7a6lfAw5T0lGvF6azKDsi4IP8Bbd6/0P
dpEt+1UkgtIbXDwHpS/w4kYt4kX6PJAo9CUgeYN7nTW591En1lpeZz91vvnse/LV
62qKrYDuW8Jlh7KXx+P1i+2peQlqXAOiPqvs4tHr/I+Ce3DOCLDqeUu6Nn8qiwxr
16rBLLtd9Mu8RNW+Tz2Z+P7GUAkztCssS7KGkZA0ZvMv1ADJp8svaN7G82JeJIfr
MpDYzNJ2JttYdja8m+8Ej2DoZJANjJGB0wRODMZx9nysbDHatJY47w6ti/Pjozoc
puxCYTgjOm3lXSPjpk1xEDVSXn8ceGry/HjLABDPptOZQi0/yHP9J1g/hSRR9ojB
rLpFH8b0xqbVbOYESuFE7gMZSNB1s5HxLueCyDBqMawwSim2SHwpMH8rNt+bkggf
Gqsa2DngzLJI2I7kVbKZs8oHiiuCWJ749+FoNVb3XiMDSdWJoiJN5OWYwJBTbZmr
jW9jo/+dQyG4whGolbEKTTXvXggtABXJRfctZ+N/LhZOnonSEGRBT/ZdoGXm9WDR
jIuXiPbFg5rQmcxsFg6MdUYeuoj91vJuscChZSHv8Wz9cksQPJ+z8+TCg2Fdr07B
F4knwaahu8Wf/WQ/7vzdve/hqVcFc16kPEsu1XPY/UlLS/2xQvjF1FYU98XdJwqO
yuKGeL4hrMUigPi1wTkNmIU739HjIYq2nahCvzZED0OIvuejMbHIj2Y3PaKxD7yZ
AnKsotrkBP0kKWIUZIR2WeQ2W7mQ9ZPEfvDVK1rpIN5tv3zSij3bMmWdiIScXriE
C/wCG+nPdhdW7ghOdkMJ0elTajjzkZ1K1uUduU6TwsB9XvwJTHniaaJns/jpbxBb
yVXgf99xmxH8pvXAJYlcM0AQou4rybcafLpCRZtqIxWSbgJbN8i1D1ub/jWRyfLx
/axRXt/TYsl94Zc4Hn13SVfjbuEwddZKRBhjQkHeqElALmci8nZqxcUtOVr7aJKQ
6BSVNuXVQ08oW7ss8VkMX37Y8pmbcQBK9qh0wqq+6FJoaEvvgQ/9GLTX0RZx36U/
QHuQ/svjHqp0iMEHyR6w8J5s/M9KmlX2Fy5mnYo1lwVL9nS+TvNDdRXU2jJyx8eA
4tqAmA+1paf9umQhu180fYgLRVXFNWpLG3S7eCiDXd9RWbhqWxpReZ5+DYk7/GdP
FXl9L40A7faZbQagO2Fh2PB1d7Ds7tVpvSUaoUcfwPuG6nHNEuVuiTaiIjlWkgIo
O0frlkVPbQ2B4lteBBUXvVf+yJ3pM9tbqJxmX43GSxSi6LZ1AYGFI7OedGMMguiU
4ml14XbVho+Q/MAjM05Z9g==

`pragma protect end_protected
