// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
jsl2UNjIxCwBu+/KvNq8ykpIi2p/Z+K+N6t20CpdJRiZWB+5LAtzpnMsB0aYUOCg
p0y0dgaDZfCxxWkZVnlHfRaSKjc/71vhfg1mkA8Qa2x9Ow/TJyhTHKCigotyLJ6P
dbX0HKugx96qhFCxE22P2Myy6sxpZq5U693wvm5Ys88=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 86432 )
`pragma protect data_block
Wwneufyrkxdv0mAzCMV+kJfJUAVUGJtRG15ZmVgQsSBN0MKLvIqyW5I08ytBE5jd
Wdd/A80TKRBGjgc72EXkN6HWnplTHFx5aEV2U4HUHrQo7Va/yjl/CHku9MiFpct8
KqlCVv3gXPD132sZetydRFzMUXKZg+m9qJE7TNfVdUzvUAkCl1B/l5DPHG5YRRvQ
XfJuuHS+B4Zt4dX2zQNVJvlpBwiMgc48yrOXvwvINoAEylC9du2XFPpnwjmoUNmw
Iu4NwPTefY9h3+jti02ytHCHSNiHxulNUQXTjO9mdN+QOWHl0WQVMXXnkKPoblvK
kuvO/dJV5tkHiw7QEXgUi2WQJRGfDW/LsEj6fo7PMG3FsF34/GPd0k8dijQlFc/i
Ur/5UNIPK0btwvbmJCZtT0z/OR4qd3AeBWJ4Al6Q2rLMPdTTcZPUsn1YljsCMozw
eRU5ex1nipQ2YaUgmZNbWjmbale00uXWGwYbtE/l1c3nS4yygbNrwV6/0NHlAsZp
YU1JQPomWEtRBHk55P7zKpJmytGBxdgwoSzvh8BGggKBxo6PHcYP1CL19760NUA+
qIiuZ1ksFSvSAh3AmuuOfaycpZtJWW8W8WQURdBey+C31dNBUBLu7hEz/z8cmtHZ
fbtr/VazUKnTVz8i2+mXJW3LckLGgXwRikLSNSS83gmevhR68pfXexYL+DrnHF/6
4WnKLhYcQYK9LFPKEDNtJAOEsjhnO5t2jeW0Z/s8jxnOoztuzU1aWkoaZeEM33wZ
duePacFD3G67fGT7V0lBGxakhrHx3krSQjnk6eH2Ofw/IgOpvn36vFhhpK64UBGV
ntpk+JThxCuefw6PMdGxyhv3D0ktm7Sg5vrl0ShSXCeREQZF3tu/8GF2fc9uEM0D
qONGmQPwRZDw8tgBhjl9gkWaR1woyP8ZPMs+XsmAY2xagfGArPlkUEVS1srHsebb
cE+VcNILYEMFXRabAhI5cwGOxeqbNgdvZUOEg7Qj6g5ooAyonZkMzta/uRtP6o7b
i5KA9ZhN3GVkWIGKvnhYUqBxf1/PYvfxaEmMj5lGZe+S1yCZW+iSLd0eM07FsfGP
ZQsjD/TPkBhBGLj4eOFj9UOKjMemvzQuBeDhiuQmk1Mr8sOOdZYexKlV8AuXdU7h
ZzdTKAKH4pClH2Y+UszOWP4I/2zvIlCqZsAT3hyaoaAozkpTEel/ZDQvCfEr245C
Btxx3nOjuB8HdW3EwzmbdjJDXw6hMFVH1psN2VXSGXDcUuGeR4rplrLWpeOinwaJ
jnqNCgCjWjSPaqOiUgJc53gH0u4uAsCJxGLK3tEAkUeNgcjjI0YD1y0v01b3ODzQ
zvCutQGGB4jj4l0eDn6iLQymc47bS8gxdaL5gZZ5dy0MVT+o2vGeW7c585qtDXcT
NNfKoU6y5MK2Ypkxat9UbKFGxvMiHUV9NuPw2AIdxTmThDtpeTLyzcPX1AlQ4txh
q0E80EOcZz4TYHXQ7xU3IgMa615VrpCNoGpD1C111sK2BbMtbsObqyFXh84EbRn/
mtjCH+e/dO3g/asCdEvYZcFIUFUEE/Bs8+vqfPT8hChhTaBnke7QXlUAljcgro9l
eieWU/Z/ENG8ObUpVMSPSyJjV9bM9CPMs0LlCvlglImcm8D6FDqrFndd7bwltaC6
S7ZqGiz4Wii53NoBPnNLtJunBdNQWuhtgq1TbRgv37ANePkU1y4lCHAYSNiFvUz4
0vlqVBZHs+nDJA+iarYzi4xnJ4bqHG/prpCaXbT8uLcbhOkFJxMJ2tA50KsArHjX
MX8DKyz77htRJF7wt9bx9kfywXMELUYwvEnxT+hb2t4c7mhDf9304+fo1I7lwOLL
2+qb7WFJM1kJ+mf4PdZCI2jTUV83WXuBnEEIHU7K86wPS3Fk/De+Xpxl09WsGdPo
yZ0u1/GaPYMxLOTX2jxyXg4n85MAj7twDh9CFzcxDF+RgP/VN7GvCqX79kgRW38T
ZYzUaf/VKm/NojVuRlTiGWfEb1YwVaGkyxnYl87lzNFtY0XcZwifD6GGIsivJlSh
7Jp6vUDepcjQNUzQQ6ere3SOH/qjNQK3UX3ejNUe5oXGr91qjTwLdZSBZSdkK7e7
c+y1IE1uip66QbBYy/QsSGMS3bKnWN2EVX4E7MvxvmMsaH7Ptnq3fLKZEwpy13dY
iZhjNTRwrx1x/caaSfOcbRJxEk3wfHl7QYKaA1UsaM+OyNOykM+L02di3YUSiaLZ
iQeu0/Y+uzD6s0pEnMyX7XPaXSqJIlnLf5a/F4CXsOa8+UZkRjC97MZbINUCgXgU
WAfAexLLG5uMVb1s/1lFiBPsv4I7CEJtBxRmXx+UC0OCXo1wqRqRAryYYx8VwnTp
IfVW/ppC9KihnrHKsmDLCO7nBSNZh5MN1zxeoN/FSEYW6YpBa8jhpFo7E21r6VDs
tdge8A3/VVpH92rof9THWfx/bG0zYN8FHtoPw/QW6fKCIdDJ4kgGwwk7iCyDtwle
M1r4/q9FFLEH3EIHfBD1aHDTZ8ytxeJBkYjYp5BbRpXx19wJCSEbpCp8bnNP3EZy
KhTMYncRlzkuubsUjh0oBiTQZGQ+ekjh7jJEDJaCjxsajE3bQykZLUHjwOTmD4li
fvPTXMTFM4W49NsTPvI2tfNczcSTIPlIAHM5RW0Lotdu9sgF9aYDw+T6dsyg8j9p
uZfxbT9oJDCHLQkKjx3RkFAdyqXO9JqKQNDrPVPqe1y8KtdRO7NxtjflpbnS7axo
0BmfrqPl7M/gx4YfLOimBhcfmzl5DRgl0BBID0Wr0lqirmfWel4W5m1bBWvtttKB
yEWoXFwC4MV8PwY5yJGhvFW9m0MZzo+VdCfysYKXGpzy6uRJRwKlx62PES/TowZy
qfIRJq63CVnaVpgvBHOnUjAsBU04Osnw1AWt6bQf52KtdoGfpcyD0Sj1SK6S6kwD
QZJ8PY7nFkhWvsVw+OMJrEYTqC+j+fCV0arZpONDrV0LBjA4BqoTO/d121XN/E5/
PYaocB1zAiujPtkvxUwhS2KUDelGH6cHLjzhVkMIpqo2n/j4OK8crn0QO0z1fc+i
adUdrt9nS2wrkmAWUZT982CnODGgsSVtnKAY2ga7IibbLpe/PTPYFeeU2GbdbwOg
GOy2ln1I0tL8H71u1zmfgAUW8Na07fSQPnYlmvNI3xmPrPWrmGn8RiXL7ubsgy/9
MdsG3J98RyRsnbtG9YNJJyAotauvAuMgeq8efygGWqCnhpjte9YSOsXGaeRiMPWf
3SnKtKkKvK93OYZkEtIlIWZd7TWtRCvrvF2ZWHxgh52fJsAbO1xjbDMIMlhChLJM
7TdibGeW6gXSheT4UmcuizP4zlqZjRRKdRWvyXDQW1jHM6AYcIX7dM5koBgAiT2T
U3UMyizlRsmfYZUjQAn/p73ThQ4+74In3dBQG7yQmu/8sH9BJbGq2oqtt4LHqv6j
RkCQG9kipeqGVF5dx3qv3GylYljzHntzBvzkbILZca/IK0ZCewLupsfP45dY67Wa
ro94EXYVwc5wOLuclIDPSkc2Z8cZbF3+zlcxKut0Gtr0lFuojCt8Lp/loU9PQbum
W0440SZYmGdxTKkxTV8Lhi4tlgoLx4cKK6N0w0KcvxjrmXRUuP4RAO+p1xHKfDNJ
UhbUmNvrnryYAjMPKwhOyRT8ErZkBNm294QmrLU/g/Pwa48Pxj2l9voFmbWNbBwb
SwR51L03KymUlqIYevJvTYjn8JayJS22JtWBQMJgs9kNa2IfQ0vjLfkgJX6vtXm9
6pIxZXsytwIw4kFAFL/hCDXf0cinQ05wOlHDpYNd0La1ohWSQtyfc2822nGdlZcX
BTAPtHOde669vl+6Ci/1WJS/vSHUZLACHkqVUz2IsYhtZ2GiuiVeAqLON4WRPppK
nga6t/Ew5VSjAgKLJwu8OX5VrlA5YTplQIDhnaObddWJqdnuZeNqenxzM6vo2ylC
k54V7uZm/LlBPbVbgZ2mPabfXxG7xrMNYE5Nn6RVtRKuIoYk9XL5ceP3790Z411y
xtYaZ90hYVgkorqvvPP/h95oL7nBzjZWyfGSdIaoZuC1fs20Zjjnm2Qok2pur+z+
6B5wPwVvXBHinlgZ3v9ZDFiRgFwhyJndv1kvZJW8KAEJVr6ZPJ9tuQdJ9PgRY9dI
G5UyeSbbSOtRWuqxNE/zXEo4jJXj/KVidRjxX3gEYQk1crMv3wyvH/94iajpEupx
LvqBt82Rsi0wLgxkK1FNOaQYUad0BqSiWoA7+LjM6HIcXeQeqE30P04dCgSmlAK0
xYCXzKXvE2uA8OQUauRDAbCKRxy7SCRaWiTSyxp0H7ss/3/0yGI7kg2d5gXb91R8
JdIoclsdkD931fYOR4RkR+tMNIw7fOat4V2Bfcr6zmBFiinpIAPGupbCR9V1U6E4
gLk3MsYXik4Eb1tGnDKLsO2Jk80cOzFGBTewEeGhsOVN1sJ3PKZ55cvLaNHC6re2
zCMpvRdYEr6rG2S07B7XrkLMuHJwBvQOgWTkPxNpidoQR/3oJCGldm+fcQSelS39
492UxAyZACDG6UaleBdTaj6DxpaUjewH4BkOIX+hoipZcWagdjnnfSA8c6RpoJ8y
QyMCIUTB4DNGts61ozF07sBek4t9diNr1Xc6Wyi/mD8e+NVHMXlpJilMuMsFI14N
ukRXOC/pDIL0DApbst3VzJi7jc/s8OCs2N1m1+ryiFI7MdulNHq9elLsHvcVMSAc
lZ0tlMOourWmdc1yOlLeThvh51K7y/7jmXHpyMFTX0KulM74idX+soahOnCeOmRE
REHc2PL+2tnQkj/V/Xh2QmNPT22p0Ap79zkcdGrRvLypmN0kJM3LTCCWYwuBH9uy
z3ibCg9VnliO0YblsPOoehrZsxJIBUY8bepxJz+NWfZ48o9OslxyfVY/di5SHaKA
spwHNvF7aZ0Vh+8gEhnyLqfOZYpDmE0qESZOxIIBFQT8xKCG1HUMcIGiDCEFUODv
xAE1OnhvtghsJg/JLMFU4oWEyuZPeCUEjxieBA+KTpXUEuHq5HFRIVKfdXoLVVl6
emRIxxiLQbOE2Yq1OddsR8rHx/s4Piu/KjazYwrSYgE+cKixv7VFtnF9839Q4Ryc
w3PQDY2s4ka3J16iOp94a4AFcxzJWjEq45RVpWa/WbwNgput7AWqPZPHOXDPyJe7
p/yzTo4ADyURUCumvDO87Ei5CNJ1jIa2t4i0z9mBBsebOaF+poP/TippYROvCc7G
3EyTHFTHuwoJWDa/mp8DmQfmUuEc34Dvpbz/75tXKDKxsjT5i5mDqrVP6eLcAl/A
oitUw7dIhqp33YF38nDXTZ41fbaDCFLTKlIw6W235PJX5uHlk/OqTcyolrOMSy95
P5sOZDQOiSeFtdoXg+P4gKOVuU0nTt8Q5+gV84a7qpjZLeGbSUVFxW7CPraolVHO
4lUnuadlF/5W/BnYcDdUzvZoov/v9tyiJwf9utsj1fiCMlyOD2B85wqiplG9xZlv
QZGtj9OkGtWB3+DaKHgsH5YyEoG7x0nAS7e42Tx4J+BemIiQcbSAAiY9YxnnWlCj
lod7TfyOECsShZ9uVFmB1Et/Ovj3AGAZSDGl2ExfDTUbeRlAmYRTCAobNqSIaJpW
k80OFN1ukE/SdaqwaRwUS18E2+YAt/VedpqbYC00IvXi0u8+ByaRqyPRt2rKW43X
/hyLNcLlSbeRs2CfBZRVvSCkwZVNaEQVI8lfM8Fz+GWe1v+ur1awcz919amBzHw7
ADx2VxF1H8G2OxjXLHNNKJ2GNokhPNQz/owO+ZjoYTIUJne/2D094yY1bAM9o84/
6GpQUS7IGdmMLlUB4gC7caanCIwwVJh1o0WJBfIsCj6zCfC/2xEBYo3mK2/o76qx
Uflmqt0SNyg/uBg0s4ktZdkrD8BCfkaBWGKwKZy+1nqi9roE8WywewH02Lw0K15X
ggs3v+f+hraB8vMlI8mlygxcv/30GicRYyVhQoX8EstsFLVuhvwLUVPTx50U00QR
SZHTk6kY0JOjT/9EGqZdAd/qM9QUld+hDP1i41NwsS6GFOtv3AlSCIfFef5R4SQZ
npV6mDGmSeeZnxc3FMmpz7gv5TG4tgNzqCuIAKFPEBxVTDgwTrCLrKrtySXIMc7B
21HSokSN3hp1BVs+Ws0etvdSwJ6OFBSGHr/POU8uiIhC83fXNIHrxjeSJKFvBgBn
7Ec2xmPjcbB9JymAYS95XDS/XtqpJDY9UfpNm68Bh2VShMVW21RNKGOPhC31WZTe
XbPcezJmS8pe+hDr8BzRzoDjBxdxHO4IVhIjb731qnHLD9rZHhyrnCeAq9JYMCNu
l4DO47DlSEhUGHJyEEyAVk1eh2jXRSdU0d5SaX5VimLCSd2t7O+adc7QN/68ZiPJ
wThmLGScl43XqkGOh7DE0VyFhVSCwgp4agooo0s14uePaJOamx92VOFKVpHIAUKw
jQbaN8D6usvRrdnwBJCVPMCM3sILFNTl95Dc0y/aHXzVw5z0txN1l3NOct1CSPdC
CZkBXejS02sqtLmxiw21GXZTtx52QnPAtxxcF8KGQFj4vCvPCFF6NgRy5kkCDge6
56FvQS0mqSIe/VkUJ/cdmgUsFrBmLM0LcaYVKCRBo/Mk53ZdZSdxZdhQS33qHyzw
6qFf3ZZQTdwaeqhF2Xl/DMepbYndPSwG9kWYsHs4R4qejF9h5VZiu80OL8Lth00T
1cR2y58R5Gv1sWaClGvMGJwJUd+oUvOmvWGlqgNJdaQwIPwAAJ4MlMxOL6SJeK9U
c1ISMpJpGECInXU6f+lwS+Chh4wBTfGiX7tjoOoL91OIzsi/y8nrFSf6hrg4+2ic
BVEcQKutW7H/NwfhfoMHxpQIGt+lqF27Xklo3pJRo+eI/8n27bPMsXC/svf/TTjL
UB3J4UB04x74XD5h6cXNPS0r03lqjREguoJRQEY7/Sd8RlkfiH7c0GjUsLgyIL7n
hHBHXH5roW2QzMmx8GumXItwU60If2svGwtAEamOTP5k7CUwcJ+521kfr+GVl5Rf
W73LreOYjSUHC96Yx3Q9xvPussxK53pnVhPIoZhKp1Ao3wA+PzZ/3nsCHHHMXGR4
o2YgXgBnAG20wPCZAcKYx7q5QsCD/J96M4DUz9JM9MZWZdKekmaa0batCCjsdeE7
lMXIz2TbPvTObs1pm5mRL07au9xc6aiDpj6ugUlcSqQ42PL5/VYVrnzlSy4FSBcl
lV4Mm+Q/qOHarN1szKQ2jpLg+4hK2NWV+qCaynax+Eqjz5A+rE+DC1ecKYBWIesY
pqawiuAGYwkkggzx2mo9EBXDDShy8xq0AzD6a7/ui9GkG0zsDYwa209NhnilbguG
SfJliGhXgb4aF9GCnztJ8kxVnO4TUQ9Ol7OIKpiYQ2lgnXM6N6iH4XRORKseAKQG
Oxv+7IHtldw2r7eXYHCyddHp74h6KL2ysTRdQGCQNjOXKrXKkCu7pxDYixa2EDHL
dLnPtYAiEG5ASUX+EOxEufyKUAAN+HGuouxoO+qFS0LMTpeyVJmsAL0Uoeiplwwt
yyBIoZDn7TCOupN1zjxjEAKH/UP2ox/P+5xV9BxU1NU11t7kREOOCHpqve6gOFOH
hZU9hx1XCSMPtBRn18bdsU1cOrlwdw66IwIxkz1jINq0GfM4tdOEnXndaL9prJzF
P4R9ofpK9qNNNupdVewtFapLYA4o9brXAl7KZHI+fvM19G3fJmLIIf/B6OhTNKmU
RtgSBb3ZCSZTyKlWz4SLqwGszbk1mM6FTlW0Jq4a0RNx+p/6xkkHVrLYVnLGM2r7
wHWUrpfnb0TKD2hU++tSo4pQZvY/e1sPBjJxiynSKzX6BoC5SZ723dhxC8bAaKgL
jahKn/SO62chd2EnCT2xSKhfxGKbMB1YVTdbDe3hNUS87GRp8YmQKXC633a8fGtz
jsFJQbhEewKS7V/h7AEWxqAYeBJHUNS1gl7DS28GAv8bBaZR2fGWoEMVqXX+LNqi
024/IhOau/POgcCagm6t2wIfPr34eR+72vfitrgnU6B91AA/S7jbOL/Y98arBl22
2cWZIbl5YamM7hjLUP3CDZt4UNpNTVb21x09xeLsb7hGbO14g4FE1ah1Ae9oKHYH
1Pmqn1C5cQ7nKtDt+ExbswoXDlR1RdbifxCWy+ds6aBIdDPNgQ0PuDboVZsoGG7r
IVzz4la+RFVnAZaEJMIVW/x7k/sVZQlPpp5PTtJ46n4KaJaPS+SkcL4AQTDTxfSf
qsoS0C8A1nJ4UYCWJbpl6DXpE/k22KTT63gsiUbArImoGobX22+bgKvktsfR6RHK
ZmZkarfeko66UMxdlU6QNynrfFa/X4CWjIRNgwBBjSWNkqqU2VM0X9pk9AAd0eZK
ZkdBJMDLS+2f6uHasiW6MZaxfTRyAap1QhAAuZ1zOi82nigsglvsYX052XrI4YKD
Mal5hsF8QjUhGhoMK+LYEoh2ptA47QkSk1b3ZDCHUqihaUtkYUgtRKRyJkwleFxr
16LsLXDPN+Ift/D2DR7rghWGL1ZnaSW9MHwsb2rwEYMhpY1YUqxUuGx4BvfYw+Ig
1pvOljRbsoUYxyon3U6p7X5ed+uTopxi1qwSP6+5n44OKWhFHaQC4jOJ7CtWxMb3
/5p9YnpOPBfDMb8Gl47pX4uG3j4pTZfxvFbNrar72aGEqr1x+QQWL8ATKd6Q70ec
okCs7eutUspkuvynvCIg/w/lHS1d4/WeUMUlfno6tLwu+GABrZ+4uW6BsQ33EoJH
o/QxFyTEcR6ha+f7tC6FPym7K6fN325Qm9sugypkLekLyGngrVckZd+U9EOi9G09
1fFWKQJxPZ9r4zXKgKLjX/QUjEo4359d1/iULi/5RACCZFIoyqwFNILGym06BhSt
SMv7BQqWjAZQgwb44oJZuWUz9MGaFiT5cpoeSKy78RHLWvD9p4fvGoTqqZua7WeT
fS6aqqaWJgE+nAgzDAZ82DdgdBzvRx4EgYP03dZoAv2u2679Jluke5OnfzjznaNu
mAkB3KqyIrC365ZKjR5LpparJnF3FZcOxaHPQ/1oGISsgchThH7cJyx9lYV8Rkyx
ib4MxdSP7yIT/KGOpTsRnznnY60OMWikjZ2o43ktjynZjAB8fVhh8c6/z5NHfid0
Eg4utvq5vk4zpOkdNG2JaP2kM698Q/Z9c/cko7yANC98YZG8oyG4mwcpfmYTKQ79
+X8Pnb/mvBPXpbFO3adh+ktS8ZYDJ8ztq67wjl1YnG/djJ4fdy6NN6USlj98LTDW
H38NAWaHD2L5MmSacY2ju/NmRQ/ElJ03bNxl8Uzi2ZMMpHHlfK8Ou17a9s2JGQ0k
vHK57KOrU3q3usEEqSiisa7QxQOxKADMeXYx8wVqokDyQM8JQsx7HIJa5gOG/5vE
zH0l58WInYbxT7msIJ+XslOY9hFuXYkKC6qbk1QsBkbAtJq6rq+RjBi+wuUVUqej
IflKP0aBfaDmPNYV1VQ10NnsMxMbU6I0VSOZ2oqR6IgsJYG6NpK+qe1/oRVEQZh2
JDAWfSechZrZM2JLe8g535tWfcITDNEvKPi7Er4AyucLopDueybGXTVQ2RfVithc
zQuAodarUHMWgIJ5pNUum4IvOgXp+aXOZfBlPaDfA32U6fGX83l4RcdXOHeCyO9U
f6gLHBt4YYWvzymuWYZuWC3f0vL9yGeXGGc8T5/piLZh7hQPcQgC/DqBrQ28A4Yj
eKDy1POTYJ4Wgwr6y3J/ic4Q1xpo0IJA7nh+SxWeyLm9mZINA4jZUMsnCM1AZrLN
b/4enofmZG/AX644VBayjSbdK+T7BW/Foh4TnY4v/6MWexpdC+nihFY/iDnJgciT
xiUStCz3J1os0hNyeI79mDMyFPFnVw58a4xgjVYjkVuwa/+AM27UyBHd45vXeGlT
yzrl6QA5R7P9uYXJe52GMieCfp3RZ6eMmZlJdxuC9ikv1yikowjIo6Ngj0FqrzXO
xxyy+x+frEWOhXzlwue2jEQq90gStswfCJlHcfBOq7F6OODwUBakWzsxqFoPsFhB
zQPxT9hTZHcbuAB/VYcM3lDuY9oFQKauatIwi064WxXBvqRFJRSjS7jg2YzklHSV
NOG80aPxydU04JW0mle/JpOA1Vbtd2uVN67e4+Dhyc3IT/cthEPDMMx1wuMWkME1
4pXY3/dVncOxbTc8xSR1lM2z6HUzE+c3xP3WpvFBxQ4z+9TIwF+HS/rz4tPwCM28
8aDtXqQtNNVX4mTv8Tc3TD6IvryviX0MXmUsi81g0Do0SUIUawYuAKEpGsfxwttK
IelqIXzf60K53yMe+6Tr2Fp38bRs+O2p5F8Py+O47jnFm6mnrZUKX8ASGOhYpjxH
yzj/8TOIPTrSdZxWe4a5e6iWSovkTxC+DW/fmgyPBsq6hCOxnH2RQ0MTE1Z0kMU5
q8rnbgnMIfFKKdeJSibfOh7UsqXQ/WMQL40PyaicA8mTUs53pXSnLRb1Hdkr3Kkr
XA6j9eJHDxj0r/IwMLskWK84z88n3y6vPQ1L8W/Ki/4nkPrE/e6RAtPxtSFEgTuP
R30HBqJrby2W+xYnEmFpwa2Mz7d94Wj/DBdQSGrBU4K/NvgrjQFkNBJ9HYK2fg6q
9m5U6E7nEzNhDNta+VXClqeFdBDMvcajcEGQRZMdI2DrIdsUVRgu9hi2qIl/ZmHQ
bnCGS5/2guR02jq1YPCZ6W1Z37WVuiXr9FIkXYHSKcF1cLAS0RDtDHAWVM06ZiIN
3JCCbF4Z3+cNRel692RKkB8TGrp94YwbO/1Bex8R6FUD6in0Da1O2NmNnO1XmY3M
u8RQSPbixB140y9EhbrtYEK92PQqfyoXZwutOk5g5PYQLQqDzLN1BPGR4laC9zd2
KDUC98X0jltEDZXEJW/7B71vrMc0S+rZ7DH1hGT3WNF0NyRxaAShnMkVqBF0IVA2
RWR/a8PhJb0vjWJxDaJfcYKylsKggFREAB0CgrsAh8RYSi6zolPB9wgaZQfTkkM5
pWAy/Ndectdt/bpW56Tze91KI7PyPX1XXNBLaavf0ha9F9QmdGSNpd13tOvCHtJb
13iL0LOFoWbcipHuF6WLojLFMdKupUou14cm1OANdYwb7Ohpt9lHdmRM4G+bnGtT
Mk4JsAhYP1b0cdXt5Px1QjkQWNal7e0QuHqlcfsiUmfttsaU5RvmWbo56EtGVR9E
LRmuu6KKz5L6u8XqoXPr5gj2Nz+XEP5v7tLIKq/Ey5eOVuH1mw7bxo5CQkN6xoJZ
8I9OnLtVvRJG+AO+wH+7Tg6c6stzISFi5v5AHAuJ+KwhznylFLYewPNprOTlE0zp
9TDr8t2hIl116hVVt9dmZQSHJupdQ0VnJCzKFxupdw6lJva3vtplwls3Cu71MTOC
ArROa9ibHUf/zSgNN8kZlaFn7U3jFoth/+zNl6OAHUQzoPqQ3d50JHGYXNJT+75c
Wd3Ospj6452wEhYf0euVLfwfmIsCdHIdZlsfcydfycI8Hwjn8w5LidLZIRmvvD08
rcfnIPWhsPPu51m02KmeeuL74wl8n1nOag8klPVSR53bjBPzPE7TF1d2Xxa6EmNp
lF7i986LHoKK208+HvIby/gevgRH8gmcW21JICyeOZ2p1/podzs/0LBxEl6TE105
Qg3exmB6YhXji71TFjaYFD4vrncGkLCr5/jXM9rE8UMzKNfeQcaT+nSbYK3suqgA
YVxL/RGUpuWc5jhT1pKnXuDBGm0coSFQhFEyWjk5ag4Vk6c6sP+w8i/VWcx3rSOC
Essi8S5kt4LRISZFZSf1lvnMHLQ3nfaHy9PCFz4Z0hb3cLLma6/FDi2h8Ag4Y2o8
vtrrOaJcIJQE2U1RQuU6u6nej8eYag8Ntmk+G+jcTSu/Xhk9AML5cZr7U6RR+Nst
ChHZda6kXaZVIZLLE6dq1g78RY6/JX0EWZOuy2KFYuRQpHYOU2UzeoOLCz7jtkMi
DudANM9OLzfJi6FAHW/XjGKeLsDyugE76dIDl8H9blVCFiI1z5jp9ZvlwGKUA4YA
KJ3B3POiCNJpqqBZrhiWWM/sKmiDiduZZB/EBOjQr+iLbaRpcLB8Ar+lii6BDewQ
3GDvhzTAlgO0hWmqiI0bxsI+ptGLILifn5KGAZgh90Rdkuh9CxsaGosmWOTNhscQ
jPKEfD6/OVMYXwwSirc8p4edw9mLgNX0KzV2zAaG1ETK1OY7QEl+EQaLooYKLiah
IoyT1vdH/GQssld7Z2JpVWPJMyIYi0fOWr2grZSJ6eqwHVy4VjinOWtGJ7cuSF94
z/YvwCbZiCYDbUy/vRihmkClmGuvN+HypZxQVSuby0xwknbX8XebM38GfXPvUmfJ
zUcF1y8D5a4SYXNZI0N8mlXUSGavo+kY0S8/grk4FfGMMEN4guiJ0wkLAfOinvkp
/Vjr6hKFYdL+J2FLJ36/4aZ/ThS90zIJikLXRS5uQ26DnpFUzGbDqfdkHDHTLnVz
NEpPRrodOtd1NtcZQYyU34DyV7RGx/SsUPvX6FzNFeH73Vwn8zQ6WWaAs4hpX2Fw
/N8eUbofIXyMGSCW9B378DqFRzVY7uH6zZx21l4SYqXy7lXfVaTGfB04fvyCj03+
TSlq3osO5h6DScRMy4gL/wOPGeRn3YfIlbU4Y/8moKnxhcXSrfVTdDmW0s+j2uHv
Ow0S09eZmKtV6WMFlESMGu0SfgxyOd/k7Y8yd+/J1oPhNThJMrNbeodEYsusuJuX
o+9t7rUMxSPpOcxT2y6crYRPXsSHEhtV90jMF5SOR13iqVOuLzq1C/JPo2DYz74h
e9nM4zn/VpJVVbAO5WDjBsHqZBc8jmbFt7TlQcVq3iZcRH/nJmzwsu2IvOi1DkB/
IIBN+1cgElNqXISQ503AwNyOSc5lTHAR4k2rHuUKt2QlRO0TLUGp6h4p8yQ5WLKO
gOC8pFVsYYTg0NwN5zK31B+T8T7kHcd9US25huhmR147lg4d+dFaG7uD35eMLiZ/
oxIdaCOMQBitWMN+DM0Zeh+Ty88ZBp7pLG1austCcrZnSx28dWkRVmhMa/yCdejz
ZjSYVcFJWwcW0JQ9TbVou0b+B2EkolxJAG+aB8mfsYm94PKUQhd2+rfv7ts4FQG5
oJqVE1Owv0gjHynskXXcmZNXIHmD0V+fUIMRSA3fb0eyhonVkt5mYRNAJc6vYJ8l
et2cVd8zYvH0yPdOOY+HfKE61Muu+WUWerF4A7Bt/d2qVUkgfyuBqctnWemBUazS
GG078JcoAcCh21GotaZGu9lP3qW46B8ykuqasi9isVk1JF3AfFG52P/VBLVSuSDi
zok6uXyThz4E2V1lWoaAd1LEbxbWzm52gmgldUXHNUtmEdmW4xEOrXGz2H5Bv2Yc
eeYylwESG3QoqpjNYJW/FRvUm030zlLz0E22isfi57Dwq/mT1zjEP6hDjWZhQh8Q
SKeha3/aTmkHCHmtjpcMAy4AAvOZnz7WAq32J4C2n2xxvKZ1LM+XnLkhonvDsmA8
u9EbxIZaZmbf0RsHJGwRAZAJE4BGiJQqCmu7p+tu4nEmT2IfUC1ny/eWRCKZ+3cN
18oaxTNWRo6+PDnwSvVzKCVKZ3Eqe6UhPZ3O5/Jir9yogRSVyqLN90onxbZ8n5C7
wHj+VYa7grc2Ve80+2nu1rkD7AaJxOptO3j2E0uiXLQQdlbnnzhJgdx7sQUKE33Y
LeMCuyRNBQUq82Bed/7DbSQ0yZqQaFsAlCGKPckq+cY3wcah1FBO+sRnynO+wnaj
k/ysjVaQHj1f1OUkHCHjhZDdH9s1Jl4YXo8MnvYNDASOqsfblh0nq9jWqZIbrHhK
hDzsay33cNpsCo9Apu0IHD3gtpdKIhJbJn0yvNVjt6mkSVMle56o/7msJgIZrJZf
0k6lRbRbvvg+WpKvsIfjECA5pInZaXQF2kop2XVIVWSO7tsWmO8DIow4M3d4e7Gy
/4qoqqc0EXkur5hPSdgjKCePwmLu1CIm98Z8HZnlD+OrZmcpHQJ+ozR8EgM0l42h
iE3TsXngGxtOESQrv9b6YW9zMvuS19qdRKklRi1JNuoAnbWWq5/zMMDACUNVCgtC
RKHjLACxdiDkTVJRRHT5uxjKPYjq5GvwQiD5PjNiEgXp2cINzuImQ4hy3RKYLvyu
oXHoPhhA4vjtrVtSMOrtXreNj+PG4CSa72ILTNMufZWL9TLMIlXdBohZlSdN527D
eOgls+M1e50fHjeStjV9WfKdeU4HHq1s/Q4ckSKk7KXV9wtvzxXzPUfkRSn+V+Z3
2eZoDDlHYtensW0ACgglY2pJoiZ+TO0ih9c7u5DUDtF+khaY9dJhiosdUlpugriT
2Ggh0JGZblfzEUl8e3QFaiBsq6LSMsAyqHZCSNfzMC/GryOc8imKl5nnWeuurxBx
65jlXw0AgKAnZUfc7SuDaKRuDkk0IOehwcoHUhW3u8oy/VXlNbjKKLdiqLBZSvhY
viyEIs6TxpJ8LcFfY+diDc5AL1a0h4qlJAdsxz3c9lGSdnKFkEcop6RIRHwWt/Pp
lqFkBxRSMmNJXLqBL6KwAmU5FbiwkL6a7AZKwXIk5W5ZYrKp52KTkyvQ3hQUg1T6
O6iOMcHJw+sPzs+sfhO4XHX8mYBi3L6E/3SgUA6H3s+6BSIaBUFNBslRu3hVXRaj
D4Thv3G28K4/Udui/n7jmMATooKI+q4RNeOAYfiH94SchZ5W5yAc74F4Y4F6xC3t
7/hxkRSuro+2NtEM5UezLBJaNoNmeTIZYE73zLq2qCWo1IsefYt3BCpuB2AROW9F
0MBf30wKo3dSbAfI29D6/4pkbEkXnPrHyaVLwxzAVblKennxdK7bGbNcMJu4abH+
EHr8rv+337imEBzbizjK/tBrBVZh3cGt1yUWiSBKbyIvUh+2sXG3T7MJasRpjEsU
K4rIuBnHzQODjT7XcSnHpeE5xbFO5rNUiat/pGRGxLm11VLfuAgda2HrkPnD48fK
t9s7Kxt1v9ZM/H4bJJCfkihJjJgoP39tMk7T6+hs5PLBvbysYX1UGj77pt4Oitgd
1w2HKjMLh6hMXiOquZN4ApKnaMo+LA1hnk4Q7OUJJCezg/E3UwW+mXvc/lqM9k2R
+btDljJi5gzHKo3QgRrojYuQxZAbkQZ78wHCTZ6DwKgd1SOXfZC4bxG/G5wpxxw6
fVmR9e0cvlIe3WkWofNxx9Ac9cN4J5eup0h5KBeTEzRrXvMPVhmjuDbuJW0lbLI7
wwLEakVuJ39oVlZxNyWE9DQDvzCfL48s/w/wxAvNQVfgI8PKl96fvd+fK2DKwpfN
jPd5HlPuQE/hXpLQNx32u0B4OsRy2TNypgvYvcFUDMG2Vlfz8oo/dHgWFUsio6+G
WHAJV/y68Pt2heLvIVLmG9uyzpa800EHx18ElrBhkkrVHQ9w6nftShuYkxZzUk3D
Ye5Zz9k59VMXC6EkMC0rAVDBWTpLu+t+OH73VHdwbXpBvB/q+TUZP8PSKJrYy4sn
aqmdJasZnEjDAxsX0vWNiJSnMVkokj0WI2fncnMaKFv3LyG91/v9YAsch+OpkVxZ
oBkVjske/Ck87BB/4fupPfknOXvdWPsZVPCJs4F1ta9WZoBg2IT+uWne2MWQKI3j
ADjxyGYT57xEZr9J/M3JQvdBJ8/qrTrzJrMJ/RtKMJzz1+9dTzUt+u956j+WOqQO
U6RBTBttMX4N20CI/0GtFTKEPoyDEZ68LrEYQJOdnSyXTEIZoA+lmA4rpcdUix0L
tu/jjxmaPlwElpiLlCpehGAiQcU2YZgtykd2yCk8+EX2Q3x1b3WlyjzaKPtWn/+5
1Yc88lITyb05P9m6AwrpByMePiN6qEYYZFJP2mhkRyeUM0xi46TOKWHmL1YDE+88
2iQ3he7emPaK0PUCMeLwHHLCCHvG2qGhylQRMwhwFOTbIIvwWUIqBASDjSw8KTCE
GFD8UXRa3o4IbswT3PaD8j0P9I4KECC4ArieqE1u0FM3shU17eIcQ87I/F7qEsKl
Q4RL6ulZGRokO0iSv3zr1+5eX3WdTaGcYaIjp3qmmMOAUN311IQSEggYJWPqO3Py
CTfWVmNZBV3ZkY/ZOIHJNzr2QwfoZ0A9K7a1Nz64KfArZuXEu1mUFnRT71efcE2l
5op9Qa6LEY8DJ6xxPRMOXYAzTMdoOFgNmOvElWaMBGFRUGFE28eB77b7eOotTh0u
BZf8pNGtt+FBKL9WAMYfuX2/HvehhXzMM3qhG34bw8vYqqowqan4taDGmBCOeyuB
bMiQde0YID2JXotpV/EKYENFx8UVgYZ00gEb4sll6bpXRXsRMiHBTBMCveIRwnCQ
mGjvpvn4vSC+0TlzV81K1TRfb6NiM1E3puqK0cc/N5Os9MgcsOrGmfPJZx0/+SwI
iHYFm6o1QrsCnJREZG0bd8QWPMm65XbPwEYYa6EP1VSd5aOvBW8dh+OWNRDE1+z9
pd1saN19tEusCEmiIGiFKroJFkSzbRtSDaLftew0P8za+u0kMsXZKbLHO1gBmHiJ
ZUogPaNmgjlPwFRuAs65s26qV8FVpxrzt0OyBGL5yd0gQ/Si/N+FlGlQYq1UA/Kw
+gX6AQP0h0gJqwz5TOcmZKi9OdpUdVOpMH3PMgtJIcXAU6D4Vx5nyKPCiBGcJL9O
KidsdfU8UW0ge0wG6ft3lNnogHHSBYoFJgvlFkHG4a7s1OQkjb2qbpDOfOk0OWyZ
l13wdJfbg+Is4EbIyV0iD9knQTVgZko5fvbUEAJ8OxSgmGifP/EO9iO2M+HmrSKK
h2Te+0p4N8IoBT/JjWwvX4rLb4gKkWQO7KFE7T6CYZfwM/0MVQWfX6NBiUr1J2tY
Kr9pAyodqCfofs2ysBFUJZxqJmNGk+ICwmgO10HMXDtW2ES9KNMX/BthmJauCPHd
qSMAXVFxR63VzJvper7JC1CC6wA+8keqsC+YTLzER1JoiVq3yJzAHGf11fc3+nC/
Nb/1sHmra4nwoBp/i/eENFwCsq2ekBVKcJ5rNdzfv0U237CMv5TUOLMb8gS1wNfy
i6u/WCuNwQ7Y2CoSt10EYBXa80Cx7PAKrKma73CVY3HfcLEJ5l1nYjUjygUqa0QG
j5ir/zPs1/OMgfAAL1t7sHlzNe0Ygj/znKAWJwXIyWI6x7iSZpYscRW6316y9+RD
ctphKNYvXs0eN2HXhExmIjl1gwNe9OBg4KD5o8LKAFbjzKi6Kek/Z1haeAL+u3cv
fMHgtYWSnSLM7Jk2Ilxf+lZxoCvLEULEdrDnY9BBbltLxPQdXfTTHBSNf0b8OZhj
nJsNdGoVfppctR9SmmPpv/+M85uAJVDcuRXRXsxyh0hXcgUyT7OFreY9tUgnJ0sG
pM9/66RMnBNKjSAgZ/dv1YaWC2pXrHPOmi6eEWJUobgMMCb/SmFPuAjt7b6UEevk
DrwJubBUi6mwbX+9AcVvTGNUgKio3On3j09pjwFeQFraeKwhMNzWoeoW5IrDMjc/
eLPqwl3gvrnOKqKCcZMeA9LnpzLrswpPvPXlnUVY36B4T94bAujAxaCip8Qu5904
kHS7NIa7JVKip5C630F2orDt+Ot7G6Lbjop8kJi7vU6tU27Rs1QI+TX3srfnI7yo
yEeEc7VZSJGp633gB2pvxeHzs03tpLSqE6wlilzYKgQf79K9zPy5ADaBqRoNbz31
WS1IQZ0Xfd91PWaqEMkRbA3NdLudBKXVvCJ5dTMU/V3DuZFL1/7WiGceuBtUuqdO
ab/xCAGBxZMp/NkyQAnHtbt3a3x1gYr5c9kmmZM0CBgTAC2DcOtK0jkIdm0UVpCr
x0JgQ/FsbiPu+vVERyOKJHLMYGzedEImVZNkZVRgVlf1PicfbHVKJ+ZCxRKd+mqo
9ddq6+6cT1W4TxMx/+DLtVxDPfWr7AbAzSfmtuWliAWiYx/5Bh1M1m+Al/daxR/7
GKefZloO+Zx+Dr4YBYPo5qxS0inue3WoF0InmJi1qdqvy96Fw3/R4GXvvsafzatf
XnOaYK2hh1t4LfRcXMS3cJMGfTWlxnh30kRT8niZNYTYBXdw84EVo+yJ1vnPG2j1
fzZgZW2LYA8KaSNTaUnBNuvVrD7pwblmqATN42e/2gqIpchKulSrgXMEjz80XW/O
XSvVmnyBz4hO2AQHuci4DlNapjOJY5WSL3KFeTCaQ+qQyDuBb9sT95Fy24LHUbED
BxGINAWXcKfrDBFiF2SNyGaHYcdnj7W7DMHqQWwiYGoleJCuEnjhzbrQ74TFHe5r
QJ/As6OZBiFFZK0Tehum0bN6lDqy0SaJasAbsjX/u61xDOqrv+2NxTNGOQeXmeuq
wO2ovEBPhcPQADZYB3bmcenFN6OZBFtQsbWtlB/3SfMtoWORjnUlXd/7GRwKS9So
PvQrT9PHG7PJCfozmTgb+feaFFoTvW4vYQ32pTHO2ciFJqUZ0JBXX443hvqksBpG
yj6ZUYzRBz0zHNTPPQ8js1CvHiVKVpxkTEejlZTCycZoic3zFEjAWDoIYbHKSuDd
WYI795xdVFXonpBJsUL4n8AJGno8gRJeXB9DsNVa/5DRyXuntvauIAm6+zB4Q+KJ
u74tddRcLPpM2WHluwrh1SIy7T7A0VEFc5IfNxoqZWmx29wdpF4D7DsuXuYOlmb7
oZSsYK585WqXxzO/Tr0hzEsI+0QR0GZ990jz5XAg95jbivZSx6QRI49n+pDQ9xGn
2dfc33HqSNXOu/gm2IS7J1EBJyduKkY789p+YzihrsqZelTLOYc2vohSdObno/y1
0H6d4EZ+9A8ohxoguhklRpuNjJ7E7HSHjeLISvdBiSl6RQbpbimZXRuumaeP5FnG
wQXr2ykKjgDgowdEKt1rKUIMl0k+F4c3TzMN9FEFth2GCDupeADwOFyiGqq/SKWf
W6p7hiGAEgKBA8BjU5N/yCj4LMXyfNPPYk42P+VbzSwgXdAYGHVonoMfo1N/Tuu1
d//seGtrNJlVkV2cex0r+DqlowCA0OSessddO/AJlMQvkZ1N+sOpNExfEJw0Kd9N
0ZLIrihCdVNfGxn8y9LHNfoPyVUz1131m5d/VyqqI8f2uK7F4/lDBBIsDkm5RUWr
fTwRl7V4pb0ebJChLLES6xosybvnqDaGz0m9HjmlvGXKpFXfjEipVCBhPIxiutyX
5Gv0p6IvWhFX8e7dpDz2CQmorB1Q7OwcoiE0RMly9eV4r8s9RZRUDblpujd2XAI2
kiLANcasfwsU3qN2kqP/abokC8dOLXvZPete+zVoze0To+bVaPjdkldzI4k9dq4C
Tlw4KQ7TU7hp2AY4IVlsGN78Nn9DFpQ2Zgkx2EX9PR7LWibKlc9vhmRWqjeJdIrX
awCs6FcI1PcGc/e2mCAJ8e7ezG+vI20uvn6z36h0uYw3xvf1lEoidKb+KpsaT4Ku
v9KUUm5JaKtf0LQvEzjRbR1QUloVYM+aZgop085DyGvfYAwmhJvWFWfNyXi74MLf
k6jlwwKMuIbhbENKmdCN2HcvySBcvgTlF/sUN4nSAOlx2W+cGjuqnD/MZhfz0Bdt
+ns7YYfDms8arQROay+PvJhHD5JKXPhm3j8Gg0ec/hxsrXjj7JlACERqvrL/rIvp
B/Zecn2L4owlW4z8o3zPqc4lnzXpFYZG1RHFMPTfqbSSUAoscbBImnxt6hiOHna+
/NHJXUAGyPZ2I0Yxf4mFD5AP1u58lSPHn/3NYTigxlAEwZvp2WpE67yc9TWD6gpA
HnBI6GNKrqzGBacqC3uZErrcFBC29g2KyvCdI8fDSHgSwKFIv7E/16SMZn+C1e5u
YIOpWUylI2Daicz6vRXwngr+0GOPtKftnwXjCmMSUsRfzkySiQpUH1mEeVFmWhyG
B3WkShY8Fet2wq0D9wvIsUuQodR3MCav/yychXLcfK0hKecXzPsrYwm80Sqa/tx+
vrshbLU1k85nQuqY30k0nqoSIePlKep2Y/wz4YIgVIfk3NNZ3qydjwXGFq8zgmml
tR+VLp5dHv5r+m0tcuOZ8K6FEK2V+ytM2WiXb7DRu+dpZVnYeYi6wH7wqjL4L/Po
SUw/r1kHgvHnnmhoDc+5It9No0CCbCBnGnROZKs4au7zCG96am2TlNFxpI9DvLh0
h3IrATHw+AVgsvB7bsx5mccKRBW9QQHI3Ue+quCUhEFHiz2ld8sg/Bku/MQaUBVZ
akw+3QAmWALFHdod3ft8kwi8dhDMyFitdKx/pcZdXwRcXqFqUYRvsP6xpvur/GNf
jcUg4S6pxQpZaQsn/+fsy/wEX4iaLRM8N5NG/Rp6FczAqHvsVSVkbs47nrNfWOYo
pfkQZGl5P/ePn8GNDaTHkJG1dj5TlIl9wlyz6j1URGYgVGsEI8AzPWkkzHy9InjQ
ImsAnnIhIvEDtz6KJMSeOMAsDmpQoYT2iFRh3HepoZ4hFtiaZC/HsxHQOuHjf9uP
RksGRXXoXzk8RM3YhzGIN4qVi3UCRZi8SEub6NqnFFH1dJOlotLeOgLcD8v1p4rw
Inh6IvGTAoeqV/OcEBgZGZvfM0FcUW7aCE2bxL2CM6NOR44BnN+8icHqF02fiYoP
bJUfyU1uXTXbhX3V2nK/Kq2B1eEG1a/OvHubqyVskGdEWKOlLiaJ3nw6LsPYTiGp
H/gbsKIsCvRmVKW6WqIzcNugN7afRGa6aRkchSX3Quij/dF+CeJesSL0nbu4qWZu
+qvQ+9y0e2xpRFd7vUAf8WrGfDquRYxA8bX1OVEW6VZ/nhfKiFkYFGqBDy7cOCq3
HhAgIGJ9zRfAEpISBzP6VuEW6hWxdKFeUfTmQv2xXKcB6fHgItbBvd9/fgqC8u0j
KbiZx+U/GEw8ogEcLESjUD7mPnPkweqG0mSljBamn+5cGAubMOIuEp6u9frs4D3x
hQcRagz6b/D+QC8Vpr7gRfLiAh2c/lwdY7XbI27YvDKMhNxMxrDT/scuZTjdNlIO
6546uN3RU9s1R4Rnv8DMGigfJWcZKR52LSqqA8C+runEZaZZ/lXZfk2BRCHQJ5Wd
VLPCe/TWRPhHAoMKY567to3YkfI2ou/vdNTlURkgqvqJNcuE7zwxBXTqIJB3rJFu
9PnYcN/tqi1ac1Ctp7f4dSbMjW0SCrzZZh0ZrHsquJ9FEM8fcedRv7y3C1ExGyPs
ZWk/kyD3YbpeiTgpdWKk4920tCYUjLess+iRyqvGd1ymxKI/ycheYwLJQDsaWuRV
dXbuorZQaQA4midznNzLfaw8zrY6ht0bJauExJHF/Bukpz364GR+jKOljYVynLzW
30P1frlnSCYcL0HPQ/a0lnYKL/DbBEeAi6CO5ULHf+0HFpZ9JgQrfZDU1myc8v4r
vCwf1wfz9q/qtUqYxMkN5/2ijTIwDFd2oHtyVl9XzjYjPrSHGKZ+0EiF1nh6wCZ7
xQH8bZBWrioJ99WoXkI8fhzLArQp1xq5JVeK2m+swJK9SE0byLSq/nx1RZ1V6JAr
kNqode8Wfc6+mk/mN2BgSXZNo8BWg1yng1Tf3f07Ra/T+Se+Cea5jcDx2wEn60p3
99eEj7kV5XS4Cok79Ux7CJEqS+UYrQWqRSyQ756zudENOiUPVhPqoN+kGsBFtADZ
Z30XQ4yC4d8Bn4nXiGL+ugTFQ1ke3LVVgueJ7WwZc+omTOSHcbJM7C/EnIZkm/c+
MeZXJOhAuKYILbSLi/xJxh7SrmdX5WyccXWlVqVa1o5E6AYwTLH9g4RTj+KC9NUZ
1FCxHuFzZbygTxiAoZ2ZX9qw5LUk9vns+t2DEfWf7AX8J+flf6Qf8X0QDyuMHvf8
PZeJdKTyF5ob75YJypBNiPEDoU5NHjeS/hfRYacr9MVuzRIjDrspnULA0HRrpN1I
DBYu5JRJwcPv6b0LtPPCpO7MPNW59yxSEVfya3D0rjVCMawAe0bIAKlOhfxE3LNw
RX/ulIZ0CfE5VGl09TzEkcOygmrGdFfIHtWO8KABAotyKLk/CrjvDSMWTzBR6cp8
ra1dQCRjxeenGSgwd/VZd59uXg4i2XdriZXWjBsyq5i8SbpshvyRK0W+fj2OxN5a
d66El5IB+LsOIehB3Mp/iuWRzwe5CmNdImHB+sx+JobESw3TY5pbci7Tx8oRYAJZ
D86PWzGybCY8QvadDS/URhDJYVQyvWOqVA4bAQ43+oyJvCJikiFFOGMkb5y3wyyv
BBau7PKQ9r9XF50RWuuibr3hsf3ApW4Z85KE+N0tAtMlZd6ahdUgYEiq6/B1ZJLE
0cFjce/JvkhKLpm4OcbaSbtaENQDRuISrddFUZgRiG3JjBNn0GPDDkHjwlcZ6Dsl
5Vgmj4QhF190zslsF8OLm+b4IU54kmYcik+g+Nshve9c/KXREDZrNsoQmJQCRMpM
RZ4FMJz7RgVQ8VuNHUCCSPFckBrGOasxuIyuFeEgAWvbWrjNfv1eS0TGqK1Tnq+z
iRBjsgMjH+yN/DSMLOgwBF4jyrn+dTX6Q41nr0NErUqffJpS40Lx1MWJqax5eBXg
OhxvU7cASEEIxL8dMezmB2cguekEywaeGA/0etcpyAXAE6GL1Z8rXuf5E2zR7FsD
xdii7gM1BIc0z02XbfscaM78gQIokGOfsXG4Uds+cmUXM3ALexrCBWaXqhtRC1fM
b513RFIzpwWKnjBfJQtqtlYbxoORUJ9pBooDC2eVm5KT7IJji8QCyurv1JCdhKhg
L7GL6N22SZJCw8fgZ1PZAqjFFFZsBc3IKj7lK2Tenrzveo3uZx5Sb44JyyDtTsNU
8qIqwIbfWeqiRceBFDqG8OpQmjx17ZqISdhtIiq10M/hO1YionA2sbwGuSaHkQvA
1NdgJhaXDWUiG5o+gzJoVP7oaig/TY2TXyoZqFN2N7JuqTbNUcI8Vm11TbUEf2MQ
FwfQGOneTmW4XzXu6DNlww//3tPBVi8dlYxncoTLmY6Llei8Tie5/lwvSuMnIn/C
gvX4w9Gpdso07U6/BkvvHLdsSJRoqnLh49u2N+Ul6vTsTOq7Oa9YJOkXZjxOK7YM
4j0wGYd5PaIei8VtK8/hHWTdB+xInBK1XVVX240Tf4pdMGNw2ZMrxS0wD9ggRgbQ
b39xspxlOWXjhGIOylkea3C2q6LmNubV12Ybp5KjruUBpTo0290j+cwGs5d0vCBY
oqOeHSckcCRBLL2HS1hkkkPA4KxyFpPGtWPk3Piu6t+nJfkOoeEZeizRt+ohzrPT
trFZEB8QZR8wR/eskIvJYE06voBAWB9iEU135eiOxOGHRht2Rbh3/yfh8SWlhbji
M+IlLBmWKfHcNfKzXzgiZw8AXMSIrrsBxQJMHAABsIl2llWKsUKEImS4R2Ve++Kf
T1pRqoLM79rc4eAV0tRYkUUT1KeBjSt3hdeW8l7vEBzWDXdEFNe3F/BjJPh82sOy
5pqU7A9UGNjWFPrWZBl+SmhuPVtfO+yPWA8MGv49eu6UJ+oy6XerRDw0GqwVr99D
tTLTE+NQk9d5zKVRP1eejDD9ZUgBTqsr/Cz/eyEGKrVV2YCg60j4U6IEcACox0LW
ejr+6qi4xdMr82JpYKB3iPhz1u7T+JkKbtoIG9QjCwv9Psq4PlMbEi3hT8tIBNtU
DqRlRJHTmB07xw71Wmnmkw1QS2r9q3TybJAp0fhZLBymYtUrHBqk8ce07R3sGppB
ErtEwO5Yl3XAAvCB9F7PF2krBkw0TJOqjwPRvM9VHt/ueo8WFfpP7+VDC+4VIsGn
XDzdkwuvgTulGi3HoxEWVMfi7lPw6lC6XyCc8INo3G6m4P+Ctl9UeEOUlCWzuW0x
FahUggKiYp3w4upvr2WCRKrTDjft3MwTurd2+uLZs+huGNou5eL2wIMUGk4G+Ioh
QvgqVE0bRcxeun41DO7v63b826dQELfSFNiv1diyeewV7cbfR1eNPFWDn68i7xmF
NOS8op8MqTLFgXe8h0KdJPxryySkoETFPB7k1Z3z1+GTaFecjk/IWCXHWgSTWC9K
roJoFHqFqxAwvTHfMgfQvfkUL2bYsyWyQt53KAy4fg+30777O3Z7sH4YrErreQCZ
527SZyf6AFg59+K8oRbFLCjLA13j1RznOLp8rzDDqlq37BK3NthIKMGmqZpumGoY
Rxgeo8/71179NObFXmkM/gsEzN0A8bCEY85kZyB1Fb3i7AfZwAlf3opFh5UWDImU
GpWEnm0bbHiRhnmpc+GNdZqqC7zhYXw51UPrwHuszck6tu22nML9bpILlm51S4IJ
vFvn8CG+NYZIqSbfF2x32YREMQazCSjJ3WtB8mUWOLsn7+mcwGoiaUmL5sRREZWi
8nZWLqUnGexFJjzO6KRCJw9rldnRXw8UfmkKky6fhYQzT+hKyfnCgMJtKBgNnY5r
UViye9k1hF+x6Y5kso2XbKvd64y+xT1POqQCS802mEi5Oh4phIPmnJ4MCZq2faAK
zRjyAE1YvZ2mGOPxnAvZRZYgA4TIconiRoAHYGrvB1hgX4uQ03Sex5u3YnFipwxK
yvFpTW6wgyP5RSoW3zeSCbvwzCR/iw78VT3PnCcso9OmOIoXTfUzIoHnlBSPWFWM
95zo9HcqqOdmh38epYA6GKAGEBPMFhY5hxipwAwvaB7/6xMgTVLiCedaX2uhn3ly
173muy57q9abrhHnL5xhsygv/f9lffT7TgmFUEIX4N7kV3+p6A2QKAAsnTSacZVc
tnZyvNeqTIj+UWMND7sCuFdgBsAZyN/QVgdpN4OEMnO7sNyaO0Pdav1p/BYH9H56
p6hSDU0TyOsR8r564MLfiMUGmpMIIwREAGURnfiAeTz5YUaHu3Fwc/aaESe1Jg1w
cXztpVrmpeIjO5uMivvMJu5USk9jJKhZHJN/WBqYG3nodGJeOA/HBU8BiXvZqVS9
Pa73ghivghazbypmh25Z3QDK4UuaMa7zI1f7mT42aKXo+q7bCBOF5BrUVfqAb1L7
OOtlWQ8vQG11ZEK9Jdn4G5sTWSzAmpVEkE/reTCgVSj/gGvvqNBlXDuzwyb7gwDN
AH6cOL28mZdhfqHXqbSN8IddrW5h2juJNTkm39QLZZTF8P9kAgKrD2+0n7Y9UNp5
DfYHmx3FBQIjzL1cHozX2MyleGj1F7ukaF9fAaHmWxmOjGpMG/k00GKyC+yK13M9
SzOufLIPktloosJ0iScKYJVmVdVe+tKRHLZX/53423/X3I/hAXOo8SO6RkRvkJey
LI88IiQlVVX2nxLWxLbMRroY9UILT6geAJJJmC3AY7UOpaIULzpxi71FRHxRDMS9
slp2FS5Qw7txaUZbA+rl5SDJMqbZF37rOaFvopIiE4AUPGJbnlmYMwyIhgd4cuIJ
1H/7MCuXX3W9kr0Qy4mJITr73DZfMeCsc9whYBbZTrEs4ONVDc0zrimGmZs/vlpj
PT5J5tZcz+6Lz+sd4ialT3E0kRV+BkhN89BN25y92cbJ3e4fCfVzriXKgeTchwad
lQ9Auu0eLD2auwIwxOJ+0HOsOJ13m8+X3ByIv6LZR5RtwjnaoQomgbgH/+K8QEMQ
54Gk5dAoJgUyL8UdQtOQHVx0JJbhF4LCqpIl+HwwWyVSIUkc32tYhn8qPTCeZ6FU
ciWxRmT902Dw7NfhOu+Zq1X1MDiKDD9IHFT4m8BCEE9RokIc9kyPQzHdbA56ieCB
gRRT33drqWMuBqoZnx7I7C3aAeOjLnRDEpdDDo9q3S2NyU/1YLrk8HI5Lcs7nGEp
Ptv4flbmZ3hysHsBZVM7G8hmWuRoehEI9o0CzEwWSJsv4/BI77i9S7JzWQsjtQrJ
C0J0lZEgCaXuxXzwOrUWnegOIn5c7lp5uXk66pSxOLvKPZY6uhU+5yV24/auCMgr
SLddAVPLpE/w+UE7ZiaMAZkSwcyDJ+5p3OSb6+aSYKlvLbX+fJ7iKaytq9rvxEur
hdgrkLfG0L/g+lNqKGNu4GXHNgmTH8/KEprVbdMPCD7aIFoKTctkxX84sdVOHQm2
xPR3qjz0DW2lGX/kSag+AU0PGpO8dLcf9OqmDHWK7+IQqieLtZevbD5oLl05cNm8
EjRQZImaZQyL9K0kYdznFACM3h+uJzsnhYDGXV/W72T62kh4aWy3QVx4R5+AfqWP
Rzlv8rwmdWB2CtKpkY3RRPOk9Dpy3lqt/FDEZFLYy+0xGTWNC3kM7vZwLkK03kaF
Fxt+3D3Xx71xiITYLQnNl5T1jUES/khULfnRslgzXTq2OCPbu9I8rB7Ej/Ia36gn
qTHos9sY+V+rO7DLHNXVAj54PIQHeuQkxp3VgMxJ+lVP2McHLTblZ/3PUgLRs/ZG
PnUvk7XxiziUXgtehErWqdw+oq8/dyof7soU9dUBpUxA4/GWj7HlaCSQ+uBX4BVB
mK/LiYhtsZQKbNn88UhkGH/+EEA+yaQjPtew/cSC+6gmctpKGVTP0MZaMirU0TR9
tbO20f9aFBaa9ko1BzR2zfOUxvsz8788LMLk4TXX6bou6t0tO9nNQf0o5Qoc3J7i
fcy9RfaZLVKuW7QVtwxhVXKshhey8GnDsv6pQRwsa4A5NJDvAY/PKX1Mk4HFdcVu
s5UB5Jdw4/hGSwkZNax/5H2ldsiBFm32vEpLZW7Z4DTD+4J0wFlrV0tztT1ft8uA
WtAbFW/Sv7GPmIdZOIW0iQHpPrxemmeZGUfgoSlDO+71RQrNCsMUsajVYp91/4h0
6zuvsgJHkGMqaFgNfXgWpSZ2WaE8knsH8HP+zhaQLYgxAGRcyTQZuz62G+v4mmZE
hnvY0eIX8rR2lSOSNtNl5HnNYJqJda3Fj9KpAtJ0mf+CKXgNBTgPJVgk29jhonUL
plh6dEte4ePm63CCcGhgUjxH45BaOknjMWmG6rI+heAEvbhY4sp3ARSusG8CpcUT
qN2B2QnmiULtkJgMg9S0OAbVjZP2WLxbm+Q0s6/tgSL57Pc/nDVukvqBO4w7aSjb
wac5JfiezDk28TXP4KH/HLRGADRnzjgA12uZL0T4fTfphuRPot//gCcumEvrboo7
wGWmW6TyHspxbIZyYWrAQaMTq+fH57b8LGSxyvMxitT9pKuvOS+xu/fdR0serQH5
TLWyiP3avETt3GZ58UrAzX+mTkApJxVI4t3+pWJft2K3OoUgVAX9/ZTmfFTStWzx
o9G9RNGn3y301Z4YqYi4NiZWb019sbkBxiAVJ7PdZkWGDztV30wDdz7oajcVFUtq
bSofIHlopNZ9KqAgHxtL5rJzLzNbNKMT9CPJlQfeqiplFl9lPPrii3hEv6eledNv
jK5Q9gSnglm1DWp8UmmMbLtEEVFZYiHYWvZ54TxQrIecyopTTiLxexvzO5UlXvaS
L+bT/OgcjGF7vM7OnBjGW038lBZbl/F9raS+/r0McdA0/9nu8JYqBrTP6XKj8Fiw
bRkCHeO9Zt5RnwcjWx6We7FlXi+7RKDRwIq9j5mbcYge3/tFephZljQ9G4C11wQR
fiSkeZLXVRO1XQFqgolb2rk2kb+hE3wi/oQIg2uHMfvX5MXaQuuolKuFPjit19s1
36CDzEizXw/MVnZ9k73Ly2dlJrfO6PuEzzvh89YVx3ZGjAh6CRQAhWzfX6Pxng6T
VEMXdRXjrm33o/TBzwOiA/1xqbmkVd3jX+pqgxxllbVYSYLRD4rgegJ6AVpWfCh4
3X1TBqzStT1MqEJ7DbuVWrnb4/aG715mQcVa9MB5AEP6TmIBCFNjbkHq9S3ZgP9Q
5jNjMuMe/3InUWMPebpL9HDOavo5FJ/dtzkT4Pl3iwHA/y6vG7NBBpTgDUBDyAKv
5mv7MyXk0F6611/KDI0b63G/7sIfOnMR0LHmW5Vg9fRuCixTVWP4QobCUpyiANH8
D6jcMuGZ9I1k6YlhDWqGZ9reCHj7PDAm+3zB34D6dWTdzPz0C/oAO3JOKL4wdHEV
b+2/JvezMPaXYeqQs+g1nmnfvtLoRc55WWK/jYI18L2JOgWwAHxFhcL6WBMULsWN
9PmS5wq7SQ8Efkw9L1iQ4xiXDN57sQBkvrkwklhXRZa/a4ZHLnZBlfwobOiQyC95
RKhmyqjpZJbENPjxkkLPjv84B6E7ifvCdszioLe/QsoX3srxm9UuHndO7TJRhD+n
uDv1kQFZXnbSSKTI5UHzhpkpKjZfg5nhdARtKKbDMrvMIkYaSvpOjGjR8Fl6h2wz
NdH0yYBk6Q/yIXE/TbH+pWa1xpSPXkXpG87p6Pja0OkMwXdBlNXi4uy5HCmDk7Ag
F8hyfGY2R3cUc8e4tOJOLM6Q/vdA7CULFaaHobnowgafnYmhb4WF3R7g5tidl62k
eTY+oBoOmmv9ITsrF7gKMOr2IzhoYVE8o+qcS2qoQev3hlPV5wekbme9cJ7FkVAj
SJ5a5O8E0Gan9C43Q/57s8or+5OIvVWbqGPhXfkD+yeegB1IS3+unGrZkdl4LWjR
ACeFaA4OXD0slRCketpHjK3ac+9dvos/4WAztTdlz/liyVp1+/qeQZcSpndnGpUI
B6tF5rRBe/lzM7uaf8HHebXoJ24Cocew0bWq6FbzbE5xAdvB4EIK7TqJ+BNu7UHG
nPd3pTGJPVV+jgbUhHqCMs5chLKSMYHKlirgQv+wW1734u/mgERj/NeCasuVB2um
0RNpdXDDlybEYab3p1M+iN8DOc7bMYCNqfxbTr3a5shtc3b/8LLPkhrNL7av5Trq
j1wxyHrpaVw3p1T+dxOIwgQNxS8riToaidqVMz+LRLPODEeCeu5lzgzsK00A63/L
boLckpVyUnM/u20vDlhznMhEeUD34EZwyzh/NtLzM4TOHBcWYg3j8J8yHq+fRGSd
XSEHEL/vImCBUsUX4Nv9pJVQ42GRouMx6BqhK+8JlYCpX+LEhlEVYMgf//KYZvrE
z0jk6Cggnl0SgljmzCpIeuDau/khs9wTtHRu+nUjCwJ+p7ONyCmi54FiR06NkaQY
5SvKTHyAJ+droDdv1B+koAkF+wZvgF6gx4cNUpnwjlFHzF9F2PV4nNNNNNJpxGgx
rSWgD3LO16Kh8FwPmeXnyKdMqyWO7CAlh+KBTlWKrZ9xUjFx5QX8C0nobx6qA4qC
WWnhxeFAzQAWYI+ztSvbGMJiWoVL/bQDFMCgNYFOlyIWoMMSc5wXe2AKzWYpLmvC
r5tfaH3dbNYdAe2gndaYO0R+eAuglRalasoj3lkvnD3Firnnqvc2ZYJVD8LrY5Ws
5XZCiIL3p5g+5V5C7+H2Qj0h+c4fs2cbi2Oz0FhrgM8l+FYacHpIjUlg/u2HIvCC
fIIIEZatQ+YE0ngsrjr9j4zO7ez942/o5aulFPg4utBK9aLDioqrYT8lWalBPk1T
vez0nRKeTmvUfuWJ3HsAQM6duhPyiX0wmI+jyYPn4rTlBDTDy5ut/6xzvzGvToAp
a9rDgIolcgH4ra38j4JCF9my6Ca9QZ5QU+8IbUc+VUnomfrkn4p47oKbUbeeM7Bi
coqq/kgWUdFfNfmCEgVwsFxHbTficGQR62Qt3imPB3kyZimfmsnPNaAdaux2zMmz
NtpKqbUkev4VB5HouEJx7xmubrOTbqpNwjhBrQg66CZj1+L0lON1tRsRU8No5LRF
EZkb9D1Xd231iQrGB5VoHiAg0ORVn3vk7DYqrDaWuD+QvT+XeT1XM3gxLG76jLd5
qrXHCdDLmC3QkutR6Gg2IvU4vdnSrVl9XmOAKpOBhY8SLl30ISk+y+wxewOnoNj7
8Qph/PP5FYHYsuIB+jvNZYTQoTvV5w5l7AArs0HFwgOo2AzxplY5n8XDKKW+4Sw1
ZOw2pILgf+e90ZMm/eiE+Kleccxz1nuGQT6p0iVzQv0ovJupaC2orGwArUqVFFYt
aNGkfHCW3V0VSgd/2eI1zdkPbXdH/CGbpCWWCZbW44kPk0+VtTqFeY9zzHYdTnGN
85ECOGvrGDr8ldqS1bDOS+ExhSWwrTXpOLH9PZGvP5kvmkbJ4yO5SOt0CLjFkAy7
Mxc/Aj8u0spuJKaxFv/RfLF/R1lXuO1sr2BVK2DjYLIi+DJb4g0MXalM/1AMK1NX
OrhCIqOYuRX+pYP7ZDMyHZ11UxYtx9T0PHuMzxjHXl4l7UemXbXdgAki6ZXH9Zxx
SX/ptu1I6XDXmVLtQ4Au6GMXruaFdvyhlZx7K4xBx2HXV3BRZYaQrGkC/Qg9BGA+
AHsYhhgin0ibI6XklpUUVZPjp+PtT78kg4YjnIb//U2FoKpRyEwQhc9M181A9L1+
ajfZjFlXry00UknIuRgLllTrJTujhwn0qSouxgxB2Y9FsZliDuaBvfiayYPyZM2F
kaV+4EaROFLoyyvzDlcYT0id4NSgWdGu5qmsCJOzlugJfYX5AOKfKDLagfOdGJL6
2DNZ3gbYWXv1wd1hpJH539YgblZWQxCJm3NpzTmP91NA97CgIgSSfQeBRXYPbAMX
yge+l87T/4bCSk19zWIMYBby+EwKzL4ZBh0lu5YK7DyFChCNLOJi/KBBA/njqgCr
FH+cW7O2+xLVSmACcZUc/yr3uWbp1utbLwJALqx+tCwKIGwk7YjNeSIpWI9h05Ht
kKCN2XY5phLilmToxQZRL5TD52d2cIfeuikaT4AJmFWaPgXQW36ELJ2Ms54Y2MFK
TCzZG9VK1lcN/ymBgIi6K6mQXE58Ol/66E5OhdslKzoDPsajjESgwgZNut5rHTAu
rcY2Ky68rPiU0haxQw8iGc74jsrEN2W1oEmZdi4udNnLor1hYIBH87qorZjLtVHh
qGH/qpvxUa+fxUBaCKyVqqsE3UAmoLm30EgRGi8vGVlqWsbrg++4kGeFNmvDZGRM
JuWA5BQnlQyTyqG2rYzsn0ZHBFagQiUc/w/lCxT/8tiqJpMijEo/IfGtg87/u8hE
fDsCqaXQOVpkyl9+jON8l/C3wV65Czd1LO/8I8+NeBUWt3n4uaB7XlV5ZeghFxAE
Vwsmo6U2xXwKL6t7XQSVb3ehC25Q/HYmJAyC4wcQl3BRv9He9IDt//GZA2A85OUB
3Q3AJZkUTv70gkCqjmctwlN+F+tR9wh0WpUcgEFH4Z/BAV7Pc+SYX0y+AlaUzwXu
p1s8ZNUuz8hlc+Fra6pDIjh6fTyYw8IvbguE/CIqCcTcpI98RFX30JDyp1lFa6vo
kW3iWDZBOM8f3gSIoXXzJmCiZv58RezhUiqV/rj2k/7h7Zzjg8nyWb5eSuunYi8L
uot87aZ2wmp7plaJSIpwVeR5jvwOB9E3h1yWhcgHt7lHqSIFd1tb2ynhgtlilNEQ
U9sPG7begCOVxkvar0NDaYws7fFoR5z47qnoGvSIG3PCuRveulh8opRN+GN+V2NI
X44C9zdlophLiEbqqU6rsI/Q7t3JYsQAc5Ldis+wBROursetcYDBGRz+hUkk6chf
gDXHhKYnptOJ6kuj7viMUDkcnGoWqhKVuE+dF0Fe3KkBMd1CaxXIhW4StpULGHxE
k4cfSnPA62WvEpHQYMhlW3jjLWwfU3xVtcl4nV4aVIqa6vOwEHcuud40JYRpIyTb
dNFED3bkx0AkpkQhl5qIfeOZuKb+4zKITOzFtOqk0TpDaRBT703Nz/tXr3FPHDU0
tAuazn5Gg1sahzJ0LHX7LpTYqKJv0mgBEtTpN6QifTQhYrZQQMUQUpYAAqZ8YJMy
SfU1jeCxnVMIWkStcxxy0Urta5FVBJ0PrH41oQ/2/2kG7d6akiYKrB47Qg/kPys6
7fufmzh5yk1jBIwyMO7TrsE4gMnfOy0fqjSC/U39CGFEgraB5yLW9PT9h+5uF6gt
3UifQXOQT3C8V3TitmcchSK/PRXmBPXYghZqeuN7m54S0H0mByr7vqCg5gZw38lG
TH1cd4iVhG4K2c8Mn6pyC4QwGqYhsl/uBXcZ/VKEz5KurPtUeJt2mfC+3gZV0KS3
jiLU8D0ENDIEM5YhjJof6BV8/C7VdsUijUhhFk8bEmdBRtLrVUkWYyGfvaSbU76Q
hnaMqDZlEc37zX58waSyC4ksI9rkmjcOjjIVSWmD3pDc1/hpPuHubDVav9Dcf5OH
U1MJ2ITd71kfh2J/qrJ8h/FsmDpq0chpQcrMaNCoYiga2NwjCoaw59KQViIbAaEm
bNbzh6TssTrggpkQU0q9QuZ0Kvsds3j7dz4HfIN6JNYbr0bOa8YMFeCPiax+Cy6V
yKr6XC4oRT3CaxnWcHgFXgseMuhjsfFbw2X0asrezC+Q9oycVW3JrM0KTUwCadPn
JGH7jtIuMm9RkPYCYSGTND1n47Hqx8Y5Op0NQ1ExNwEqnm3nkvd4ROv0/OLKsJKm
/BRU4+xkmZCvuO1de83oHv1cFHeLSMSeK+iZGY0zrTjCF2Sz9NNpqtwZRZvM01kf
IWuyHS9AoE8JyAl6nLMRqpnPJKtjeDEfZmJGxg9/N4sWs0F8H2WDZNJKLGXJzAKG
JGwjEjs7i/nGKpSMrO6CNO7aGcz2UqH1S7nnSaT9vAqMYV63ojIZPGWTTXGYnK8f
H0Vd8yIsbKEkvc+Gr0FKUH3Vkspr5i734G4c4qTVwgUNtyFg1i8QfdzZ6G0RNXZO
sM+8mp2As9OFJvG8Nbu0BG9hgVDqx8dYPEaOqvaQBvReKC51+/B/BrJt6hQN2iIK
4g/rPTFXDptUyuMzWMlV94zw0kp3BdE5HFsAv/MBqEfFItRgj62oLPjy2n+vwgRl
6rOQT9PgPKK/ca39kablKH9gzR50mbzAgY8nVdHT96gTtA1IChJlNqlsCLude8nu
7T9XokjvNQf5CaQx/ylF70IFaFjvIcYFgd/ZjaqAdchM6pKGBdBSbanL+Xde7lWu
aBxKJO5gAc1D62YDmi2TnZUEIpKQfxMAeEO1gaw8bb6xLnSZ2qxI/222SlKzUeiQ
Jywu3+xmDlbvXbmNkJlRJ9amv+ouDfuhJbXz7q6Z/wx7xHnhPWnMD8lObQp03IfB
grwNcazi07XnGrzZto7+B9L8luvIr7rS4hRPJ7f9Kzo8Nsk0xvElFAUA2ukvrnLu
Ola2cP9NxYthS2upKRYSEL0EExRYSFF80wFQ6yRKuIBay8bk2ae2tKEDVYXOM5ZN
Vtvn5+cKkJm3yqYt/zujcnX4Yv7SXszAnfJ5NCrH4K4iXno5S17hcwwV0iSyUM/S
RArNeOy9dvCINPKjnrS3wskAaW74PZansQdUHksnLVx5lZ45oJQ5YZcJ1LCjuppU
oPX4WqtR6cV2tvKzQ4hnwsRt8pa+DA+PCTfpWwz0jnyLN5vw14axo+UHdL/ZbL5i
9HhBdrZvrOqsNANK7KtvwbE0MjC0cJthyekHyGqIa+sYWTvNXuCSKbypJUSKzH/H
J76VlLxZku8jYCWpgiwQCvYrMPLjlqnq678JJRXrl+olc474MWS6Kv7RraLjcx23
rKJyCWBUUI76tfeMnWSTq3LqBGpyuhUpocR+zplcipS3W+7uxbxs+CWE1pgYKun/
ZrNbBCRAqC9SQqK7FI+CKSG4xAbAGMInPEa3v7NXNJULfiJhYgjyld4TrEASeRPQ
uqd2XbDREvvgMC4WfB0u5PxIAjm7P8I+JPEzQ9XVoQdsPwzWUDIXM5RV//7cur7e
2x9I3JilTTcFwRAH46k/8orNKQH6T24x6Ev8QuMO8fva5ms83YXM+OMdOW4rDVrU
ZdmWHBDjHxwX83sR+CbZ0ePE2Zi3UC19YekNy3Igo8VcW3cn9mwwGEAEuIZYP4jC
WGmLLBXPhL7IR6YRmPQOGFKPj2rgxarrsY735flxvDSnDAuqZ0OP2ED4NN/NgXGe
8mwhOz7s5bp0unsVsrcetWR1Lm3py0/+NP2mH76NNGlnqTEYcalTIqvGdkfc7NhS
Ui/ykqtuFGUGO+5jDq6QE0u/jdbFUjQ41zYfLe8He6OVDytlRk4pWOLX1sMtnS/B
rFaIXlc0Vwh1vm5KTHfHzWS/rrJr+Oj5NZj8JiR2obG5M+26PgAPIiHoCw74VgXs
/o/s+cdf+yvwYRbSnH71lIl8lk2l7c55xHUnx7lS5yRKn88MWviX7SC+nOCP+BRF
YPrlg276yVLXFqoEZ/4SY1ZxxmzFzlQTHDQhfMiZ6WeZi4ZMqWWJemwywHJJWnva
Bnegrgtvsf5GXaAfo9XX/YJj1mN4p6YtnOr/y/03/ohjexKNf64NAGt12/PLxsKl
KxyCAYcK/JGNb02JGgwtApEPwivFU4umu5V26SLVzosrABy596QN76aPMeBx1AjD
S286Dxm4IruuppkcrN/6cxh5uYpBQYCf6OJXzGkyfXvg8rdQQ/dhtzJGT+L6wlKE
HGh+0juPELUKpBxpiz+cVobU/D+A8bngM89ktStJwPrg2Sjq6QeJ7wZ9dQJesDix
thWhs3QqLyRrhO0ofPVOrpQysaD8b36+yJDE8zls0tYJe5L2KnIMIYExJqzkiL3k
XmQ9HjWv/+HpjRxh/L1aCb3hw0ArGG2amswOn/ZRpXzX74tOUAkiNAfvffHKDO2T
KkWQH4VGEJJ0X6woZUXXE2sqcbArRqfoXSuaNxul/LwP9CSJfDpJhYCsLFrDxquU
RA3otDzLuuIh48c9Uzms8h/5giga6Q8REFlR1X04Ii9As/gD5tn4eB6qDtHUBcWK
m7ODobz3+uowpvb8Afjfw7EOfC2qA4UZDv7BZuE2uTKbE3/ZorIw85UQq0TkekAj
Ctm8B0Lo7C7rn/jHB63bYFjOJe7pTxZEZKCH3PjlqgXdbZTiC/a3lB52wT2xb/At
TzaC8fM9mIqk6yMfA5uw2k6xsQM+r71ld3n/YeHuejy27+tTbma9utwcjTSNqrNB
+pu10tz+/DRrZFPVE111OCLtMyRXsBHfkvMAaGmbeAfsbeGL2jNf1A5e10q76I3E
DL0qpijErXghpVMxC/Up/ngkHiD+wNLI4SudoicI3HunZqScb51hHmJrEY+x1ahN
cLGkh7heg8l+jwSCeKDf5XMwRwZV2lwBMl0dAUWP8Y9Y5EEurZhKM5w2gFQ23BL2
Av33usyIlayxOnwVb+GXd3HczchLu4K6/Z9bpVVfIj8ZbPyYPidrqaD7rjFen3pg
F6hJQmfENptz8A6F+vZQBmd6KyBaTscULo1Pj8DVVtpudmWOkg7ZNtBCsO8qsj1j
2mnGbPqeWWQ0sx3fYxpPL8Uw7sXPvLWEJgXHS6ym+/ThDPZqwNrQDPw0AGKHFGsg
QMAAMbjPRMBDH9xNmV+fVhOH99acw3F889uUUvGkpAGbcEClPhyadjWEFg0kM2ea
EybmKekmCnnLXX57vbBUAM+4fwbndWuYQi1FMN+JgWvhJR9u7v51UO9zQmfjNEFj
FN41zwmYbDY1kKXMfh9cR9ikOLYE77ZKJLs2l6iuvogDVQcIFnhk7TTHwdP26qot
9RsYSdPuGc3NqbFmdePVjMsY89cCE+ab+HwSSq1cnJyO2AVHoFk0GDMIlafWY/T+
4Kh/qENaThqTLeUURRr4OIqkD747nlqM+XDOG50MrzwB9rP4FFAhBRPrX1mG9pJG
VQOo+DpOoxxU5UehuahlZqrEvqsb8ofB9RkNMwiLtYZapu5dkS9CA7Z2HFhnElbt
MiLgqV7P/23IgnkdZUR9Gmoxx/mr7w8X5Q7N3tGk3u/oE2cZOUlYpZMkQeA0zpMP
fqLZHgavtxnV26M4cmOKtANoylXrqLKoMuV7osMxTMvWCZvj/vdBDFY85YzeVnod
WrkVxNqBV7EIAA3QZxS2Uu4VJ4qgBMWSnq4gKIh9s3UKIIC05jC/GSB68pjC7Dja
6VA6ig+A+mDdJuGiPTpl6oLalrmWWB509nPW9aMKO7csCFbPpOznaQP37xo7koIj
carWA6MWZUMGsIFXDWGsI6gahm60ZKnvCA10V6xfDo44hraXDssCLIbgxPmNpTtO
UooVeqT22UNOshlhM26CvOA8v0yfh53P9PNrB0DnPraPue1usZxyyO1In7ON2gV5
SgyRiA6pRZFkaUkhMOTNB0YtQ9Fjv8e4+TMPyQN8MJY4/npecMqJeZUQCH914uln
2Dx/e/n6DDNhoHCLLau9R3rHzBDshxHf5URlOnlj+AQMl6jZINZQ0Bt8ADxvFXaJ
9btgiy9VACn4w2sD463y7LtOJpJuopVot8ys9H+gA9WRt9alj32acgVhcrJE9rxp
icBx2kyrwHTwcmUattIXTpO2vEJdscskYt9j9skNXTbrmtW5ljRuMKx/s2T5RcbB
2tUejztCt9cf+Uf3FwMp9ghwhL/suz8M5EZOY15Fo/LUaaboslbCArhQXK2qqsDZ
Uw2Vwfj7Id2BJx53iJw/nNQWJ/zN72BXPZoAFXVTaImMWMxOMkpR+3k4PalCmCLe
7FprvYp1GAgSxsnwEGULcQVlYDSIPav7VQ5FtV+YU5nSnD+41H/8P7KtQ3GDMat9
yIecdSVZivKxUINiPZfeFM/nuajcKK/vLWufeS4lb4tPRkgZ7PMzH8Kdr6rQe/cj
6as2uOkyH4uO77Bf3XDhKt+adHkYn3WdsIap+UpdIRH/dN/EU86Tjx9Hyl20FUmb
xUk6QhSE188I8pOPFnTcrQlzpX7RRhcvjDNXic8X8AJolKPVgF3q6JWJWLjJHR9/
N8ZxHXiHTwJ++cA9k9w/pLKBo2wKYdDs3nhpeR5HcukLYJVl0v82awzMgRaRYV6N
AeVxVgdOpd9RyNA+zo4z2kpWNkyxp1cAZn6Gh2qrIob70R+RiuG8JXlORFwcy3+k
0NPCRv7l3SWIXhwOmVrbs5P27OW4Skca0V12jwygKG1qa/xUCQ7t0iPbZVkcpcGr
eZYAQFkyBIOtSeMy40ihrk2bwFcWxQUqb3zDX9HUIzosnJTPHzLPwCv0fDuenn1Y
HmgbdYiFODqbQHaZf7F/JfhSpCnJMnqIn0tmlHpsZK039tTEaR7UFD5nsyaABsi1
nL7uirMegG0O7hFm+Dtypjypy8CWUkyUa6ZLnVAWMgJ9R77o+BloLVQFAMl9IsP/
8reG4p1NOUfvZRYaUfD0qP09W49CsF0ec3vbzWftZnd5psGUEZcHfsQZcJZ+pLY+
meANGg8spZSGCmyRgmoI4jIp2gnfhPaWz448afUScFcbT+v+C3Ijy0JxRNixzUZq
YCgpT71a9+r7KxEU/tLy9G1WSfXtMY9UDyWiYxZuhMFCSqZc1wrShi52At0WFNcv
gzvD4VTQ96c82B7f01rBky/p10gG4gUBbGxi/hV+QVf4qHFRi4ZaghTXM8wbUKFF
hTt7woGgy+FHiFD9E4pEQ+GboslekHD3rj4Kvmz0WQeQfH72M37QuVdDvNik6cL+
qF9iStqEnJ1KBioxkHw1EvIJ54wfGmXhIcrTwweeUJg8crqnf3Wlo0V5t0So2z82
sz5Hr/rhBgxgCF0mjl6SZW0MWooU8AuGQ5v/hfi7G0zlnOB36foyu4NKyDH90faM
2pfA4exXEBvMNWfP1IuhBVxV1YVrgl7h9eOUyz8EVDabpUwC4lzyz97QSVNXWPBP
eau0gn4Q70ztaqUaEbEBJhwGbzxCsksLwH7GyKC4Iyj2BtxoXAAkIMMycf4u4av4
2F0QHjGYdTFucRo01ZT+hXHsOx0/YAWcsdKyKlTEjdpckQYl7sfDfxF6V6T0eWyW
uSGdllFm9N/Mympip8f4P3WbVwoESOsFb6lgKydY+p+G+N3BnlL83O5PfKOevcKI
FSXTOQ38YTd+T1ztAu+Qtim6rJCE4gv49YlX32K143jDa3wloeCsiTErTrhm3lUc
1p9yjRhre7KRqV6IZfdIK6judpuQJVxSdZqQEbc0ZtGjUFRLJnTx7T7xSIhtWuvJ
w0bfknNU1uFxYLuBtYQ/95LznCudZ9aJi5cIW6aKs474EycGrIrpiX+1X9P5W89r
RAGBIkAiqlwDwKXCY6rHRxBEl71wFVQiZ/usy34cjwIr8FnkprCne3ShPhy4Fg2N
icx0ww3XIrTO7BuuelMSN3eTEyh0l37+GGihr3KecygHcMzAi+y1/2V2GJR3dVqs
xa1cBs3DsCvcMEmaN+LsulV+USeD+JjNJnWK9DPrlX2G7GY0BSbHmuIdY8iJfA0g
FVzkVF7+ALw32wc2lZYLxw/671l+hs5eqW0Hwv84aDN6aciWHlpiQ4hpPtF+fzVt
fWhhVpDFVRjpNMSAkAgeX2FPD6cBxhit9hYIQi4TVmhLDxuPExnSqyv2lUg4kYFs
3yks+s944VX/6WKvfeJHtgg9P2kR5/Ha8cu9Lt/9iIxWRXdSRMnQxDgy2vDhuYTB
5wWyZUCYVD04WslgDJx2hJVWSb0gXhUdkXOlioJb/jzzKJ6XLOkwRErm5vcqyGrs
hF0Pv+IfC4VaikP5ZuYymvp4JdI2gfcWvDXi6rw79rCfZstFN1EofPf8kZoybe9a
ztsz0i7aUaDDxOI1NgESVB46PyoKRqE411aWb/rxVQhKFW5eXsxf0FfSKJgwni/d
bb/Y1jQ3rKNMQEx1CYKYWS5KcE2DqG2Z9fE+1R5IAOaA5fCskcGqvPsDEzi4+I9S
iCHgS0+C2X1uXiGCwzIRb7rCbas7HLckb6VArf772rR7bE1c6eoJigQka6ZYPGev
fMIPJnwSAj331SVx9ObFMcZS1eWeKH82xC+SYYIemrFQqQ435NiTcG4Jq8XtZ25Q
D5SZJ2N1ROXuhA6WFOaMxoIj6R7QzvkqDII3iTmtwQ7AN4tHmD7RkVeaJKMx88Nx
jXwpyE6F82pLSF8K5HQvjzMaNgXe0GJPyDHukWGwjIjKhA+wThijxlDempD/o4QA
N4O6u7YjPUtBJBsq1Ktt9xeM7TI1rEFuhCmlBRlMf7H9W93mqNd1yEloPnd+BvUi
LU5h2JfgvUc/SRkr6RmUDxNMQSrMtCmiWEdijxrDfyb4yexQsCDjHcvoc2aWJ4z1
M/qNhLh2tEaN6r+WJRimf9fMDQ/ecODbA4g1Um674r3D8JcRNrYpPu4Is+1sIs9r
fiK0hi2v/v4f3XyTuXrFlqJPH28EJ6Yv8M/ZPdoQ+XHJldiWe5oabqLTz6tTxZhn
FvlkSo3DsEM1e/WkVy8uZL3cMvl8S9Sk8oer9MMiU4cpUx7hTKQIbSx063wVa+qz
1PNtaGV5qxnNMLltnGwUdmhJH1Rze0nXkfc/wpzBRj5OriF45YymQOePBTU5cOfl
Z3hjLjBJPNpO/j3+3+NvznIGxHnqNHIHLfhXyFPViR+ujj5fkMvNC8RDBr6+P80Q
6nQM8WAU8tZ/J25wSpCfyKQMHabtDI/oGy0At6Efk5JYhkMFouvos+Alpa60YhWy
z5VGgx8P6+htweDimUI5tGUIlGlb4bY3wVWO9soWAL11lLJoYRsu/K3q+EvepoYJ
zrevWRbBuhxewQX4f66IacCq8kclDIJqbufNPluy5W2pKUu3hupW8a15o4IqDBco
VKMX/063dkINECZQNjC2RReOzY4+VhtuOwmn8s/L4QVSSahrHyhaRcYZk/v1Ie78
QWxCRhWC/rVGVK8oCupC1n3aycViy6msHgXt3CKGAokqVSq0iijLrFCAOV4yf70v
BEy2T1g5/SIBj5lRX4WAtBqhxxEspI/IAsGyWNxE1J627Zcl0mOu33ltx5j0Dmk2
KYFaSDDKlbh3xIMlifbZ2a6E/E23XMpekydIdpLogTvNX1AVjbtiNqTc6lQYXrhv
P49/Fx8z2kK/yeiAmKh8H3YCeKcsbOCTDj59FJnae6S3nxnaGqhEwbyZ54kzHM41
Pr5r/B2tCvzrXNcljuuUPURIwT+gbY6gnKTULKVLj9RJ4fLg/Ng93NMeNeftRBFZ
9Ncd0LVF/Nvr3BLpnTL8ugC3b63exi98bR1BvoJz5+QXVtXIZdZJv186tFkG/BPQ
BnNveKU6+SeC1E9NjdOffGz0+OPBY5L76aJvkLbOoDL2Msj5mBdLP98i9BgQdcP6
Q4/wM5EfPKzvuf8NLi9/S5xL8Wyo264jTcLlO0gdmY4OJO1zagZZoC0MBqhJnJTJ
+KX94WANboKnl4mg+i3WhgGKwSqkHJTCv3g7hSKsh75GipGfMqL+7uq7wDrbhtuE
CbRo3J99qFwYEykLsMJbifpHVLPaySsp0+vVC6xcaosmdOr93MHuPVjUE3g4HjO9
ZpW/AskD4AZNGCVrIobYL5LeWQq6k1FNeU7CHZ478d9gqntLUeO04uhiqJG8zCoK
Aj+PXjokk9VQ6oJdcB/c+aHJ8UMoAy6V4R6cuTKI90+rkDbMjCCCKQ7rpY3Ml/TZ
iAQW2yEztUqLV6589BJi4Kkfp53Eo2xLgfMn5Pa3pnNVazPBX98RGyL5gzA07/Xg
AaD9me/6Q7IfgU1GZJWPJo254jBV0XFPUFjq3FaeAJoo5QYGwLpCIu6nKKCyb6pS
187HoJfHEOptgJB4dyXmQ/pePJdZGZF1j4QDRfn17avqEFvFyZ7FpNSKu5rbrvhj
T4z75YOnq61qQNaNPGjTHnurUzJS3tFq+5vxz+8bLZoCFG1znIPWIOT6ef1YLBAF
ARpevQxGk5Of4HYY6qfiE2GuBWCHXHD/N05K5Q5S0u73QDsSm05jrREwJkpQBCUM
bZeYYZXeU+fFXgIYcGcTQ6/fVPLOZ6Y/S6N3v/EPfo6f5xZnKTKX6N2Wbkj2G1tf
Wq8rEuv1PxP7NPvzg/wf3n8ZQH+uELTedGQvRY3LoqlrQkatbSadya7H+4qGB997
O6HHYZR2BvJxtRJR07Tq0dAl55RsX0BJp8EzLpLT5YD7tCoUZT1sLtKQebeZ4Dtg
QDtBIoNgzgFt7+e5fnaB+uwhH8dxw3KfZ9ByI13JAzPTobXJuc008XfezCPWiskO
xfPSwIGsfjjFeIXwaSF0hCtrTGRtweUH3gJtu7P9BdutbkWv4ckmL3MGqumV+LHc
qFAS8lJYFQA6KVgb5wQDvUVem57pULlvufvqk3Kvbn3F0kI43o6YWFiuooei7Z9j
55udkilqsbXir11euOqYP4vOjQd3zwFw3Y9lR1lf7WFsqKknVqy/IJ5bs0lM1AAN
2rndk2yRmLe7gSQXwI91HzNt4rXhAZBQlmcZNfb6w4OTrA18/dB+VZhKSqErGGzi
lVZm3Kk8fDxMjU5umVmqsHUAjG8eD86D+O+pkOtrXteQg+WOLoOe/rRy5zjJxasi
76ax34vurqco0eJeetVmwyWSZ6pQAiQfwfXq3JHrjRuI3VPfa2Ciy0dv76ZkC+uR
WaMbogCuGmj5Xaf8cKt1TWns/XTrPYrKTZhBdsz6PpC/+K/fCAeWbR+oRBoakA3E
0dV+aht0mqApZQXnPOu73YVkBhXbQKwZnhd28Ldh0++N2tEfDfgeZwuSDrkQAG7h
aPDhXo0Ki94dR2q4rRXZbw++isn4jHvHnK4GoMW9jQeIbGPIBM32vliWx4G6IL27
toL0qKKQ5dYMaJ0cFZAmF3YMUSRBaRlQMbZ8VwIAE28HtW7tRHas/qQ/iGGBg+mo
BmyVMvVrWV8zDNo3Nntx/2DwN+e/oMyc00vC4tY/tlkF/SQYPQhBHshLHd+5TkdD
DZfczOpYE30ELI7Hp0kQ9Id5n5yiNtFdG/82lkS1vI4yU74R+JlrO1NkwQIAUMkA
nKLzBIxx3U9T980SOVD/1h+OJ81I29+xNr1CZMe2L+0RCqdsfmYODFCHvEqfygHV
msIN84pufPUU24osD+f5gz4af++IEtHcP3oGKf4Sj2FpBAjHgHwtX16YNjDyHyMf
qWtwab7zgMHeH+GiAsimEkQ7ZupLYUl0VrVMfEJ8Zhjg693pAiIRd/2WKTwAeW0K
L7Z6hYUY7nGFpkBLlPeDE4cDqpzjay2jJ8w3RvETkWaKrF0Cu4o/lPbiqtgH+5gz
bFMPdy5LCgLCty1mtPZxiO+IhTOr29cuj+2vHD3JmH9mpkvoTdiFRkh1uglGfFEa
NvY5e7rySGXDnBSczGoCw/tbmz0teXmn9hkoojBzNkK0v9kM4c3ErWSnNtf2kTwn
rdUrre0X7mJugAXv5H0x7n5rO0qHfa4HiOWX93fAqy6E9ePUTp5Cr/qCRPMehJ0z
+jBuj9cbD5yYBq2T1nLWItjsO4md4ZQ10VT4e4n5lMIqhCIqTMxdmnxCWvsTsKVA
r8HJpGTdBrkOTwEIapQX0A0k17EsORowE9LHZUjtIKU2WhigWYW+2KdvIsBIu4eU
+OZrrHsQm2QVSWmBS5WVay+Rorqpb8CRXfEOgV+trwoeJztUB75gN6xJNI48ZGk3
nn9szDKjIseLDhU8SQyo4ZnqEB239hy8rJzRT1M0utUqbBpmIZH8VZjGf2Oj0V1d
B1xKlVtf6QYxAWW81suJK10JzrYhF1DYBlH60N0EJjaobCajskHE58iCnd35mfAX
U3idcuKtLBV2Cw3jhOw0+G55+UQv0fDPGHi4X6byE7XYq7J7FPoQChK7bvGk/bt9
NYEnGROuvZ/+LRG80YDYbPBIhf70hymprOU8kNId4MZdWifGIeuOTZHxpW0HeoUR
KUXu6CNwuJKhBczNLIt9eyupdKThz889qw4eml0NLFAFNiDca4Ro6LHz0hKgDVTb
TSuj9/l4hS730Z2PcDyfhZYcEGRlG6VYV4bdGBU6g04r/hppXWZ7YLf8gp9ZN8Tb
K8UdXfrK487ETLS7W+Yxz8jRnCZ301jb4k51ZCo9bCEXdIo2SACqEe/GyLewAPt2
4U6QvAdYLQpQth/dRRzsf131XeQmr2RtU3KmUXYcn7YBAHls5tBxH3gNdcJTxfbm
/QNAkiYpQbeYLJZM7rEQNRO0BQ2ZDlzgo2xrTBWa5u3rFUgfZLgLyKN0HOmW2A7l
l4Ef021bW6L46+QnbK/Nj0k/9EQHIm5NQsC4RVZgOGUyI7xarxZ7lohx8sw/w8vX
Rb8tzbpFbYD0YpDsEgDDy+tqVdJ+Cihy2F1YFdUS0rLne/XF2JdEH0EQYLWpMrbt
Fc2Xkqpw/rFEL3z5l6pLjA0ApJP2NbR/WxN3OfEKImNQ+XAxSJnKmVY1Ilvz57EV
US0rNKoiW7DJ6z+69chIFvE+lJZ6f2JUkhe/rDDTRJq/Pc7TCyymvV6M2sBvbVvq
nhXCyUtbv0UTRdwXpMhJePiRPHyrReF73tFrXqwWTwI0k5JirQC+iDYlejgDkNgw
lEp+qNGGsjuu4CqDAVyqpHC/fukFjtoTU5AWxmsTwhwiA/uHDTQozQi6sZwp3Z8p
MRtaGlap0M/OAhNixDmhfTQhCV4PMsqkw6LnYxd/rRbUs4i2NsHnofq0wKJAVauL
b0MyQIN3iB+16nkvdm8CzmoHNUUS+eWfa+QST7hQ32sZwj4S3PNT1A5BP1+4EPmZ
c/x4Z4bIDWnCk5HoSiVlbQoiUQw5KV9FBi6TsCYosh/KbgXOVZHhUF5yMC8CvADk
lCgT/zoCvBA7Wndp8X1j5bP00PHjjs0NSVfyL2qr/u9ZfqR4f08bRiNjft8TJuI4
4GE3GvIjUh+jAtV9NMHzyMyUkM8a3D80j19chKiq9XJSG/ELtsD4FRBED9eYRMR/
98jaCQsFVoMNhFjrXDDok8SXft5wUBJeGwKfAyGk8hisezlnadlvjGJuU2RAfY+l
DtWLKn9Q7aNoewV6wX6ynUQ7ngI+6DM6AcAixSD7UqJHtD6cJmKOa6LKsMD45qFW
nFKtIIOhmUeDUvHJWczD0Qp5Ayb42IHruvQlavT1UK+foq080QPGky9FgZofR7V6
PDPHsLTN0I5L5tV+CH0kfwzuSyuqK+TeUm929h4d7ZJBYGFED589HRWBaCgaVagI
/fnUB8zoygjQG0FFS7e9aM6o/T3r6yFYvBPZTerQ3RjsxHVsXVBOgNQiAiuCbcKV
jRo3gTxyxW3v91615KJOf5tOBcsYbT5AjycP2qt1gjMJI9HPe9dnpKdmz4vyRBDy
xHmnpbhB29MZ8yVQuyl0SylaQqBv4RAg1/b6KlKg5ohZgPlTbq6cEiCYkFtkvYQz
WxkhmP44ofIxHWZ7r0EBBrmKsP/OQhE35NeiGkZPFe4261Na8EY1pQ9v52Wen/sG
YRrK+kpN08vQEUwtbGedzr7jXu4d9f39cHd2kGkbVAqz9McRp3xjrzlzAn/NNRNs
8LK/OkS3iwKxoWvfQIIeu4jUtw3KsJQqMEdbjMYy47OsYYTHVV3Ny0tOd581+SV/
7nzzcoQvyWdEkblBvZhDj9/jHzeoUQg9jxghkGxiUj4fdzX8y0pyxdn/WVdiENwn
2l7e65LU2jU9gRmHS/gx6XJjmM9ldPkkcKzcDKaH4xxo53AkOSQTBlBbKqIpI5qC
3Isx/jees7RUevfDlUvYVYOuuqwI8X78lGVr/wByiS4i3RPGugYMLIy6ksYiqjBF
lx234ZdDADIaCG08AbQCQKXN/hs793jtvhBmkHjtM862jF3DpHoQUv6R1/LIBt+H
JSRYgrR3SC/bTmm30OAfByiY4MgulGQf6T6arU6cvAGlpY1s0Ilgwi26fwIp/J3j
6x19F5MxsNz2jWYqbruz3ba6fn1rt3jG2iiU467LQQT1OFgpPrBR4tLZCUoLaHe7
c51aXtuuIRtyKrxI1ipCdhvPo9o2zcRzVt+BMGBABAHOPkYHSLHO6Q9Pzf2kkxCD
hEOFry5dSnsUvImMlF01ZkPa4ytjA2ft81ymWs/OmVEfDyPnCiYyUCUdZWiaLSvy
7wc0bkyw/aKsY00+0C70z/HpdEpo++S83DXYOoRKFan1Nlx6IKNN9R4N00SdM9fb
jhMc5HA1wuD9lG4XDCjpLoeTL/P1EDdbMWIj/6UH6JDmp9oOzizSLLyk9FyxWfsg
D2+9B+HYeYsimms5+0KByMS9MMG/REfeG/vdpbf64U52e4eahaFlOF7L5KX8YK1v
1nbzCXtkOGPGkur8zNB0MHp+JVAfj5byegqwX1OuLiZoX7wDCVMt22ryM7TMLjIP
KjxVgGyhmJXRVDnmsZjjerZHdinzyiqJjpNQPsYNs5LHc2/2ZF+NX7Zdjp4rJLuM
e69WJvG94XSTPNjIXig/QLcbmciHzTPlq13HnJyuAi7H/oKgx76ralApQCF3iBgX
ABaG8Kb7B9kljZeGLAB1tuiv/JVFmCy0EWDUywSkM4e5AkK7OkjCm2ZlFtkkQqxf
p1EnICZm9tbLwcRs0rHhRSOnB9gxPIaa41DeQGgUIZeptAxMmm5HjATUR3b1+m6z
kMW1ouwjImkLGvMx0VcbV9vAVJiUnrMdlQ07oKHueuOEAWUbMOLq2NxCkVqwf0Ys
1Srq6mSIyzpQTv4d0xgwhYQkbiS7/RB8KDVpOEVxkDXTxt/QwhqAZKHgExrHvxgm
JsMxRGaM5NrBV8p2ThiGn0WDOKMept//0yQSQXU5Sd5NCiOk9jKOjZRAG6jrGKxC
LRm2uiOpsmNgxt4AOeDDh7tOa+PEmHFwYVbpHnskJygew01UkrEaz8r47AToVZAs
mg/ZTiVJiTm00DqaMpYQezpD8gvhMhthojBr3i7c0vGmbLt3C47vp6pXzU2iiZci
Vc4qE64QVcmM8sDoahkuMJyv9F/e42/JCvQilayejVZ3kqUQHPp4SouAXxFd42rf
FdNnNzLVU4Djpm9AR5OPoorjpx6cCZSr+2DZa5yZBC01j3L4kOqZ9LD2jKdDXXpA
cg8lKBmUs8iLk1qM9VES3/Y/XTBxBEJ9lE9Nl5VLJLpPHVAja679KS3yj2vdD7Ap
OMN1moI1KoGMyRxpinvMlhQ5BmDWzS0KfAxeFSlH4vfAeDWdJ3DDCsZOMT8jEmym
/0ENpoyZ6qLH3+hYSK/bhCU4zkGVOgNwdl791HIYkgnvMjPa1csYg/BRzfmUhNoU
xP/xIsf43HMFZrdLI3Jl/RjtKWcJtcmgT0QrWHQN1+pII0+FKLLmoTBG+b9xKJcS
RekmNLxYBwEXjG/Af3rfxnLwuvJlS56veZRbKPuHWGR/7TEwRM7m73sWQi+Ia3Wg
XL5bjH6Ekh6Za36oA8TOFAJoywpoFvnQ6fSgGocggmWI2wC6I4z/Su3OBb7yuptE
hnLcaMh8vLocI3NIV7Rjjlqka5QbJCapr0N1uqqoM8ZdzPBbsFlh8dWsAVBfY7vb
DhVzud7VgJBWcNHFIfpKv5mJUg1AGzak7r4AZvwBh+LWFlsIPVQbgRWbMkVzm7Y8
XEygEQAjmgw+voybValR7G6g6nvfAxznj5UCM9t5WFY4w3BvxEHcAMjMNC2SUHxw
UtjEY36LFag524EdpCKbELtOEjoJfQ4JfYJZ3TNjWtY0//tjNgIE3KcINbDaI9dB
CJTjOtYKgQRz5RGChUITd93flontCEyeK7bOmxR6mGQrnuBE1BX6Av8AZLD2ZooM
75XfUBWfYEoF73aROgqk3FQ4hBdAlYXhrMi3qN+8UBXeGYEvyGFyR5/6sX1iH1a8
8F59mRGK9vMcoadqz20qGalPGwEpSwPP8l7q3aiCauoIQihR4K8CdOJNel7cgq5E
zvs6D1qQOJwMlog37w9oeu1x3wYMV19//O1VpDpqM1Al676y/SuZ+QUCvVB9eNWK
CTA39OP8QW79Qjqgw45btdVWlvNKsIAO8VwxLoAhwgLkecK5tvQFcGwYR83HdCBw
967G3m1jw0f0+TeXwdkC50lMpWNpF+8hNBzuVBqDIFpDSmfLF9cJku8KC9/OHuFo
Go4kcIAyKJbxgcvhL7/9Vk0znUeE/fEcKZtfbN0RBuyX3TGsRTUE+y8S0pBEF0J0
+u2g/+JzIsp4w4wLCyZcLXMRNF1qY8b8WPr7o7JglOVJPJC7mcNaotBrZHeZE/Aj
b6ogr+QQNaj6uYJI2D9vtPTiNE9ovWp7VUPxtY3HDV3ledwDj8w913jkRyid5/Zo
GN4DsRRLVPkFDuDMTaUd+8Z0pxonisvaAG3N6nwUibak4B9iqOmlPbCGGGvtGChu
RnC8FnSwiDmZycDYOJgZQ7LncWdW3ffK6KAijIem6zwI3k71uYiogqg6ozWR7TNi
2XKPUFmYKrRr50xQpq9MEpYDyJJqKzNsrQY7mbkt7AOMjUm2oeYJ4D57WbTwR3IP
/WQjpqelribwJA1T4evb7Mo5MYQo1TOTucgZRRVV6KMbyZ/QDLl5tXxkx1eFWTCH
N5WTbZGwQTbav93wQaJ4/GMjDz7g/MS4rrUyL3uPq4zrbSe+dsOgeHl7adyfuW5u
2MuH9RieGSK8W1kOyXqoUwE4aVB5KqzoY6sBY7pAQ1CE0m9UpMV5Xwus60g5wu5v
v7991P7paEUhTRkNEFDgaQWMBrPJAOFJpaWGbzz0Bl85YWHB+skWntd5vhfyCJH5
ZIQcl7bueSS2c3k6uKiLNmUzbDlsatIv7S6cyyR1xknqGzweLqbocVP3le40sz3N
5yv3d3o6QK4Fw7ugeG9k7iCTCQuPEwkY3cxfbvSvtZRkaFGW83TVFRCJyIemPfi0
Sg3Y89iMIbeYtVNWNQZCXsAHHwEJWTjmassqAK0PA+hBELwx9yUboitTIvAAlfRB
emXs0/BQ9/d6ufVKzOHaxwsELThyEXiZS4kJbEtk0K4oXrrVqa3fb+SROKSO4qwm
Jay9cE1yjvWy8oW0k6W1ZzePR9ct4XBzF6CXlRh/Unl+3/sLAI0FsKLDVt91YLKY
v7rhTa8Kv1v+HhkJAcTa8aMJHkWzMe6cPNYGUEV+uJPVNp0CkLlHHZ3dvAM9kKAf
Xxi8tlrhdLz2AfBVm47uO+LLtrxn2XuH33KD4iajV7rmZwnQodG+MkPOqmWMK/H1
Xo3CEvMC0sUi9gU9dqJU3+Yvy+Na0oWYQNpOrg0sgjxsf5vW7B5eDeTOr+TTu2IJ
GZSvBVtfYr3ostn9F2o10iFkdg75AgLnt1FOQ0wQH648rILBZK39gPTLYtNoAiz+
X8YncWe+9mKu6v8OYkXFafdLl2MFghqQ5Q/h1Cc8HritK0uwN1qeZLprXQs38Hmb
dYPEmtLQTvKtxJpt/hnZQtvJFcd8mYp4/lpf/5Grk8dzBgH69n1+yAB7ZKmFI4U+
9fhQMqdKyYzm370dcH3rU9sqwenEx+FH/v8bS4RU8iv9nxpcSxCkRq+P+ZSdWCZX
Zzte0wFcNojqlMaT2PAamOpWyiDWaJ+aba4OX7Cf/d3EECRyO/6TwPEls90BeXFL
ej8xwklr43S4ow40l+d6ystpyzq2WVmToEoeSbDlEMPP17LLmn7AF9YqDiVhoU8R
EsbRk/pDv/zuiHYR6GzS2ZyZySYKYO4V3p7EvsWh3sBrddeAyfOqWQtPhlCb2ETR
Q+OgWhftF6EX8AT/RjjBHCnfgPEesN0YoV9A5hyfcK2TN/40hAo22ZDQOZTNBZR/
6tt2clR5ekgHXiz2RMJgLkfbE+Vg5VVyP2o98EdH7Lxns7BLFTP9chGQ6jZPeKRu
vaKDWcZ1YBLP07RpIus9MDxBZksSjzhUSzPO40Mv7WeGBTnxDUMeZBQPEH6hXxGQ
6KIRsjYdxCUKS5Y/ZgCpblpPh0roEXsUUlFoNpNMoUsGmquRI9cZzlXZzAOY9pI4
dyj1N8vbXn8C9kbdfn0W7n2Mn6ApezUW6bxlwwAx2MuqiLJXuz5WKWnmDa4DGnL0
ybuK2EJL0h9VAhiVBs08HpprMisgWPc4xPpV5ZbaaHbXpmocrS3JBs9ZzZoaMECw
JkMISMaY+QnoIwgtsuKeGQF+X9DK+PDt4/OM2ryMs/Lj1wYrCXZHGT5i0Pw2nUCb
xHZT3Ie3+y69cnxq5xR6FXDGcWdGUaMlegiFrjh9y3aV8H01Q2IZcmsicvOZ9BcF
SQFDQRIvZ3WOkB5+4dsYdTQSdrqLYc5rzrGLDDc72hSNqGIZmUi57E2BnfxkmlTD
AJZWUspWkqQ/xnUH7ISY0hBwiunt9Aei4CeCWICufBtOe6DlINaIs9vxTI48Pw5Y
UaaeACVMX97cumpMtoyk2725tcCOoo35LRw2eDR5y8luDbqEyVzw5TniuqzHedf5
Pa0HAilOlJ7uDPTw05Oa0iuZJ75GT+9nmr4zH/nBRQAxpazgUwm56Mjc5hgvioc2
B2db4+2jWZCWlAWRIZXIYrl+QKAwL3fVeElwAYMeHO8A/ST8L4dtOde1cHHP+mlp
b9yqbgtNgbjwzYqWKFtSknr/ocvVNZuLY0WsWQG/8u4n+iOHWrUeUVHv2A7HVTsg
Z0w1wD63tfLFjFdz1GB4UqYTOwAc9nUhiiso47gHhk1Z6GM70rG+COgjqNeIuaw0
EYxPkqn4QVmIBu+FmMP5wjgL8UtxNpkUyQQdlBiD548hztlw2sOH5C5SrBhM7Csl
e42jRXzI94LqsahIQQIBizAN0dSaqPUPuJoYlqIRbH3e1JywkY4iIy/7Sm/nmAoW
+/GNUERH2HAFMgggKN/AZOHrZCA5jT+1nOXcwU0KSlZtzWwCwNmLwQgslQneb7BX
g7cE9QKKjueB+62eqeeAxb4DFVNflRwPMSOi0B9zVgoD8OFB+qlb+FN+fkXrTYad
Dgf4Zk3ZS/qH40Y6UF5sKCIAuJSCNiUnVp2n2s9T+9Yxs6WUriv8jG0DE8aoXX1w
qb1236jJXw3WOZEbgHGuZsBmwvVRV5+FJpcs1xkdFnTz1Yc5KriHDjgZONRXnY7k
F1BbeF2LSn5NHfc5sPukwlcUSFG/0VJTImy62mAOP7TgH9Sa0Sj2L2Gg6ghqgbo8
G9WKkD0oTTgZzClZ4rRse95wej3dabUtvZ4CQMjBdHwKM2eK4NT9i0JveeFS3rBY
a5dpMdhJC3RPr6H9FimZMDgEwP2UlUOWA1sT8YYe1DNqUmqOqW4n2mKLw5jzpgUI
mz4J7DCRiYTL5H4sQ2Gx8nJ4wXIWvO0Kkx/6azqZoRDdPB+sa0YVVNusfzRi3QFc
0o3Ta7HkESjhX4Yc4yIlv9ZrGhLNJ/ju1KphdZbekn/f3Ei2+GUvnt2IqGjj/SGC
YjuIKAjulDs5Q4ygfgvrcu97egt1MKBw/7mz/Nd3yVEoX/YnsFSnExYUWaGLkEgA
02tVh7XGmao4K8SSdKQ/v6aGj/+uDXfnSlRqoEqGSk9twnIuSMWQpe9QNnGBxrWL
Mz2LLSEx8xi6vic5K9tXry/Y6vpmNf+irRy+XmA0MlL8k+5Lb4qg9Co5j5rydlPT
70nmEYlcfRYrDE5Y5sBLnmMPNn+8a+MxkRuUv0P8A5dOmD2jboVo6XWHuMejLua5
Q+xi/Y4DHP71r0h9i27P9PCjFar0nAUjx36h7YnLpcx8v8jLnBv2A/NBoXKM37UG
Ta0rk8/mKyryaWRTvruPdh9u4FL19A+/tNjdGzOIoxz3e4zDHyZW2t66HOXIa8GW
5qgoh7DDGyxHIvb/M3k0NK1kEtj9IX9Ig3Trto9egkuAyHurKd4Qjk38DIuhTkVp
KvnWhbbPLzAQpmhGOpoZJ/tz01qmS5rpYIpXcFHWrNu3rS7GoD0XM3LMsHeutxrl
QHwQI4hgx79ckwIQwOd5ESr63nNn/iePmMk2L+4jXB5P6yhak4Ia925FwhojV/3j
AN838XhGHUr3Bt1LvrYNTHyKHIVTwLRciWLSMkejjo9kPLcllOewOP34R6uJceUC
ko13x1Ca4+3LfGxHYZiNfZawoo+uYd4UC5ZaezJeSoyOYiwVCb8pJzny5TzsYgrG
c5cdxvjOdfsIuN9sd4XrtqpisyaISCfFeOtZiGB27yOZhxC5HAltrZfeswXIBiO8
sXhmbRdeo/V5fw4emAOxe2MSV7YZ3y/RomBx2obXDhgHTYUDE7Z1OEMXlu4kR7ut
OglgXOZ+6ZJHJyxPn3J8PyY/l9N5fJWtWixLDEfScuO1rexUZvtJeReUMKZuITE7
zDCjj4CuiBFV2khw0n8DNXr8iuvgUhw7VZSxT+ookJ9gAJ2HP1M2P4mEfWUZJX1V
ytfVJMBIGSfFUG3UTxLzqPylJ2epaAnRadvuoCYhQVdDER7ThbXLzK4zoESbVeG+
/746GqywwZsO4i4OIqN5qtbAvtbG2WfYxb0/9YCH7B48/o+fTRxP1dlgOGyjNFYe
NHKaS18gEXA2Z6DB1025RPgvPjX1m7bHO9NkZsiMpR2dFEsmNcBW/Q+E2JH9y59V
474Ft69s1myf1KOzOyIvpf4QSNfZeashFP98xb98+yYgAcHv3wNEaq6Rw5KHjvoI
hA9XB7jvEzltxtF+Ck8U1K9CvN1ObjYQawM2qazfWehtQJlzAOMo0eMbPUoHiCGd
c4BK22L1oRQPEBJVk8o2e99nuSl/EPx13HSLYCq7r6cmMN1IaBUmsSlvVtZvbnl7
DImOyZYpoJ/UXPJvlx1Rz6QIyY2DpuPTvZX1f2f0I7wwayMAIPNhtOKE76+LV5PF
TLApTRhtvg8fNM0V/xgsGQYNvknNP6HyPYdiVRSLiPQ035i8LvNugb5vqB9AKEXk
c4zBYdkwTJvr2vqTEAc1gJa0nJaj4dHpkfrOmJoUNyil4y9w0uHsB3M80W+P5TqV
mh+wqsmPM9AiDCWg/7r+EDrBOSXyVz7CLeSSuFITl1fpl0okJz0O6wNo6chu89Ce
6j/VPT+Fqk4KcfNOsDHA91FJ7OlRnGuWTiZmhdV8D6+qR/mZlSyKJDXyrfFN3fcL
A2Xyf3gcOMAqJs3Gig0iyU4OtLWdSizvpIhyrKDsnzVrdOIZuXRccC5FGvaiPRwc
iag1Bg95irLjpEzA1ArFdoW+6lpEvDoC4A4tEy5qRKBWJaI+aDG/64w0G8Lxq4Tb
YGuL3FhqjqbsrUaHwQ7HFzjxOj6PTOuvWT3Mu2nohcWiusRqshbv/GeNPfQ4r4A/
sUBfT+0JtnO5QZ8MwxdyCnGDGosS7zdSyv6FQhYyVF62zy9737uv/6wECmgxgYJg
FI9VVqYSWiRqtbd4jWOcn/9/G3LJBXu5ZoFCuQUudaqYnFQUuHKl+HwHRl0qCDWd
taJVlKC0o3c60rumv9D67BQVqP8JMrmaBVK2G+Wnv7NO+8GctlFu/yVFeAGqnTqZ
mva+AjEbmtLWCOpyKk3Z5DLUKSfbwh9rF8YpO4UT6KaCT+Wsx6swV4UL8M24iH5m
RwJnBbWELlxS0ReemwL/cAsrds3LnKuB6mPjrhk5NdLz8RmMYwLJ1hbGbMUXaejw
QEJ0poTKZwB39LEqWI67zbQ0RE00ooPGJjSBRiVFn8xfaxnkMei8a6it9+8Exrbd
jEmKbP5ACcIWljnwwJ6zu1UlajIX88cwWgm46tVA8JmhDlL+EBbF+c/hzQyRIzqe
gBrcntPoTS/KJssc1zYOUqzBVE3wSmkvS/LsZ5yJnKUGaExahU0K654h7n9XkF5m
EWW/XiaMcghbHl2bfNyp3bt2lwiTnB8qF8NScVGym+1DiBdgwtIb4ntWvVbmJROC
VQyehdwFGrOJqOkohOQGNaET4wLKZyvXdPuShfzdnVsMaX/ZurDrMvk8Bu55Oyfp
PZOg+TtQi6ZL3l7MJq/xNH6YvP3cVLX2vFC3zcm6HflZmoHPaSosjJ2NeI26tWV6
7rwK3f2tWtFxoT7URuKJuU5Sk6+bng+bjGa/rPMcVIMGdQuQTAMd9ItjUqC/5nEl
sDaaZcZCeLWEGcXvQKj+tadi1g+PZNGhUDdMVkvFu41CsHQRAW+EMUJh+c6G77pL
JciHOHiGg2ZRz10m69nZ+w31bhPkRGUxbYXeJ5J924jIjU2wZ50c77smTWSluLOt
/Zasgfh1u74bLiOSdP5mSjnkPyA8pyH++KojkeGyaFY95ZzcrYR/OpxeuzIoisiT
ysdYtXKEd0jt7Hw4GRSPtTnrKTqNPNaMAk7bSwJXSNOpqKlJORMx9JusN8POTQxx
reMRt9lJJGlmEwDZ+SF4QGh4GwGBQVvRTgY+tm1LFLW5Sgm33HrKslXO71hErCG8
8iyfNAjBYp04kiM+XNimuuIhrMU0PPymx28GsXVoclqYyoFju0SftLRkrrxh4NI9
wCN3wpG7x2dmMFr1Il+u6LKHf8yiWYCgghi0kCvM4xtHLlIOX4rkxMdJ6vafqhcz
vcfoV4CK2oBUGZQSjEL0+YxmGTquS3WbFg+l9xGpazwI5Q/0A7txasf4I8hEGe0H
ecRA4q63DYfOSGOPaTzfW/h+8aQhWlIIMnyNDUVCImIsLT9a6ZcWRpxykWNGQL8o
ps9zhZNMKuqLgmnC+pZHAmCzIzcNS8xtLgrVYopnSKSHqKMeJuhLrRhoweDhzIp9
z9YwIzGe4T9/vOX0MqbtK4yyVtP+jah6+vhBLgwUWmo1gGW7nD6u3XjEt5ZoznCu
eEK0f5rZv+rxNUsdi5Gad1qAOLUxi4VbefZRDCJA8Jk7XDXyeT6PDsxsfh4yYL51
chCQIq1vTTjMvUnI8C2rskVh0ly5O3IbMBWSfQbYqqzde6u9QabyuW/crf2eA1Cd
djDxnIDRa1z120EuTK0sdjeer1VL/+h2X8nMlLHL9D6E/+JTYAnWe8zqUhSDOA9N
rAYwAW2t57xybJsc27190LfqUVpfgXfnRpCJYJAnLwNuEqad6bWim9kG3Fsw7IoO
P0r1enDlr9CyX6+E5zMHIPp1BB7oipNsBAm6rkNj2rfwWbnoAbJujOeaZxEZhub5
Ktcs2qBUj4CZNMpk/iwufEmUfXr1zQA+lTLcxKABqLnS+Z7RmOhXZwrcby3GOGae
We6ZhdaJsvpcAHQU6rHCnFi/+fhYyYcD5rpkq8KP0llZzbyDPLa2lnLpOyyQaNHG
oS28VyjzoAPlwJFF4j6ujSN6FpMC3q8FZKC4YrVNTcY//uHVSEGTBzVxs/dGF181
YsMz3PrzBbVHJGKR93rs7t1Fqp//FUtP5TooQhsZ7HEeQDCnyVFStQ7gBjtDPhU0
0pqsraua9h3gOc1joVcZYfzAcSmGA2Y0Sw7MYooaTd2tmEQ7PophpPYFPCcwR+C1
x4A2/2/6YAe2YjOGqjzKNNrcsd45zqmfY6siWB/LwWKYdiCOgc6nUTMMkeMChqbx
mID1VSt3l4HYK/LRVwvntIXo7ipYWkScYnziPVC7FnwnKDIjm8gqxkPFQvswbUOy
9Duzp0TG2GFXt1Ic27HeqFvuGp1xk9xP5NpSyXTPLYlBa/cYgvmOa+pE3vrff9UB
gx1WNoDxI1fvPNlZubuveEUfbTI3zzbddF3zW5QZq5YXC6nB+/UsGlXzdd4dgmn8
E+ReNDI6EzJF/bH1PHZpg57HaXQQHWuxIl+2SHPERtINlSsbOYDBCQthLz4E86GM
FCv3TLu0WwuM0HMv/NNdmSkPfMcLn3LjW+fwe2sT9OVvab6BQfe5xgpzSsucdLXV
2jq7zcKqeAdErdbWH8gx4QV7LbAZLDF7nt8wXuB5mOW0BHXlwHscHatQux2waxTg
WyMtr01PL/5nkIsJBIRUDA5RKVTmPI2Q0GWr6yjbDF2Kv5VR9Tpc3jwBjj6ft2g5
0c6YpeDCmZrwKNw+XIG7KCAnwoffSIoHav3uQ8w7thFetj/oLxhwQVsapQGRryHr
pFC5RTiCrohva7lrAU0+ndArzuaxfw+ASJAMs00A7MVJ8KwuVJV0ycXc7FViD/xj
2rn/ZtcaTk65api1PNQOWUO2aVmiMWt2IQQPmGsmtI0d36SbKE/OGYw0JaC1FmLT
96TDHnNQDzn2W40+h7xsJa4uaQUm4tznMz1SatLBOmNO/s3zA6tk3/MJnUvu1ONv
kS4qnBd/mPa24IssfihnEbbfyaKwwhgliTDVGooB3y38wfuITioPb9c9oSiIPlPg
fWpA+0W5WvXM03UAAiSl0BRelGoBoijbR0bYkK2s7Zp/AQ5jy+C4PNAWJSdMAyBQ
tQhkl+gVBGZyLm4CeEVgY/I8Z8rF9a9zOS1ZCzpvPMdYNGQLc25lgCubAPyka1aa
gpp2qwfWwfVyXtjGgeuxcVyidQ6Q+MQEfhzdWFITrJl40gUYbYf3HpV9SloAPUdV
u7CeabI5t5GCMmcF+mOPcNdFkRQ/qjkVPFUMelAs1fGJoRTR8yaudIAr+xNZXEfy
tdoWMuIZ72FOoPWWKTHqDM5TzU0OzQaz+0TvqJ5+Z5amdDQgxCsbKXzN2x24DAd+
cNw1E8xLsE3dOrwJ/4/lC5z+kmzyI0IWGAzaw4yg9XJbQkzzBbnu6M1W6MeydxdI
x/McS1+stNSkuTujSQ9O+1XxPy4yGUgrkUmGgOJNXFHzybM/UUgGjLeE2MGTpBrZ
tOTbx5hM31LvLEyIumwR+2nfVTZodhMWgNStcoMIacxWiKp/m0+zYKu0xvdu9Tda
n0BFSffTANSWr3STzbkLGWnaFPznVOc96+tDcTnjrKWsZHreXupMx3HVTXJcjBoG
3St2egZHMRYE58+KpUAgEbdvIaUavPabZjDKGooRN8JHZKLZ2HCJ5CM4rs1ZpBEK
18QMXopESiWAlqVPI5Ia/PBW3qHnNSrlqXecQG+TpRcLzWdy1HK+cnSDdjTQ1wDL
00KyYSF60nKpvtfBsxTWm48Vy9241Pi8crNp8+fwN70b334nCML6LN2ANlR8z1vK
O5v9DFCqO5FqcTK1UVGxZoH5EOiLfu0eU0MtQtFHwEitFANpO+f+V+orzNROWyK8
GhsgwTo6R3A8R+FsCYh2epf1UayIyFx8g400BFlIAKDBjk6RykMvNREP0m8uwsPK
idPdAvZkdkjzk2eY1OOnAcEqRupe70RJDFQPrpu1nWgyRjc66TSyfJ5jbA9PpZv5
23ye28cIMl2TncbH+2qrOr8oKjXn1iEJO44rWUWTADR0yxsIPbnvidhdQ8VwoWEw
CGJrr+Bg2R1aUF62n+9GQjH1g81yvY6HmpXENFq2VtoUtYsVWpFJ5Y1JtmUsmWJn
6vbCS+9fJRXpdWn5Wx7pU4Q+3FwrmZJg6fUQ5lK/Knhwwe/TthtgqGFs3SJHPlYt
zU26IpxLYAclznpKQV86hhDoaWqTucWpf6WgSb6tHUCOGLiy2xIMJVF80XitnUuB
SGe5JigfYfjm+JiB5k6uhaS0k7rUFIPWYeK97GHle/zmsrCJGte7auJmu8iJIwxo
nYzjPNNLf05iecmQtm2jPSq/j6nymmZKq6YaIC+rwaJOR6Tfu/fwe6ZOfrGBvAaf
Xad0Rnj69VjBwbbn/1SsXED9qmLHojzI/giqgKcr18sWuFYEI5XmAuWTX30YzE0q
fz0mvBn3F+zPSNHaNncgcxDvR64vZqeutoP9puZNOlZbCP0n+g7PU9wCAZXKj0Bj
sx5s9G7bTix9dQ1X54yGrwmD+7mITTjQJ/Nyl0WvNWZgjv2xn5zWS3wZGBSoV/w1
QkaqIYgkidULT7xsQY4QVdfO08rromGTRdDv6pBlZTlTRk0yUmhXZPFAphemX5z3
UDo1unj4GRIodp7f3XIsBfVVVrLe0pPv4wF52OhQkWivtaYAUQVjZS4tu6AU0zLd
RHJXxf0/s4CZLsL6XZ55gRohuHiv8NhciO+1Fb3WD7Begt/sD/1d5XwsobJFmuw5
OAN1/+q/q7EJ1X8C7tcklQepgITYYRhO6wtGt+4ox8tHPh/70z0iRwiGyGdXL1+2
LVwixK51/Mtxgi/eOMucwZ+5keTv52s8qWhC27gsRpoNcuUOuSxYfS9Kfphddt11
Yvl5c50pO8Y6t25IsC0B0Sf+PUw9Vdpcv3tDhSA1qPd3iLFJSTzDurUlU1DDZPn7
zLz307SirSa8Ybj5VcLnyiBm2Ezs3V+Ie55g+wqv4L5vSSOZYhqP83x7I46Hz1lt
ttbr2vKGCFlxBZexnqT44w4VWPERKT7V8HcGhT0PQpe25rQeMIdYq0og6jFrKHPY
+21irZjhpHfMb0UUD5Bf9c0W878w7ZOTVyT7XvQkUkFH0xxLs3zeVNdwB141IG5K
FdQnGJt26NiM8Zm681q2dB39VI/HQfz6CyslqHltaYOzjPOZ1bybHT6XLtzL7gfk
JHhh0F2HafG/Ye9iJXHKBfKmKAxTaWHY2pEWf5MWoTg9vZvFHeAbbUebwrZkh6cN
HEPM7OkGT56+Xwqj8AZnl8KxnZ6GgVkKy+QcEno/sBx1aQYrC9vxiIV5Qc12+O7r
jO1437ZGYjfB6xGqiE3M3iILiHfPBRAk5HC9qGLCSf27/+VS2/SQp6qN+KkTcRWB
CRTTVgtVfWV2/vI1TzrKNDLhbK6K3UuEM1iX4O6CWi0TNdZ2RhWycIqbCGDwmhkR
9Ch2Xx0g8WdkNQJHj8yvQKXWVM3XTuuaD94Id6DvbftIKEW0h+hn253Cx5eoNUWT
rDxKgBjz5vWfDOGCSmj2K9+hoVnypzKv0Ngqw1kuEiOyPe6OtZEf92e38PEfUcXO
3Im2aLjv/EyWgwfliPX1XwMDOJyvbiAVC2RISOs09rBvInFx+QDy+tKUmGgt9fYv
7LJu7YQZ6UltWcvReo6S3aZUn5OFMcD6A3B5BK3lJQsVbn1UfuvwGkAZ3BCXw5PG
dmy2A1I8RYbnK6eFYW50EMvRUt09eWyaiGg4G5uNqpLHE601NU3Si+8a3qrUbNYx
dN7gm09X4HOywihGz7Vu9xpgHzJh7VkAs0pjQURuoXgBM5ASMKJ9ZNKItaEy90AC
3rgX6dnoPtqB6MebJnsp71JraB+/sb3RI/org9IIHFsfIyFA2l5vREnY/kD5ZmkR
mB/fLVUzwpTX4qUNGMGCNTsV66/0/Lo8pfZuUkca/WFn/d/0PZDBgajXgMTLccUU
odDRLJm827bfspk6uaKpyPJd/X2erPYNT4PqwQPdbz8ShO2Xf6L/73X037RIo9u+
n559sTG30TjVwHjPX89liiR226mkJhOEskdZulXBxZ6XHH9OdwK1BowQW0ef/154
YMIhgtoTkEp/neKEyZDc6CgZorJ4O3K3DfAlkBTgo4psy+sQnozLp2ZBHP8TflLv
CvHhFkAu0fbh0oV1We+jhvrylpIssW5o78GpjOwWQN98rF8nEjWr5zyYTP6etDxZ
/M6EJYGI/grj1/CmlA/q76iNJxfdoJd6Lulys2zYzcQXPm1GWjLMUnxdEvhFClyr
cAobT4VuBJUooxUZu+D8DDvg2z8CFmlULhB8lF06WKjp82Wo3j5M8srM2XFvCgUT
EVETv2K8aA2rKECMO59LDC746H69VP5H2yqvF4FiPyIHjgt0BbEpK81FT+IdZVMB
sFK4zxsz9z/WVW9xZZF5UKyQcumtsJVE8WfGyluRMhsiMEFCdNbNFJoJbcol4M6y
7CT+eiwMoo23uakOEEO4stbp7oRWGbW7Q6Xf9iTHza54jVan0ip5qEa+ez5vsm/P
DORYiKoD53K1AjwttPu2cCNI76dF+4/v8RM9Sztz5hQAYGGAg6WtBnpBEq6NLQGs
14EY1w+9IOODyHxzthAwFIisAeX0hPiDq6H5xEFu8GNezgzM9ehfCyddq5qwUq2C
X3uVUcV6Ptfo3yubed0RQO/IVuf29PEr+6zdDSvabLa60JaICzx2GnZYR7Nqj1++
cRdxEn3/uidK3NS8BkEKijhshlK5tUoSdyvLi6Ydy4a/8vsUiiFRlC930n+2IVPy
NdRgUwMWvJ1yzkK/pHHrsboDPlubNI37mh8sPuXkxUWfNXXXK8+vUxcow5b78WgR
p08zO7fkiqoDlgkxtCBenkPnY0RcATr352Jc7QRdoh/MuKQo+4QGzLOguSGEPSAh
IbQmveoVxW+0cwS/ITCd8YZaWFesXHi7brGdeMwonEtkHU+Xeecwvv3NU4bQFqyB
05xvdTlmWPW42P+2wj2H9VpglIQ1l6fOtb5rVP0cpx70IpO/s0Immb/dlvmCddgT
iF61L7XPLqgmmX+3hcpG5n7GWyMRYMdqo6tJOYeLloahqPWgP3X9MVELoR+DcN+R
R/w5XDQm++ul6HqBv1gJ6vNMFpyPqZk2of2E85zw5fzXqGbuwIPd9pFkt+MijCVW
fdwGjsVDyTd3dC5U+X9arVNhaBtrnOL0GvhN4ztBKNROJXq1WF3aU7klR9iKaLMx
jTokpvuvySd+Cfs0IrUCyrswv6pr0BVE9cPZqsQ0Pbz/UIn65rmmr9Y3MZk6prGv
P3NjvZDESTduL1bh6ENSp5QW8PZKhPwh89rwnbN0UjNez0si50F4Pjul9E/1m4Ct
CkIYaZg1BjhFhcP5VP88t4CFatBqspdzcyjP7venxQCoVCtEbgXuJDV/RkpJwxLs
TJNFb8OkIvuDR06WZNip78nRZ61Ryg7AU1VGMe74g3JamotlVEJ+U2jIvBJMjpWe
7X0kTgWI0YoGYYXJ9TuLC4+6nH9WdKSxtthpOAADr0JboUx6QWlLOTKrPFhcX+pS
tg8wF4fAzxLmhmv7smFpCEGZZxZqu0Y/jeXYaheRDKrQ4IecBZnTjJU0+NzUNLLk
+QdJ7rhIEsfK3wTPvN67NXQf1h1ZNEc4ChzczxfwHv5/24aYDw5Fz/BJtVdSf6pV
mwY1MlYuMFbyr/UDXOMKtLYa5TLN7GUUYkmbY3sE1adci5aY2JLa9gUhTlFDHUkL
/JemzKAxhqrOXxgSNDiYMqx71WqvUlnRozdW1/EwI8Ltayr/5S/SyYjwH8L/jGBg
mFyiSFqtlnuDKwjSCpEw2H0fRY+8ZcLkgphJPyx+TSCUbhdHGmFnyH18MLtcGeLf
xF96RBNiTIkPxWbvP/0BmkhdlkK4c4LKTKoRl0YzM7I0al6g6N7ZLiQXZINtV4zq
D4pEcBp7NDFlWAqtazHvj+abMimBx/7TNZiOLTLsOZLURim2N8RPCGmFCiJEl7Lh
InreCbBD9F9vL27aZWCZzDJbGtwauTi8z8tAQKg1YNkhLZjt0RjhIH7gnJnQIEHK
LK158ASg85jRQdqG6fyobI++jfFUlkpUx+qgjxi0yTGbxGKvO1C58XLSKqK4knUP
plbI+TGG7GgBA6D5ot/lKiZLGsT+LeJoHWncNd+uOtJXCkh0OefciyBf1qSamzYe
3cqQmu8qLoMzOAxwVWzssnUXXIGGIoVc0+ccP4HeorEAQhWvtvnFoX+fTIOue2Mz
nOpXrNczPh91FozBH48l7Efo8b6XCcqWRmsRnztRs+dOh21CYYijmU0ILZzTjawO
h89rUZv0BGmw3irSt8KaGgq8jLDKlP4eHpL3OmEDqPYDhivYk0x0Bt6MF8eZWukU
GGXRcdqxjgm0QcQn53j6Fadsc77eHGa0hpqBSic5VK3YOLcV0Hc8wSEhTJFbQNYV
QChfTZFSpGKKmX4Dn7qgcP+RQLSr7NApGAuoUyW3WRKk+pWbhy/Nsy8PRyNmttRw
dFx0jwnD2Fi9UPcYMJfDyYy0/wxkwVvHg6vZ/klQ32f8juyriiwVmEeDy0X7rs0b
QpNF3AZL6noWSHy0WuC8T8qjymQjokS7Sm0cxcxC+rzFLb+ws3K9aaz48bu7jOv2
UyIAgAON1hw8XKIsuEihqBYVeEJZj4xD9j+AzSI75PBvSJyflT/VAh8g88RyRAFa
bkhIdA/hR/4Samz7oiM58T+Hi7Armwup779gic7A7RsUL/e0C+Ig1OGOBDjSCZkO
Czrcrc/Dv7FhlD0sYF17hzUWcLDKxYebNOpnoRaImWIAtnb2ZGyJV7k5l9LZtMdo
jvCN8ON4EmZfZUZIlTSIxHGhPwx4s6zJJ/ZAx513QO/0fusKC25q4NB7/ZFzKMie
yV03qGvNYuiHFolPukddUV7Opx4dkDU4uNZRou9qRgYFVvpD0451lmGKUJvRbSgu
Cyq01Ie1c1DCYX3YIuR37bJgJq8D+n4vj03Ky441MzXKu5d6Bfnk4ygTMN8KSX37
lRDUTfR/KKHAszxeH3bL9y+wM4E+q4Ma7KoKVPyyY7gTXhB5TE2mCGPfOXJI0IAU
ejX+veipYZEr621orAwOwcfLx6T7IPmmtLsDUT30K3WfHIL9x3eGf3RQ73+gT+Q8
5D5iyY0HI5Y1Yg/eWXQHqja0xyNe42i3yvsik/Uj9BTpw4GrSbqM5mOZTFny06Sh
IEZgoz9bsSohG15MyifLCW5oLnnoH7tNC8XZli4n1vOSStKCPR10RBAm9I23MQtD
o/fccYEPDQjpsF+jIwPhJKGHcUOuzYNSXeGCjPVl26I37nv/4zscwZbxcBWLnPlX
haQ0zjZsPqkwTZ9qCJyGV40wJTBWqPxqwIP8QQ9hUlvZznDto0LjxGxblEuDdt8n
QFJgQt59wXSgv+CW9rx0BeAQtiovd92jXvROfFDYhHdUmCLm1ywV4ZFwHSzuySq0
ZqXCBYew3y63CbNgSH6epDwHF6loJVn79tHByu4U6/6Qrpj1DTrGgwucuERj2KXh
aSnetTifJ3ICphEnb/6pruGPyS/3DqSX7HoYN0fxrqzrDiLuk70q9uVa5s5zH3l4
DyTR0pw/IOQqAeZjj/mv8uWGOrkBH1Q87Yk5q9uWlS45t9L3/pTtuHN1d92GbaNv
82MpE2WUwSDk+kp+fsKtHce86m3Oky3gCJIuwksqvKvDLe92qPholGTrcs4TIlzs
/TlViiAkydFli+1/KAgfugUPBywtX6YnUqG8wOgD2hshFhftHn8nT5LruZNpiKcQ
5H4yVNqexwlryEXNqxzYET+Dw3fJu1fBrxZYQ+zx37q5b2oVQGspVRpbmHPuq2f8
WRAfvS0PQpi7sahQhi6V67wGoBQnf5rwbgTc/MRv+U1xxWVqesfc32WnLyLAtmet
xjAP4wBKG1+F3AjZEzypIPj5PXZR8scgc4e6BYYb6R632XQ7ClRUN8nWmCANZ6ss
KkSTN3dwWBa7cQ3S8RGllUO3WPTtRDiR0bOE2dWkkKHg3TIPSvnC1NjTkyoKIh3q
nOn5wtdsiOx53G6IgzFcZbyODZuVATL0qVgBZbkAc2l/JYDhPQ4LYcoHcJ74fbRI
NQ99S6WeTWthAs260Q7ZC0hTC7C1uYSQ0NlXcAdKbjriWvLmddhtwpNlS+O00ae/
DKhWcByYJ4L4hqAW/OS5NzzMsWc8xVfr7gpDInIJs9PQuRj1UNCgP/yLoCl6sL5S
uTnDB9XvxG9VXlJ0/7pO3EEWjIwswqmRDCY9UJjYP8m2em5fJFh+gU55P2y1t/E1
q9NKw06/r8fQ7fo1cHfIQPDsEEgaTYWp3p9lf+IY/Ei3eZLCHWUY1wqp+S1PNyB9
RvalQ/X93vORr/+G4uDfnD9ZVqsWWWoLqELrinS+c6esZ1OuZ+DOg2SAElH1zkD6
T2LXEsH20USpkwoWeCmoBMTF4XzXX7jsUkTvKCFO4G9WTD0dqqLrgwvxL7m6G8iS
r7VQ2SVSoicg6Kgjr99pyBVM5HIANHPfJXmhRNg4Bp7XhQfiL7TIYoIpQBCRCYRn
u8NMEupcLBc7Mn3jSqn4TX8cOewh1VwO0JtbWdr3KxUTHmH7kkN5TBLamSaE5J9r
LmGxuPk71bnuPtzhVmQlP/k6jzhTsYgcJkBIcYycm53K3zkIA6qa4jhigLv3kS1R
EYJhFfG7uxeFaoWMxJLjOnYvCgyevcwdzVixFSXJVmevhqwLgCAhosHIIxS6dWTU
DIbtXnHtPXYoT0h17J1yxG+rBKVuKH786Dym3lTchzivSbn+FfflPkLQrp+dhju+
7/dR3BrHr1n7ee03N1q6d2t809Hs2iICXxaTs8VvrUAOuLAnbVBf93IyssytZY2W
SG0DwSrx6WCfhPlLMfoWfb8WMyeFsELxMysTwI7KI1mqh5zMqNm7KTiaxhAywurS
ufbE4hilq9XnmYjA2K3cgzEtKrb0wZMYeSPILcwdj8puaoVVqrS6vJXg5L8d2dTD
QhkQ01BVgOVQVDM5wSGskfymha+n3w0p0EU6yBMP3R0/Y+Uj9gTccc8sXAAer51A
lJ9/H3fP/0ij+i9ShHPmFLBl1GJe7TuSnYRgu/G9nfuuSvvVbZSfO1OnH0RKktCU
//SFhACEB0w644she/fUAplPeGaIpWbV6oo6siRpY0L0lWHmxe16exYdLhzQWCDW
OHm7JX3MLggs5GRoTFnJmbDgjy0yKR/BhbC5cmYHVJHxrPy0L1xCNOns9xmhW3jj
EHOsEu9zj/g+YLlEY18ueiMugER4YzaVRA/9triBzu6/t1rTNhRP8sWXPUAf/gjc
rMPtbpU7GTBfHljs6pDYBVC5AuUtsFAy4nrWVLxzxgMmNuA3Cec7YcQwIRhWEnFG
K7W5ZErKiQ0cTcCXgaXD3BZ0+CVToFRTUrEpBRioNrAHJlVXEA7s5spqsKHlx8mU
9eT78s9y2WHRRFqp23NOcgiYLsh8RdNywmyjEqrrihxCh690SViR1yw8cjM7+LKN
R1fwZHfwlhMS8cvE/oGSCcLlPmw20JjACbRikIav77JtbtFg3QOFr8KQdBlVCGpa
8WY6XucBhSZjdcYZJsuoY5NM5xbPU0mutoMtGf8piqrjvfLEV+3d9XeOFwTB82oa
YSgPqEYD3M/1t11tELNFhYaD8xC7FJJE5UDrZOazxczE/OZ5hkRIdRFVZGCvYyjq
g/Z3MX11qxdVT5oupm6FkUfqK8tZ9GXRofADtaUqDjo5f2Per/SCJe54rhC8pU3z
4VCGW7N6Vs/5SbkseBavL5xc+EW8kaIDKhZvc3Zz/V5YO1aloC2JCJuN5x3AD2Pp
Ts8XRNpDj3H/mPJf0IbIMPDUlcsM5mUnnMp/cK29VMEsi7kr9uWB55N9H2V0w3Tl
9+TqFkLE1hmkwcF+viQYgDnzzynB7M2A4cwlbNOYLWfx3wZiNCffvGlfxPEQw8Sy
Vy/mmkre+5sDRGIzE4f54EN2RpdTwZW3VsezRIvQPN9rsOmRhVWDF0jDFm+Ifdnc
NhalepRm6y/MTj/wy1tt6rrEUC4gYyl629m4cz2Kwf6jSWjTEUxCedOXKOK4JOxp
mAzmcTxjz5vEyTh9kPJHsFQazuSFmPmjBNHOvFm5Knd04UlhPBHOxEZI36NAKaiA
dUbIPBZ8+7IXFSN5FBz8W2FBkYy2QDcJlaVQrroVBILsDIoQWu7m5G0ay//6LLmY
nEL33LKlnNfk+32/MtjL20GQ3ZgbR0M1H3aiSnors36pCIMSZKHgISi1zbd6pVdc
ejHK9jN/HPB0p57CAh1kAKOnncCSlbI0Q4eA0rfBaDD6wHNchIZIbYijyAv3dy8Y
/63jYhsKomxJd941+nXrtc0fGi7HMMOWvMUtTD32slsZBqM5svU8Tle13ch/kgQF
+szGuaP4BTcQFkMPovdf5zLZovAlNJi+FGW+g9uL4VMgJOS0EbmGvtKO3t2uaNXh
9SqfHdnWpJjoLOdxK/LixdCCS86PIG9yPslme8BikB3g8YjeCnTOPTIOv93lPNbW
ysDIabyX+a5PhXBKPa3623VrmtMzU6HZibDnyw/pBAs53x7BYE1Is1jnFyk6oiSo
d8GKgvf+Y7zDiPUTFl3mJdZ6hQL2CS0w7iMu33svyyPfRnGEwHe75nqj+Rqg99fD
QIzRZa5C17bSl7GRpxHSt4Wu63dB4vXRGNtMMpXdwmfC7RBrc0Oz+PhJ/nMPFmoj
yi92k7LETyrHNK73NNwdoH72tm/ibFSs85NHFlrdt+cX4CTQpSAn5qf/ekr4V0QC
IgfGAlrSjBchQheEleD4JEwkxgkJ6bNidsAlR4e1UA+UmpQl05W5v933TWlBSdD1
KNTSV9E4nxazeMgHKRx90CY61FeX252WGIgzJxWFtYt6TvRmSIoU7SOwheuoFu1b
Qd48SYPNZXnSfpRFwMEnanZs4kBGXRCH4Fyr9e7OimO47e7UnQ/7NbXwS6ToNcFu
/zo7cn6QReVWjc/c65VEiHMHdcXVWjIDJvvQfevysOjKawYBaFVkfVJ0PcCQ6Uua
LxfqIrYEsmBc+eGIl1WhjzvuJS6+b3RANkyo6jw1a94NdpPx8Wn+zfNzFoZBryb1
LNatjcvGh6in2qclgfPokk4JTOoOgxmXUdg6ReTpUWOd9AomZkTFZNCKiSiwYtnc
EtsZ1KYQFlPLvXxzXIP6tTj6PyCGqRhh6Zu3KBSoKzUn73s5HMtI+RYCfZLZwj+6
RaMr5fDJSskUmr6J+8HgsqF9aRF5p8xhxmaz8YwLIxYdwTAZacX5auGUY0zyBNUN
kLD+j5sQ7tOcAz4H+3d8VATRrC0zwRdGYLps4GgLxLXF1mWB4DOXuITNlCgntvcX
x2vgCcpn0oBIrXJhI/gPMiRcGoOe7m6exwf4PBtke8ikElKLg4oj+G9JYCwurDyS
94MPhZoajcRe3NU2Qb8e591Qvr/eps6KwIHk5V6oSomHq5uXUf9NVfaYJrnYKo7Z
WOVKgmUfbfy6SCOqOfVgVMq0mOKoVcHRPl3PHb2zfC7oMZk+16BzGhhfrp3n+a+J
Wx0FIfw9yFx+uEZnNPht7ko24QYFEkkra/6fa4WWz0T57TgA7R6szibm08665VFl
jVDBi7JUzJ5c6N91Ft6ugCdHZlg1YAT3omkPjTOln1G9DZiWBATwQrP9QxdW2f9/
27L9mvzBVrWoM0P7Y/DnZRXgZqrbGe+S9Bw9Vx2qHcS7a5frfvXG6Dshyl0oo3mb
iuUu9H8AkACIE1GLU60h0hE9c23D9GthY/ZJjk+rUibyDJklmM9Rgy8z/0GlQjm0
rBUqHksXCx+ouSa6CBgQFWAML+Qe4V9MOxDe8XQx7ufWFI8pDUJy0oxkzVLkAXp2
en8i95ZUSzuVabf8iM1kN8ap8lw+Ov9J1HdHADGnZkoh1Sl72PLlzHOlSlkekhIq
OU+x6S1grW00/p5lzjN6WG1ysoW9NU6bjg/e8n1OVUvsRc8ecmt6vi7JVXhtXghN
5FcAgVzZp3GWmqLtmFzS7XsB/T+4b5xsYfVMkOHGSFUZ32RuoR2VtfqKrN7sgcTn
xx2RVICi+2hJCywLlwZgRfUwbzNiODowdaZr3i9Og/MbZSE+ZEADUtMI5x/9RHji
uJ5FrgIFyhxv3mUNPvdGowzZ9k7H+k3B4es7L8z1lWi1TfFMTbdaXtvYgY4hC+uS
WXJE/uxgGt3+MbIeYHd+jivzwQX6n57AzcfhNpz9fLljPnZhqlVwblP3mHr8VRdB
/jMxB3og0m7dBuiUy3C1hSwijbi51eruykRPD+KSFRr8Q05pj+J/Xu9DrufH9a9x
PX86uZlbmspnd66myGoZ+HXSuhcC9AO4D3GP/Zosmr3mIAvQ38qCRavT7UaTMnSC
FAQjMMvcTPEfuDgrtW5rbAL0n3aadKwwMGmccddOBNmKdV5Fy12qHlSCObzgJ1uF
m+0RIunEpmpkc57jyoynRQEFedxPoJXPsJTCqeSb5FrXkgOiK6t0CSwa2mEPxvZf
NFhUMbgdpQN84L3VPnddwmM9alX0uqhTwX/mwAYdd20ur5Ku1u2WW/qZL7174UqG
tBl1sQf867AlXFo8B9WNE34/bQXUV4kurYsdLq2BrDuk3SXZ8yWSY5gbDluHl16A
UDJpEuo3ah2SP08PSn0ZYS7PDmIDR21p9MQJizdwzuR4JVKnno11rL/FXWfHHO8+
fNR/bY296oLZa8DMfpqNWdDVqox2Q0GXiMXCOt900fCq9EDT7/+fOCxt9WBw9U7j
l9OFVs/rCYyaC5MApdljMG7k3e09bGA4sl0ERfn/hPlUJ71ioZ/XdeWegvpmXDP7
/zYYHFo6/W+l5BH6dDdb02702pxrt1qTE//cLzGD/FCt+qKSw4wTPrbh7+MztBtA
CdVh+XfZ0/Q3ada49Ocl7rthEh+MAYYxC/domMZ0UvGsdZDMG/FL/o+6VLlU2R+e
2uq1vxPUmqf6uTXbsiVl+Cz5htWD09jt519BY4zKFHJyUrI7i4IQgx76tPseLiaV
FMehWFZWxhTxf75wj4ibauFGcLF+He0FN7nNFSORV2prUeSYJ5OtcBUidmXrtbHA
wpDbAnfYX6GLdXsjkMulaVCAZ+ZHrvzdgPvTnG6CbiX+JlOk4usKU8/1UH68IBOt
O9zJ2+zGE8aR8l64Uu2ycJp6iyrp9gjB9TJS0knKSP+NdIvMnG83227XPDX61RNB
Q3ZRKNopyfXKv4VWjVXfXDAOxpaRmpb4Pj7HDCmHrs/V2o/7dgcNhFm+c22XYfVi
q1+Y3ovaAZs4hwqV/mxB5N8XiWkcDtXn3ixa5Nnx+mZevGZhQp6ikO+uFDqlllhE
TsgA3n+BMaeOls5T0PCyJVjUb6r40p3x8xdH46Ig/aAJPwB96hmL/N73YXNJF8kU
8pf+yJRDCc2vFRhF9fLE7Oe9n1g5oYV3tAbZ5PSasPbLReCuEqDz81BSVgqie2il
qPGeWkMutBadSB6AFj/qq8W9tD+2BuBrnwXg9RZQqbwNI45c0lGoy0nRhmnZgyT2
Ehp2OzBLiynQkjDbA9ajFrzbo92rv8LRNEJ3U0AIiMww4byU41X16sRjyE5zyDYC
RRBnGbwBQjzB9nykrN6KRoQSWPlQg3UbfH/gtM8F4b15Hn0XD0wmhx05CKF2svkL
DyvvU1nr4HdtG8I9dslzBUDSTB/NoYl5cb9hmn6gKB8AuWUC/0pbbrBIv1ucX/8A
ZSVcT9WTVYw3zmn8y/Xy16POV71+qE7zfn7Hw6V6t59GkzjRi1CWfipNn8/PpuJR
e/LsvTTx+vDhSvAtVqeHqQ7IFNYNBi5PjDkbxeqKPM80Q1+s7Pb/eDogcuyQteZ5
2tXB5AiMR1YotPy/dbxVNfMIPLKGn82+AxnlbWyAvVxA9bqGaGuqHpSyaqycVdjF
mtu9e6rtQBXKaA8P1goFDQH6B9RmmBiiaJrxQc2PxHUgeo2ok/7y5Da4Cxmkr34K
3kLF7N2Pqrkv2U4MZ/dC4nSN0YGJQgIJ4rapbf8mrvOfmqwXmv7EXXlUB35IRaz6
5mmHPXa1YmB8d29FNlNKjo+sl0dlkUBLhZO8JkOTz6mmC1+i2wZZMO5vZ9+8M1b2
+Pt5NeS6UursH2rkSfTjyqsP8l2rhLlP47do7KgAgzfT0RlaaeAGaBPJaMXNTOEB
MkcTWxFGLyyAkx45GzJ3ad0vLZMLS6U3FE0LGz/0YFtuhMu0DKnVBwbphOszGIQm
6lxm0Kk3dM/siPFhxfQcLtYlzaUhGbRTdP4IHRRx51MHKv7VbQKNO4WmoiLwzGst
UNPWo5656/LR6iHMGYlZTCDGkErUeEVXzbxAG463nvvm+Lf0go0FRESr+ko1seC0
/9QwPAzO2AwnybGillpsU++nxtTML+1SHDVS5GCkYXCIPct87u5UlZGmCIMEx3eT
R1PnTmpqYHIRrb4t6il5I9Ovz4fPyUJU7nGou/xfi2Hm3lzGvyaqwn0vR3eSI33K
XK47Gl1lGLMc7ZM8+xljIYpphtS/+b80cuh6M+82CtUsSvr9DRBLTbXEOdEyWxtJ
ye6CR/glDkPtkfXVeKTqc+UB6Wc+mX610RTwE65MIiVL//jUeU9C/0FjVEDXUA+G
5+i0cEqgGqvZJMSneSwUxQxZ9h0L1+1kExldRV50rdZWl82TrFrd39ennKuH2iC2
kMDCVnHOAXzKnErxVsbrHrbJXc9zhemaq10yRP2lBdRF7nMdJhoc25MBWjs2l4Wc
2NjRGIqKJ97AWjr+mwwSl49jv86w5zZ5edoh1llMXOhWD45SVVIaGV1E3LR2CrYe
1EU9UJm8eZyuJlb/oU6qtPzFfhX81sY3KWvhGGHvZAxH3yUpfNtl3O6pFUxO13Dd
jsQtm67hPwu0ZAbj/IOhsQm5WA6e9Y6olhP5xoJRdGKKxYR90R9xUvuCx4AyDTYa
ryLxB2QFAolUtbCIN/jyEEgntNF3TP3srMDHuapMq952gJ/psafhrK5c5Qf+UftG
70fQR/hsPV7GQZ0T7NHxYiXPhB36UMHBvc+ulRv77/sLyxf0MByuSm0mNYrvJbMp
LjXYSpsPylkbmmAm1Yhss8xeCWt6Z1Fj3qeVu2RbEeGVj0FQexxuQ7cmlNKbWypW
mfI/IepRIpC5uPfV4NXtRPZxIfrMyy8EeaHDp4V+udpDSuTk5opMNk7aiu3oM5cF
1PAs80rxus8XnWU3VB+XFQV7bZdnB1QojF/9VIQgjvXq0oDEmjcIfVa+cB56S5ia
l00nGDOEXupmYOVcHEnH1tg24VALUYlfIfWnX2NYtoma7btkOWEzcYTbTYjwcKXi
QwsYjtNeX9lCGcOQNcqO92pnfOdi2j0jk2kGM+mDuyOrKH8MGaAoFOm1u3UzzUJc
1di90cQG+jYK1NbxdTZxO+yomuvtdJau+zhYUMO1E0zFrFTuqX2L5KH9Dj7HO0EZ
TaN2LFhHzv9tQLUe23X28vwZiK/uxmDtTVwFS/wVARX2ueP9vPkQA6NECR2+nse6
GvNZ+emIi9HMvgrXfHwKZzls1IsJvdrn4X/j2Ggp2suJxjPdX1aLOq5SqB9FHCaa
5tJJqjdQHA+Hxk6wd7wnznUWgpgq6Lt29xJJCLaNw1uQntYs7DGfte4BozgyLkEH
EV0FdffaJtq3I/aMHeWhaBzl/mtz3r4J9ihr0uQq+/VeFUrw0DUQCPtbP5vcz1GY
qohC+baswJCnFZcXFbQ9H6zHdP81oR0KVmQM4OxiJsvsuJczXN/2o/7EUTm7n7hp
/chz19eoSUN5GyF7/+dnKaq2gBPW8d4xEmqGyc0f+90kjPxFS3B6PnsBLM58S2uD
phrBNkn/RzxZ1a6ck4h8ZzjoDwgz4ozE+fMyEnvBe5xaR3rRTT+YnYDegTl09R9x
BKO4Gtl3PrOV2YyQYKXT8ukCiQO6oAAMLu4p/89clk4OoW0t4ddJyPcqsVrIbleL
l5KbSXCoTJVRVE9QdUjeRXJYIkNTGbQq8gOyCu5A+IjoxnWNjyQ4gn7O2ti7QlN6
ZAk31+tPa0UXbQYhctw8khXzpr+XL0PvlwoVEF5NtTC7nfxsCImRVltNtmkDlvPy
IYYhR0OoaOwAgXDjfRQB9f7QgMCn4ihhe5mfS7CpEMw4Uy53jRnqfs8DaK1OvJIR
RNcTfQCRYSh4nRlmbcXFxng7Hj1qgHLd1ONHA1HtdDdGRgYMhnijftMpDOJTlwEa
8ub5wHcnV/ekvpajrlTuZr2MUPhjrTvIc1KHvG5bI6k/LGad9l90v0vzIwrTeQn2
J3b/AjKeBD0CzP8L+bjXgtbAgY+TMgwi40zYqUHZhyRH7GUWRcSBVTTNMwjxo3Ij
vqm45KArL00zsTsKM7IpIvnZbemmIGUNTvkaESIsEYyocAFCKskhm8e4BuoDz5GT
aFYV5jodj79yDF/bqymsHCMlaLbu8mpgNsmRkxO5r1x37atvc/SjNe+jT45HqZ/u
zq7+7/rUdAWKmT2CeGEtI3RFmzdGnD57A23aSvNzTFo5EtJTCxrie3SeqGTY18Ce
3Nr908/ImpJTnD1ZHoiSkisBc7TbMi/m14DJQsKdmwL6yY06QDj5zoae7j/gd9OA
Q79QguBkeRiSFvTVuzanLX6N/M09Q1CvkaOVaLwwLfoK+5qyHQF2IIoCzUYnlu2s
eFDrZnYtqj5HOOalFxc0rJdb+XwpHhvGxAy+nXWX/+KBUrOG5e7FOez0nK3R4JDL
tzKoVwmdHojOcbHxCnMUqZhAX22yeUghcRUqDbowWJvXEjzfltSx6MznHapbnCWb
rYASH9w3Adv8MhInNoqYX6JwzAHUOrVdlsNMNN+i0m1dvH0iZg5AhE77VAECPvny
JD8eFrrDAnv++6U5zL1Qcuo/K1PmGflC1r93apOgFc2Gn1Fr5zy0oFyHsjvdujOt
J61a5FhirQVbb6FV623ZWOefPksjjXcflp8DV5Tp9tnsXIDFFIySdDeYjUXmaeXz
3+7SchSa4f9bukh9i/AdLvMs2z2PtUmUzCc+A4nk/WDPbMol+3iNbyHYjCRcwZZr
CJmZv3u1Ib1K2qgp8lpcyJXohI7oj5NmShy6h5uV8BSBuNgYtQCnxB31t53FTCMZ
7KMYGp2+3XzIZqm4XJSltcVKwncctpxL4GSt5aIHmU2xmoBVtWbI7z0ooSfPKLZG
qDyyrPrquRyJtMGfXJwiTJSgkmyj9/hxpvrBzcPpRNx0crH516rGCw/tj1OZlGmj
yOLLH6t+upY0aWseCG8t1DZnpK3gmpwjZRftehZLglHl2vjSeVtu39421GCLAYvK
BaWLH4TvFNw/5CqsDzH5IKa5MLX2QicIf+1y2QwxCUxTYZnRdSrgb+jY0Wmk7Gi6
yeLzrVW2oMhpvaZOgAcAU2mXhEUOpvpwU3Dn0ONzxCXLaDZLbfj5eD4TUEVXgMOz
8WDI7jR8iDyzL1B2C0Gs/0hJWge6iJmOFRgAqMt9piFNsFtzb+ZR07/kO7G5k6ae
VQrNEQzIXZAqT6CwoD35uMB8NF+UXvZxOtjbtjRhMQKP5dKmfi9d/KUA3sMBCZt0
rRjFBFdI3jVTkIqB1rQThTmkHcTCwcSRxX3/KpjD5ELHRYjTUwTUC9Ok68X6AL6r
Je+R1cFFSOhHMTZVJRveO70+hTXkZ7NzhJ4PoSjV6VYIFmVPYKxhtbANhOZerImj
B/5w5MxiWrl6pa/RK6wrbVyVa3SoHnNKmy0LCczTtn5chNKn68Z8QGvcZ41oJlNU
IOzL+MO4GU6zkfcY4Se4VjY4LjnvRZ3rPzuHq42V7rv+lYzvqO25ToTwwneTTPVy
KzB4qSu9hSRHZ4IXpXL/bgzIMxIi1B/SbHkztsRkhat19ywPj9MjbJ8gJw5Otf1f
bwwzjcv1M2jq8DkF7S8VFS1ACq2czJSwV72RZqHKMuJjQd6dCMBQhMoFB+tsCzog
YQxs6LNlaj2j8UijhDfY1fEUrl4maMjcbOQu4EIjyD8aQkWV1qBOs3MaiJSjOuKq
KnXUDGVe2RauId93Iy16AG/hByxIkyN1Ct9+nuCIBEuJwfg9mrllNGWBk6wUlxvR
flBY0mghrN81+xhAJQ0YCzG7JfEnm+GHafnwCg+6bUFnfRDpJ10NHdBrEOOx3lv5
jZ3SsfsszxChy0uaXJEpZodgUEBcs8ejMqIjWdjguruGgpbkl7er1eltP+e92a4z
DBN+2rg+NToIEyKqMVtNhs3tnI+CLo1ARkGkjJTMsA7NG+zyOzLpkZ9zL1v2UZsT
nUfWIDYfEQ2/PslzqnXA8MGXKo7zqzI+lKNELUFxOcwfW0w1yzw97Q3v5CPMczA1
sV622RFD8T9hQK66X82v8ZylgDSrpdW1clwtCHOzRTs7CURcSsLJzaFvwifjSvQg
OdJho8G8JL4O+VS2+EmWazxyv5jFS3ifzWDf8mb+bJbkkWyPkw/tmTB1jV0f+4mS
Emm+TSEQMY+rwZKRs/d0edLf9l1jwdotqJb09yu1BHnAWWuXBcdxpquEDtkXacko
Ny4imeBmAgm0GBNJnnX8wR98TGnTCVaLtAd7ySzy/Ux3NacAcL9VBxozUyF1+XWC
RZDR0UiuX2orjA72iVOWm1ejEiOXCaJOiRvXYkNPppHEzUIsuQ04/YdTo2xPy8ke
ZXaUuR/mMKxxPCsPDlIOn+b2CA84uWmq+5S0aS6ESXlbb2cJH9QXgFFzFjU+zq1F
n20MtYiYrZY4TS+fIMKA/XOMge+9O7pu8kmdd4gLYQvuFaEbfdHrB+NVmuzSJl+j
k8zZStTywpGz1pLglSxOjkkTl231W2i1VRAsf5DT5oBmPTAvH1C0vFpXW2umSzEQ
B3bMKICLlE23MGPIESLQllIqp2gZFDj1e8tknWubLhL3NGelZ6KTyJ81Fmpxm7cQ
LqxFUQtadNsQEtuleT/f7PlXBjWpCg8LX1Ff8TKSeA5TVsJyIN1kpDcBT/pBZqpG
ChE5m1WaMTIEfyB4VLV9j+2bTzTVibnOsBKQUp5pNGQOoGr7OPEuWjbjMsa96YfQ
0WR/EXvQlRwGB9Oru/21rhHTUgStFdpPXmmEdCmsmsGYt2w626KBpSSgYefoGMv/
uK4rSbjc39vsc6OzJkDrq2f9p54chbEpEeWb/fs8LIKOHRCFyU2ME02OJfQerR2a
yaBsiP2RxfXK3trD+QxfbKzEg8MCLwRIZc0zi9Jg/y/3ZaXhihstwru4aN3uY4RF
jamE98VpJoaTKirjzwO8kQY895p+PKTzj6m9muhY2/iiTpAGUP+AIHJMJsdh1Lsn
KNc3QmSAvXkCYtkO6NeQzdAENwXmnkJCeJiSfXFpPMmRaHDXMjwo5jQA/nk/dxgu
rMckTDqWUjgJR96/XJQO8SVO74QtFbEnaaueL7nQoM+Fz84Wmsew/l+4QM3HJYbR
obl0LBiF0GGapDwf74UnGG8MSntUIU3vGIlTyXwp90tlYUwhYu4wknfzIL0YlCd8
8wE90o3HneVjPH/zEwdLwv8g5za1FlMJvEDZZj00JwgGcjwsKDOvLGnPtbo40aIJ
Eoxbpio4sxt0uBKtibyzjIay2UB3ekPDf9IYzNUfFy+NfVKeY6nDkIH9RDY7YJ8C
J1ga9C/zLojEyY5Xely/FDwpZIyIcPKRJ2q8TxtjCioLLYdx+RSdRh95NA0H/vUP
IjpbEi8n9Cp9XxGpLQI8OILpC1lS9sdF0MpObhy7pfYSV01nosyAIBhJO/kJ2ZrJ
axBMmFwYlnbp8EqNIbslR3rQLt3jd0voYSMcZVO59bD8eHDpN2H0mtkGMG6UKWth
izRrckre/xzWmbYHj6rNMFqBfwo8b4MOdIOOvRmaCoPkgk5DUb30+JjSegcD4k6+
3jpep854kFE9w/mBti9snTh7MV6xrqwmkoEv4nVmHnW9q4s69xF1yBCCar09vdH3
IQbICG4Om7uJ/eX64TXqHPs2nZjVUzyhdGFLf+lNpwUSodFxqqQfnb4qfvc0b1nW
ifTGmoGo+Pe0z6OLx66sFUi5U6Dg0CiBIHy43Lns6phdKMJiFdL9x60X1tehkTvb
e/ogBz+3nuBd5vsHTlbONfx6t9M+qbT9LTybkXLBEMW9/mTaoQNOVfa8biZRJprN
zkO2OHZNPpKUroruIO9ercXj0PExaYiGpGIT4/7mcq6WWGWW0H/dDlmgSMlMNupD
HVR29oISDMMFC4gZ9MOSv5ungd92eKPR1lzP34geQNOmX1786m9p5aJV91r0YZ7e
LQCipOhLqYswywP74t4FZ5pSGNVJQO64mbOSy7VUHq6+pDRPpZI85M9nXq0YthCb
zLO1XQKlGw4cWYnJny19XTRZNLREgzVDKSbzUUK90rjDlEP4e9bIZ+xmudgYkjU8
7+A2T3TV3cWcmSCf+QVgOEpPkB5XCv1R2ivdd3/V3Qsk/lRiuPR4aHhoIO+xtTkC
OEl0LniVyiCg8HN1GnjCNMA3a05UJjPK7d3JjE7MuolpsqVqewla7FKVJaY1C+kA
rEvDD+im/CJITJ6Ok2jUS/7kzZiHPOV8Q6GlykENKjphfxEQ4GKLZItLEXSIndk4
9oztPBInvQ58jyXy8Vzq7t0080Up0z1D0m9YWHr0irXdt5V5KdI6iprOHoCSjCDt
My7aEAXgMSC3FC53+EnFU8QTn+jmBoYJzYdWqmJKjjIMwZFEYJnCBelzJWI3st+F
tAsfdiS8uBH25QWd3NKiUwRiwxN3Ecx+sH5yGn2uJsvCGemCHy/yDPapbzV3JFgD
EY4meMnBQgJf7WClHkK6UADjIs1Z3uBUF1YnIUwOcIF/o9ZtkJSfqAxa2svTvqKx
CZQSxtXxNdHZX05WnRoQrBesuwgwn0BtmpBsCSWmeC/jlcIOXSkrb46RMH4PRTns
YIt+GfoyCpB3kRUc/APt4YU3t/y0fc5hwicEGBa4GA+FzgR0vhZ9w13fcojY0M7C
OgkRwSgMLDbkwI6juqITIYxakfVBUwYJmjsbw0Op7LFmGssVcfWS8nRxYZS2H/Tv
rDxdfB/1oRMjgcPbiXS9nlOBmIyxGgI8yCNd5mxQ+gjwyJZjLtXDFOpAd3/pHOoL
NQu9an0PtoycCjiV+26Reyh5SZJEOCXyOJJ4Ad5UZ+kaLJ5qk8g/ByWKD5joiv7p
MoIS8vbaRexTSqxI/iA0PIDtQ9wuYLHlWrp9I/MUqdRLS+UXbaM0s9G4ORDhF8FX
xZJhxlWY490/3KyFRoSs3XBdTn7Fey33J82u+gMDoRPkelqqTegnw36NOvg1ugDu
Al/DPUJdIMFeuWgRiTfZyw8d0kuB45cVOjb/yOJ6lHDttWhjwHZw9KwzMzwYrJqA
UnjpbKQI7u5qcwa6ISHpc3wG6XYv176L2obmWXJxapdH5dIupm5Pv6AFV5rkuXiX
etbvaF2zJBt7ZngWzopn9UKaM4H/MD57KfSms5SDRuwY5309hiltnW3DgH2pF1Li
YwbYzYezE/kpQ6AUw1KVHrI+7pcszvjUSXQHwvqIQTIVgl5xyj8sBMi1d1P3Kzek
Avm38fxy+Z7QFZih7/gHVEmyZbHtX5FpUP6jKEdzUMyQVaNvczUDxfKSrzCFmCPU
xjrC9JhZxp8mpYD+NIi6JSuY1Lw2qU61w3jfZTqeIaJ0KVimTqfAYnfogMho4bfz
pRBxQmjIVpWRBh8yRbmjJp0dK8XMVU8UUvHFCVbKfNJI3v/NIWlvPJRu7srJMb6a
3ON/D4PvS5B6C8QsSvC9hMv6yaPeR8QHdA3NY3/6euWkRGuDBA++31IJru8LinxA
8n9VaLJ30DunxARG1HI0i/QAeg6zbMzShIPpBSSUHahnayaiz34UE2k7vgWQYEXe
vq1ERT2MtwO65ckOmRjm1Ypq7pNtPFX12hKklYGU1YxG/Td3OkWlp0gTu3U2kK/w
Lkpc3KA451XeYrag2iqB5bczgXm/cEJBhsYkuOc5QNRyVjP/gvMuIkQmrLASX2Kn
uHg0k9mqVtEqQBbP3bDa1+yi5/vev7dBXPTOJMCxHrLJyC/8xXOeXCBeS0E5jM5x
FfuTZCvz/gik2nwEqDDCJRjo2V98QG3FmMJLGusihd5z82CczJlaGRTsVlcRrN6V
1VwgtYoTcnIKxa2qlK2rNbiEC5piUurKBDctUZbo2S3iDgVvWvPINux2hzD4KnkX
zDTLPb24zYuOm5TUbcHmVm2NVWYhiQ1MDnljF3P2ibh0TI1jHgZw9MxTLrTFPI9n
P+D8ERyxqCDUmMaRfVWKaBqWNKdth5fy3ObXuUun2PjzDrZIvYox5ah+sLvoiBzp
TxgIOCGxmVSpSBJX424Iiyll8i1TK4db9fVjmy40WDrUrzA/9FArI1rgn3f+IcYE
r5HcP9T6IQZP3nRc4qh+PJrHvLUoaSWyJmUSTfNIbArZufY+e9rVDa2Nnw84Y7ag
UImm7DtwASAea2iWh5qCRVOXDqJBQNxMN24D2zxM4ucDe9iSxc6FUZCp1svnTR+a
oyQOxN0QxbR0xCbKn4PJ4cg1IzKjUciNmsvGb8+/srzohHf9m8nge1gTvMvHiFD+
dRyIwNVrC/SdLDrcEv1yAU+hOCG2ePDc90LPucSY7Uwgha0J87P3AY39JYjoYa9n
TaJrSXqKGIxXiwyldDSsVpvih202xAk8/OWX/aqFgRwIquhWSxq3v3K86ScqS7tk
px3hCQeAczLF57hZev9hz3DQYUIABFN/zlp2a8YpQTF88dniz7LJt1oN3F9QEX61
RWUXDOzmx3GGxRlKtW5U7F6LJ7FImw/U/jw66mGoIb9A7O3ScEWjJNuqDyynEkFv
3hUCvrw0BrBQts+OQ21/PLfQvE6fwOMWDcAaJd9TrOGg94MhIvhZH5/KQFZ7Df1n
gZOhp26lcYLlr0HKF+hnz4P3TZS14RJTvUGVEO8CJspB18nVNinQSNgucHkwgzHx
nUPk1dD9Hlw5lMFujA1SC0algzdt5Aa+k4AQAxY8yiiQ19d6JM7tIZHbJjRSHl5y
9hAp9NooDPpBSaQpZkurU55rPjZdV5anfZKYhvKr44yEIgaPXYD/Xeg+u6LLScio
Tko1u27vwT08rORdxt637E58E/j6I7lGRRT8zP4ZIUgekP/wxexdWEbauQ518lWq
74OTbntKQwC2VefsP/TTlm4m73K8dC1cR8rhAfvdRO5nH+CWVlfywm4ZyB3hskaF
Btrgs3+UvU6j8Ot0DUNTiKKVHHyzw3IcL2ZlDdl+acxvtIbDtKLNg+t/9f2YpEBj
rp6qwEyI/CquuCey1ClDD29N7NTH9VghCOp24BJWuyiiL8KSN+H+wq2CZy0mlR+H
0NdhDhbF5R0or6LsO8ctnoxo2gkjHvyhMCoLBrKUrFushxfdmC+ZJObV/b8yV+cE
0YOG8PtAovqfw6QTIUVtSvVKUCr5137nfg66nmkx9nGFM3w8SQ9Deum+xVs5Twq6
orCoJBUZN9xXbwCUFkjX5T/pE2QyifvJAJTM8qXo7RcgKaKgIzR9OBsM8iFe9qdK
SnQIigi34y3AQa1pO/UCipUiUldK4m+EzoYmkpeI2Uq3tB6WZBxyY0QyYyEhS2Bn
vmI9JM4w2rF/BCA8c6mVWsWYspgXIKPD2EzXLQodYsARtqacDNuWeacxlzszN9Za
psjopykM6PjaZeUOIsVniZFe54oYy5ZM4x/loxTsG2hrb8139+xgGsVsUX6pbZis
oVRprNQusYBRscV2n8B0I5VKXFBe9KM5/mfgCUkXfoNwLeh0wf8OqHwdn7Dv9kuA
ocHALMLIx8WnLfaCbPmaaI/pcii8COUksw44PsmKK+xtwxs9OPtLSKfd4W0sTc8g
f6th/XDKML9S92FIhlL5y4qDlWr4SwZg6ptXaQQHoQyjcXExN/o1ZEaZxXUTwnCp
ACGmruyaf6xcS0qlTY+IQTAQ8uTOHlCJFvjKnGZI0+BO+Lfyu7wgxl6q+wgXDZPy
VcXyTtl8sxBMjnB+zWt9eT7KAJw/1LGYGeE1yLT/Kbde0kB8MwbLHrkEXFVe05ci
bDow08MUCKcN9AQAqfXxuQPUMi1igT7N3JwoWft3feSs+vFStowTJUlIQ3GYbzF0
uT1ITJnvjd2MbzEo2sTL3MX01gTbSGqREK/MtjwSOYI8GQx8XH70d6xFfqlmYykZ
ZQD0Bd/CVE1i8rA2Wf/qfaaombmYDnuwhcw4/cJ/3M3Y3Rwn+TDxhkFiRBytBfTt
s7kvoxr69McZVT8cLtHP/pDpJNXwv55UUWfNENO4SAvAbh6dXwuMVrgPVi/joQ9Z
9HNIT/kgGT4XqxqgybXEnhbNWyDcdpV6Kv38kAcrdy+NYJRNFjQJXVfmK0IYd03j
9ooy8m0ByFxWQR7xaTYwYDCiO44xphxB8BjqMm26H7G5IytIXEsm/TNtwEtrhQVc
2ebZbn7+iDP6RrncM6s6eyJq5OA22vVArNxg9Q3+7VxOWxgI36vCqrCpvr00Tr02
Hqs6CilVZwWY1+ICTt6ofNvE6BYNoNHzSjyTzXR7k6D/FbUoP82glx/8N6xJNdRk
xzsUIDgE+2gMZORJosofMcNuGUAha3yClCVWqShuny8FDxvnVf/8pzDfHlEnlMRw
UDO3UvzkRXIGMxfPkgcKPqNUFS3jEe6NATBwUlKFosSsKs61kk4tYWSNorYrtMU8
mjgFihQUQDydK3vFIXQP89CqRCj117TGyAo8dHv91bhK6w3SuhmsacmkaPX7vL0X
UkSQyzF3M0YlagXhGLUcN/I2ENmYh9cLJA60kgOkwvjxiwYjbZxmO//qJbx7XHTj
zYVh7W3cBM+hD+1HTrYHzMq/46lt+/EUtbgyDavcXks4hNeO5tOOq48w56WhZ9Rg
fo4HITbwC+SaJid6jcnXZCbuk6GFxYG6tvDvyFMLp40+3bzpFZ56yUAJimtbFBTs
LPACzxfBoQ9CbfPaCct4Xilvf9uqmkQ6lahFaRIBhcCgd8TAVB027mmRC9Ymvov/
Bv6caxF0fzXE9M/oSNYVmL4I9mpxOiHymoxvk4BKzEG2obWyGPHp+fWBxEP9dQ6O
VtYgz3tEgrF2r71XO5g1eg4Tg09mI0RNVH+YSN3/hCYTcnWmdYve3OOsmWNawuay
CeFklJlIjIN00mH4WsUo/jjgbcRARpCIvzlwxypNXBXjLWn8w3u/jAtU8G8PctlD
U62St9LR0T0pM8AbNMSgyHTl2ondFfFt9+0hHx76jpmNmPKq6VSMYmCR4ZKFteGy
rYkWYERGT+fmixiP9BgZ0tUKpU0VPahWVhKUmHMFqC9CnayLUMddht2cDqCFcf1i
IKNTKPXqA2f1r76nYTzMc2YveSF1rPdawmq2U0Lj8J8CgVanUkbbnVfv98ELHnSZ
iF5Aeo9+xj/vs6v2iJU++/4dZgVGGWVKSSn9ZHGGVkrbph9PQiR3ODafdQnX5V/4
5bNQL2sUjZbjUqOtp4iab/Wv7CPOGpBzAx5yS0cSg19ka80zm5q2Y7BmWcAim2C8
H0Vbeja+FLsUZOX5P2Cx4U2tFFoolSbcF2FVLzH+DJDlvib7S5vD7d2UsaxdqDG4
g4fjdwiMuWQpLyKCFl+kM2uzJ3vOCG2ME4YgrcYJRS4xRyq4nbomudNd6UaQJ/dQ
+FE+gmfnbuozXLEK/KVfG2Q/RZqMfHDHeQKLTm4Gy9nW7KvyM1Tn4tzmHrc4BzZB
lIH8ynypCTgPI43Ap985fjS41KWGNuxeJwDjfhIMQolpZcCtFXYgYCD8Kf81ffw4
M9yZ1rbsID8HwCOqb022+qvNr9E68+tLAKnwAb44zYfg40LvdTtgVPrG4KFo+DZ9
mMOp0AwTiep2lqauAdbnOGRKYu6MmxHPkGrm/4ihGLln92VE7jWxWmQ4lJyqPa6O
4aBnNKaYyl+tJqmuSxXa0G+NiUJyOvuBacn+Ox0BaZDWB6NgNPShaY0pvS1L3RSx
b2wgdWOm39qtazyTuZjM9er8SkcwS4xv7CWIgFYLHR2rS0f3ylr3dO6HxzEs6C+6
I+qj4g/ZogPMapny7y5UeYm3ZJA3elcVGy0xp9ptrXFugY5TltNM+13uJuAx4Y94
Dd5kvPSZ0CAFdhgha6+m99B2Y0stEY5bB47SrP5AOIs32HINDS3/6iq3/JXMIA6F
5qUoIUw7FAbokwRXxM6hGzkgIzckhF6uQmFTgBUTown20hI7t4UTKgFqkHZZtsu5
2yfGND/UMzdNKXg5wTlGT86r4RDT8Q5SmCcPlRhfkyClXlPzp8G68lcSjnBvzZxu
SJHyaTz6mwQApyzbOTD7K6gW65RMpC0EGpp1nVudPFlLszhlz9LoDpmJECPSxnb/
j8rsgfbMqXkIRTyUM/XWWRqDT7pwREavV2XTUS2BiJB92y3HD+v3PeM/4EXB6hbH
R55Y/SRwWZ3aizm4YB5Fvqg1jg7/u5JnpaCf4QZ+pHc/fC9xchr2NBbMeG/YMqTx
VHDdbFR1244UgQbrKUHuRXWwUQ7sRH3yDZy8yLjStYqJjyw9BGxmfKxzOJunxDE+
6OEnkwe0dZ+C7uA0o1vC4KnA181qUbWf/u2vKmFeOyUEwPXDuxeFbN5lw5FxNPmB
MqMaTAsNcZgD7uvK4BA+nmFQNsWD8NSDp3kQZyHNJpfjxH8Tofz+z073tGP2XJJ0
R3rY4muqmGiyGhoYXffiy4FEGOw0u41/1Lfybx/4tNw5hCR/aGUxz722d+lKufdW
woaxEKbf7dLot1toi3quMGMqXobt8OECW1KoWV5poxPl4cJjvvXPTBr32uAlK0RQ
+pyLlNjFFIhVT+3R+fvl/7kxs/NIVNAKY13K7KySLmOqoTqf5qOHr5ZU8wfqVrwB
mpy4zi74r4syvJMhuO9nxxd1kMidCkISi2yPjBRxJ08LLAO0NuiiHSbaVz5xclcM
Y9mN+w/smxrIkwoW7uf4kMBy6KjwtGllGLx4K2hrruHarbCHlQkOs6k/7L1o3nM0
n2ekQDdDj7uH5YcUt1BEY5Lwb7b4kTUyq4u2WHhpFgT4K9vWpq2OTsKfnjvBJdbE
o3S+GL0mPXZ49zdltyEDAqRyq7sAr+PL3CJVs0P0+qjnw8EfBBxIWo3Eh0SXv7jp
MbKvRhRyg+NT8gPfbmiCi7P5gfI8IOmhXKIjLE7nitY0DgHHHLAlid+8E363Sx8F
beXtJ71ixIVtoX8//fha6cDao1Ba15qGX54dTIZ85e3O8sPBC3NYzJki+brriCpI
QhU9kCjNeajJ+L9OVMqJ9hV35F6MaV+bfxasDlYaaTjl1zeLKHDcIsOA/BciaFbE
LvFhbbAyQiQ2VUQJEVwGt0WlHa8eojiqL3JrPz3mTgt32G5Tx/o/1Y9bQZdbxz3R
CCDBtmZzfIYfV9tzFHdJqY8FdMf+s8JEobjLVva7er0gqx3Iffsec1eg0pmwbSmF
hR3bD0A9rQSoQiDgQ6xqVfs8jV42dk3INe5w0yMpPZ6aVMHuU4rdpaO6+fNRIvGM
JgEb5lTby0pStozc9xFCKqPO2ognsUXYetgqfTfNovaVoaqLtHfT0uzDGhIbEyGF
CF8CAY4C+sVVkb3/2dD+MIU8QZJryG+Lh9tg6xrWQlgXskYD3umZyW4UwCxwxUH8
6yGAVuuTo8cT3neovxzZwx6e9YVLH6aYSYY1I51pODH/+vDIylgMFSPfZPpXEzi4
kPcxIQkGlJn2yFGP6ENd5q+ZP1vdwPbPQyUaVca+VyAAYRhp0rsJlgjwcAlkQLbx
XFN5dVaLOu1Sh3rKbke83TA9f0npzdJ6th7gqOCH64X+zgPNG1Qt4QAcrakJowV3
e/tOChYTYQHgm53l07jIOYTdXhIZq68hW7iqfrBNTBRUrTt+n9ddH4Nx4E5bjB9D
PFqyUx26syE45+Cjp+Cu9qPnUTAbBYQI6RYO5ZeAqZfPBHqWuuiiHJjVTJLCzKBd
ufPRDog8FX+WHqMSKWjhpyuQ55pcBZQMdqsLIVNQUpRVKRsBOgRRIl4mh+VAAOJ0
9Qt2wi9dGtuWPpAzqHLvSvUZ1hZAuVf6OtBGrAbiTmcOvBNvZnK2E2dwQirB2f3X
1STIYwHr53mIK4NqX2Jw3rJ55/7aF+qb9Q/IzOL+bqlYCtjwSPrNBj9MSCboXaI+
W1lcTK7XS8CIBXQYswv2f1elz140hRNaTV1E4P5ULdbdtaEMSjvTmd3x3JPG1RBm
2Wdu5qUjvtfGHEXEVXOpYe2pfH8RBIlDziXxzbTSkotgK6sUxnRcy6mv8Fq6+ErY
gZgVNSzilMa9gsEcqRrqLDdi2056228QG1eKCbmPjVdYngcnnRAXF2K86j7nDZqa
6hIVX2V0QKDqiTnKVYm8rDSMIlUDShmf/VoTb6z/MAmgk9LNMc85h3ehDJ4f5It+
WbpTOGJhDNg42lqq4kCFRjo2hrmmCcvHfx0qtSA1FrSWKy/19zOwl3sknJPyumOQ
FpHELqmMxFvfvkSBH4KqQKraZOo2ZvepFM9bfP8mcJxZ/GGj54OO/CT4WO4dCeEp
oMbtWtGtpFg+22mWPqv4i8SZ3ex707mPfQ4kcwwY+8BbCi4hPbmI5tabfGlnQOSB
uAPR85LoRg+/TBfkOrDgAsT7dLDl9G5Eup0P5sPJqmEhVnBSIDSZk7QY3zDRjLYn
/P9faqAsmdqKWpB6+aFuwv3H+EU9o8ElNN8StEmtuOpB/9b4D9ec9KiNfFQIydjM
cB47s2p7rP87LizTRP4hJQgqeZj8n/sfJqI2KAfnmlZL48uLRMPi/W4aK6V5bmCD
kTu+Bj2fHR5heZ8D10eY0fkVwBsHBQ614JWq6UykrSvsrQfANt0W6p+Y6qltpF7C
JRbAqXnRbelk5OCg+jTS+Oi4u8sib0Ga9nGqbfyc7/Dhsl8AoYKgJJmqXGrxYrdt
GqIM5WVJttdPVPvypz5UVBfwLiYnh4V61FEpgLsCKtGAiGAHQwlshHfrTV0yi3iK
ktN27nHNHpihLhp7O3BPrBQV1+X+TP10/unCcNJ8dCFwMow6I8zkkGcewLrUcoE6
57sjwLODxc6DdvM0JnzC/ZbRp9RFLS11CqeDZzDTa1sjleKKyLhD15EAH9hq8ZKx
up+PqiJcriJqxd4nqfbH+o64t0CG+sODx+tZcvsTnTlWjFVW95cUXgDetncPbsNE
bz+mh+L6qtEb/c5iHWS+DIT3Ge8K9FFvyQzxYY96i+KTxxRl8onCQ02UCzMdB0AA
t7cPwzHix6wtin2/4Y/X2BXWh+aB1zQtf6/Rg/CbLW+r/TZeG0wN/T+nBcTgDdZj
c7Hg/p6bci3Uc9TUrkE0MD5G3IXLsj9GqO/TMFeqUKfL8BuNCqwYK8UPDGTxl7Yt
hjYp6qRYzv3Rc2ZGWgrlnVxdrNwXUyRp3/8JvIdlzpJ4e4dOYjEn+YO4FTM6t+qr
xZZ3+DK0f/e8xVzJ4vo8C/nx3LyQ15UWPp5Vwj7MCa1reEYrzkfS9QpT9HlkMZte
5IQR53V5gKZu7GFtbyZAf3X8nLWTqzHb4ZT4V0H/pPhxsaIM7Yb9PpXvLliEB0BJ
u+EH0PiO4bPXyaTIMThBzS93cgkU8tK8j9QzG8y1CYx27DHuARuO8xK0lWLQUoSg
LhhMsbuDRxkX18BKqknDC2TVP41hp8tJaLCs9FlfIu1TolWDGrmEJlgUreJtJslY
sT51XQVGLaLaQJyjIQOS51RGReJn8CgCPWxgu3eaNR13sDGby19rq3b8zvXyYZqX
roh7t3Z8fRrIpY8gEndOrQwNi5CoKUKSSq8E9BxI01GboKyM7QOktFJYElCrmwxB
7l2rCAu8QsWX1GSQw5USgi+KgG5NCTfFdlNv5J1xmh7gXwuzZ690jZSh9Z/ioCbT
R/XmCiFzkYMoK/l56R8yTvKB3XdA9cgz/3G31KX4IP9utv9SKZ2vNTk8UQq01RDl
j1F7tT/W8aFZmQdTVfwbB0ZS9J1uQCKVxsNiANlxx/8CsVk27kVt4NRG3c4i+neC
5tljWn1Az/GqL2yQPFcmUUQP1mT+uPhgvh5ymdSd8O1t2LaaFae9LtVXOngteKWb
RSrzidMxT5jyW8qiQauXS/aXLX73L5w46Vfi1qrvyrgzNE9Y1BlMmmAvcPxSrSTi
2EdSNaMrCXhoefANabLGjQ+sqT67rIB5qiJm7CqpqBz3uqNM3NR02N1s8xlz35Aa
jODSZ7wHuuwna7OW0Gu8yJFG3AwMTOwiyzNl/UyZ7k+isCax5zDTeOJ2hhHdP2ka
fHauKWHPThpLtLI7zdCpEkA3QFEXFacNzXMVwkA+YEBmiLCEQQ6ReGU0nJyKQqdD
Poc4CTHV2aBZrsWZighqYL0CJu3AtQ116ybR7213c80QjP/ORMGuDGu3dXVLkkro
qI4sOUTJdMtuZCiNUBelEOBfGDtferC6pxppJWeBl4SS8jfVtJ1LRsfwO0TtCeGE
zBmHcVcnE4WkyrOZElltHV4aITt9WHKThjzEY3+VFrARB4wDg+kvTIFbx3UwtuFn
sywXH32NYl8UX1ZcuzgM9hmTrpxOFAUB/P0a9UAViGJNAxGz8keKytvtSYyfMxY2
nPbqta7slSIIujZKyHn1tZjw/qSc9Xy9YLt8mPLkGD/qvSiFuygpWBgsZkLiQMlo
DKE1Ff/R/KSVEqDacwCUPFGt2Am8GeLIzYAvPmprOWql2TOxAquvrqaIFZNF64fL
Uq1HO1s2e8pWuTw2w+t8xoMfb+mxG+dgOKS1zq8XxviTH0sPfE2ahBVpv2FDPzjj
doJQEIZl1jKfyA+xj24ywU+DEBKQsBUJjxbUnBZOJ8sN3YIA2du8wIU0Vf2jIJSR
Jio81hJcpNlW9rJnA2NuNBNtTJdcW6VCTBwy2tezxabz3faOZk4KAf1vlRz0Tmhk
rpPr4OLWldCJZTDvMBl7vfsV9XF49SR4lx4X/kdmWUJOInk+ZnT+Vdb7It/5KzjO
oICOw16c0VXoT7cB8ES6Y3pOwkA04GppPHUivLN+WQUDFGyR19swY6LSzHyPF8+H
j08UGZazQWDqOntc547wPZ4jQxZShfGVxiT/3Z4ngyGsra2wff7AXP5jG8Y8BUZo
ljTnbz/oeImX8K+h4k/KoaQSZ7VTWYqkJN6vITLxHW/8zC1WRebp1fGGfmk81Yr5
uIvZB4knxYLVI6P3XGQlGJ34RmbKnEXw/oUKeTjhXFHKpMwjj2o4yGOYNRUWiHZe
MzIEUSNJyaLBSRnEUa6WsiIpRZSf4s3tnNmoa/MVtIjaWdCpT0DF+Nv4NQAbIu+p
3KWbI6veyFtLzjgQuPSZaCElo2SWbGyjGXeSDvzrKT7rah3JHf/GUZ/wvZZv/J4C
1pmJ4yti3FfObVicwY8/8JOGOBRN1Sv7C7bTgkTjL7KMAUACiL5CJDQ8dMKgU21S
fVtgJmGujFKHmmc6y9UO0bHZfY5s81fSvDknwTikkTdRurVlEjHXlJ10MMA/Xr9f
tgrwSauWBQLvuaYKaEJH8kMQvCZ2VGdrSs7G00AMoinZVJlfDi4NtbHeAUkjWe8z
iLOK6OZfNKUxvz8htankuCypTPKw5GkaYkavGGDpu6jCXFSJj33RUrQnFeqDyG9u
IYzngZ3Vmcvs8m4K3RuQUtJqHPDN5Ih63iqdv+8NpP7Rx5DuWmgn6lFJlw2t1tOZ
9kcf7JSpUL+owxclERgJf/KL57Ur/LxUu74wsLUK8C02plEtHqOGp7ESCN+tdOVp
32pYmtJHUg1HvCZAN6sW+WN+K2NzUw4Pa/1UfqcjXlbJy8lqBfqgOumfAVGjeX0g
wweaSmE7TlTgTW4oePtm5yxswVb59+MqMNOOUvute5VO4XMXIzZ5FRDxtynUOAOY
WpFpatkSYu31fOVD8g2a4/dCD2RAQgg/esnsjSLOcaFrTlXD10Ite+DWQHx2B9Ee
MRe/S2rj+Tw3Y+X588e0NJrz2d5Asmb0saka6SaG3Dt7JP4OCilg4Pf3DqICyTnT
FcFtbNsccr+Mfm5ZJUe1cnHk9VtRClLpqVm9EaVMNfxPToLDOeMxKYqPWpNjLiWH
358m71wUtrb31NfaJnL5Y8kFGspcks+frHtDGVf+T6FYa+zR9keGZtwAzOs1VO4N
P2LpPbA1JgZiLXrp1hT1AnhLTsqUWydgz9FbBbJeIiGuQ5+1Ic8ILamM06ne/5g2
8q6LkVruvcON6LVfHvaCQfiqwG53sLrWb4ZrOPBFZC12e2yuRaj398mUOy1e7Khb
6iKn7oyCmPQ+TIxhYZ/7cmZe18prsjD6RKjLN5YZQLfEnOHDDw66SJnYQXHafEA6
AUG8jlY5XQv5u6bLCYuJ9/zLFo2r9y/Jm5ROIb7ehPJn8GtGnO3ZbEVbWdfB8zls
syWuywPOBcGojnuAs/SHIn2iEPLa2E5ZqqFV+3inLC9QonY86S9rB3QHWcvJY0Ua
GuKxh3RrG+XLoAtnDp6QBZwIitcdImxTsmT04rMQhQ7nio2fa0LRIzeneyYxVQNh
jBiidrSsmqCMLgfXdRoqn9YPMrsQmoSnqKhET4wNNZJUNDJF8l+xEmNGNr9Z7K7F
grF6bAepemo5sVL3heSeaN2qtoXISsOPUEyBi64Khi0dkwlpLE8cm94DDZXtxXxf
A1JSnu+Hid8hVMRtv++7w6ESHOyfn6ubZM6k9yfbta9VPPKsHRNOyHT7YlLxjk1I
j+Zc4hC0x+0Mv6+1mgI7BvnmkU+jXG+flrMesbj4rv24IHxvXNygwsD7Zfe/wgtc
olvDkvbLnfA2zeJ+x9MkbzUsjYJgis7dlYB4eFAVWFBjEWTLhAJKpyHCprUN8UP8
o16aPJbIYNab/0JCtnTAymHVkIHVlfG5VPA+woSlNdTa+YXwhk6fliNwyT8phojR
jUFTBnpoi72SIQEgLSZB+vpKodMkNQTJJ4lR0NPFaar2wq89Cedw7Eh4qLvYC+Ug
w8y/imB1pvqg14yiO5Wm6XEgGezPWff+nWJhTWKt7uB9jWa59R2T0d5Vkke44J/6
yNthznkfRmrXRqhWhcy0kcJmkdJf9bNVvCc5JihiGjpnPXbxW+/JOoA+4gdSamVO
XIqZbiU7cuDr1oLAZwH3cBIREPuvilZ7PzY3y98kRV7Sabn8I0a9XqrtYyO2rAp5
Y5BoA+0i0irTF7ZXC42VwRW8BwkncEQ9hEKvx0HPXGvwn+76dRccU9ZANHIZiQoM
ghKvZ6DrvTAjljYpSCYih2XlhZqkV0uoN2psoVf5YNrFiGepakvcxtOp12BYfRfL
M2WZmxF55yntAQd4HNjtnjOmVj9/gdfFbhxlWZ9xJva2ZoJftQAXgboCD9Ebgw27
b0yRbVB5uYSew8oO2rg7ij7NRAtxTcVa/rbUuUIOfWlq64CZDL79+NQ+v1O1vxpc
EnreEyQKH3VLSefMGgrWaTXV6ZqSY8JbUtHAxWCycRkRkiMtF7lUGcSHSutVRbfC
pTlF76OkmLVMRQcneVMv9LhKfujpNGfY+Wc43CKcHHylM5LtajqnPNSbDQa0/JB2
Jp/0t0NlqEoBGMUsOjWaQxjZPMXwyCYW9X65PZ2eYz5GE5zByyGIJ3Sdd/WdvZCv
Vm3n5FnNXs3D12Rwxu+4C6ZTqDNcZzekp20uJ83AiaWjA9q7glnoSNmvBxw9rrFz
Mgm+h00S60VMpKdl8RezvHOhjnhCY1n7jzH8QgJu+Sb3kprASdJX/ejPUmqgJPyf
EDjFaHKSVIfOhoNHuZs8QpIxT+HnjIT9t/aI72CBliIAPZB0CGS/n8r4u7UHj6e3
iWT8LpLjwCc/0+D+mPPEq+39IDJUCG7vzX0Okn50qAmAj+paYo7SmJpAyn/dHy+Y
4MA4IjkfMREyV03SKxgyIrcsjssV/eQpGdj3CgSW/OQfEbBNGPfiyky5RZ8oZb+c
Jt44AUyo1yOE4hNNnhh7xexd6KoY+EQiFaJQwSLAW7ngaqJhZEgNyTbL4J1CnQ7d
NOs6Br84WFjaGHdSadGrcg1YcZZEYBVFf5JCLA7Gjcr1CzmZf+LjzdlORjcN0MvE
nCZN63+ui9Km/uTDViYaAUzHEZOkW+c6/6wGIV5As7cQ/oxKepDHO4GN4nwa7Xn3
uCIVaO7CHmdLWXBUqWmQL2k3SP8F1OthJX53GNNmIb/ZOSNvMW5wg5eRL1m2KlSP
Kj3hqczBixskoYZbwFGOBh9U7T9PegU2ZFfoaH5i+KXuFQpnZLwOuQApAM/iN6XZ
ZJU8sx2byHGMUmOzdb1+DSQKUi+zOdA8JP6ckmXHK6uxZxK8W0v7e4fhZnlcZSt6
PPYf0exWOtewdG0t/kQ8GLoZFZbayCGqi3FmTetxe/QNRQOc5MN51z9dV31VBUrF
i/lJG/pF8l0BFZuekmE7UBEKeeoczjFJtt8ufrB7UfmxoVpdU7vMTS8AZitHolLd
wL10Bk0pvipSrl9z54h5qBgRPlQVJxCUfH2u3ig1qEuNOcmdRrpM1yEUah0Xqx2Q
9trvYjIgVL2xEXdygLgXk41F95gJXiieFU8Cr7Ph0jaaMw4YyXXe4Fu5powrE+yq
dt9p/SR3xTY7RZPmNgCBz+kI/oNFXZ8GXCYzqPp/JWXU3Gb4wO+0U2ugGXpoxIQG
cpCvgOAHi6Jc3OrsBPXZKfYpH2KlVNILKGn9n13Eb+Jq40kc4GehusC5JAElNUlh
GFkAxYxLGPexDUOJ5q1AZD8lOov1TDmXQ0G/2fRRVMbwg4eAkZyijusD1fBDV+Q6
y8axTTLyMnkYiLPYN6rdVcmkz3GhhmWBASzMtfwwY9CHqzX26Wh0I5TbQkMb0MyZ
kbDMekSfVaL6/xtptIycd5/MnJUeWk0FKaK26GSzNiY8g81YWNjqVllg1bwAc1ll
qp7V6ZPUCjv1soPYTNXhw01tfiSmrAOtk4JPedE+xcDJ1XSsRRpEy06x5JEf5UF2
DUuNOiZX6YtbNs1CzV1V1scHhUWeDNnGU/31cXdM74O0dDChUhPzK8rETGT1gfni
t6f1z5NR9jm3gfHxEdrrEsEI0nmt4wexEj7kzb+cWkY6Lkh3nRV/W/T/kAG/R63R
42DRze4oz0s0MVoqNdIR/3K0VYzuq/yDe+7QqajbjRJvqDQ52KdTN9BGFRmefg6q
gloY8uuJ+5OKNh0VmJuJlC9PYDB6jIzPjpf90t8DXKXso4q8yyIAvEWdsf7XB8+d
3Uc7Ep8ehm41RjWu97Pw+1DFisQmwZejGktY/Dee2uKFcmhJSoQ5TWB6YEKWdFs+
BVDRPB9x/W/+yC0yOlVgdEVuZdRREjV66cZK8RFtLmAWqB/8Fy+pngnVPAsx3GM8
ny4WcHauyGuEJBzCWRGS41zuTVnIDjKWmtP1KcO5Tv5XPWTE9h1LsRsCX3g63UcM
ow7nMLyq7u6Iygn04wC3z+5WiZklub+xf1QOEDmlDWnM1eHcCYkSI7bFe8Nup+Mi
IPB0Mza4vcHGQI0gIj80JAY6C2dEgZIUEOjAPtmmoy1lJqO+B59zlTdDxY/s30W8
NSgIUAhSbZcZ0DOeAd3eQwA2jGFDd3LwNyPXejcB69o9ry0Q8yEyNagqpWQjvI8k
4jdt2fF9X88OIq3v2pJkZO5o1eoR2BiTr3THkPHxaL3ZvRs0sk4OoAqrZz1tPt8h
Muunmju+pmjSmnFPAjmhjGG6dsPDe1y9D//VfBfi1qjY7CMT8P5OkHFcX1uENrQ4
qMezSxQS6Xw6l53OofmI6rJArN440t8/oFTy3SGuc+4pPrtIuPhPYdWiQZqB9mIO
iMUFxMyemXgBet4M54oH0bVNJ7NmoD+6g3b7+YbcKbWy5gqHOj1pguHJio/m7rs4
/YXHorjNt39gkMgi2oXtetiVtaW9iUa439HhFx1QnksgRARqYYSkpSYhSjZWoIry
4h3t3+LmtaqObB6ojmcDj0vRM8UYlSXzxgfyX+zmoKhHJu5fiuhhgtENv/HfiBlh
O6CruNU0HKjD/YEq74dU/Z8a0rp2jls+5Hu6ftdPcBocpRDpxbCI2QNn7ErxbPv2
5qkb/BiR/NJRBFaObJUlXk8ucyPw1i4UzgBFWyljkwzJ6W769QcegFqwnU1gx772
Pq7OnlqD/2nUeuPRNhl6RmlAV3cnE4E/N0WbASLtbYJzdhCGq6LzXVkGQzA94ph2
cdB83qkdtlfHPqJfeG2E8VEN4a8nZBEh6fsIWh1I4kYn0xTWsT63JfGQgT0QPosU
IM93mfaABEfVktfaRoofhmfHABxjPqoyBXx2jnAsKZPHO6YHBXRjkhPCxNcxvVr/
Qo40yGOFlvv0bqh4PESBRgDyK3jUENY27zyh9nuRNNoQqJKzO9vfV40aanXPrWCj
gW9EdBmR41pUIgeTZYX5LS9ip9OlcwhpAMkpcpDpv7rUhsxGOU8mgQsabJpX/x+c
sul79PwT8v12MFH1EQ5ZyInqWAId/xniO1ByY2mjCAvoRlJy+AvDF4mO8ei36ncZ
7Uk0sFEcoNPMxxPs14vQPMwGeugTP44BSSo3XPx8x6gQZKi/IDEeW0OQcijwa03J
ESg0hhGuGdpxN3YY8x4fnfVQisB81wxYVRDRWhpsAGqBH7JsVSzGXFJrFzJZ5QfI
tcQmaMVejG8W4V4e37TZyDk6GDJAR8TVEoNkOO8dOAikLnoDs3AQ3e5Ug7B58Kj7
atKkBJ0aTq/6U/v7bKmOTORBZUKmUCjwgEwKLXvzu8r47/LROZ8sNLy0omM8KBMN
dWUbj9fxC3mnKu+iIysISu8PzJHpJ6zu9XT56IcYVdyfWWr0jMecDFwPYypYCOXk
16Wo0GUrPbgKj/9leX6WdXRXFF8yrwu69sbVfPtZcjjJPpoepMG/6tW2oxK0Ddmq
FxxiyEktmxRmtAVkK21d18vWesIn3twkV0CxI/QGoSHAaYkQjUqmqatz1YjbKWCd
atV4gqzfhih3Rv9Kb9bdT9SRQB4a0TAux87lZQPXb2eU4ojRxhbdVZRgRcoT2JWl
yvuthfGyNCq0EYHa9SH6o4odak2XpdqCWOfql+qXbsEKfc/YtbrbCCCKO8CTo/8L
WNhtBRiD4MfzsXxTSAUhOZZG3F65hOOJe5E3HtPTZCH/jbyikOiIl1NYhyB5dPdU
eT1xG7OKvwVFbIyBeGh7KcXjyP28bWvrAiIzbWznvBu7E1zgrDcNz7fjQfMMIkYH
LPu25rIsodFbjv7eQoWOkR5EZrB4bL9FmM0BXp8EW6p2mrgQzsPW62ndUmeOcOMF
TtGffCgBLfFPL5fntmpi7K8SoPkOeHW8xo26m4OELZooXJaKJXlxb1e5khGQahgk
0UW5Pcu4hH1Q9o8+D773ctggDcS9JqhMmV0iJIeLTiq+4Ka3kS/wObIjXKrg3dSj
/12v8VAvReITY8D9txTu5Q//NHaKMadzkbntyeldhObqYy1P3fZ/sI2e1g4PPbs8
u3KAGxoz7Ta5ziSQgaBPqWtbORVaX301UzXt9HIt3zuUfoEDwuGaebevAz0swZYp
CcUJOMzhnpHiGFa8iBVp8zIylGW4vPS0kmYSgrzpmh7sD+IVMDO39MPzHMm9m9TE
sZIAFRBNti0kfCVfqWprDILvOoJbjqql7dZ2DQ1nHymM0c9OU8NjwMg5LhSsm+Vx
vbZmIPRDj7oeAGb4gZa42U6JWUpW3JEAvacwUeqL9AWmFINKzhVIGAwJhTzwS9U/
9ryduEK/75H0ak4Q1XRN4YPbiBLD2+fq09inZWzMCMpx6Tgm1RWzSQvA+qmdNK2l
Z74v7pp0gIACp+gv1xEI3DfoouLpubkN2AbUQUFWK/npQjzaZSBkWZz64lcZqlRV
1hdr3RDbvlCKerIf9bDieNF1MYXvtpeW2fG9ioh4vW1TJs7XYaK7QJHCBt2SqVWg
afyI8zYmbn+S1k96agmwHN8OKB2BhwXY//nx3qcewJMW4ZbcBVfGjSA8yO+VyoUX
uC600im2ZrZ2KBLrmgkgpmhEz+WU4bMAjqrEh1VHxQAYM6ee56hgyaPEdlwPgo6F
Ce37H7cOmLpyk2LUr0fgoznaIbw3MN7L+XoTbcJxugh7ayLDWi/nfwE/GgDaAz3j
zx/DZXHDRQ+crdnPkDyxjzVx0x2WGvZPJeUCwYLa05FrXBc7DQNc9i01JpJT4nPc
05rfGgnsdw4h5StOFkl1gr9HgsVbl9T/BnwwxGTPfRJv02WbTiTejgw0633/PeiR
O3vQLIYYNPwI+ka1lamSlOv2KskGY08YdOwVq37HvdQOiY/v5TPXeRi1kdbe+Daz
MF3Hb3KsRLQr7Icl8sQCc1uR6RpOIY1YEE6GaigyqtRRk3JYv6fTphug+ZhqNb7V
7kwqqhQXPbRz3XvJKdmK5kcH7onjOCuS1pHZttJHl9Ysh90dAX4vuu2DO5Z5kOfv
nuTcKTEqCdeukD9DRPTlLKxnxwTYakIRY5VnlGeQWCrZ2Ln5MrHeV5n/39pGMZkR
+7dlm0o/vbYg9sNsZ0opmLkm5uha038LNvSlAKsMyBs7gX//f9FEgRAQcLal2PNb
SYACVOWxfNG1V8En5VgF1FkrwQqK8bGyTH8IWR6FbaQ402E0EAirybMPD48IBNyu
UmbLt+mHVwwM+puA3dfABWdgXYS//4cRWvt99aaAmLz3gYumayPcVUJblrD1+boV
Qbds5UKFBOkXQGt5JQsSqCdu1RxAJ8m9lS7SFGtOYnKTwlr7S7t+G7OPGO9iOJTo
De5fJrwvxvQk9D6yGgC+S06l4Xe25EMuDfI6qBdDakOblRBZQQ514BsLkAq4hx2f
9jxciL4I6Z+CQsh42QUQY3d0dlweQIa+D7BbWh/5hMdjq6nCwH2GadgOoCJIRIAr
RDbQyxZYFd+RI9PK6CkHG7FxXeJPmEHyNP94naXVRVOCx4fjLpJ7S5wV2UkucCvf
EsfZkCSXqCETvAz4sWFWkXWjHqSVD0l8YpC/pEs4OSSExPoRzVPt1CSPFrG0xMmK
JWR6yS+yvji/qHTy9AP4Er5r66gi/BMWMfRfXN8tcp6xGLLMGoWQ+7rHwD3H6l53
tIzjPAH54vSoqOBevHVIVGXe8IXwRgEq+eLvh6FW3FvkdUvBx+ZdwQ15rxp3OvSd
spwV/IGsMcD8Y/dz3CkwjD+q84IXaFPo+sxoB5Gqv/cHpl8RziA0gDs5kX7NrIj7
u/4zrh99MjTjHSTRHfsmo+Qh4mb+soBQ80zJ2df+EeWTJ5Nx3oTJMX84EsIxQ/r0
q123zDYPJu+J8Da/KaopgS2G51yNZbkvnK1bNMNcowxLYEmrFqZxDCahfPlIcOo8
Eml4X7aIBelBtW7UmQXqgaNSGrF5mqamD+2zeXlBcrIXIQgnLsmKbe75t/t1xERW
EoiLkg+Z18dBOE6m61wAqW9jHrMEL0AaR/sDqsbtuCxX3QFfGfhciC/XbctRcdLm
m0MKA1uI9cQgoimJgLIe+tSB+l65XOM1eTq5+ymB8TSbOVk4nHCTdeVU5lzvfIw6
PMysaRbVnrcRd2jc3xhbkN6To8TMogXZvt+/DTOExdVKEB/RI2AudaC+KPxZ3vTw
0XsTAYNQRY56x7I+wd78aL0RfryzF/F6g5W93vCEE7Rz9NfsC6HHmd1WssLcWH0W
yaDDVP2Cu6sOkAnZwd5NZ4CQcePnOeyZgGVlMHmREPkfVHa32K/Flvop2t+4to/7
SzwnKj0LB2NDCoLanAHJtfJB6C70zgs5fmtuXxiPo/Y7AZ+u6ftFFjh+Iiq0PrSI
6lw7HOrhMnrPP5NNkzQeUt9h4zdlZ2B9hziTOh7qGr9Kb8ZNv7EsmRJ+VS0oRNHd
RBXHNMnPYpfCsd58ARl86W1tc7UE7AfClU8Y9XNFReusFndnBBysqFfCyvWe70ou
35xOYzSyJA/bc1QChViVjAEBJeTcYGqfYKjBt+VY6AHTwJlz6znQF6QmysY0bHiq
zKJU8+HSMylHC5FLw/emR2q6oc9A9/eN7f29k9inNF2/GBp/8Xhe3SXmdQQ4/M1S
LrYUhrItQBzYkP5HGBpTTSYrsGGa7rF5O0HalFRdXhUOeCpjb/Oknw+UIYxogFLQ
Di0ADuzAmpvYGwXIKspIHYCbsUMmNlCm8ShwlCgf0IHp8f+W4PtY/mZAmMR/ljp1
JpykBfozDI2e0uWvYRdsvGiqOt+NoaM+Vb7CzPvNuqHrpE9bXP230f/zqD+tUcR7
771D9Nc56pNt31yg10N1DdKwS/5Q2AAwzCVzNqkJSnb35aSKefvxJzHu+Ku8o8o0
7vg0+hNq/kRXPMj63+YChQajkBr99QBR1eas1dI9z+XXEIg7M9oDrjNuxtsgmvog
VrzN12Or+q5ROpuZSWbfJvLdhtXJhpnZjXLXnqCB3h17opYByTwSWZysTNfdZ95P
WzaUtAP9fQvxUsBl5yKXlimIdWBJt+cGLuMsJRVmx8MpHNwv3aw8Dvuym3Z5CASl
NzvkHhHeDWq0OH+Kp5A0olrgL5I4SY9neYAyHM0R7fAKj6bDqXH1IingcVazgUwF
yzhfwEnBERD2X0jQTIBUtQdJlfwTUbqemj4OnJjfpuuysRq9ftolw+sDanROF+8n
/sEvowL8hXBhy3SBjbKBIOw6bfxiHw9i7Ly8WS8J2/ooNX76Rl8DT+12PUFre6HJ
5bfMOdFNiiwJYpk9zVyGNN9hO5r4RyDE7KxlB4vrv0eVouKWuPALormhbmKV6IzH
hR31V6M3SmJ88Asz+lqFA6rkcEPMJHk6lPp8tVZE0BT0AUV4ryOV57YpOQ9lJ3NA
N82482rGA1Nb+dvdaKgb2APJK73Kmb4GFSLUcIUYtI1HevSxx6kvXnYI9eZgkjuX
CqA8pvVmpn2REvToMSx1pyoxlIcvSZlMKkXTYBGgfXAVgnY09afvThLPEs9B0MBu
wMthQxJauOvR1xlT5kCjJMUuOPxQifzDfcNghfW10x4FQkiXciACXzPP+5Uo2dti
Z35vwXePdXvFbNqkyT7BQ0r1tAQdlMnnxGk78+ufbW+8dvN4jqX03DZIGbrWq1mo
fwwYiY0v+kZQ+DVz1L5WmASN5Vh12nQa8DURRG4Q54rhYcqlRckkNOXgp25X3V1N
EQKgtcIONVkAakjYBcg6bZWfEYUMNLGv2gv5FPtKS2enHBSbF86N5dTyEJfeZIj3
031W+jPu8qG4dsuvn+lu8pYmuXooieM2J3ovlNre2PzaOkA2cQKrhgY252Guyf5K
F3GXvpJO0cBzQy0BSSBC8ydYSjPsgwLIPyM6LjiF+Kx34v9CHbadtCnm1hRFUnul
UwFOiuFlsCp2M/CZpN4aZ9yb7TyYDNCi17ddl1S+UiQriPSXPBecagTsbOX2d+VK
JP45iRXwfIJo1l047GgpzWyNbBP6T4Tk2yhVwf1QoPud4VRMFPPyB9LhgIitQbeY
MwUYTAtzEdcwCeKRMZq4Ic8HZRHq3Kodez9r3/r9rJgeo9IfagEn7AS5HDHweS4e
LGSwI1AyljnrLzRhTf26VLq7PiLL4THhTg6XyFr57iu8unsJYxMYKYGoQdykM42H
BRu+aIEXe3++D0PYaCJ3fpRh0AIIMMMjGJR25qiMIOr5i0Zoe/S8x6N1gC8pXNNz
eS2Wc7Uo8CkAvWW90uGWnetq24ySDZrhgx0B9q3iqQhlIPE6GeexLts4+HPYhT57
fOZEcCsWxQDaIQTWLK1Q8OA6dJsBpBFsSGUWhLFfdIqKJhYTlbeXBjQQhA60PjtJ
ieuZmpGFcr+hKcN+qn0tKJ1QmoWwzYpKMmUg7Zzjv3kAP5KwCsi/ZxazK6gaGpVV
erB8Nb8rT+Icu072C+QjTqf4wDUNTaDig18QN+symEZ5TWBc34UkcxllQ3c6Nr/y
DI4fKe8ZKijghi6wA4sKTYUder/WQu/CrM5NKs/e9GphWRGEQCwU7dGI+/cNyNyI
3MiT/Cwm1SOPeBqwMfPVlG58jx74P9g8v/j0EDzhKmgE4r2COBm/fUfa/Q76RDxc
CdMRZFHII7Y51mjo0t20CkUYm0ms0hJ6W+KB5TOyvoTPzK39ENwUnWelgCc/c6yx
reMmBHjQbTGcWFdC8Hh0vWm9BlJET4O3UuO9ebbMu9Z2Q1AprJ/AN+TwzHCS9EsS
LscAUzfNiy80C08uNoJyZTXZGeepkNVkjL/NTVdKVw+FEIpPExSBznkRdhdmFDjT
uIZUA/w2jtjZjtCnFPFSi/AwnT5Ug016WbM8Kt8GP9o/kxrd4D+brvz46jT/S3ye
neIwQ7q+aaRJ+6FhT1an7k8ag7JeBLmeZz0mr+qAAOHx0pWqNZu6pBZoxdq+F3ZJ
497s4l1i6NDg19vBTP1jcNdv/pYHrDYrWTHmZGmHi2YL9puT5wdpTp57sTTyOm20
+JGuKCWy+NW2Cyj5QG3k32rUvkVM4+K99Xv96rEOg65YJkMdGkfc9z7H8TIrjy7T
IxlVvxceu/SWY+flS34EJoeo0+cYl208KoSVBLFzhdL3FmC/UZRMmyAQjqBHdZTV
VqetNLIeE4LFYQVicSlvjVBMCFShZYp/vMMR9t3t7Ckrl/Nsh+f9ufgf/4P9oXT7
Ok3qmD8kRdnf5549PJMwP5BRzxnjyk6FgF+y5SKi9qjMUJe5Etiyl9gwvvv6i7Sp
YrOXS9vYJCRDhqb6vEnV4mctdDOo1FsT4GvBcOHlkesma81dqwc3VQ+BUmIJCZQ2
XZ63xp4ScMzI6ACW3H3V8+DwMKegTj6gfaJ7nsvllj2Wby9UZ7HKG36kbZDOJUaU
WZnB8ddcL15Odm12fiBBQO+1nanfdB65Agxbtug3Kl+4nk8Sd+r+D5Sx42nAIlK2
D8CSjfw/rTDpV/d4d5R1VOv9d1PaO1hi+3R7vITSL/a33JTPR8vtb+8oSZzFGFSY
Udzaa6beqM/RQE4WvalP+co3UOAHoNSd5yfKQwjSefdcQ4lp2L0tN/9rWVhLno8J
ad9GgdD9x65278qDFxVa2EWLvxevVtH5Ar1YpGK8pyOsPwMkM+IT8Usa+c/dETs1
u50axlbUJnaSG/E5R1hPx/RBXCGDkVeQjhGguOQJE5VdklqOI20vVvvjIvMzqrkp
xiHw8QRBL4HT0RFFFzQmzZZcNqcaGw0SzN6IvmIsNfV6TZzgQMw/tSnM/bs9zwRt
3owHpSmmVW2cwyBN8sUrkaOTEVsnwCqWpGKJJqH6IpL0ii21GwULsz94DpYQoZXv
42+OQ+xzjyYQHicc4+C2NWpxF+/YzM9A9P5ahPoDOBKPa9EMFwGsfkid1gne2vqG
Bz2A0JCnUu1pJK9BQ+i+W1WV/ToT2CFJDtk8oulnqrkiyWgqp//NmdTtIaQP9LHn
XVALJhGnT/NxqBTznjEF8zSgACkLxDXjmd3jNwwp2wnE/sUeF94+8sL+hDXK33rw
4hGW4J/aCHu/dQdHRj6tDuc0/WtnxIFKxxETkopxooIfy6LHNGzgCj5VYGcaV22k
1B82xSXbdbPmxUR/H6UJL9F9yweSzm/BN7Y5ig1KTDt7WEo0KqPGS/j1MTRgH1w+
XGRbC5bz0aB66kBHCsjNOKNp49V2gg+Wf9GhuAiBCpJ9Z6Z1opngVn8jfpqr3xnP
yMPGoLXbll8Qca7qLlKDg5nVDFXN8pge9tYQzbabzeg9WlwOVYrfgqZi+wHYZAra
BFBFVyUHA/xvC79DlmxkG88ivOokSP9rf1zMMcBJS8B1fiKnHm9VYrBhXbCL4M4T
SXCdV/tgv+23j34rhkFae2BkILHx+4FRfvRAwodwA1N0l7FHr6N2qclYVKoCexPD
ajEV8c2Kd92qsir+7ylJcakLRzF6paxNXSgrM7vJkFjUatcSMeerTTgaPJW6yNd8
2VWeJ7FlZNKPR6Hu68Emhc5VMi/rA8OLVp7oJu2vlZeDw0W7FGabRuDlkvnboD2L
flhUIPZWzsFx5k3U1PyhwDXdqgSQvVrKtkyuhlKzMVscgA9X1GkY4JX+l18cGWRJ
vDV3yEd4ZGSzP2dwTwddbEybH4amXnSoriRSYQDbAA+BNsGsiIUerByNdLX3fT3H
EyZIGiVeYdSZpOugDOY1HJ45fEOmVD+/o17kgOgntpTGrKin0+YVgmDrC1exnJlX
WD2c7dNHDBu8JWK5fMvCzsb1v7eBBoBPPrFiV191wvvZcggPk/uCSdyitFOZtb2I
S0nrcGbPGTDfcNzS3funnpxSI0dC3gOBSejMynvq4TlFK/K3eZivf2hQLqYb3HpQ
HPj+pFwDcAWyNeqZnzxjCs2bFuSYIT5koeUEcT/1X1k2oG5+PXeq8nRZxkXtohDP
cknX9SxPYdi1MIzXpf1UeyIyyR6A9fstSskQZyLH2dimkI1eM8q8a7FVMtKCRMJM
F71hWO0XjOSWFxMLr4hEaNsqXhLm8Ucuz9vlpti/qh6CQqeJ5Xf+S/IB7ic+EDyG
BLeH5a1pNydusCxHOBEaHzFTFgGuBkweAA3BCsO/chJOchgeeMU5Rnfxe60ntOQo
ZI5bf5OAiTezHdpSJBjUEChwbozGqrg8yChsJnVmDcY9vIzY1Um+Y2Rj6NM5Rz3Y
J7lUebhRRhvkgXsteEPQcp4OKL9VKttrQB3q6Tc65K42NseFh4JA7oUwvPw62Q/P
sypnrHN0e0GK/K9HQQ5J/RYlGxYtuJxJWRbyrnG/R4x9kUB1WCComkXXyshCOTj2
RlGqjsgV1d5+df3eywY4v0dTfxos/oruaTrXIcFVA8/i/mmyyoXtE3klfJbLcPaJ
9RwJiM8Ch0HWnD7JAFFctAL1FnoMFJz7nIqbBeP0M23LhUuiPlSEkrRqOAkQSrMV
1In6Uhxjy1ZPoLlVmXtHNnDClHHzPiV/z1tjrW9pSgXOWvRjs+ltce1Lz4bytGZP
xHSEtBSwhH/TD9Vjm+OsOMKu498n/ox+0oUNrhoGFelDmogZDH4mKuiqL0ORYJ3n
CGDVc3XHwk1LIxx/+6jKEf4gpEawMjy+FO7FYIctqQNdG89cgpj82yNo6K91zir7
8ZAr97m7+3McTB63jN7R/WFYSsfZ4qFRme650Ts2rdfHU69b8e+4sb+P83/F2TV8
MwWO+GqR2/fsDk870WoHlbxw8wgWtuvUlM27iGfM34FhhyGZW0hCBkxgiVzJU3at
OuDwugp9q8DuGIaaVvU2Eeth68Wg+iv2x9kI5lMPz5hFp4xF7WdVPf6GPHC7Co6V
7OgYRzJX0LwzjQ2sc2C3Td5LMMiLnTdf0WrH8f5/WaD4epkSC+RTZ4jC1UpM2m3Q
+eqTaRi+uNEFKFeEhXOrHuOg9XpGHatYD5apWG6KuXzyRBjeZePmvkMz2PGmD0io
sSGc70lKSrVvbi8snRMwKzIRDceY9fEo7hx+8vqKp7u7n+YWL3v/bzEj5NUTWDMB
Z4Wf8n+PKK0o/ZPNTf7yUi/mfJPRnpOt6L5gz0ramOnW+0hAKZTKuQFtw5g0oN73
sh9Z5WEOPXSg9VWp32de+1e0XCY4MKnefDJQpQz8WhTaerfXLhjL9/42nMb6lggz
ILfORK2pB9uhao4iGMQTHH23NAReybcC1hAJoZhUXEc5XcQ/NV4s1VI31aaKllfF
LjjabgEyDedKm2mrwsTgifE1NGrijWPxfe3lmOkAeCzBQhwvKcXtm60wReJjbDRM
g+3/P76I4pNljxAOTtwmluQgBk+VdDruyrRs5fshbFYjxQ+qVgXJWEJI3SuuzZ4f
rpFghABYQ4WHe4NU3HpNiDYGDNqWFmGWMbLfsji3fxG71z2gBKgpIpfrVCvk12oh
SK7J8lqjdllCDsv5SSHq5Aoy2N0f1BCOJC7QZ7hhw7ACxinNTekW0zYf2f5ebZz2
bN5dK5oZfW8h3/iz/1rGP/kO561IFWZcNT+pqNDldsmk1G0COY+3ElnsG/V43Jxi
vxQ0xPlq9IYgsxU+PWLXkbJzRlePWhOSCbZinqMFibMQ3x0in2wv+EvJbRdIwj8K
dGIf+E/qNWzxjR38Q5zSME3hV32i2anuLP840tsH5+Xg2w+dbCrmxOuCETkdxN+i
YwtJhMClleyhy1SjiWFEyFPin+cklFdrNN/yaROEsbZ1p7dGAZ+NpSnsdjAYb5by
/fLb0idjiK2T0XMfXFtKCfu3esQJyXaM4jLK5TNuITw1GdOLuNTKFpazcsZ5oT+k
AXx/xIvgs+XSxgl28IvHYdSCqm7fntuLJ9Ooiv8sG3fIZpEvLS1avrCSNCk0IlBu
5KtMRa1kX1QtQxEzloh36t99uNt+AljdvEcz0d5RD22N8OxspuTGKYiDvZkotc7+
ISBO7fkJPMQvZ/wn1GaBJfl8YBr2JijXiSsl+ERoQQKC1/qbJLQV/Qn5qnvm+BgD
gX/4avbtzTUctaIPqBQx3c3iU5AmY4IZWhtZcT4YhQ5ANf5Yll3WYClgP5jqVsaT
XatKroC1icxD/2XS6hq9gtw12EknhgM/cQdQqq+HEzD0Q046IKx4xYR/ori8Fp6w
FbCffdKUFX2QLJMbGoxZZUtK0/g9jEC3zlYQ9ePJ3bakxX9elNY3y6murov7MEJw
2E7+bip5DgEOUh3V+E3cDxBc6USWWED/PhP1aSuZ73ynmVBIAH5QRcaI3tnpQ7ew
FHH3uhPhz9wjIe1gvIQWxsgUffjtIcog+cSEVhYkab8dR4Q9epkboXmEB6hxiraS
lHonk8ghElxBE4yy9nk8sAs2MF2smM9SaP0rc/TAf6FLXt9m3+llvJCdm1/O2S3S
FqbIEuvx9t+F+nLLBgZbKn8X6uCoJ1PuGO6dph6dLWqdaPLYmrBpznte9oOvhWdE
Ee54xaxfD5W5yp58ah0ZERzTrDjVZ9vDewgjc3zQNvCe0FEKlxvTA6xxZ9tctQoR
tp6iWp1debq/6vLsrGOr9CkNEKOgPj6LgycIX5ZsMvNmvUYg5ge/45pdqhA665mX
pwmIUq8NgtTo55SomH7KcOxohROqWkvbjBWAB81/CNMTgjyHVUzdzYliNiLNpYFz
3v7xglsYTCliqMSGkMMvnRPw/GDl3HUhhsBz5AwojfXvFchmgsCRCf/r4tWiy2+5
nEDkjMPEC7FcN0Vr5jrhENknAVcGlzlTxT6d6qvxh/FpmylPeO0W4G+VJy+eHbiM
lWoa7Ap7eGHBtT7xsiKxKvuDtwcLlrpYN5YPwiqtYpdtzEWv8DOncNqaV68Zt1fR
Tl3ThjDGY0BCu7YtPajSnmh4MGYdnd05Vm0Tv6RiDm3zZSSUQbqTSS1HQDymLzNW
Pjqy65vRHaSaGlH0oV0Nkgr69n7pcmEGRe4noI3a+2/9e280ac2yWfU74kGknUWL
790y1pr4uuaOwi4xX/ddLqGOUTA7UtXUqn2R9b4LE1AcFreuV9yWxlML6lrahbPP
E2u6lEST5Ga9FbcEpcuUwIykscINvXg7sHnVuoD6Lf7qh00N+c6PYr2SYvBQQIw8
7/F/P4O18RGYSU2tLVlMv0aiczKpecAqfonJczFc+AtLyZButqpPolKUW5/Ig4Ov
reD6Oq2NA51Bew7LfcwU5uoIw6838gwSwb7ZZdNsaSrWAPq8TSwWlLfGavy0LzE2
d52VUwtPatrpCRu5KToosVBwipIBZWvmj97C1lbAJqdTdk7K4b0XbtFADu25Ji2Z
tdte4Z5UZIxIcHul5bRnGyiQ7clrv6jS9GRJ+B/BrUn4eQqBLxsXhsJjvYCLbWJL
PLTwB9DXiRwXZQso45oUk87SKZ70/BZXQ9aEt/c/k889XB4ZWUiw/ZBflsGCSvHp
qf4ZuXmF/+eJz9/p8w2u+SGkzAf4YdQ/0GAcPld1Ai18HAuha/HKsG0yjIoXqTok
9054asjBklNQ+V/+FB0l839mo1m6WylOu5EAhXLnbCAZftPeEDMEiov/EbloZYa9
c9QOV89vBmdoLydOIap1OkA5sPIORtkcVpZvspH0fSm2DEBL/U+d3O2P3qsyQ2Kg
7aewQc7F1R6ZWCr50mTyMAY2mmoEs5RP1g5g3LERR3Jm4ugu/Vp+0oeEsUDAa5b8
WQRbI81e4gtHAhnQbI3gN8FX9awAD0nVF98piYAkGxUjgyyKX9BpykCxGb0CYotp
eoZSmyP/yVivSTN6Yo3n+7ujVbTfmuPI24Q+Rj99Ws8klb0Xyd29YGbGliSOGn+S
qKxtcrrT8DQ30UpvjuAOeLR9hgC/sj/d9eSigsuvcFxnxLOArxVnNIzezRVqO0lI
HgU9x8fBLqePAstkdDThR92pIhTdxHXzklg/hT6HClPMLAiyQRHn0E1CgF2i9PAS
fGxuhL0jWMXAXneqbgM0THdt5s8CRPcxYqyhkfLBbtC4c4qwMApLWfQ6SwD/rSoD
T3sxu8ZysSCz8DD4fSY0W7rYP9g1PrMcXmyfnU1bWGEmGLyYe6mdBASUrYW8+MNG
3cBUWa1KaaQdNjTnpBsbxBdpy0RvK7SZJpqGZhYDJgeCir7uhFdd4uy+qKzpcTqE
6YB4LdHkgFUEQoDk9zDpRbFI6+hDZbQSMb6/0AQZrfPXPnFE4y1cHSRZIgkzapQ0
VZgqiXVxaZ5/xFlc86SPKuuZ2AsUocs71QhtFsUeZZRrzYJtLruun67cmDX1hzNk
VHTANZ5wWHUY3hjhQm7ql6kybOtVUh6vk6sJweBU6L2Zr79U9xXcjCgY+D0MYjLg
OE0mV2NRqJkNgDbJZN0M/i5obDGVXUizE6YkNWj8xNGW8s1Aw8WYqgVep9NU+kcn
k9W5iqcgYVzSJEszb+XEZMmIU/XWfnRDzFShC63FxZU4Pn5d8Rw0GTZDwfsCMSrA
kGuGRvm5R7zXp0hLpG1aElydBDoT3sQIrB7aKDGjTl3LHPmDk0mu+xanHKX0sTNW
cKUkmkAFuLb5HUrAT8ltiqldUDD/hDCP6/oHY0YKKYafT6Pk8J49s0rTyd5ercY7
tMzcZ8YbQPLYQljEibG7sWNKNL9jcQKByoFspfTFZY33KjUgGvBp8JH9Ff9X14f5
bt+4QQ1Ll9iwwbQ4Ox+/1F9KRRWLnTjNS1FMzhpzU/qRfNwucIEvSKtA2phrNWXL
ApxmrRZhK0ur7Gk0EdOZKYX9lH4fhHUYBP9osOqvEz6o3kiIlI4p6g5J8aRWUMvr
MBezKnACiAcHqAebpjEb9eRC4SEVv5yqg456qG+pRdcb29H2H/U3ObO6nvHu5Svd
RIaoyyFxrXKJxU62x7lFkYzQJFCbAcAvm1w298n/5Pf7cvsal1QEs1Ag9n9pC+n/
ZtclQG1WCPbVO2HnHcurAwC5YbOYZj2It5i0lAUqxim4pziK87oZ+k8o/ISWDKBf
u/bMQdPqZbu3OP38F8gM4RjnZWAlnmz15KdLwjjn3o9IXqLUzQVA/uQ8KJyL0uin
bQK30LTnp3dzMaEgwlcujLcYAcEfk5Zwj7Dz6VBTr/xdGMIuX6kQqglmiHe3jCQ9
A837cPqNh1Tn0fvPgf4AP2dQc1FINChmTzuYCgwQd37JrRpdt6bfWW9RaP10sGol
RPIIJp3prOX9rDfhFCgMD3AR0a9lqI8C0rtxejmN0AYK2ml0qEBf/8jKwCOR7Xu1
W8LH4p7dT50XxHHxR7iv3+/DKc225g9d8CxV9Tk2yvPf09Lbw6cvjYT+M0pdNDpe
WwfaJ8vKbtMOiMPsV/YYJ5Fprw+JQwLRhEq3+Yr5DV3P7uUQFefcX5gkKHRMHvBU
09WmfFn8b/aYiXeaPGMZEdhj51p8JD14le9SUMuhMnlusSiJiVKocub6hINIAS9v
MofDJUbtlcArhHsaBMn2TvtpqkYbPDWncLHnP/KfSfaz5m8mnq/6pfsFEXtsNJa+
CypxZKhd3mHhCS/QSV5KtAIVCifSKyKUoxv0M8QWaqypjghO6I2GQ6eLraZAgj8f
i8SGWb9D8NV0UQ2qwuUiY8Ub4iAQ77WvCURFlG/RcAmit9nW9HjAmR22Uf2lFLse
dX0lVqZDhrjQGhc55qRqgt54GDT4XjMrGTdUuOw9Xqo/gIPVJsgXHE6KQA38OiIv
uuAG7eSxFQo/yrwVhcNeGlQ46TdtpcvGpn5DYJtWgtl4brLmOATYUTUueGxeHe34
5k/XYSbDxrUwa29nJJWVpSivyF+4fDGxOkf/nN85eGERlUY8N5Xl/jc5/WeP4hqv
X6x407fKKdwZsR9LA2TayTe/Oxa+JkoNjVerHGaeRQddIP11iJyM/ScFFQT9MODP
/bvF1oLSoGh2Nbf9CuVgb0xOg4bpaBV5hT1Oqi1aOr5vfOvGluUsgT9LiRsYp6yt
799+sHgO2B+6rYPaxqkJHY181TaZBs88onGJR6RURA7mPFOYUVmr5ZA0AjtxJwWe
zSi8MrMQqsAWsjDDUoZvgCPSiAD4KcAX3D8mA/kx1B29kQZ7yOfzTw51TgVc2Rou
rh/pd8z8txuu2jUQyCGx7/DWABuQ3BVjo7C10rGVXRxwiAiDxrSPxxRYaBXJp5Xk
G3aIZTWoO7B4KOH1uKTbYTV9IdjHq8GNCdddQZ+JIJ3uP/VWpB5/GYog8HrNBMgQ
fudleHxpyIvXsGYIv5Ne93Hzqc7PrQ9rU1mD8ysdgACqnf7QRmHNPb2tN4eueH/P
Pt/wZHylHEmJLJ4oDYvFDtBmheIwHMNspmWcfHOkeybDRWRMgKNw+1XKFDW4LPB5
Uhtf1SAtQC++mp0memSbTF57xm6QijyfOYi14eN+DV7gCEpCvMRRMVjZyF+7sGV9
7vfrJnk8eArFkQpdKQ/0PlsU38BE3AK9K9ag4ji3OBvszPTb9Qvew/4LrcTVJEq2
mbRSlrPcgWxmqOpb6IxQXJNXHJq6UXn0BUkcJcc0rPRzsgG7Mnw5qORPXgTOCC3b
Ex50hO4t10MmL3dqKOVhOlW8Zz88eqnndCe+TUhaPlcN9FahG+42O/qREZBfpYkD
i/m59yuXnQqcFyMOsqPQnnZ9S4S04bxoHhlCTiEtOXFuaVbjKuCxo0Oy9CEmM4aW
ly4iwp95jPoiIcGHvngEw3j7jiD6ptAMX3Dl1m8VFKyeeilSKb1U6MVV3sJSmbfD
DG2YFvu6tMJ51fOo7Z+SszeHvpih+U0IiHnfprpyDFTyWd9gWtdp01zODwwuQHab
6dENXW7OplSkkwKyj5r7vwT2hIKv6aczJv8GpSHY6dvtRk7+20n1bedh7FhISvMk
IKGtv/yxtdzjVVz2oMzRzD6ysC5LvaQS0gOhMxlwmrNlOEMzALKs5YDhS8jlD3C/
TEKymxKSRdxoEMAPrzcDbsjtJyLQr6Kn+XYBe9lHiBGI1SJzwemKRzXEYhoQ93Xj
42wuATshbp+lGjlg+q/MMk1n9UaOuHTxVmlrjzUKC/CYNHsmgX0g9UVdGvqSah05
7/s16Fp1gbGaJbrNkphyKAtie0gcfjhrWsHE7vCr1Tz1hBJaRo7nJZcBY/jq6Hsb
zGNC/iLlh59EWjSSJ30SkuYltJwQIAF8qNOECHQBTPcwrJL67UW7kS31RfoVGMf1
fklvyHg1pxpF5BAjFsvCt5A+h8bTxXN1FZOYsX6/j7QE1n/UiEIoyeR7oKO7MScJ
HLcfhT9oBIT2vPFxX52S76kkXzmD8GVlptrpnnX7VBuo3vVCKAYT9/O/RggOG/+U
0KumzAgr+qabqZnny8pz7QPAckfdRhvb2HZ+uLpMAr8FshRqBAh97H5j7sZptslr
Uxaaf8F6nCWc2b+VCZGH4gocJg+STtmHyYIj3HZetCVdT7vHuse8Qi4b4yxCVcT+
BTfYSvVzj/u/SG5dcKm3+nyzPRNOHKxTNRMyEoTSFhKz0CiHe8FfPSHp5LDajrgj
HcMzqneCZ6Syiy5iR37CXNBBBKxG1U8xNEpjPTChptXNmCHonM8wFwpd3EF61b0b
Y6s9bbhJ2YLQ7Wb6+u1MVF6dTKAc+enhA4MVKCT0uZJe0idmAsqVK/1o+2zPtnQn
gIHjKA1425BOU/8mTQ2rMwO4P0TpPPbPz7aDh+pwV3W+PRpwt8pRsf9XKE5OYRhq
QOJ4e+ODlxlX0Ol6i02lzaDacaU5O/z5NkYpFDWfLddfGG1hML0EXamVNhdJjxH2
QkS1Z7KOx9kSulwMh1SE6b492rTD/LC91JOu6OoNw5GWILfTrTFRZLyGiWiib7FX
7IK1ZWHGzqwBh2bUCPY8wNdhfbmsV8Uk3TXetnb4+jEWXBjz2yt9WoF0iBCGNkK3
KXADhJFaC13Z3e4nM7RG7daEBcMZcg0lbvfWaKEb01IXtnXhJYFuYBxkSt1gSUlD
obGowTrtW+eaqDbRPh10wUI61GdWNT1Uk51iNZNXa/NaYyLCjr+AG3g/l1lkoWGG
71wTVYEoUPdhsP8G4RjlmLf17YkUjlML2lwnyGARJK/0FCB0yR4GZT7UxFFEijlO
KGRkWRkYXTrkuo9N0pwOswmvTDlwoSbFHGHdRfk3ALbG689OAdCMuM8lMOPS2KxX
W+HiM3d5V/wj3zKzeVk1d6gFzHY2FbQXFgMdnKMu0ddiorVqgzEWc2WLlt4/FZgx
6CAt3mOm/abmgdG3+Low3fuHXR9fNLSq+xetCqAkmk2K/qGnaJKb68rHPS2KUgp6
g8Ec03uURmNL0zistdFwnKT+H5pgnE29bWASS/n9BKwTY6yzLxNYHjBC7qv3SVcP
rbNS50oyeLwsow+SeqWBcOyachhC9kneD2p9MRHeNjTmVscGeXdh9w/AwC9C/O5N
iOZUfRoL1Y5kqIr5fOg8gxaMojngqPYqS3KZehyeEASDleECEV2reWVRs6Sv+s6y
Dpc/8WvPMHTRmsdITgWdqwcwZ4zU/pl4CD4STpqISaplh9P9ylTaKhbAikcBBeEj
FeBpd0LdcybXWQgO0xCOOjlm6c+MgAzoKvUaq98zZRej0U9sldx7h6/l/Xe+qZmi
46+qpwqgKHFY0ji9meYiDDhQmnICQYssMG+QVtAoeHlnrH69KsW9dx/6xVjrBLLA
mzgwFyPDrJvmTdO8/8hI0Garsxvtdukmrky96ABxr8+aEKR+8zrDllL3/Z0XSpIo
12CwcvHpUpzgvlnonB2w3Xsl68ZEOTCyx00JO8I/wyvLdFOjIZenFSq4V8rbPkNb
qszYrOfkBuNGG55QMHjxFQVKQdeWFBsgdLl/jvcxzO4h7d1kYgjDB2YG2dJ/0gok
BbbzGglvq5R/jnbezNPzCkHcNlBvM2jlKwSzPBbdhu0+W5b3uNs4kv+p3P7CZwmO
nZKP2Y7AUzV7XQI9d5hTQFIyPFqIiPJoGoQkK9s6GnlgAT2lLUPTY+vspf2r1gAF
IJEu4NuPbTXBNqLqCqy58rKUfHK+BaqqE8Vygw43yE1SzXtbaxGyHdeu0sP7TUXv
sxbnmuv29+4qtsk06J9Gd2m/Ly/k1JUjsgBXbQF/2jvldwdpzuXp3Z6WBnV4d6EA
hxE400UlIoRD0MiLUr8/3ODnHqtH833EaCoyIQiblCJvg5ePDucHx9Ezq0nHYgad
RdH2a8td49QtHRw4Hm4PSlr3CqmlA2ogrlbQED1LoAofvhGSrmQSSsIF7+Enwnof
nfBpBcDZOYqYLCBsTPZJGHqKqTyJffMd7FEshaJu/aYhD8ZSSyzWLasC08BPYP+U
1wJcNjoTDi19/6OlJD2tqAWtQm9jNoM2kQAVRqRZfuOFj5w28k6K+JNfaX8x3UAc
bt/Eywi26nVUX/Nb31lUgrtRnrgLNMiuFBscBf4v3R5FFw7XZdJezovO4lfbVviV
YgIflL0KLDZZ1StGfYxpWR42ETWfcTHYEUsJsT8ulcWk48Py5AAySSHOPgkDeoLb
pQX4+3HTHM4VMzhwIX9ue4rHB952Yit3iGEd87RLwM5U6Azf+MPc5YzwtL5F1gKd
Wo1upVvZZ05rXFyFzosKY6m0l3y3C0H05o63m2bmiy+tDTSjYVT2fbYsrt8+N3KG
me9pVr2EeDEdVO9tu2fazgK21x15h8GywVwROZvUPrNHa9A5PA23boD7ANOJpr33
rf/XnFgNZsZntwRf5LO4x77sxIypN2OYrpOmavGWM1OSCR6siqYXX7oLtyg9+rfd
mbkhX4sg80LG4h+331GOGjQqu2tXv4mfOXSVU+CQrH/LVVBNwGErh2Y6yKeXy7bX
K4q4o+IdCN4Ceem6usUhOFq+XDcY14v83fzVPmmS8AWl4GFHCoNH0po96YAR8KFr
ky9BlpZkl6PH5976YewtGkj4bzKoqYWGNv89vWUO70beyz84UCizSHBKx/DL1+Hg
B5/WOoXDgqfi/tkE6mKiCfxQHYJ4U/wIUYe+/UMQiG2Sj/tumuRbvtmEW831D7Y4
5N21YCq/sxU26KJh1mqmWU99zqRz4ut70VHX2DdeEyoJ9grE2Uce2WArHAYjaVM8
GQUa2s+TxBVFV+2P3dh6HYEl/cVRkKq+aGAzIA2J/vmdwGFcmwdRhl+e+6oQvSGv
m4040i9VlI3mr7vSrWs9oLqHr6rt6bjN3BZnpjY4NUi2s5VEoTtm2zgDK7PtzYD2
YS+jpUPnFb6O2vW3XNsk/P2MyjtZpk55jJsjjPIfeqtbaqatjotMeHBq/XOdhU1+
7FXpt+9nsL8lEwm7eI36IQB6Wap0gzzpvZzqxe7vWBeE/Od4alDFqfGANJxyIkYN
qD8GqHK5svDbVq93iqzLPKWMuDz7RxMvTYs6hdtI17OmIyQjohQMshSkDk/33OIv
6f30xZhhl6o77Dr4BN7azJ+dJ1/sqsQ0jPKOrAA+QRzNGvjwSAzJPpkIEZZaQs4I
K+PfxiXZL60gFlWS+7ltsvPcHdh7vaZERgvrSN5l9hr8zoyRtAq5WUv0E+q8IWBj
mmNCFWftqm8QGWmU1G5wCsiqWFrhFYTaIPP1wLhpMdqLhk6k4FUZh5RXYSFPkd7z
enVWb9YD6ujcRM175eIqUSbVkP7VGgfzyOVrlRti3En156LUYsR4QJkZKxXPg0jW
X+pdyWCY2nFJzuNcj9q9NfX+WH968zvE8rkvnK9ip8IbAEhCvxD5WQA8b+z4AUIc
iOdU+aNiCZiYwi4ZOsGK0m+VCfvtrMEvrNWIOV1I1XIAMUEHYlpuRv3MSlvMy8S+
zRIFVZqiHJRlAC4JtGR8KSNMQDxvuUx0/X2ciLHfFVm25/wQD1+E1mZRlVDXwCil
G1btIN7pyy5yvOa+ojzgNAZt0bJTLx0nspL5NKBYFUUeHyxvpGD2Sw17J0djRjB8
HHIWRmp8aQYVUu/sfAqdEkLxN9vV7/3vzDO1++DdHBp7chWtb7Ec4AkmM5R0phkX
6v8rZyjGM7F9XArUmSDcF/EeBBn/WprDIGp/dnC6752IldiMQZY06jd8LlLZFqdR
GpjvMU5JirIDgkwkyMAYcc/1e6dlZGyUwlLBcAq8Qo1EmrNxiSKmOu43G7NqlUXr
D4Wf1WT+DTSHOPGu+4M0+VmkK1Hc4OzBpSbkqyz6G7ZDNPDYJ1JwC6mLUgTbJtJd
fSccirQOsd78U3h1yacKDqY6nEZYSrCPvWwUkcqSd0mESZJvTf/2PC9dbBlIFXnp
dyziMPkdQoaMi9JnxVUhOk/2ISgLF9QOp8Dimzuk/d9hRH1oZJQmZrPrg2G959bn
fvux5Xvc9N5hfCXYY8uN0JFrkGyT/90zFlq7Z35HBfsMibL+lgOdNZ3hpQUSWXo2
ybuBOuY2dYTLM+grXI3tXnlVvE4fpNKScEkhdCOsjSlRqhrGNcjRduarLI0wNV7/
JGP++cJfF5b3aebk+/Fp7RRLm/wxUAWHv2+1T1td4C02S9y/W9cDG7TxYqZOLIc6
IRyzbQ90g8MSZL9Bj+buCs/4JPQZovMvcDXrpk+SXoDLmDTTJbGG2nClBiswmYhI
Kl+A+cJ0c2wgQiM5NrOsYBg3pmhnY8jjqk9MUG8JkhbV4c3GKLnjEusegUF6VWFu
+/gf/W9CNbhsNbm3n9AKVfBZyiOLmki9rzmlAd76clfObrk4n4twnkbpE9MAvw/Y
dsBpUrAizQdcCsyf9rZrgeUPrRDcj+O0B4Fit7vjKLWuEyI1trWZ1gD3Cypxn0kY
L4O1DTaEaOOHRxxliy72wJ2/N9UJxV1vnkMSL2UG2Xgj3OhzgXNCQfbJyv+5j8ok
SyzZs37twhN3cB6p75iBH/7FYxA1IQu81zQ5i4bHHZt5xDa00vo/7vPUZxUYlSws
wbJzo3+D05aUboaYwwKEIt08UJqSIHnb54tXaKCyvMRRarYH31/rLMX5oRJtpyB+
upr8pIR0DJhN9DgCGNncAnvR4YKxPPNFjbb/Im2lSR61OqtazLk7V0wr7FPdbcJI
DZBRP34FRuI9e21M+Zy0ryk7QKMYmOxf8x8V8XsLaKQR2+o9YOabGgO1Q7qcfSt6
meOJXbcvRcgWKFuMg2n1FItVUQ/jCBBOg1Mmw8yW2DQji78Q7zcxl6mTj3KpFULS
XdJrfUU4kSt73wMsczLWHSBZWZkz96whfKK7GOsUM8MmJ5lULu+slNK6SykhZDmU
OZq1PKUxMWZla/PKr+wtNjCtrzg+1VMpeg3DB+5OYYTXm7rhy5xFxVkHQuI4aEfu
9EdQtESsAc0GFBzTcutO6mWY7ntHQHIizwKq1A+hRO3ljRDtpnxnX3Gh5CR3to2n
c7LjqL+7l0T75cMV0Xj3paA/r2xidY1m08P9T31PzWV4H9ftmzmgXNSog6v39u4f
e8OAhGBaUDjkYJsFq1CYy4LaCicqys+E1BZyv/4XVvLcXWjo5bbYwAWZSCVGClRz
vgAUKVHfu3UeOuXV4s5x8Kahs3SECEKkp//qafrQfLTeNTbiCPC82NbIrwMI2a0e
uoCXrb+O+lkGaP1mEbs+ghR2ynINcNH+2L4Qsf2nTQn53M5oJAS1Dn+ahWyiXY8Q
3Me+9qQkp9oihFZ++ptaky298kvJfWlHAepB/6v1yyo7UGAtwNL5G7qO8tJROmoe
bl93YPlgkWsohoVSXfk+5iFARTNoQwnVxCuXU+B3RQC7jrYOZAvq7Ei1h8RXixK6
oUSZ1aVJl4gEsginYOejvl9kt9t7J8Tr+wTN0kPa2+dtczRqN+G6WKnbWNlxz6Ej
hU+Ev0oUbDGmzMQ6kHCqOcDZNSBvNPeLb3MBZnVqReq0fX8BYFVUVwhVWNP6X91U
6lqhg4RdQal48KQTiP4jNBEmbGk8k2akazUaqZYyrXRU91EBgftO63UtG9tI3jLl
+W4vblTw9+psWssKM0x6VPsXrovy0rU1uinMhrToaEJdJV+lrzvGNG78LI3q/HgT
pgYY0iztm+1uXyjb9qGrU638AF8+CNWF7zVVXW2imfbztVitMo/WSLnpqIihSdvx
1CjpK0N/UTwXacX8Vhkikqf/Cvk4TjBVnM5rwmihBsC0Skqkt822t+GPbN57NtoX
TTOxcwBrDLQxlrsKaDEVmdwJN1eSqV9qmowPh0S6xIS3yof5YhenTgTPQuYZv1rg
GutKIndj2nGtxjT3ztC5U5ivgt0DTwaDufx8EzXPLsPHWcL7OLPuK6hCW5W10y5v
Ic6zAZW/RAIsvb1gFqjuxG53zqGBzGC0BjsviVS3RY43TABmfd5YXjzDOQyVbjQZ
t0WlAKp8gAAmukirNMnLSTmjJGnM/suDn6qzzcNIwlVwhH6i8GfpeUb15Suy8Azn
vSAna+J0Lo3WfOnvQUr6MVtfazz4HDzJw3q2+sI4pfpGAmPXRjioUlb3jdxs8P1B
pr1f52lfiiNf75IZ6Xg2V8J0L5RcxcqCcJL09NrhTIuWWXSCRnL+ojx1TcVl9oJb
szoIIHMjD/ucdq/HGAeTrSrGVi6hblVIghd4ZZrrpBDtkPRbj2Vea0FBVUF/AMaQ
Njk4GIB9e8aLe+ZGLXYMKCvjayKnW/jadoXj9gM7nWOyfe6Wwo2kI/0AsKBYmA5F
psvje9EyZMZ7y/Y6fJThSBY7lVqHXgIw9xkwNgzbALYs0/R9SOHb/E90TkpadoZS
ASoCK4pluG9FO4h5NAz3hwf5ABVIg5YysGyi/RKEo0f9hWtAfBQeTvJRMPut2c5x
gZHIgqftUnabzDHrxeYwvzjkhmkuNMfz92IvwIcGiAm79y7bthDSJJuS9rRksHXV
3GBLLc5QVhIXFoSlyo/vemHN5YRNCKX11zKWnb13QsX3DmMKqvrzgrnl7fvhg+Gz
k9f+agSAyPGz+jMTNe4438d94lSkSIzCc22ugccAmDayiLSxYNOtakh2aXSLSiEX
xO0QXMF/PLHw++AkIyp6gOF4Re/yqFT5ipJwMEJk5TrS+iGc2weSjKqtK1j0h4rH
I+t2W2ZVsbZB2No9I0xJXgbTQmkPcmpO1aZJ4tAvwpEKLlbRrPIO7v4tubg0XROh
fILXqEqxZP5ly7ZIfKpDH2CYKx/sbUPQvAlyQY8HH3tiz4ZQiYTsSc6eO3/k7haL
sbW+KORDNir7i6CrQFsh1JtrPBfcXhWptr6Wjop9mOqa2QIb5hWkMRPzCjwsjw6P
d6kXDCY7Wsc7iRl6ZNTPQAv5g6feqHqnhCdl+H7SPG/8DBONBlWG0qLWN9Vize5m
n0VNISomTlRKEq2jq/fE3Y7nEe/GVl2dZZiIwRpVmp0B099FG9c0G39uM/3MeSKV
qWNFnl4TjoyaCBOijJq5Z2uE1PrEv/U+WEVPn0v6JDjintQEbCPLWLNF9neZZkcp
NMdYOpkQmnAywOaC0K62eQTYFiiS+/MAA82SH3M1JXSB81/5C0ROQIoYikCgvOqW
kOAlDuV503XmlBCvng1xQBECKzwfze9BsmtwHy73iyihYn6DLeLy7K/5HYu4CGRX
cTl5kMsdR3wZzoGt+g4ouAUSQ3dB6ycAvvlr9m0eiLyducbO+RtZh4aDr6axOKtv
ZOsGMqAZgfe9iSLxSUBrcnRW1E+7pECOXNI9YBTjdFk4iZ37HhU7q5pV2krjyiYl
KHipTH184bq0NASKOJjO/neVQmU+KBwuLSC0k85F27zFGaQlypqcR9XFvcg01HFG
2u82W+acnkfXN5VDFxZ/JWUfEL/I2UE5G8wvtCv20I0toBtO9ESW7VLmBg0P+z4z
d3XrjGOGybmo7RavQdtcIIsvsUlhp7nMJAaoRKxhY5f+f9heNMuEU+SykamUp2zq
doyqLcbCfQkF+A0weEclBXYTi8tuAZdvYIipsoqOt3/GO0pdRiUaLbKpFKWXTQbp
rKRDXx2qKIeTcYutA1MEBRvJUKfNdTHfgLWWuyW0Pt0vCvFprc2ZFUY3+nPJEUO3
yGh85yy8jJO1oR39f9C/BfYTC0QIUOC60P88sS3HRJClqcot1kQOz62LltohLAXZ
HVI9I//KeATtWw47tlbjo6urec4zImtJ/Vd34vPHeffCfWoAPn1XgnQOcx/NI2ky
2ZIUGLM3OxiKvxbD3hEnpLI0qAn87oypkvhkg9/E9HOFHbnnXOIiXP1eRr7HpkL5
0FddPNpsnWWs9Yqn2sHN3qWhVUMZJmgSZvlLMiinghIeZztEACMxIxsdZD0AfAe5
LPSg+eIqjcgg+hTOQ2FaCJJHdS5Y9KB9BLYEyS/C9Q7bRE3nXgeZ+XPJIz5S0qxJ
cxcGt1C5jQoxiTJAUuFGX4JWQCNFpnWjRJ2Yb1+UU50wojAY5rkDx8SnyQ6u07mF
ShqNaKFknCMu7WcW8/UgdfPq+JYhnax92Fs+rLg+EAmSNCDOEuyCgqfw+DVoRTgm
c7uN0PDhVzZjaCtfpK0O275hmenlrJLntEGNOFmbrJ5V81+kW5AJffdlYTLyrzxN
xtqk8LXTOiCdoubMlUqvO7xWXe8ZRpb8YSL+vNvpAz1Xi75rNh96btXm1MWRQQ14
RFNn40zv1s6hTz38Kbgrfo0u9XRaNMFQxcmSfIMIio5/8phwXE9NdtDI6oeXCmF9
XNvtih5Bev+Nz1wRLzX5mxEFzJ9lnvGjy/SXg+S455WnrYxmxddfZKPK/kWNRKQx
y7EzmgZGAHsiVNYDvmMh2AKMV0SCo8XQ7RNht3g/lw/olFPYV3XrFrqsx6gvH8k5
pw8Lrh8ThEzZNKpmkg0l7UpSbuuauOfnKv4HsfHEvdyFhe9OlQ3s8c16cJWZacBs
KoN0VQPK0PT+i/TFWmnm4N1ophjDVcgZyPTqHbK/AKRPQBR5KHwpsthy7XNAJd3h
tuLEnBfBWYjqvl7hHhG+B1fturmoUXCC/t8Rob7KdF8JghiBPAhDAyJzxsfFau+i
0HoaeBKWLMtJ8rePcRstDDTB4wheTQQZckoHjs13iQEzi4n5nve0UOnV08tPir7t
J6mYWFJ4P9/Wl3BbNRTDoZs8JcEi8jejpcAKWQF1NPPSzxjQAQUsg3HfaG0mldyy
2TleZ90xaD7QvsScQz8nPAes8WDfjQcnCQrgJ+41bt4PV0B4UgBGpHamSBoHiFfc
k8wQSiy1pIqyJndh6w8eBalsB1hxXxouwMSwmh44a1xFYekeoMgeP5Nm5aifhvX7
7dbZsS2BgT5UQULIMfgNPUGvCL1T8yz0JaBOidecQLlwe4n4zEpffIZZJmN1RUfv
OE3+NZIN/MzpbRGL+IM4SGHLz0gQr9Aa/dVxJkVhd6i8tkQjRcg8OECeWCrt8C0Z
Yhq9PiylV18MdsvzV6TwtMyh+FpV1MVNx649Udjhp74AYc2HZfOVZ49Y3qMJsy6s
lVb02sKjwErSP/oLTi0G/inNCauAz7NPZ9USc/jt1fq2R30h1lesynWqLuyI+3gf
5dWGhpLbRhex1eEqzfIv5Y2d44DSNuF+5pA/dSgKFTIZ7seMkwIhZswhB8oohD92
n8rOuxLL0Ds5YRoYgQqdulgbSir/WM3x0Zg2KoB85xb1k2LJJvHEc3NzgfUq26kJ
eSBQECU+EyrWoegGeJsPAZKvRsUwjc5/JXVQkGwNBUodVSKSjOCEId3p/ToyekGm
GK2PoCs5+fBFGi8QuDvhzKEHHnr3McYvAq+VPHlIqRBEAmsHbwN0Fled/dZZC0Rm
Mcb9IB7BhEsQ7e9QuCdcno1AVDurCZXGWbTq6TUne4TyQEjI/+L7dFzMDuV4JJLY
qWp+KZXrll1X4OHpDZCkzcNdC6H02r9fDlfsuSKFRoWbAXLdUEV/lOFcE68vKB8k
lw/4xc9ojjoJbMWMXJI2G7H39KyJ+6vnH56MJv4avnYlOsbBOEQih8y7jDj4Ue4P
XbxzOzA1U6s2yqpswgHGoND8RZkT4e8nQLkTtWrklcDAmMVifum5vxMaMantm8AD
ej4R44DPGk3PPO9IOS8n+GKnBCG4D8hSkNG0zYBQ/6Q2KqoRM+ZJo2dxhHdftPhw
TRXJJYjDvjwY6/15thMoop1uqm4uXCcKPOr33RtANh3CSJw9+5bYdduL0BTPKRR8
dtxT3WB5BA6t2/R6ZgOgP2MTYO6gmWmviFEbaPxUoNXGyyUv81zaowHOUW02rTei
V6e2R7dFCTpCBmqHalmDvB6TVCoAdsync7ftMPMXe2u+a9FPlFe0USZBi82OrNhP
zbXbkuPq6eE0CiK9PeRxYAJ8A/TN0Q3Qy1mWqORUliMDh/RtbhkL0u2CVxmnz2M4
/4q7HEnkhgdDxWzkW3taB/Hwzi76s3VvT8g2/TXVePicmd5V6/zRdhmoofuHna6y
bABKJU/+6lZcB6cvSsr59AN/Bk2D8hDHhx4Ai4XbNKQ8juPxKDS2VEjgbSuZOiou
n65JEy7KZ57h/EziWwIM0AIPZp+6uQtLyzsCZeiWqxQ=

`pragma protect end_protected
