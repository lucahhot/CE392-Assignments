// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
tTgvJwdwm+HMPVslT9LaH2KV5zEc+cE7ONtP/w87cP0p7nedXdiN6Z5+7U3zwWcORpWgXnLjdxcT
Wf0COEVrvrqA8EIb6GnI+E5g1lyThfXc5I03UTD8orsg1u/WNSuBtk2AE4Fp3yi2CMtqD9aj9nCd
Cu5vuNPTCzF776GiPkK4PXe0ubbGsTCiLA04GlAgV9RkDznxPwIslYeif74/DJEhka5SLQ3iSnqN
hCaNB78mhflH/6r5tPM+sMebw1sCi12gfh1+emxzmoHyLQGwRqg1jD0u6QVXzJiu0VGgjs97VFf7
D9c+dbW5xxD57F6JTH9/dgctXVQuNvIOybJnVQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6336)
9JqIli71KGC0rhxZ/WigXewrq2HclNMlhdvUQ63UowurCEbe1dK11/EyZJc1f6O1uQ8kip5/5N43
bPO9P3P5FnYDjezaXRxFHcfZ83Cw4bi2Ci2Bc4SpQeYEBosqt91QcsV7QYsmZbm8vfkVJdWSK00q
vf11iANJ7EQTla16FXTb+p3EP+P67ln42b/k0dz1d+EGDuBTYx3J+csJEIx6UMJJcaxecSb2IU54
aaRzvMuohy2SZzAT8sMR4u6ARCnePJ00e3jCGRVPXHV9RI+UZE5dCJ5fqQMRAptt3WO5ukbXKTVZ
b13GZz+/5ypmwCqhpU6wQu5Ag1fLWgN4M/5lWHqPBNMeVfhodQQO0THADLtqfXi08Osly7R0Gc66
2Aypm26djxDmfXRokfmae9Zct+Q4HFqKRokih8+PCqGG16jfThaN+BLrfl1IdngiJsW6wy/aToHm
zNvg3FaRJAuZ7PKbHYJqcx8+cboiFOheZss0GIH98+1Dh1K26Sk4KRgXP8Lus9KVyetzl3jSYwAV
rYocq0exvIsCcfYHD80puglbgrzzXxUUvfc6qUMjV5be3HLey5JPx8/ugNxYQuacdDIRrEzZSGpS
OvPfLrJbsHBzRr0kdzjH0hn41HIJ/8uvxgrFKOCH0o3conr2f7akoauLZiYpjhHoWqYMjVQ0NAQu
qzdehGycbQLnPKxo1kviGbdB2gtTDv16pZYcsOXsrbjgI00bDvymaUNa2wXGD3IiUSX2iYWsfSvO
hI/T/+9r0ICw5wNmkLtEZML10fnEo25JJbbFibL4JhVzIkKkSuh+S5Dqryfh2FSiOhhgGvJH5R52
mZnGQweMd0en8aME4bCUoydtakzKMMuGLu2DDn1348G73AGhvB6q8OFqsu9M0ERG78cSHNSCHtJD
kyMvh7C74KfOP0hWE5tmkaielPbNCjs9k0iHmk9ChxbzdtVDfGF94pyuLH75HRkOJXdzIgcasBQf
9bhRN+scnKUCrcZO1rit5OsDlX9VsHY50t0kv7SOjqiQDyUpvXnlOTxHtofED+7vO4hZdqqTD9I7
LfouWOYTIz+tkMcht4q4b2a0QEHvKhdTRPRpYDsYtnkE+gp5s9sxMmL8rnbB0FhaEKF4pQ+YR4iO
3WwB0tctXBdpyM68VoMfXhi6/aMm0Q8aOkojpIZ1s+QoAB/1ATwFZ4HLg1nF2Qx5iLvQcTXUeC1j
d3j1orXICKsgm7Fy3eMQswOkF87HD5fu1LyEZoPaBYsUcNbMONSOGV9xxKvgU63P/MM4CKnK/Pby
DcwEpXfNwqXZveGddvt5mdW8FgPU0anXLwGa8GECYTMsl3qzVhI+IkwBGXkmgGzzDThTUen0Saz3
VPqdueV9QyUtnOqjAdoUypHmh1nC8zxOPyCn++kp2OkEyr4wgYwuDVfW4TCcH8//QiaqNPpwZ1pP
freU3R6Y313FDDhVzR/Xhrt2CByD4C/0nt1lfuc1tkZMUmHAfdmTbI8hjuRnE7Gl/J3RHPfJiIkR
/PXWVNd7QLn33p+8fdHFLKz8ujqD0MBV1QvqfK/hD0926mLkcpVrjmdHIvv7kn78W8vkGqdgfwdA
vBBiUyXTAb8/4flFK6xM9HPTGcMqxo44DJtrtGy0paU7Q6GVe1mD7Qc6ZBbGLwDsH2soOPvN5RTg
4pRhVTmYElGyq4D9SGAefpgYYTvUvRxcUqiRz8K48ETBe3muoQPJjrwHqDi/trhmK/XQt2u+aM9m
IXwcjydIdDCU7bcqGOSmdK4GXFRHUf6w+HkaeVJAgjkTJ1yQFz6ZNG88kff0kpR18/fjZLzGiqGo
yvLuIHlt/uZP3fNq5bwam3dHK1XNHMeiUdgBpshHZek24TLs9aDYw5qiMbSHJHGhTmuLeyuQHenv
/vFHrzOG7nUEHU2/PnU816Mq2uezG8FGeyQAH6YV+q0KzaoxJZp78m8ochdVJxtPdmAC6q+RzDlZ
+jD3QEgLrprTyxALcVIAMn/U/usU8Z5aQ3m+yFu2N8J6uRR8pbXmMB8b99cd9cNuOpWjPd8EnnOa
zII5mfhIfHoG1806f9nW405jCAI5X6x6AVjYDDo5ce89iyULv72yOj9QWFdcueLc+apXPZ/rFx/y
ZyJr/l2yzvVb8neFg60LxfTnJjAp91HGTrOEf6jHLpsEvP8elIK7vvGYwnAe69tFjDygfH9glwhp
cmNece3FdaMV9hY9GCR0LKPWwKRH/CdVw0V6Hr3q25ziRWc19dHNpOUlf5F8xevo32aQb0Mp/WxX
0PSbko3bwAZDmujyUF39OsjFXTmQ6h2Jx+GOlYNujjEtYVx03pwHvtocuiJLHMvjmxf+TYpPDbRR
HFXYHt/RZ9H2NbZUCJUUAW4aoJFEOnyzvT7kcQtn7eFo9yspZMcqL5tRMpBgj/KwBhYZu4V6twD0
ISyD9ZJy+6o5L139nhsf9/fNIMqiRhKTtYJIVGlxl4X4IPbeLxiE0fpuTw9V4LsWld93SIWtCfje
RaVgBa/a0wIulYi4w6AEL59kuPgy78ak0RKUbiwM1QqHgPzPHyVhN8xR4cYCC+73VzksHwfRZV+n
Qb9hhmK0uix9ZjByTJQmFzASNGLO0mVjSoMomfSp4qUrGxjA5ewRu67uPn7s2xafQ1EKuox+QTNe
I1QDk7xQg8+pgZiswcQC5MQWGE6pVQ+huJvcG/qRUNDIuzF7Au+JBKm25Ukdu2RNSo7ZMACgpPSG
FZOZ3me0qo44UjZ7FDZlUpI+dZJjNlX31AKdWUXRW8U5GOAcM27rytY6jctSR1f9pZoWpwMu4hEV
PmugwvLOOTGm+qX4bkFhUdTvtDxWtBTfX4bcSbgfY43HcbMPPVlyS3dxv3AzJZS44PopQZcST+5/
U7eB8gWRk4SArAQ2O9GEdVcurqIMtbkSOHpvryHqtz5iWZ1I9w187Sf7VjcEXQ4VXwgl9rfR5YOo
JgEy9rG9peKivhdo6j8c++ognjoO8uHUmb48MM/6FBbUJxoIG5Eq3eTxBIWhVad9h39XYfEH8eBd
dHBK0BhxT3UfzLremlC5daiGp3mySYO8hJ2X9bBVH/TBp7rftuM9UnwD+2M1RlTqoQuxeS9de+Cx
NL5qJ7FJxIuqXRTzFwIJT55/Jw4hXQ3w61ZXvNntkgVJ/C0ncW82AFwsBkFw/gcQJpzbtcdlCpV9
VJbnwS5MKGbXmJbNd2Yv0UBa3oxf8vTh2mPsk8AjPZzKeXA3A/fxbO0/hoEWkrPtBvO/RxKk/UDr
5QSPZINSi6kTQtTrAv0DgALuppHf6ZBe1l4BDyULZHR4a6ldcywnHdZPcJwmLPZfnnaMwrbP4Ex1
eWYu8Z9AiaBMracfADS8Y5aMe+CV/PGG8kDa3qY0D2yTPUz4YcD/Yb5xA8lINReok50bTajUVbJQ
uV98ZuPt7K29v4MMERM0p9/SfUG7QYGIYF5WTxlohDeRSyvOq1B1IQeprgLatFxpsg6qNWkn5yZM
CQoln4GngOPL5v0kcvbcWDZlh7R2IYFBAgGXZgjSXrNteUmtywOFAdXT32QUKO1VWZFcBgoYTH+B
zHk/P6r9c1tiUbqznWAJjOfiLZJ0mZceehXh2lPDvLZ1xos7h8BlDAH3qCSlc8gsfc+PhPkkG5QJ
ZWApCVDoF53z29tMCnhH7BwJL8C+CWx/zyQR7m+Ek6I/CeMIlwJUQ4n+cBpNoswNAQVGk46+mvSp
gEchaXgbGtJB18cw6NogmGE3HAY1H1m/VPVchi35IFBoaIfeJt+4fA6zOnavcFcxiHidf3UokVSO
xZzLpByXs+oEVwULL84RVH14gYJKpV4Zs0I63SG2no4JGAnvwrXjQDoaNW2G5wmpS6UYlEspT9f9
9xENFCsStd0gwWyzvMmBzPvRmUlViWzKI32Gb9bgIH4+pt9UigCLpADY7yv5zgLtm24uEiSwLOFp
+be54Ru2CEIXfKjeFPf/ypfNZD5BreoilDuiZmd1i+2ElbY4FCTxgqNM0oOgAUKthnJ0U1ioan+R
/9zAps6bqPKTuwVXjyET7wdYsFQnSrnQ1XasQ+4za1pdiowvN5cTMblU1Fs17Zga8YVaVQsoXG4o
7awo5+HG5QE4lkCnCpHFRgzHfqeojci/6PAR30l5I/rfaHcmHo89KPSthpHTY05UO1xoyhFyX79H
f0SXwVM+pck5enwiryavCOUNdoSxC6Y6j/Tvs56jscoDs/H6Iwfs6tVWKY6vVeO26yXCNC3bqd1J
RkVA8qrIV+zHO449/OyKSw9XGcrKcVnL0HDLWxahDDVZ3ZEz3byLO0F5q45y2qENNTyCWbCV8Bpm
f0YlYXMpVN3FOHROBxhbb4ueORWOILeyMWYMPGSTglxbAx0ATFHya7xEt6umGVowbD35exfPmXx0
aYzy5TDWkfmEBtsLj69b2w65k5XNwIp5fbQWG1kAScPHpAx0ihy8L8i+lEflRWlrH8fVbIxzCpcY
6ZCxrnY0jGUiVoLPnJaI6/uBm62iWAaPLIOwZG/yEtcIUWtMSGXhyMcZNCW3UQXf2qZcAGhbpCa+
mibMf6OM39XPhQEmEPeJbOZJu2I7OKU7YyPS5yES9WjZFyhZY0JyHw95bvCaujAUoVI9yfP2pRly
WssrW8Qkn/kyj4VOTqAeeb3uUZHGFaDSbGdcIJq0mlcKSyV9XegMpEswUndH6wITCAcsGQqEzrbf
Lcop+dXFiRoEUrQcUgaSjvzeOHp/KGVMgLbHLfrpP1F20Pbi0lomp17qUUzNOVZqNL45lk/DNg4A
+5AdCadSWBjrzHMtFnWCxeUW98Er5WN0HFA/OLR0vKpq8K2Nk0UHpftq4BX9ZnHT9TCgGE89EaO7
mRiFNg7QsPM3AEbZFUo1UOS6ypGRSSW7dDQkpfTcf+8xDc5ownjJUdCvu8ux6Z3Rcmetb7yPA214
eR2GpZ05QSkmLeIf7RxjmKlGu/ZEv4qRr6/Gd4oRPVILD/HMkr91RDtkJZxTb4GMzccBvny1mjhP
+pooHMibyB+wFVYTz0uB2ZStBxK37IC/MxtWVyA8TGItlk9egcbGGPNMlAKsck89PqAba7PgF3X7
ReXC2rBwsAisVsm1ycBAFRfV3VSXu0QC9Jbw8JFMWvTk4E5rSynyt16nbWmZ/Q88bBtNnEd7ljWL
/FmqzAfjt4w63+k27+ISlHt4eclyIhZ28DIX/Jl7h3Y09ABaTRjX06EDAgLjAo/vh0UgUok4xk5E
pSUmQT5tHR2uXUYwrmZX4oTQB2OqmfFecqkyECKTF3jReQLRXIai2+fAi3MRuzS+Tm7Q0YpePBqu
4xYymCGuXA7Bw04jEP0mCr/GyWiPvONUsPpKNNnbK8J196CiliKgyRmMJdAeRdp+/NkzDcish3a5
b/yt76xlbemKA10ztHNhE1ooUmHVR1Cx3wH4LqYIlfpKJl5KpigAa+aj2EGya1HztIvk0yyGQSbj
wXHzIbS9vXWxPCGKrGsMUmB+GMYzi8r5fAaz1ubQ7DmpUNAhQx8KHTcMnmkrvIGq3IMHfaDpRULD
ofyBU5R1cupX4yHlFta6fGJW1XsAgetrALnOOPiTN2qyxrLyotyBdDgQokf6qXpS2gUXVzj7icXY
Rj68KS+qoMTQ0kIOzMfl6DaXoLCQZ0fs4yspYYCyui8As14z+Pu1Zypaw9UyIo0CCOZQdZn4INnZ
B4uTU1rYXzyI45SS5T3te5k8nvkH396rjsW0YTSxgQZ0B7S0V7jUWgpXvL+ifgooJkqNCdAt+zI4
L5hb47BswZk8HAxgy/xFC6AbxmVsQBoGVobBa+SuY51lT/C+cZgwfo9aB4E6bAamI27LBZsCQTeW
7MB9EZF7DkZ3pdCK0TUmzt0EB8sZ9T6CPySCAd6ziBSSBhtrvt5ptf+vG0BbMdEyWxqQq6HcPfVr
kdmNibrn0KzG00qTlj6WSgLfsh+2zQWVbnKxS8hyfX+VpMM50SqSJXZfu3WeKygvfITeJGX/BuMn
ru0tekbkpggKvO4VT+6euuq9UvFoytgo0Yseplf4QsOjNclS2SQN0UZvt9ZvRidUFUFjI3UpKVBE
CNVTUO5Z3J7X9Y5fRY7FlKHX3t2/hRfA26T5CzJ5xtm7krkuBUV5jIduXGls3QM2DHH746YbGwen
i/eYmvrKcceaZsh4aW/G+f3On4eDn+DRL4RLJe3Bl+D1oUSN/fyoZbcem5wpvJ//3f21JfXc/xDw
y8yMdA/KLJo1MkixM1e97q4g9A9BancxUq2zjJNdoyZhROifz2VGX+Tj7/3QBmWCxAXRh17lwrEg
DsWu+r7ru6K+UJTyNHUDhVUuY2/H2Vz8k2A69EpEadntpTzDJeYRFJ8vsaxB6mCSiCp3vbADfNyd
8jMmmIYKMHdMr1BHazi0brCTPie0b8ALHUaKO7akzRVSBjpRzvukCdoZGCYqLBtLJ7oeH8o4Oo3N
KQ7rXES5QU151Wt2PJjUM0Tn4nGn3NTbWs5NUq2QToxyPA8NINlnCIuSYBmP+UTZKmZji3ouT4iB
sFcbaY7gnjtMl5A6WdlIpRlYE/W4pftA/XtV8FiN1rWWGQskYWnfK12Kz+bKcSwja/RMwIfWIQlA
lmp/+dDV6edUbf/zTd4CI9B8ejS6UPtX8MWkgOXwKnc3eWoT8y75mI5gWhWa0kIiEd6W1Emb+pb7
xb1q1g6hIEBoSdh7mVjzjxCX+MrYGXKe6B9IXbQZeaH0o8Rzqfy+1lKaBjDDujyk7zc7KWLKgqOo
4Xzm22lFe6LKdWvoiailXR6oR2/7J3/m28oDQ/ep1JcQHvDwwO1lhs0ionJD8hmDMzzVVjFuiIQD
Vwyf7Vfx8uFjiF2Lf2G/T7CiDKSdXTf4hEXPNBXFn+9qpWUToh60vM3dXiXhMwv3bSL6ZiWyd621
4p7uOhxNW074a+LoeGd6GSK8za94Ps20mXrooyCZGy7oNu+bPzYUG1F8Xr3bho4GZ8gV3sYBo2+2
txRjRAjlVQeI1lKg67cfyiM2R8TRsa/mL2yktWKxGRTNStOIMOOiQORj+L7h6InhB6e363EHa1Vz
12iEXE9iHG4DowJnhI4C2QEg6PR7WtL0wKF/a3sZoO16gVwEx/UmjVw/Rf4tXj5u3lKg/LPGnrLd
5n9oU3hTnfuiO6oxvUKsXGJdJkjuaaL9D50pUSBJ9nBEejMfAtOpgt+bjdFxLAofJGMrPHSAP1w9
9GoxpsRSJdKzaJ8JoO+LfIXrWZZf2b0MKq5IXOjDJvlUfWbcAbZwUFBCTREnvRLA9qVoRqVUL7iL
Q/bwdF/mg1Z4Pt3ouGwK8dlWZxfACGd8crKr0M7pveph70Jb8/I5icl3i98qiqWuDSmtrLpAXghi
o+dfr/VJu3MDqSdaBDjxm0bi4jIFqQAdEr3aw/HKBvgyQc1eLU33d4dSrpO8Egx3mSOKNiyzKdu4
/i+rE5Kwpjb32FSss4ETgDIh0h8ynT2aCbOi6saT36yA8v1xUe6Y9pZJYh+sHDCJ1jqMN1cqfcd/
KrnQZqMeLC+8j2XaAt/4LOzetnUMaBHMkeTo1i5VeI00VQxzyBhrriTD5xwIISODnRkkYJyLSfio
HegoHBH5TqgWDf8iCzkwB9Cit//l/ZHdWD1hcj/UnYanx+oErWXMqZC7hzpOnflKyhL89urEQyEk
tdnYop9+SKz1HnPbG+if9AH83ETmJnBDpuGA7k/SQW6yb/lS6PeKPjw0Uq0dzTs60O1IWXwWsVPU
vKy8d0lepgQsmmUaeQVEd+F6+gzzOfr9PLhP/x9zWZ0maR7RCxEmWipK3IqZN/AGAFmkIxXIpITq
kOlHNfHIQAmjuG/0HiFTNWFkFIL87iZK9afdJF1GJH1WpYwp+iKFHJrvMcqS2YAjXNsnfmzJwv4h
lDdjV9fmBQ9QgorSoMtKJwfT2+0G9pbVJGpiIC1uZScmpuuhKA4E9H3N476x3XYun/zts4rMSg/5
2ffHLIovHquV8eDfk0qSCS33oWeUXModCzYJGKoJdwPG/0r7kL4DX0KSeX1z7Cd6HlzV2ZYJIjRX
vkxqCzi9xjwVpQpHSzCJKe8N2QbDZNKrQKUl5j2L+5jAG/8zGiZaB5unIrefieib+oUM9nF9aa2B
Um2/opMIhxMwprK7hjSjy5i/bsyy98cni1ECDqg8DMvmuimnBaEIpDj6UXHZTcosKenfo1R5NELk
AyHZFV7gRFxwuYidcX97aQNJWymWC/TN68BKViP00C3GyKSx4nHJdxH8tv4rQwh09AZoP86KPxRx
90EQlKtSmCo2zbCLTgXukBCCqkjT3yzBH9GQ9g5Y76JXrQbnD66Y+ynwM29G2PPjtAW8u8FqFyBg
xyz3851cDTH0xuFCBB0lwnLfvNvQbxN2PElzST5tgCSpPX9KfyEyg73/WDsvjYJwm30k8vb8aBrt
SNzsTAIFMGJt
`pragma protect end_protected
