`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UpawvuYHpZzY/spItBpqnuY/iqjVnOOkES7LYZHEI/U4WLeU1X590n76wghkaS2W
Vq5kUuS6OT53byLHjn3yF8NcwfQFEJiy1/PnOM95o+VGpplXvKuR5Us6OOlytjPo
Z0SrMcIwPV+yXaoiBv15zzvUQF1FD2jc0MNyZrfEeyo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29856)
YHEfY2hs3IGjOSPW6hohi5aprmY0xqKQdM6dtpl3d0eFN+KEQc3rryw1TWK7fVYs
DaEYmoUNQD6xpJalWmqzdfzsB8iE49krA2BcrCMI5ybKkMQqOi7ZmybmzpJI/mMY
hd+dy4WmXrgdZ+rtJZWJCCZufNXGRWGIrVjTXkdgRKpo2eOAN0a1iCz0X2+Ge5X1
/eRa3eg5kkB77VjCTwZTNncJTewJ3sSwSmni8369nxK5Vte8exkWVOT3wmGwN5tN
Xh8VMG/M4cnSnL9Bpos3zQ8Cx3pjgqbFyuG9sIxYT38V3wBYXDn5c4MsIAnvHwBi
CJj8HEs44MUq+GOdtws2O5qeM8G28GuiXO8jRpygz8w8jHTm9FspzkhzL+31iFqS
eGALPu9dXuXlmB23ur15G5JwvInOnVIRhllA/l4C2lgICMar+1avfwBvw5KhS1lk
XR+8fP9nvImN55uRJdg+h0DU9CODBk/uSMcIEsnT3anlmxm3fXXfm1U/6hRxQilk
dhOrXDRv/zfPdSlUF+/Pi5MOdjaTiuB9BJJHKbYMAW4f6ZIP3OlrUNHhcLDXsxmX
i2IHDhVVCnIUS5lHLPTWkiRkfYBYuUCMscOUP8OYWeR5wvyP0QD1b9pFUpeHWQy7
/5XYtcAjTExcu/rwLGtHmL6VGXnV0rF35/qk4AOQpcn4ygcbTeu4L6u68PktKvbq
bDpScFONvtX5pVsNI2HbbJudxCGR5/8iAN0aIArX4AlM+37f6klRcQ3EZ5oNYTC+
Iaq2rR1B7K4aCY7z/PBNbADQeBIe80lb4xBGrnvCU8Bvzp0dvyTdWgc9RxGuNfOu
lj8bG/fUAZQhyjT3drzmTXHoPYWuFij4BKalpMiF8wxGYhIxHF5dkqP2ozW6yQ/u
Mj7qQ2NX+e9f84E4Yl8i9XPr3tlB2khgaS6QBYnxSaKn6FjgZAI+Qtj6/5CCVvFj
8pIFKPFouzv77sk5ajZu14xXowz2IAcx/Qqq9pV9w6/hPiIItGwSLoLVRUFVUXPr
MeIrgdTfZvcPC3eTuiehPgMJsgZgJd89OolO2UWXip9wJ4Hqti8MeVtTplxVlEFZ
jVBAUxAa19xyBhgBiSEmmFsoizj6UXeekssMIYbcpHLXDMc8TNdfGRVuNHsk3mBo
Ge+pp2GdCtcMFWCiXl0GhJ4Lvhqm60kSVjRJqThTe/FuhS2M+c5dosqw41McXmUE
quy1Xa1iASXREHXBbt6IGvFEIaewUIcokaxRtERG/yrPcPWnG5FWI9ZhBpj+ytuR
/nKbtuOHSOmupBWyCOkVS8AbK7RsrHTHrTkCvkNbkkPSwCMcMXeLMEZ0nwSnRVwg
kjgIFhXVaNo5uRkci+aF5YFW282x43ybGCT33FXbhHgI+YYo5bj7AmbbNkPEkeo6
n2LyXfHMXCQAlnBpR6/fBYamidmVf4mPYYnuvdPhhNxkb52wqYEzziLjFLmqhjSZ
wtiPH4vQwMJSY4e3BSzpmqszqmiWk2wZ4y3xA4Cb3ND2suj+BrrrzUGRdgo1m3uD
DC+ETDqHs+NZKjQvE4FZ4U+oe0ZqHEypt6EMugRfV/4NdYscdMrRfApkxPtjRaA/
QJnmzO6kdkP39vxbLBMSx4Uf3qxgfmGE3ZE78R/4DSaKMBv/Bjb/fYxYxT0VPCd9
CtfWeI0/pY2JXZpfKe2GqCNXjPHUclxLySU3bgEVEsk41Nri3c+ofHYiPCQW3aT7
GfTr957Fq+dgXb9spY9cfbdYAIA1zdGtym0Ddvm8yK5ksgWpz5OdIAkAKWttd0Ui
NXPTVoPiYwe4fhO2Mh9Mm2fGCt5xr4QCkwelv6HkGOIFsltv8rVf/bYhfOczZs8L
ytJvjoRPgZ5DDNEvXJkPqXHs/SGbXB7egWIXe5EgZMNb69vJHPSjiTE90fYKYmu0
lSJJFn+tvwVn2NX9tx51LdQqtwxNaw7lnwk2FK2BLz31SWFxfL90QbnB2H7w/O79
bPmhkSuyVSRqlvmFq9iCPNR6TNkucMEEI73B2qMy7XJgQlaN4CDgdSj4nxaWCvtw
CBmkE3goYsrPbKnMvMQOerPAXo5kRPtOf1v21VTnwAgxSnLNhZ/+Nn4vjPdjuOVX
cKDRwveYX4zZt86/WU0daguJgQiMeJYw+dULlpOYombec0yUL5U61ehGsufmrIRC
thSXnXGRCyVhQ0BeL/mw4vzTCkNoP2RqDhLeZj8weoRNqm3tRpKWDIrvqSGZWwOF
+CXbj0bTvNoZAUBhwCeov4a6V0/gxOb805UNwKgvPZgv6qKbZecs8VeN4ZEVdBCC
2zaWG9VCbkcFkiKjTohOHjLeTO7BYLtyLJXNK0wOrCS5IJdAUb/PDmtY07Jub1zu
WxA/IqOLGGFnCT3Eg6nbt68cKFPrMCo5zckoHUEQNqnRF+dG88W+8bjYRw+MPivm
iY17AZF64szGELrZgdAcy7OdRk1zXLfdb2BU2aEbpi2ArwM5lTD5dNuxCUI+f+Sp
AMa94zeZ9fefigIcagJhFECeIrFquKrraQ7Zh7JRP0fFdAw6WEN7EggFug5t5SRx
4cUcEATBoS01HDJ8dJSLfI7DF7WtdwpCmjlv4vp3B6iffg5w3ezooPXKbaZJGMGc
4JeJQHypqMdymdsfEie3MPNPShPCEkhbVpmGqFimVPzMnycrj2xPPPaH24NYnER8
q5pouLjzZmeIiUkBjMikJG7mxsRg7JllQtcnAeemTtB/TpkBU9tMFJjcl1wsb8bt
zdvITAlu0xLGNXc/ItboPs97cjxgrxV3jz9HsGkt1J4yeh/M3F2WcZ2G3SM8AMWw
PYqq0nDRzbXWEMFNecPnHV8Jw1/oK+QIZbLISZYXD2q25vlktuY3b7ZUT//AGuA6
xW7MlItFNHfqQ2F4ddC7b9Zc17/h35fRsFTg4A8qxQPtcHEPTTXYmHwa1V9rAIR5
Nsq1XduJeLDwXC3Vyebo8y5cdtpkzHwX6awubsimo911sLemmX3p6RATUigvPfsl
jI9QVV4b7Z1sOxpmQAneKJ8FBLZZ0eKE7Ox6VAUnjXG7hZMw7PkmmSUFPjR1RDI4
leL/+l3gZgJM30er5Cb6u2i0ZkD8g8pGI7y/5VJ9h4iHp/DpVqGlz0RzgwxAtJt7
3P15R8SI9363sR5V7/9HbEfwTAQZ7DTa2J8BVurL3Elx9YatPFoz8tol+qT87S3t
vXV/JONpFXpKO5ouGoACD7dmNMWJDqMW/NDFgJX3pNyupaS37xzvq9InzRXgJ+PM
hn1qk6MDdeSx0EneKPxS9AG2idcPApZY+/uKMQeE+Q3HOgT4RpYT1zdi8K5LahC8
itM8RE++hPYz7pQc8JSGaib6YJMTWZqzoY8NWcSzaOexMFVsxvLkYUqPYAvCxIIu
BsGIpUO2MmsMatkVDYhDclwTC0sooRLA0dMMCgo4sgWkDsG9J4hhS3D9hP2Kpibo
9dFQMkrzoFD5v0Cnc+EXOJr1WL4dQF1pYl3eB7sgUhjvPUn+8ClLu7D2BAjHf5d1
Xww20grRYsNEE4dZ2Ul+Gy9YMpCfUHPmZcza1yD66M1BBnRX5IU2TeBK7l8QRdBU
9YiKNXzUr/oM4r9UC/DQC+F91LiKLWEeGQKe+ZhHDV5gsq0EXbvoI2S43cW+fCan
IpM8luAaZg1OjtwSoPZbQ/Fz1hX7ZBPrGe4Z4hxCCN6elwJYmv1JmP5+6CHU7po7
4NvZ+nVTVoKpLXlLIIWntUTz3EBowmgvwkSvGKMGTjSdLGk1hmXLTDKi9y39qo7e
cQ9Mwe2F4CmlYz5ZobKGebC3iY1xylLRaQCEBr3oC/ElTeVkYwoO+k8ys8C6hwPF
C+t/zThJ1fnwg5MQx+j/j7bst4q2ZLmGt4OYLl9a0Hypo/Tck9tlPyWEKm8z95xm
WinqiOSkeuj6ILW73eu+XeemF3VExSCLbFeaATSEThYmKRyfY/Yi1jQfX7qENG4f
YmjHtfGJ9h05qWBF4vDbg8zJ2aztkN7Qq9Cm21iZvKy58jOGRa4fK3BWk8lYphc5
CUOoGsKIVATHFMUXVxQufhDr5eIg3a93FMt8I+5v0CHPisOqy8Q121vVFFuFqcV0
elAs3V80eRcMmOhXmE9eFcuAup2m1dgUf6GM/uQ2UEsZlHm2mv9Kd7kt0u3xuU7s
4veOh4xuEyCoBIDPaPeVxm2a99f8DF2ceROWocQMRAl2FSKwxrUw7SYgiCl9piMA
ja5YDqP9rmR4zMRtU8j99T4QoFvozzRTtsXQveAAkHnVAC50Gn8YaDs00Jl/9Rjd
T3LdtkUDr2jX8jC30u37UI3gjbmk7xfnXo3SVsCtYjfvMfViA6Dz49YTQsvTIm00
rr4M7EZJVgi43p01P/YsiMRTbuCNT2c46N7e+R5q22YxmLe1jJuxuRAa9PMUCrhh
eGOsic9zMWRhrl3Sbqyj+wL5oSZjYsiev6vvNYYgLYcKKmDg6k6mKEcR5K4xo7OQ
00qvahM6+ZCLMKpb/poE/QUM+zDL6iEQNTgTLRyxFRe4HGNwTldFmRs7AjLFxNcj
/9L1tqZ+cb+ZTp/8JA1xSHpHDwA4y4i4rnxhu2Whlkq9TEkVbUcne/SV3p+x7Io7
vbbsY073DZlT4bL8zVb+2pR3NDWEscKVOw0d0Lr3LbHBpN8egh/cHGw3mGxZn956
akLkHsYrEnfFi52d4TOcDqyenOI10DOcHcHBKx6WelBAayG1Ot+6IevIOX4deoG5
QmcA8/gIL/AoqJaJGg5kzJaVZXJeORLIyzOHKHs85/UJsNK+a2Xt6UY9JOqttx9k
yz3Xt5Bd7/WDtQIGV9gUSQHuX0IJEw9zGlPytecfvicwgHtuzStgyEyafKn9a785
yh0ok/qHsFcdFMYGXKt2MUQhOlAtjUI4XNUGu47iWlRvSyzsen19f0f3ILT8J65n
+qosbyQ6myl9K5kzCR9JtY9u+kbEFjAlqDqltEKfp5zwdFgX6qX+7K9mBQBYgV4E
itd1yp5ZNn3otahMItfolY1zKj1M16hTu0UxR2G4rQCG6GpgmzKokQlHMHCsSr4i
P4t0wdWBe/S6dKHM3nsy1ou+4zDMOHlkkHYz1yP5K3bRwLesRBd7hFaQOXo+VnUm
X+jAPpkLP3+hmplRlQpzoYeS3Ik+POp/oHng3SBtZdTveJqBrqSgMOW8LH7sODxE
2y0aXqvaZjIYBvo6JPfpXvq74C/3WRA7WS/ezIf7/23o/5z1TOUFbnmiARFrVDh0
00jxOrvEgl8PKZl0c5NSNWQUDIoPBadR0ipt8x1q6ImKtt4OwpSvkwC9uib0b0Dn
7TxqJ/HLUBDg7Ju3s4SBj6kdTEMVMHjTAWigCcV6bdN7Nyo8buvzvc7i2uh+hzib
XOWXBmhREDNKhepDZS7QcDuIPoHaFwD5oiqbuqduKB/kQq+GaGaJHzqmFRVifHLL
H1kLQGAwa8EdlVDoJU74a+tRR5Hq8/EBzzmLW7D3wVUwTGrEdeEPPwgpwfNDW6hY
NiGdRRFUCiG7z4h+N0rQS+GiOTEgTtVTbqMQbNDtjKV7n8QseX1nvQL+nOQCuoid
2RXSYPLrCFIn0eLvywUzVTdC/v1gOUy+q21hMZSC+OutG3sbyeVU9jRkhNhVIGJn
3zUJ8Z/Wz53Apne/TAiBwVBYsC1e2KfPKymcyvD8dVxZ3ABG5kG/MMKNOXY6Yg8S
pz5mKX7jb3/PvUaudY/l0JMSHMifDaDwRVe4xcAA1Z7R+P358XAqGdTaYYK3fdt3
1PC139RAdyTRrJoHJGjfE4mlsaSLoX+k1F3+trVFPBRPOpXSJF0/blUvPpxE7aDb
dhFLZ1DL+CuvEIuytDlhEZoafCM4vBCTMEcHFN1zgHylGdIdpvR6iseJdWAZ0Z4o
Nnu4cQycVmbEx41jeTVy3HtQpI4zgJCviAVm8guknfMrDc62vY4kKQAc28eehvtb
lDTf/EU2R3tMxH4xQmG8dOEiGsxF4ZvvNsIWn1/yLPN757Ltan60F2sOVLDvHQyM
Eoij2Cmmvc3T698gyRRG3GqkTjPimbYfG21fNmN55trckoHQdY5lIEc1nr5QbRAw
KJ2yPq6EuPv8FgEksaCfWI+Ni0TS9SRUhDr6B48Moq8h/TExxm1s6/ZpoiQHe4VV
MV9yKC2aKRIv9WXhuu7RlhZlGrNtFEqi6vbT7Ss0pzpFGYZSahgz4K96a6GSmvIi
e1xFkATGBSimEQ69o7TKCCxo2pm0I33hzJJ8ICYnrxpTiskjnol1+xUkzDJIKAcW
6g0n+/tK+inD/FFSMk6rYHVOGRFRWMYpdwMbRDKaQbTpunSwWn5xNRzFXG6QISqq
abYIIrKyUYbw7+6W++1kHRas66kS1zCv9t36e2pudVH59M8dGYdRT2ckQQ9fjyIA
9wSOvTA9c6zIp5ZbMb+iQB585x/KQjwbEjKJQcmgoTK57axXiPzitivhnyAtm3t5
e2QSus7Yb58jFPpK00AN/KTXCgwImwoV5nOstPZwYvUQ2eKaLGOY1jHfXRURtUcc
5OEc+N1b/KHFAE1aJMstGrwS6AEM90ZBLbdUL3LrYgdVLuy+F+nGYIYcWIxYmZSc
lzGJ1M3jT66wDq1quwEkEsziEcvfmEIQid1ofIKZgDxjVZcJUGB5VnfGyp753Jdj
jvvGTlnIM+ZMQ895LBZjOzV5l1tbM1qgJ3v+eA2p/fGRhRAJ5j1vrSFQGUowQJp6
Dr8yQnYpW3IWboK4qMl+yNLw5xmGOrilTqhnbCrNq1exFFyoll+bB4InnuxM/Kcw
1wPdpT0zuHJIp54klMeeDEzQX3es1jZNQ3w0aA1XCyP/jyMA8jJTRM1Cvz7tDGjX
CNwBVINv0TF5mIXMkK+v+JCBrZaZAVmwkOEcKJE8hH98/cqsg11OlLh5uE/ExMEG
Fhj2+JpJtSHUsaWNXalf82Oyk6TIZlVLwF1Eye2q7VOwDJGhdNSx3g7xTXIS9CjN
9uWdHUR4YFH2XBXySAkmIAvgS3GjNha1uqMEckVGOWdh+SibdfiNXiJZP9PN7YmI
J4JNvQHm9xerFFE0AOD6hqulAhLNu5O4/Ll4j3ZMmBetJ6AYs+HcoHT2kq6ITYjG
21p2Uw/aaWBlNkNuIXIvax5hm35XlWjyQv0V4ooKHfR+Pq9LD8i63WnyiYuAUaBV
JjPsQ8/sJlRPVLcOkWJ5mu5JRh2idNYM5MnyXlrF9PrA2Ar49CwSO7NfSQLJCXP1
HewjZAyK5PwPMn639A/vh6hu+YUCqEEGR7ZEpNlgX8ZTje8cypkZ6Wi6ghdTEk55
qkXcNV8dZTFAepiGd1v1TznEnvp8TLkglkB/3CR4VvQ9hdvb/B6yT8S0Q+PzDwb4
x1fOAGDbOwNST17pqJvpdiF3aYc4XMU+tVYahscLoBzmQUIOyHG99dD/GCmyr0YQ
XuEVCBMWWnC8+4T/Ikn+McRHCsoyL+XAdR/Arx/5dhDSvWryR8t9gh2V14o8jStu
Wbcv1lMLnL6Xb23QLqCew6++lpvGctVYfrC3/TxyqUrze2/4k7ffnYiIqSDR/XBG
ND3eBE2IEPIGvC5SbXo6Gq81NjlYhMRxPuiObnpBlKZNaSsE590IIOAfImQs3Fa7
tKXNhjKP0J+GOLe+It+sJWaiNGwum5KPNgx2/aJ899bnetmwFz7RNXTEBjCY/Mya
00qiXxwfHKkT4vX0SRy3opAparaUTy0ZYoe+BWcmuEecvZ3gRjk7pb9tdHM+wRuz
XoHnNjnSolJ183TC47ASFqoum9c+YPJhdbEmyVVZ9mP3Sv9JP24+0S563opmrkJG
2rJ0IloCHquMmfSACpBuTLIP6OkWd3v1fbpWzq43tLuss1idkRpjldktw9nqzeD+
pTyko1x0dtN6ideqG5Dj3NDwJWEXuCUtUqvTT1c8vJNJ/4AHGPXPt36ABhIDzgoo
7bBz8NLorj76kig+FeBdQkNMddDDz5oEuolHnlwIzIObJP+ajJREMgj2mdtFkJVG
yphIqfDlW8wfHAOX3tmPzobMibZq92mcgVy6JESlrsBHB+P93uHTsaGyl+8nTh7t
xkFmFI7T3+acpqYHAYD33RfDY5SGmbHmSs4Yl5Era4f4Kq/MioxkSCjRb5nnkauS
KPjonutRnaa84DYakc8Lh2zSBNir8Hg5alWJIRxDyyL95I2KV/OqQNPhztE0Qu6W
DN64vm409eTsp0CHnTOMvhtyjPRHaxXAs85qSe1j9QyU77T7gLwTEF794eWY5QDC
W4aIxBI1se9fItQJzO7R5OoIGs93IFA/102dPdXoS8t0xSzyXFnfwQoUILpL3G8D
B5q8NCe0H9fZUfYpvdKaWmFDM/xnznaACzKqFszfCEgPoo0cfYkVu+zhZMUsitgW
zz1A0vDbDD4y4AIddarQpTDvNTU+1bFzkBldCeo6dOl5baccn2LkkYrL18oVGImX
Z8LE2+k54wy848RqJab9utCWW2NzBPebIMG7gRffPPUKCCyTzS8nT9VutQJxo9cd
ozJbnT6H/kDqb51qn4XQTAM+wBppUdKRtepx5vFWOZYF4JUPhoZBZMTrtCtWr+Ks
oV2bkJ985wSyjM/2jJg0p5qW/AGpem9O7guo5hX2NTMNxmvzVl7R0YPBdYTRQItt
XpnWF6stgMF7tgi66Lu+INUaj8S9qaSSB6RB/jGySMZRBUDyBimMS19MSAvHe66h
AmTSB3+r5S8R2Cbhp4+deFpMK2MKRV4ZB75P2iLLp9aR02kLRLRj0OmCDoummoIK
Y/fHC8d+wOvpWJKapdQ7lb/GYy4V8PHYYKLtx+oNCQifIbo3u+CFxXUDZxkfaRpx
X5O7/Ir1/SoP8f5HOOuG2t6QKog9KX43QUcrNeJuGwlNzY8tOTNSHq16ASgn1tYC
oLOFfCWBVaxKcWoutZyHwKgJA/40Tv5OqqPu8W6YSZctcMAV8zwfrMZBbslzkTGt
jv0xzhH53heecHXZyQ0i3A91xpAFTjLu3osyMRJp3YLa3dk1f8TJz+jpXAqP1/Qt
7I+jGlmzvU8bs0Lkn1eYQ25tz1j0Tjepn7iyhVS/AKPjEfSsxuN/HLkkTANT5jMf
sDz2Z6aPIscwxO8XXjKuF3bdX9T0Y0LtDk9A3fXHPdfODrMWlpKIqsu5HPYTT9Qx
TSWUAEF9yA9VsTnziMggdjY6K0DQTY2A4YkNkBk39oBUZQidJ2Tlzttqfkt3y2/J
V4OyEX+yjDkrWu7grcluNwpA4OGmg1CMW9KieZz3UBK9SCufVA+jOEVc3vKJ/uSh
It4GCjC3gyLY/FBIJwcIAvbkPUNulx2/GI2hhuuc9vbWYMienROTuoiAQWVqp6U+
3huZl3SgkbXKvV3jQ4B+X/gPBmJW4rqiJmCshSDtqvQBTeBUBnlt8HMDCct/wwTI
f0shaTYVU3+LpmJH0kIkdcaoej3sslr7AENz7eV+ZRYTOJRA0ZViP4B+nSyCBTs6
i2FPBWKmXbo5jEUqJ9Rk97I+IqQsvJvby1wqxnuAGYgN4t+UQlz5jshBC3gc8ptf
Zfvtsapqr9lfWv4gQuh5sfGuyYSV+ImhXce0sSA5zVx+Fh3BFWteRRX58eCTRw5N
JeS00uhwR35zwgz0hSFGhMM5mY/pQch4dXyiGTKE59aR/m8mJJxQ9LOXHZL4oEp/
7x8E7il1bKefy66f5n2uVjJ0P0yvRwp4+UagyfJiaCsSrPJEUxW4J5ieCMN4fPNs
M8zwi0RpYqvJQLR3K1sDCJr98BHUL+3rAp1wBza6EInSToEvFqxscURLOvUFWLLh
v5Wo1NzykuaUrdJ7rOPe9vqkZAwMABz+McBhr+AtG1nocgm4GHWmcSYptiXEZZOl
716Qqnetd84vQZ8iJxLzQ9UtrAonVXUWOK9ZUbzQO33ZUouZolKxID4x+13DtEY1
HTbENxK+BrsruI8gtwnEWSAW5NVg1n6WTgOftKxFSoS2QPRqJSDFEbLr0A58HAZO
PCy2cd9Wiw4iioETy9/j+sfk1Vd2CFTq0AS1cIofEePq1CyjlF4K+1RTYXzslje0
W3MzxQOLLeZmhQkiL0w/FCl2yUAJr4xsPxk3KL1Y4fibhe3bj8yq3X5xf/hkmSck
8p8Q2BWxJosi4qUDGy6JRKOqqxmJNJW56i7/mLp+ohhvyG6iIV2pec8+siOInBpS
gzKQVEGxmxCytYKbqK/TcQpqLz42fedlVLDtXf+pH4DFp/NYabo9aFzWAnqYv634
ZOv+2fHe+nl5vuN1DNybuq4hyz9jLuR+UttxTj6QtqSglr22FI7AOnjnkuSPCzoi
p7UwmIA6xPJ5N7t38W/L6g68+H4UG49AE+12DcTwDCO/VlPwFm7oQSMUMWA/yNmx
BQ5NUJEjtemEixb5vok3+xTCcGcrC/KOiic9qgOkFRAMblxddhVzEjIKGkBXZdj/
1E/X1v2QPb8LCvPG1PD4FLcVfmBaGkD9uRmEoetNqXyw0mg38+fTf3uyQIYz8GMn
PUxruonhgljbXO8U5Lnne+EsR3SR/mAjMCGYJG0tiA+tLdu9Q7t0eOoms7R5yxyE
tp6HmjTo9eY7Lcvu9o/GR/oR6W+ZKN06nWUAB7du0sJEd5nq2Q+H5bezViCo/o0u
4Mm1TI6Avyt110yDTthkL/agZakLaGUpE5UHYvNzU5w4WaeFREX5wxOe89/es/JB
qp7Opsxvhx8TAEESVl++7x6hvLU0lwBa07Po7P5sIvtlzlJAwuWJrujKTEzbIvXL
l2OamquxWqfsfRogIcQ20s4tRuaJKRUCTcSBrbCOqn4nR/iO6JpEwIQfPhdFUMTr
cNOUpcWir0DueE0FDka8T2TncnW/+Sp1VPyAGICYpySVjqmXPDNatsV3KT/O5KI6
h7VTF8Mr8Uc/ci+80M7sr5Mvv5LMCurlN7nmZadfhlUK2nEeXPzcu7O6FvSCi76R
7681mNjP0TDRIUQ5/05nXsO4f2evWWBQL3g0UWvLfg6be8e8oNqJj/MSb38RgrBV
niay+lkwY3ftyeMWb+DHmqijZ51f0Og6Fm4KyP4VAoQFMFb6FCQiiSmNJQES4Uui
x5FT6nAS2aj7YzCflTtTSOffywCYKeYEQvOOfFBa2wYFrytuYnEGlCBzDRoWUy3p
q8NOJ1SRY50QQoIZcNnY7xzjWvIR6eA/d7CsEH1Mozckxgem2y42CDWdZX7q0adr
LBlXZbUUux/eHHN//4c135uMyXb9r8VU6yER5yqHNN8OjW1alHkrzxl/tQUrPkEf
wDHJ3wdcQ9RH46lD0YPLujWk35aDgAYC3yEx8s2U5nWIx2PDl2ZGzXcEPHHrqL3/
KWu0WIE3zsbGU6f3TpXTgqzr7uVdTG0MmcKFUA1dz/70lYkndcW5C8P+jkLUZw8y
TdqrmTvzyjWaons3VrEIITYTgI8vesp19d7Mn4BYE6+9TTs+7tf+3CLwAJI4ua8k
BKp0wrc1AewnZlTQ9xczQ3SNPADSqrfZJuxrVFw2YLOvET4mMcnJho+ms22pjbEJ
iO/aJlMGuC2L13atvmSPS6EoMYKSXSX8eZFJS8fw5tp4ATJAcT/+KhF0A3u5yuBT
OpbEh836+Fu6Qi8r+v+6DAKlnpjis/ZB2zlPsC4nBGTrlPj7VBLNRt9se/9geR1T
R+XYhgdcQcPX2Gc593jsRUDXdJ5tQXXNIgoL3u5bCJ8BW2dbQyXrcpfOQF9Si2SU
w+JNzylnKhvRQVdFY34e0Dc2YvaObuantlI9b0u0F8xLCkzPRWHaS/3hAyr1XOQT
SynbZyA8u963SPpeC+HOq/xHpX38N4u/vceRW2ztYqo9YEi8rJ5KYTLrJ/ljKzA8
K76t3yrjRn6IlpQsLQxYgP9BEssMrBdVz7MxlUPSOdF5ipqnffxruTvVlm4e8Emq
wwMZr8+sa2bK84jnBL76XSUHKsLtrpV7Vvjq6OBxiaaoZ0CaVWYbKvS3Ub/ImcjB
Ac6Zrcm5rLEy5V95buxX4mlUviuH08gWjKcTqH54mxhMb9sZCTDGTdVi1U8Qofdb
4kge8O9Jjdw7sT8BYEYTQpPCGkdFqEsQXENaB/d8XK+c6MaWPWNgp/LL0eyGXtCj
W4WOaMsPEloAMJ4hd860n0lqSeveElxMi3rrnNkLnhP6InKkluPBmR7o+XolZrkX
v9Nc2vHR9yyzvPNOvOGgaZ1j6EDkNtcLLG2f+XyO5S5o/GajjvFn98ib67B3v2FU
v4E9OM9/2wkCqtN8zf4CfuDIiBTaRfuSgzA4SpjTYKF2lVFsjpmnUh/zTaMekxzj
d5nEXwzPKxmrTW7TEodHw9HPzhSYLZq/EebTyhXPalmeBPK6PTjzosPLRF8N15Ja
0v8o/8wV3c7B2pdqlUncMYiE5USB/bPr3GlEKB2gafcb5Gc/fVC84Wxp9xrZeG7u
KHtFC3HD+VrydN8r04fjAdRg0vBIiRlB+a9AGBs4hVeYu8VIINgTMEDdnPulclB8
jWZs8dphDBrPn5hLcjaSCmYCM+HK5jggWlczWgKaBhyInBcyqQu35/VZxRR17dFl
JiI4ulODy61SmOeLoA8HIPpynO/14uxV5++dtm3W54dOFVePp3dn7xpSrguECdil
J4e92CWp2FlN+XXlZiYi+5p2ouTIAt0UZLzMFqefy83oz9D9HlIQMXKDwoI59OlU
JaiURoyuiL65azZ9CNprgtrD8dfY1zwt2NYGfcB1ADUCANwfLtUL6QJT2WtnTP8W
+DYL92DzIZOG9cJmpF3IvExFM5egdpYH6yiQxiW3G+DIeIkgw52HoZGgN9fEqal0
MmGGhQFfyhPRSjwqQC1if3j+62aJ6fRJGSZGxwT1q2SxWi205D0LiNM9H3/44iuo
Pjp6B7h9NRsFht+VfSpsF1Wmg3kAL98R1p4jgCsciwjQSSIS6m0aTqaEP2ZNYy5g
HzDTFvtcqYxRS74MWzw+j45z3EE3RJQEjeSvhgRHFOH4pNS8zqgkwx2P8V6k5KEv
WvWNqvTYL0jbNrbs8+L+wKfFefZAigEr6BBkCs3c9MUbPjFUelv7OWR4j26FtgbL
WE//LldzRMJDspMMc6x8yvNggHP1Gqmik5kWCE/2vYW6yVraEFuGYkFkg9/Z6MUO
B72zNsB/9FZZq0tiQ/J/6zkkrKoAtsgsyGhB1jNkT+5vhN6T5jcaHV9uFHAoxvPr
fCEBo+th+KusaRGNLVgLCoYMA3pNnYVRgVCtqzs7jWpmJseaH1gf6JeC0g3FeyOe
M5nZpKEYZhGm3DFspvJgG2T8zVURrNkYMEVvFYCiaDTkDRk+2d3SGnQ+fXNLmTpc
LYXsln5mPycRdjX1vodcOzJaBR7d2tant/AiP9/pD8NYs2nXpBQlqojghbNFJC6l
TbnQv3DjU02zvNLRuW1hvRq19AoRRn/PfeJBdxKzX6fPM1YArmeWzCvKFef+edvX
z+SO7J/ENLxFjJa1jg9SAQJhdWEo4/p/mLPnjjx9598dyYJh+chip7uXh4mQ6+v3
FhA7HEdLNMc9/gJ504u7IrTuo0gmBLFdbZFYyoHUKuW+6fH0PXtVvypIB03hFkAp
jTzaQ5a902t+C2b/4a63m4WYzH/4PYnCRaPGwifYOhQ3nPXssdNH37y/ANDUawXj
iahTUv8OhGOAEcSDXWciakA6bbxj1Wrs71bt2VAJGnSUtgYNDpTO3jLDapR18FDM
4ia02hQHs1uKRkLA97xvZNVciFxvaDJJA2lJd8jS/B58jgUEcUM/dhHMnhTzEbbk
rq+Ur0lHRyWJ7BGphu7J6uvCRlxKCZT29lM5P/zz4lTrdnaOmiUCgVmRXVtKMDwG
DBykxRIob++C5fN/uVMyroT5kM29Vbjyji8iicLvf0WlEZvx+C0xvJGcNHEQ4SeJ
zHld0zyngKBhmmN7CtNPZM3PU+t+2L4LGSANuE0jOV/3IFRVUbEMx0lrSwXrrbTR
l3y0yfAwjU4/oYoWl/Z9bEYxBA2ukcbbwwzjo+i4Oq8wtawN1lSVs1TMEREQcuYA
qw7vYirgRFF19NJwyp0Ha0ygetO67gtpYyUmBzwlQmmvDsnU3d7DccYzO7MP+vIL
g8VqOgorRhABvnCYcmXQPmQkgrCeMOIrRb9ggJzs28ClKiA7wCopV+TXrGrZyOhq
sAe+8wSpMPDvhzfoY5CZ0Pg7R/UEycb3DiJ8/xeLyCM2tHnTJN/X5aQC9N+mM8zR
58jSK2zaHpvNDbVDT84yQsqSslcl6xKMjFhqH5KXPXGlIts+1gCZWojn2OQBrPT8
pEUB+OvowNzZMW61kgfE5i9fLGEbOtnHjHHUEOM3+wt6mj9rSuOa0xIWu3gnYrtX
cD7XpAayACMlPaoBQshPPiydYoglFB2Q6mNlKv8z7aD1i9NOrX9FEbuRA1JsAe+h
Oe7HKpYqf8ZbdcRF3EdwNwvQyV/cdMdhk1rqsUd9AdAN/zeP/Veoe61tRv4ItrNG
QBj2sS4U+9VGYd8dKsuIEcPUY5qtI9CYQN8CH7ym8rXdcTwdy9DBduhyeRFW7F1E
k7KsAgAM10xw7WJCJOQE9wIZ2PpoUGhPy3VLz+jNCcb03mdtIfrN+cJeBzbCTBNx
Ng15KLbeC0Rc2bwx+zC5cDFI8qIc0MvSOoAWRcHHLn2zPbiBxudnhZD2CA7dSfP+
BjaRXJyToLn4gXVZ/ZyVLKrq5ZHWqKvsi/92DLJ6ksBzusa8bbV+PxWIXfyZOWV8
vywkWdL2eyjsdwcA43w2KizB+b2Feyx2xnLWZCz/i5TeI8grTASm5ltLgrJM1QjA
cjuEBtGom7ovQHza6vj5aW1pON7qkeHM2lBp7vTRHex1afqjjaMiLmBVPg9RTlPd
lFEUy6UqzPjg/vrWiZQ5y3HYkXGDrWFrIZj9wSNXGQNzQvMd99MLUDGlOoz7whtk
FoKh1V6l8KEky5JQdBL/YTplfADXuzFBxArgcUR+q2cDSX6OYa0LNMGZ0KdBUztL
DYh1LSmEPKqw3yNTDhwea9KqD3KdQQUufGrMpB0T4jyVqA2dtenCb0kzHWcLAPfR
Jku5Vha6R8NMDSC3RQSDjwkbidOm/nsA/98mEu2eN5LuAZn7s1v8eIcWbwu2SlL1
Laq3NM4moPGMZXhK7w7YtoLUlQdsc+VqIAtl3iIIiHWld8yp9R8CwuxySYS6hw+O
7N7RGj62D4AFDrNtlq6aCYb3JuEYYJgf19RgIIlvp0ueqPovewAJhLc95AtdgTQr
f6ADJ4X8TQxmtB6dsZGmqeyCdCkwDKCLZAdQGnisryaRbAsesU5gQZZy88qJt9tm
lonUYmbBuvNrWqHyvnKqCaz9RtTa+tRYvTXZPNqpZPuTrV1GDExnqyXZoJgZKuFA
Q9D4/XnC8AesgwQFr69b22WbyWO3YDaR8pCKGBCo2U2pkR1ESevZCwmbmbGY6/hX
PzWOyJuYVs5cJpNoX/YcDUFF8/0KiTDH7Oehq2eIoEw49wfYJBlityF2oEHDa/0q
EB1f50jDlBYvZGC1tjJ45AWma+phF18Tr8OtQbsM2333NcJp1DWNFQ8nVcbOPvEt
oNJ2anwQoslCDDdBtNe7v1r8jjyKKGnXxDgLgscMscQOgvRPieu/leCNqwaPIykH
8/Y1lLEDqMC+QeQ8XtOp69RAP4kSugoYjnfz105p3GWhJwDHJqN0sosQ4xHFo9QP
B+EMjWAS7rZtRTJuXzYppYsAPnZD4VoYTMDhfg1H/64yyVxfBvHp+KpBc65CIcPu
nvrEtqgwlhjWTh+y1ZUbtUv6CRSrrRXtRdSxf5DL2aDJstIF3UEJpy+qYlT/Aduu
yhj40SNVM5T5/EsjsyK/iFVMokYfBQpHewqbbXHoAS+/O5gVs+WtwaC78vKPAdGb
YxhcgkdBU+zB2jP457Ujqf0SFRkUNZZy/Gnp9LKa2B2Hk59qW0Am8w8kriEpQr5L
EE7IUglMUq3YJeZGHhw5tgKEDdGOIMdv556SjmV5cOu9iDVSPXP7t1RHw1ie4fCe
a4l4o5RlW7uHfT+SHJZXco9ZNTYJtRooNn2pkFKdSyKXjx5hCQdHNyGxBcbhktpF
JzqwIEIyMK9IlbPL+sczPYFC82XAvr1nYaBuxBknANLabOmlIwTHpO+szfcYCewV
p++tXQ21y2rmKADsfEtyaTgAAQH/JXmdmqBzjwXXwD2o8DHyHbrmLeDo+U6ztOTP
H3G68B6AVvM5XdugNEcrXHTTOtBDwudNiUMbwxUOb8rpELzLDxOoDYskpdQDxykw
0MgzXpLwHwCK4Ui20omQkp4CDxnYO9oGJ3NlhjvKyyGTGjgZAOtLk4S2H75bd+Nn
2BOl5ZoqAiCfN+rvWKGuBUQmKXQBDLOJMgT3gz7A0sMLQeYBJdYx+NZexefCy5ss
wSOLz8r7dAg7ms0XffspdyRGlvrBSDb1nzrr4C6ODEChwki3NvBloR0C4ZiBc4Bg
mAMpKzZ1nDE0XAvXiSaD/kI0LtP0EcG/ljQffIpNELuX3u3Yw4sF9A4NkrYhpn7C
udMBk48rj7Rlhh/i+lhhDA84qS2Zly3vxnsCT4pxOqt98teZtWB6nSOgI7Bsubv/
Y8p+cKSjnKunaF3bY//xpDM4hKtul5hbNprXBSzN2ZKxZIh6vMxpuAHpX5Gs0N4V
Dngt8ca8TvPb0OFpglU9bBPF6qFEBUShXe1lluQ9G1Dyh9TwOJ7dPKd0RDuUNuEX
ApwqMXblKdloRszeSOzMI1YtVunHJKw86Z1UULQZHOncXXQx++vPYhs8As27ffSI
lSoIkhlyKx0v5v4nz3j5hD+pSwTUT/jBM+gZSMV8OZ1j8P4QoG122N5cdIc6jeGc
cBFFFzJ67rTLmR1zZV9ORE/3qYnnuQOEUjl+Y3VdF8d0j5lgLdWkYsQuRWeoEbtg
ZAKHhh2XFzZLqPRsHHOygME1Yqik5ELg4LSqBlenHkMqGWjav/fxXGH7pI1aPVFJ
IJi96g/jTdfoMd/jfckU6f9JHORl9g5ASfxvBK0668j7cP403NPPnQ+nuRsvhO6j
8c+POADAhmJ98w8fV63k3G3n8wVqIUl+UjdI8/peIh/MlMYEm3w6tF3PlScy3ckG
T55rYc/42GLFFxfKpuNobU1FaQPyFOke295f1Z3F99A1KDKU2Zo5leAf9ZWjvEMH
0x1L86jY51rcUbOHhgCOhiRUluAG2LXSZyOZxitHbM6YLOMGXO5fK0GIxqXl3fDW
HJLSLQeZxWyHmBvhKNKCWGSJalJLAPFvRpomm09f7LgZVr72dL8cVVL1hc3kxCOZ
BfLML6R5dbZxDSjNX3PF3+OjbOJ9RyYZPR/C0KZBfiYXMGXugLSxqzYWP+xSW/rB
sklQcYWGB6mxRt2tOsAeHJ+K+ca8eByazJ3VHxVdLXJzSDMzNevdeQRGq/TxJGRB
han+goe1miJfve1TFOLwHeklqFdKq/p42960gkX/5AYoDPxUB/D1XGKinfWsLZxc
yIPmEanzqY/ZPEcCA7tzBdThRNpaVDRZv8njx/0247FOcjD9+t2ow5YgJ9zRdbbi
S3Jej02Pl4PMWC4S+gaYiLRzv1VruaJpIE1Fa4Cbhme8QsDxC2lPWy3s9zB7mpoM
kjyfNq2q4qZLqXeQN8x1PzPShYHMckhCZaYbXpBtxdbCco5UR9mLeB1aHoS47I+/
wk9eksM3jki16GTau8Ctzy7ziQSXFqBPMYuHV9e9p81yM0Tf74pPTnEd6KXv5Aj4
TzfpkWsbzTdEzOTEZ4+1uoMp5eIQOaHar7kX6ZNFmW43xcDVjTtoApr+RAO4LAig
PAxcy4UbKmzI801i5+jITJC00AsZk0FCx+hL2SnwWFFGdHbdTOPfjc+otIHAPHXW
O4xOGkgOI3QADo6x+Evwcknai/rm5nzzR6SzYyZ3do9s3bAqTn7b/+wXsrsUw87h
uhguMigkyfIC/cZutDCuTDQr9rk5FuqKBBgbDb+IsXoaWlFle8CXvvuXRG9R/84E
tdtNm+JBNbMrUZu1m+2bcWflm1zTYD6c7ZqMvkpRG0VSI1OhOQLXK/dnEhOmkZSb
StQgLkz+Pvsihy0yWlQMpaZ5tUs+k4BX8Eu5AeZFEx3qLMXzMbVKvniJgUxlokB8
+lan5rQud96Xs+DSnPY9fZslrYmwqvQKAUWhpFfzk1tiWpItmsYWOh+KCFoLaKor
6vg9p9A/l/L9H3zLbbw0JIXELQ3TTI33alhn+D7zvvHxqkPSkaiMGINRvQfQoyJG
kWoJ9CuA2Z61Obi6akwsuBlMWNkYY5+1Aw98tCqVw6uK0yN7GOuxqL+Ng978WCoC
w2WqW0M02j7cq8Bjrfwrn4VtjOKxqtl72r5mDneK4iYeteCSvw2MPS9+3w7DQi7w
crV90oXe+y5XMqQ8zFhGeXf16IZiJamAJHJUpIU34TKaNTerVDW+s9tIoGUizT1x
xJ/qpCDBRToVlyE0Z+WvvYxWzC0H5zPT6yXBPdT9iDjpjeYgoHSDo2OPbfyf36M6
uL2EsxfUYq5YTydfqEO+cm3sBi8wixwtdXoaH+RveT5zHbwfWHwtZMPOE2W5Uw0/
Prh3Cyi4fttVMI3tTJVkR/YVsjcFkmYLUSbOW7GLGn5EglbSL/lOPMl2KcY/01HM
7I0qkOl2AHOHh51ZjWgetmD+EaU06mS4Dn14WD3nblCOd3FubVuL2XQXZLqSaNoM
jTNm7pIFvX5uVTyRestiJkSm+OZBgvq8yfn0Wd8LGffLDf+jV3rTPk+DPWPFOfjp
h9WDO3IPBhY2y+fOXY+g4S1vLvASXwveekJe0gCuAr51kO+ulksdaQuJ1RNplmej
s9mQE87t0Y2PcOJkqbWUqNSsM6Nsguoi5cQ+ptsDFnaybpx241kvCNuV6YrUvOQG
gCFUgzqmAkQ4D5s4E9yGmw1K4sWEBeprRu/COXm3bXvmWAyLvKhwm5yLVmOUX8HX
ZJTrvjjGUP8vkwSv65+YvxP/eYiqVUNR3vkWiAjNbixU3KpRO2AiD9bYAZo9VYgM
W27JCJeacJfMy9GA2RAbn6sVhNZcbh6yKmWFpFs9LPDR/8YdSr8lwQB74rX1vw44
98f6HMtm0EMA6uBHSRWtm6mIkSqO9mvn1MrHsfwbFl35MdOcTwUViLGP8GqS+8oN
6F4hIr2YEgwGewOP+l9Gdt444dM9QI6Zcf0z6vFxBkakpd7/IndrY/vT5f3iaeYW
PHWAzC/cYyOB2EQLjjO56Te1/mXZtMRwaqPqVcIPmaTdBa3ebKzUpTgz24H4Js/e
xDGxa/0mOrxL3iKfA3JDobec92aQz0Ukd48uwhPuBuwm9liPV3gYQ/vWZ5s/bCIm
x5SxOlY8x3sVy7PAkI/K/Jnjcvrj50RTbyrJ8Cqdcb4xrHdc4A3WoM1RjRf1D/4N
s10WNvQgx8LQEYXV7vYMBFFKMtAvjABi+H1RBh3HhW6n3crskNYnYDbI6cdAFr9w
MH/N8y55WZ4w74wtp4x/pHGGQY4wEPxZG4M6aFLzWCaadYL+bU+o0Li5Nc34oC0P
VZzvKW27HNd89146oB5ysQFdXFNXZbDmOdhYhxZuRdKq9WfvDKXEyc5VffxFGyem
HQ+DSf4fVYipdP/FYXbvUpKmlHTy6r0l2IkP06Uk+Fgxzdx3gC1otrId2DPrRGMH
wuz7cKIHeRCM5uMr85FbTJx/fFDeqWyOYwE3KxEA17Eq+k84wNLdAqVMJGuNpbfj
/qUslsoMF0lTP4vKRrxiGdpv1yq5NxxM+k9DzzByBIX9B8qqedl2fKR/9dskg/0h
PwI3rXjDuzyMsQn2w9kaYDnf4L/t4/+muGfL8ROJfZZJp0IG0kKCqKhrHfepNbox
OiFcO4MIZTC9CJ5/jP8fDQdBDhozlSDtrpyFx2Ke9JMpKvlXl9r/qwBUjr2qGl9R
5Ck5yZCBhnBjbSFRMMJNafQZTHtRaRk/6eek8msQHJh7gIjd3WZ6iXqwNFRJjFk1
nx3H9MbQumcOnYYYUV/8S/vRxZVGI2unt5qI190yEI1IVD1IOfur/ibufZ8AiqtT
yv1UmY8Pa7p8ReofB81hYHDdZXte+xTbjsvCAub4mSgZFs7jqkREndkCL66DK2r+
6ogDEpLBSM+ho71v7cl+c7joCncKrlNhfOs/jGP2NT9RwvNYiLtc647Pke3DTxnn
f8ZdQeUE7usrEpLpYICFuOjj4bLv5iiaNR5878P79DiQQGB4Q+I6ZMHHvCqQH6id
u8WHWFBFrALEa/0Ty7DTSxrDanPxYly7Qojy1ltig0+MACrpd5ivknkKzYv1/11c
NXOr9TCbCIhPa40HYf8gyIvpVsEq9TYNq0homuu0jPbUAYj61Fb7obWpsp44ruVF
qp9j2LJCjsHG6ZH3T5oDoCtOdX+zL63O/YdWQcBjkgQi9y+C+fsiZ8SyHTnT+Fr0
ypjlywJuOKiwo27ss3Znj1gYj6NDyMV0KEfpLuzWf+eqyfDWzwa9Oh5EhwPxjFBP
BZZ1xKhFD1XHQRPnCDa5Cf1Bg2UB+NeMjhZd84pRnSwDeyYh0Ks9aLcTZkvoQLxo
2gJgd4bLbZzJ5XM425u+aPva7XPdZwQlzksHiFLzGyGvQX0ulQWV7KoHnVm7pc5s
1eY6mU7Y9dME5ETcB0ufEtwnvYv29P854TrywAr6uGhQd1dpqtN3t4HkKELMOzfV
Ec7TK/suF5714AEOEGYEbcADtGTo4N4fkyFB+34ZgedOvgYf3judnWdyXV5MoEYt
yrgTKHRIwpRCwmbuTH5zMPUsDDn84bu543+UU0d/3ULmVLBGWZXh89lzIqiQHjfh
Z9DSsded3UMgyMW287X089de7sqBmuYyT/VT7pbHzwXpRuAv/S21LtHd1MzfSRoJ
zesQoS55RhFhZloN/ZFlyQq4V6IDEP7/n9zHavZX3p1rc2tJ3sazABW3yY9aX2BO
ngvON0gznEOt+9+CCWUtM4dqg26bsQ1N2tLifJ12PU6qfS5wzZnLTI8a7/hiH9M9
HAakNvqNpzsopXhSz5uZAkVbRMcXbT7hGDi4+HnkKh2/ypQrd0+nHEUJ0kHPs/M5
y5ayiHFj/GogNQGo3RfYy7Bejw6JSdCKKOwtdYiOCWy+dt7s0uQHaVcoo0tcAb7z
pBN+VyMc/wxi1msAObaP3of6KowMngWnWZk/3in1hRA3D14cXnbb8ufzPawcmKmx
7xbu7dhrj0YmraKVsLfBrnTUCM6NDiPBfKOCgnrMfIDXLh0kRSe/T9MjTWyDoQfm
HVJn5zlMM0bD2mhiYWaSvT/Ldbmsm6SdiYWYvvj5PMcutkJlFcFs+3mVCGREsJAW
UhVEOT0PLjcAb6AQv8WNoxtZB6Uevw+N0ywwLkK1imU3ZWRDI3kggxuNCICJKcVO
Y9l06EY5Fwf3/Jr8n7cKsXE7tP7BazJbXxVwI/wuYUdnJ96Zc868K4UpGIq+mQsx
6ZKUQjmH8NQ9C7nxF61BRSqdGrVKxiLyCtaae4R1sw/e6XhWPP1RcOGH70dXKOfQ
aWFaFuStz7w/qkvp7opTIxzs7TD7WLQMqi29/uSvUY32MVPDSqUZ5Rx7nheYGtTf
JWVWAz8WbfoMnfTStnjwfAZ3lTV/AIsqJms7W5OGYIASM7hao/JKMh0pkaMBg1oH
bZbxtws/IbHgfwlxvmjI7zcjsKhFKgLDyCLvC0VH4fLvSbnbN69+EzT8ZWAQLQhT
Q52yzahhgm/MqOgzaDsZo/0HFt1u/WJP1PSvVQVucZUeN1zrLLsZshIwWn8QdIVj
sHtaiZWV5vK53fdOdgM018g3V5Vldx/yaKfQpS5z4ZvyJjlMhuQfNfXZsRHk+YiW
pSZUqmJgKHVSCjGcmh9vWKkkEwQmX0jiTvLcb/fWxLwqZwzVWjdTOJ0pIqc6rzJB
i/pOMGt42UYl4FbEvE7n9+IBUd191nVRLNdqGt0kEEl3h8pdOtimKV0MHDkFVQwN
aE8RQCbClWRj4S742GJ05xxsGRwgZZETAPlBRBTTjwaKUEsi64lcWqEeH4vBJE2Q
iDVAjn0qQaNBt2miw2E/9IfdXLRM4YYWAPTGk3aAzy84uYdx6U8n/X71ZW3irT0E
6qIIapg5eH3c5TZq57Ex5LJJVnRY0IsebdOIriqtRHqv9EJ5oiOAXv/J3pxIZu4Z
0duW9jbAa2NMXTP8nduGF74iJmQDmHQRBY4bEr/mMCvvzd00eDTCdZ7en3Twht7j
4iS1tG4YPU9WPnN97llJyZj1fnxca+GhrMOqbX7irpEYy70IFs/DbGPaTKsim8XE
qCKVSWlyG8D24goPWEfT3yGlYaO3LJhucyf7W4ilOC0qJe4a4oqNxcyBhe477PgJ
pUJv308vucByu2khj1ZZpMdi3jPjkXInrfKBGcCm0dP1oP9EP3f+OqoUg7AsS2Sh
xKXiIDKVmrtwRxK3PZ4c/b3E9L5EBsbfrAcRhtblXJcW3rwQDfmnLklmYw+p++dm
l6D7fTKnuyBphAnlaweQRXmnS94K4uB3tFSN79P/lsb+Z8FMEpXkuVRT0XrEyzoL
OCYKN81T8X3/iUWcqkeu8ReXj2+xObkNNTsNkHdklHiIYi5iBDLwRdjtFGX/irDL
TCw6xVxUzWe5TvbyaHec7GQ2eorLFHTI91CpThFUZsLAryg11DQO9UglMI/DB/xS
owTyZyPx2l9BOSApreeWFDSLPXI9ynbRS1fk594ycA5jn6P6g6hkBH38VwOrCdBN
u8TVXQudJbVjEnDliaS/sU/o9LupiYz3QO6A6qcqReBxsOZLAuHzVIdRorbjjTbo
eUyZ1cjC/mAgMuRR6aO0FfLOn0XSPmrgwKTvNL5CMRhl2exnA8c6RlxivWCiTwlZ
SC9j8hQFP7Qt2i1DiX1aJHN1BPsr9xmnbxAKmfCVt0S6U3u9GbydYCDBDUPvempy
dYxi56CF7c8S9sRGgV/QS/YH+446gUvliGkzG7ty4RhsO2ZttOLQC1lZLPSWDNkS
ju/od5McXTKC+m+cC5KLmAYS1fGT+ICj5q3rCAS1SBspbaSCqfYKFMrAwJYks0ac
K7EkGsCHOYcPhLbjqSdvIcmDPbTnYFVKGGfbFzGTrdWjqjD2RjMOiq/gju4VTm0q
I+5/IdFuEHDT0eWCbk1qRrh0yOYuRT4ScgnRzTeKIarK8kBJm8g22YPD/Yk/LJh9
8QZn42mrDY/CbxAYK/T9G1jyLrRj0EwpQJ99Csg0fnm2WO80jnpHS7+4PpyfGGMm
K4E1fjmf6YWmfIlQxWK3eSIHaAG86MPIOqemPvOjudAYXPcjudOjNVxwnABUfs0t
dSSWmgIH3jrnGjacZRgSzVEk1uTQjdCma5fxtB96SoJtMmL3RQ1aUcSvOw7i6p7m
pq8i16aFe7YFiVSUCyBpWumFqX2o99wCRI79TKeUBB8TobzEO4AFmcCtd1Gz4QFz
Jqc7stJtpVqxcuoStCuTq2SXJPEdDugiabxBRMgN/G1CbDx3fkwC3dOIKuAWSFo3
vO3i58bJF4hjVG3p31FNnb4TkSSljzLhDWGmTKnLZDTVxfqdKLKVY4Ij6y6+syVG
p4uVNgozDLAYx7fjZvB+s2aBHamj3mcakVK2ldIXGpAEejWO52F18bazVboWUB44
qQTk3t9thd+830QggvXs+LXf+BUGT3pjeq3pgp9NSkbjiPv/HkYcephGautpevVY
m9UCaCILS7sxTS9t7KHLMuQgoh4SCTUCeDGpsBFo/xxnMOIEJtrjuXtvPSTuRhE/
xZreBqo6HO9Mkd7m4PDdaq6Ey+3OXrA6Hg8Tu9LxT/hKvcn9BNhXS136SrCH67AJ
iOgAdHC5hsuUFy1rbTmHISo+QdBklTeKM6+LTndBEOkgeLBTaVxlSP0gpShODznB
nYbWmN4lbCff3J9UZpdaq5L1HlY4v5VefQf/ntcbEEfCJiKWgE12AbNGzZzD0f+H
w8ZMMRiy6St6JwWSg0u8anb/htLTBbAKuMfy0LqxLVvc85UnD5eCoHA0rNJxn8El
2sPgRKywpoaV0Wgwhp/jOSBRLrKiXudv80RsNS8eG7x+XVz56bgfVv2aye2cqead
TVc9QfS24gCRM1R2Kskz2S0ah2CaYkdDdoIC3M+uVd7AplER6q5DNKhJMmswH4fa
mge7eaaklijx8uBY+EU4oUeGCxHGd68VJ1oTdNJdxHiLVCHsId5VN3S7847R3WaV
u9vEl4JiuJeHvDnoTcZc6S5NES3hQ1mAjbhLUkPALVPaQ9OSxsM49DPCIUnvq7lu
HRiBT+kawe9+M4x3G73J6xbJk2bznBkzesDinGO1iuUHbR+d7S9w02qhAprLv+Uh
nI4HyRyvqw76j7wjB0YkSQFdtEghPiG9oPfrSkld/KH3m05ZwPoOuXyvbOVipmlB
y+Hjmrz2pTVpLOs+Zbqx5qxplr7BxDyvWsstqIs2RZ8O8wPpD684usgFTTMriIG5
h4CV9jWsACxBPxp/zVCdrM1oEi1Mw1sOEUOWmA59Xxd1ZzPM7No1vbVg7JPGA4Tp
Qc9vNQpPiIBlR2dd336S1KT13FRovpY91YkwJmIQmhXFHcfuijhg8/1mwZFQi1xD
4yMujnKVRBv6CUYda/9DEI8d9/EfsfzLfaXxVBqkjszVFpL32tQ02BYRu4kY5xln
kW+bZdcJuRgVuQ39jr56VMrEMhGYGAHuNgr20sYQK1yzGx9zSSCCjwbTbBzLxTdN
7fFd7LVUfwDsjh8CrCTLEDapubeh/za1sZ4Yt4ltrrfiuKUSKZ5vceDZl/CV5LJv
CYiwiUnBVYf4Vm5H/LisSkJIoHJgHe8HaQe203KSoE/AnmYxspPA/TTqKdWmu3qj
nDqtUEv6h+jyuAKNhfcS5pl3oOEv9D2xpfxKLmyB0AgCADuY7TakpXAS9WJd3qbt
QX5mXAvKGI04a8hDRwrDRb/W3Y9bCWqYHEUQepwjNRaMgulobWgxSYtZHRYVuoBQ
H+V77lAr2sChuuaboHZ6UfgAESlZuXn0oUFovgXUxhdok/ACXNZ0ll9ZVJKnYwVv
UFaZjvHIGqZ+o2mqgCT08k217JeYMY1m4xE+mKZIOU3qRuOITNQqHk+FhNGdnK4B
wudOsRXAV+NdfSLIKtI26O1ejMInTlVLs2HD80hA0OP2NDGlHsrW/6KG+CGQDhRr
7Ekq+XpsIYGn+YH1Gf9WPiganLMeZXMZTFHd3LHEo5CwC0BpOkOU7GNiTkQc+8h2
vsMNSY9XEvjR2KbPMPJHLEQpkl5h8Tr1w4bPk8gNK+G5d3tSRYxRXIuRhRAgXQnE
No2WhHbhL8OYqDdYfRJls3QJ885bksbZSKiYL4DE7jcucDTkzV9dG9e/vUnBYQow
xmuWhcijp+NH9nCA99Hwp2axH8JxhzLxWYq0sSXifCQOKH5i1822q2NUE254iRXi
pzBKhth5cmbtJ8aesABXHuN+JwZ9/oJaRYRK7kEu4NrQGgumqTA8CmlkxExiXtXA
F5V/mllEENO6C4T1UXcmP3/6FANoJ9Wy4JH0EeaJCA6TCTBlk1b+aXeDFgecrw6C
OEcZYHtbYXvfyg4YstTQHy2/VwrI07hsNK0Qx1C6NHkdm0nSAiyexgwfkQXnfjwh
wMMgxaYM9CMWzYWdMG3+rbPlL+uaIielE6KVEGGtnQQqQpndHAs4wiXL9ak4BfSa
HU0m4RymjjsPaFnm9JYqUpn/ra8dPi87jL5CH1ywY6IuSZ6JV/I9V6GnKYWIkh+l
OtVvXOttfRLLnFMF7VYf1s3il7G3uWM7lWtN+ht4V6bi53byGiHov/vtt87JIk48
QbFiscsOvy+UQFTUTe1JOapDr7BM99OTSMzvP4+jctanxHiAtYCrNNNRGJ3SzkCL
SNLjQVafa19OUIiwtngKA563Z3G8hjFt2HXPAu0R46tVrMvpuLDpUISZx8rESAqJ
JZyNIWCRQVs8M39l3LCvmw991KZEX4uY2cu4phBSAwzDlsH0bk0137anW4LNIjOk
Keh63egB63CWoP2O3NFgce4dgsL73WQOGHuHcLG1CxwDg5fqVZPHsZ0hz1fqW09C
nzfCS6i9JngLmT05lHkaa4DAAtuDucbkdrqhNgkUBX574pBTnrmWojdAFLeQWUDQ
XcoQFY68wAul14bu+iaCq/Q6Cc3QN2mBGG73/I1bkzukyAitON1UpvfHqha2J9BO
YX8qUTwnPaIKSzWp29N3YEHWwPwQwAlghwdUq+Y0HJKZyMsrLiT+6qEl85PIpVLY
Ukn9Z2AqklYmIkRUMfK2Mgyl4qDWIMBuxmEkT8Svq3+XirMqL+MeANND6W/3teqj
WRVDRHtr3Zw0HdGfjXxicgiVtb2kPeGf7l4h4YIcRdUUJGSsqMI1/qVTgfDogodJ
SedKQ9NJmNgfjQPA454SZYgUZ5HuCysHT/lrCL1X+cLqAkHpFpM5PWcTO2SuTgRI
E+iCUly+hMzNqrN8OVUnh/dgujmGh9HowPSAAjMRlnvvnmtAaWHQ5RJpElzo+7hn
ZsK26Nfb/3G2Kv11HIa/tk0Z9om8sjbf3oOz87l1aaVYXniLWrfUOWVTnoD8WcAS
tP+nulj8gNuKs73W2FpJ7fdsKhogLJFAQMu041fJU/Qx1MdUlzl/KTklj3irWS1U
pKoaOSip0SdFSGpgSp+2upAMu8nx+iWchvCED3T0rxfyH8JMCQJrSaV1HMd1QOIv
knwn1JEmoT5JAswSnXGqA1KisCMf15CtAuc0ARFzFXDA/DZ8EItYMAWy1Jo4xByS
OTAfKlkuXplAECJ6wRCsXLrC4gCtNNSZ8CdpmPBVPXkGAljqGOHqSGkRUBZS+kdu
+3kg/OyASb1mN972jIkeuoE75GEiw6knbk7O5mgUNxUPzPx2kImWuT2S1qNx6yh2
2L0uZ09wxwie+yJ3RVqPMP6IykjNteAbzMK04m2DISqe0pp/hVPtFYb8S6A6/KqJ
BQ3Ab5iwM5EcYukdhtWv0uH+1QEFoaOdgzXe+3AbbWPtISz7UJz1lxMY6sbF8myP
z99mNSZbgdesqezhRUjrEI49X/c79ubfsZ9gDBJPG3NljcpLZyD5yhxDWV3i55Gr
zVLcuh+70KBV94Oc2fzYj15u98nPMFF0jmDd8Kvx9heKUB/ZNPyn5wNFyJI1Kx5f
vVbx1lxsA8AE6cDCW8I9hz/p+XGLYmIUl6hB1+ggva034dJpo8PtxuYlKrTUmdBp
WMKJI0Sf9vrRjKiInaxkbAg/mGdqmfEjqPzPiQ8JOVdqJVFVKHDaoIhpZKm51QWq
nrkgYT8UyrZvZ6R45RG552IlOqmL1Gl8yCGzCBD9m2PpWvD0iyrzM/1Hf4vhAt4n
S9ChiJHibf5WwCDD1R2fYTMagvA0KZq3SM3gYpcZOVSeooM/bbxvU6Zb9iLer50R
0DhwCi/UKhMiGI9ZAxYWbdQsP9jDbSst2eyq+8BgrssZ9GbWZqlwobvhC8zCYQlg
26qF35ADKjYrkqNV1YvPcY775/hu/fbhHnf5B5LnhZ6Sev1VREA7uOmOesJRzR45
QERjY3xdGfY0YmpLL2NwQVJs8mO7CmG9J6T21ScmdrhB/tz5yztJ0qn/nmxWmDsT
lp6xTp2MNxK2o2HRQ51YrIV/um/LoPPbkfuNtZIzw05n9/MXkkNrXoYEnoGBuNsi
NBX9nStNGAyUaCeN1LIG7YQEwC+sO+etTvwb1RZnjvPK621EyNSbuJWJUW4sp/5G
Aatpb2tPSVtuKuM2K5PoiJyxIc7KQuGaLzVmVGvOLzTaPWiInoYPs1zm1oA6LNXj
CDczV3rIkhjGvZLM0Nh9X83/gKbUut+x/CtBBwjySNydafOXvmfPVcU4mx5C3gRX
A3xdxZZQviyT1Ij+kCp8rw9MqAH9mJSSLbGcbjRl11q62vA8nt7g0ZYpj3SxZyp9
Zz8liI8ZDK30ULSngX+OBp6Ue9dQ+1oyInLHT8c5gweCrBI4XEjjbZeaoCz1tiGU
RPjYTZ+pQRTHsae6xAJKsz6iHZM3sTRd3Zas8wjYVwnQsXEcuYpyF58TRpwiYViL
kXpwa3hwsM/fD8nQDVOKHvzNdESEtx2JAp70mH0jIyiLdJ9hn2cOCUF7trFTKpFF
UaEzR4jKx/6tmUBnLjwRvPzxXynGa3IOlLRBjlydwR42wUUDADHRD0KzNTRe28F8
dXRd6AjHglefScDaIGVz4ByfAVJLqWMCzuxbSaAgaXySCfMaBv9qbgVKjrOxCvNm
kTF9eg+OjnO/H00IxX789QhkBY2lbgHhFip3Dqb56lm0bngolLr7zU8jZKm8wUK/
USTHCzB8wUYKv1l02U2ZRptDHzFzlsk8SvYf8J1COd70y6tC36Ppd47gcJWzTlb6
ixL8qCYuaCj8D+8c4CJyHmWmRWG4oACA25OMrZLS9KjZch8ifw2WvpditWxjSNQ2
rUVWL4pNDup8vOHzxDihEYi6Vy9j8VKtyoKQKD7oyj/NVmtukFSfi+2XPkvaI5jU
BrlcSNmjFiGPZ3oHPpoQWsF2Gn738Mwoj92hkoAo7xQA9tOHErogk4gWORK93idV
uiLd6cFG0rcUXYiwUcP/H6V17DM/LOj49XBx60jGvxSnRdDs7SKl2BWeSPCzaA8J
QeNoX5VwMwQX6yQYNhfaFA9ELvd6CQUw5F5kKYMI6Ad13spHsST+Lmdugj9XzBot
ZiZFHTTf2yRYZgm8zNBsGzsR+77D7SP70ihNzbgzdowjRVxw8QO537zNdme9HOgT
G2HlmXhf2h9J7SmWz+MGavhpMwkUzfy0Aqt146vCgG+sDW5oTIZN+D1WdidtpqFy
NsJVYicQXPiXrw0AHZqRYSQHcop2RyQZ9ybphlgLrbeqZWb7l+kpZKSGdCcWwbpy
nCo/8z22RVPeREER//s5l0SBYy/KPCnC3TvSVly353+bnu8Km1fdCIFtYFdyjmrt
M6Oz9BwHyz9R3xbaoF7UF1+q99mW+um0+Vq/CdWfjyEMXY6LHc3QDG31UiU217oM
GHFbrI/Xs3/NIoL48lUvbKb59saAX2f1T+enksYy8NZs2k9Y3YoUN5GfdrBJ/3wp
bj8C3UokxYOKuuzwUqKnLXAYL1WhPorzrQcMhwjywbSraV0gYMrGutP+Cf2lCa18
AyUdPtb/iyGMhUfXE2LJsnt2JKIIEJmPqvw6l3kP6IWrZaKGdZ1meUhXmi28sfaO
eIZlm9NLVOVMfaWr0GJr5kAvrpgNpPnKS/H/O1yf+LRR/Y+h6h55RkmxowdcFeVS
JB3Ke6FswS0mw80qKFHh8DNCHLDHpxYX0QXyTW0L1svHeDKOCKKJmrjFRwQR6fjE
ESzyeM966gl9nE2TQAoSh6CHLZBR7CepZ7Fq6ZdbeoZjYWuc7IfSJE8bQu/3EQE0
mAEeXKMEuUbSlkxudjAylTJ6FDJgbFgTSLEqSpPg6xgvVtwL+0Ooy8Y66D7E/tqI
gQvYhtK12pr27Iezn/MbZ10dCNEgO2I2Db8wU++f4wyG4RROePnizBsY2CLobrpQ
TqOGKdv1OCcMTgpfE5SLyviKsYfsfW3zG6oxGOQ6qO6hblE3FC0Jxhia5gIR2uZ2
kl6ZnpiG/6S7xraUJ2O4JxCTAlAXOPu5M7XZ6goEPfRg+gCEH7Ijc/G9T08yRiSy
OAmu972zGAI+2zmEWQy/h8uVPZRb5ReYeGbWvOp5shrWUiDmIOth2zA/BZlnKwX+
CiarOL9P46XXkwQqd+yVRf5QX0s2tfnA/TxxkeSE0IRHmW5SZInpxEl0hho7cRaf
hDrE+McYsycUzwaXRWyEBX7FTcrxz72Yv7PR11yHJcR6qppDrN+VKXYVYsWLXsYM
siA3Qw//4vbB6l9zw53xH+elTEWrjc33wOrXTciddag6ztJgMw4fjN8ob7jwYU/H
NXZvPjxGganwR+rdEr5tb0ambqHz2eWJDiluYfzQ8vjNor+ReSLTtVYsI2NqNzEb
ZXC7qAUVcwZZIK7yi/KkVWsUp1qGfwSDMZ5Mh9SkNRIAzNKDzXJ0UVxSN4SQWs0Z
nnbCM6j5nSB+FKvV5AoZ/wsGK64/U7zFUsj77OWi9ftPxGD+Ya80SYyxJYZNOaAz
AUWwyOSUt84TICin/9LEU7e3lPFORMqo9548NtRrB4TJ6VArxAlUrM98LslhF7b7
mb2WEkfjhu6PNhI5aDOWtE+0RPBd38WqmmmVGB+fwmq8HFKnKmE7AQwK8EFNCy1V
cBwVLNlKU96coZhJEN2edug9ct81oeOIpZ2pwTotB9TVGp/kuONNv/hK6ywPQwIg
8LcP7Pj+5CYmWFjMHfId+WizRMsYXJZemKUC74qsK83IJmiEWvW32cQo6J3MQ++5
We+7nUZJH0fbBGgoAirLK1JQfs8okwmP6Y8qlR2jifEFcYO1oEuRiVdgcLRNc5ZP
zN49WyRJaVGow/bw0XdqPhR339p8dtaLmbtt8S7MX3puP3lpAlSky5Y/rF7+EcYm
YZSU2xjDo5RuU1kiF7FF7rBvd8wB+NNfYnovz2pxyMEqtl2Vum7cbE11EmGFZ7bm
lF6jRn7nC1egv/X6+1My60dH8Gb1GzolgNqxGOG0nv3IVEH2g3v02uqWSDp7ISqC
jpKvoQRjUAa3E9q/7TkdZ1hCxgkEJwJH5u+AMxUU/rO7kmIM27hs6JmPE2ExXs+d
Wv9TjKtKeW4fztVvracRKjNW7J7+PoDvUosrjLMiJEiPnq1xnqTGcYi5rOBBH9r4
mfQpWjWYI66zPhreB6ZWp+JGlTxitB5jUzW+1eHwX8qX09wt/S7uQ9bR0Ak0AkXW
hO4vYCJ2ka36DRtEk6dtLNH8L1XuXfZ78Y53zVZqtcnHywO3XEMRt1kTyUcpYOZv
YogTrRlMas3BYbFU8O1IwVvx/zLgd7Mwfrfo13h4yRyWKb8RUkzc7+gydrbCk8vL
chL55PTQl61zbc+Vi8W37erl+Afn42GagGQRZuLv2tK53DnFclYlrKz+b10ZIVgA
tS0GEF6024BJwp6wsTwomXs72czQUNt3ZtrcNDx5iRDmi/31RlWJTiGwY7SThlvv
HutQrQOYLpe0iHyZ3CEmIgmALVfLx7U2deVp/DvFRQSjzyHn1JhZG2L3pWtZbQKw
wHWKSzR8/d0mjhMDo/3V/4kyftFJH+bloFvf5LTN/AeYu72YOhY+rLs3CRzL1SGE
miegQrPXIWnVwS/1yv52TtKWC9VYxoyINdkjpF/+f3O6McCHy+f0yNOqM6BljAYh
Mn1oVDZk5onVHgjdT10rR0KdH3EzTHkT1GxLfOz+ElqIqIEC1OPgcORS9JbD7k8o
FmmmphfvJ+wdPt85BnBi+LkTt1JIPJ5fJCVv/y2AAaY2S0ahHAlpTXk4ccw+eQfJ
vfn/9JsTMm7T8NhdFG6PF/yZYekjctWn2eNX5qtg6T6fp4OORUFYPC+1lG1Qc6Jt
QfySnYZ6dmpPE2smN66d9Ovy6pML9N/mTpVcpcViMLAZ9EqZyTwbHmw9zsHGFJ9t
vcLTpDNYAEcpIbyoeRR6q1NGeTLGqdlWNNZbKeSSAAj/58P61NKBaPdB/o4aJFul
74QHriYSp0IJoVR28wxf3BVJWH5q+QeLqfZse5HxF70z9FJ5AsW4aUgEYZqHgR/G
O31Fgs9AUnSl7io4n4Fa1vSGDwgjbQ61f2SPA/JLKtgSko0PZ8wZ7GjuaZ4SP3Ld
0nun8Ko6EOL/wO3cqABqp50oSs8OiYdoF4gtuxxhj4mq0aVYP0ImMNqgqPBR+XEG
V/FmsiWB1cQnACHVnvG72KOHDUlJ800NZRynPlIU2/oML9OLqhj0QSi0jIyXS0PB
5xqYsErQoyhFUgw5ma6buzEMP+1+Uf/VWgpGxRBBqb3hw2wj1LRzjYBiM76qyYKz
rUcyrd+cqU0Cii9K25Wf7XtC6OtwpXHaqcNPc0F9ZchWsyLObvpo1yurAGYtBc2Z
EmhJe1NkKrW6+AvRtNyrtVicWu1FNyhB4JZdcj01YwP8kk95dftAaqqkETLTIB+o
i8OREyDNZZ9AXDMU2PDYTyjZuEVIB0+NWdVOK46EPj5ZIJkwGSggqnE8jHFtvHkl
qPSha3gdDgtGr36YYjbWZukmKdpIKtfBYts98JRp3mHxFE59kykluQk16uZIjiF3
Jq9mHGoIqINcAFzfPE3+R/aIq4a4jwPsBCC+lmAR4IVQgiVDHoNZLZyA1XA7O98e
GiF82qdDgxJvfSQVRNmBJEIpvOzyLed9lyAJfW4w893ae9dAk7m3U0yajpbRAdX6
9UF8vi+2EBys9de8U+cL9wIjpGDkmD9gBVH2WC+zySqvzEbXvzF+0vNCGULX2+r8
Vbx9p5PRFNF5NgGwrNLqi0N4T40HRThMJLUDhtR+DOevipLdumZwZRkAzO8KZiSl
gA9rZaWGLUbNuF7wkL5xjkun03vxAmLqziHRrdbwkSx5F3sL9oQXmExshBEmW4k8
264fDCNn0cn4ktBiR3djHK5aO2gBPQVIbyJCZUUh7Z2f2fHb/x8sNWAhVM/0/fkM
i/TjV0FwtkHdseNWh0VcuJ80vPwb3sdU5gHvmyjLaqsxHfDxwkXsqgizspbumK7U
zXc8juDEsZLvz5z4bFEXIN29J5zT06sb4rKhcCRnXhJSATIdDjTJW2dgx+IoRhV/
p11ek4v0yU4zPx/6lpnOR8iR88zd3I+h1OH0NJS5PLoN+LS824GOkebL9PXe9LBP
A7UMSEpEUgSRYdqcvMRIrVYvAz3wOMOpAMtKm35Sp0Fd4BKhFhPfEahOPRLVIbYW
wYtuYgB1AyNu376XT3m9F0TIeHSrjqIcKKl5fqpWeZpbxsY16Crj+xZn5LaJCgmi
xWR3/pjcD45u6hJ6UMy1/zgP3XBOyxCg3KsIfqX1KViUCRLoOnHLSGYdusgFNhop
tQDPK9yr2ERrI4nRE1EwBiaALHZ25ZFNuXF/uKjemBofMn7UDEGX0cNVkoSCPC6u
XvOIQpm2lUs68Zh9bMzuP6fmR66IHsquPGZAyFq/PrBC8hgXEV9C2XdZ1S962/KG
+FKH3MEmv/B/c8g/HfOsauvn1M3txqT84RiwElRj42TBQnI+uBUPZ3xZ2zO2zryy
BM+XXLw7v53oBFEG0ppn3eXu/xA4wnOmUKiRsf5/wUoD5kBPydZ4x38hJHrPfvB8
7z8z2uWeMt1yKD0xOX0LJRFjvU/pYAgxc97GayeG80OBSCIokJcVNfBRsNFfKED1
BCrXgN15hLAVKI3k8KU+ENSVSZkBm80zyKej8xUyggjXEmtDjbEK2cvXPCHmJN1p
blbFiNJ4w2XPGaM3n830uta0fdgiVuWtwgtIhE6dYc9r288ZY3a1Bq0Jko3HzFDp
A6dKkBf7FRKHPajYUamvHLBtjWSeGvEHDgsfvOVcgb85M0bGfOOIVKCxtwNkoKUD
Sl8wLJHPnO0klwpxyucjWB8YMHh92olziQAPDNhEPqaIw9Sk2jQzg9dxonePliJs
fjcONrG7Dwy8C/pqOBWgQP/aNcL3rcfABbdkcYR0ioJ1Ml7gBnaMUDfY1Ezk8/He
dhVdi6S3sZ+vqlqGWB3OMQCo0bGiJC7cAli1orDuAmsnceYv1M3exXchJ0Kcq0Bm
mP11H6WvyJ5PzNyhI0KWhg3wen3B1CFeuNm04HSf2IKYICPfjXben+Dj2OHKkKGW
uD/PlioNNDKUFZGgKDWy0j3CEAGKr9mGX/DERKedXG3eGE+pQRxFY4IWGjAz8Jjf
4IlBO/UFwC8lgGsCvFBebnyZ9FKvrePWufbPzIcxq2Dmjw7LjkWYotfGJ7dkeJo8
+rkoiUFq0obM1So4lTCCZaWE1RodRa+EXH/z9GVVXnj5XNc16i9KYNtWt35xZ7n4
XQ1WZgnLjO1UI4HVxHNs3M6EGgQVBhfJf5WYPk45x37BcZM1TueLLdVFXdB8OT9N
nTJYMn937sgq09cgbrJjLH98JyLSmvMXDsDcMAT5h0zbBwucvLRNPL763V9HhJsV
A52WiqFiUDFOq7NZWGGh0YJwYf+jyPOOENmqslXXPM2mOOsenBGhLapg6SyVZHc5
IAwhkeWs1GyZbN3J2Q9rmcrXwwdB4A3UetEKRBE3DxxCKM+xaeX+UJHAjSr7PXt9
3oxRtFAglSA9BgfdhjDvakyAYlBxjBE/67ukVcR1S+Fnv52Q7TcNupCW4F0tMdFP
sK6XA11EgruAv7e+mfbyHy4yp8U9H3SBWWJXIHbfPuCBJcs82mpfD8RZ+9i0F96x
nF6JnRpKIS6XquqleFaFjO8qh9AXBtJzaNchnpU2eFyqx9O/yuSc+hfLHYg8/W7i
Aw7Re2SdvFwX5ah4hwAs076u1rJgCIAw39hoERHGWQIbAqAzFXXjVJcpXbJ3dddw
D+IN+7N7C17BBob796QIpo8aEKl8BvUwZv8vMoDY5Hk+GnxARD5rGO86tOjk3m/D
En3a1Ey8zRqrNTPThTWFH9TDltPaBiS1ven6bnyGAZP5Z6ib5jQHomllY57P7Ta9
1nWwYKcR/VwlcscOQLf6Gsc/Zn2Mg5ZZeavOJrRm6QeDB9h5BF69+06gL3WTz1tG
UfvKeTwSYr1RA8qcdQNB9bIXg/Qjzy3mt9+kHCHpu6l4yV/5poL55rfpZIoebiKV
2IAQ9DkrNq6fEFCgjgV4xpalyEfqpuQcDLVpWnJZj6CJAM32iABV2EuYxrP/EHjy
rGBT8jRJCRBZdXzv+boz9veSFpEeDRRgfj739iQr98KH3lkn/wdARPkHG27Uft1t
EcNxVWQWyjMly9Zn1mHXiN79+QoC05FRQDUYIWI6IxPL6xbfRgEk/sJh9eBWbIdN
QXRjI8H3b2ttgNZxOwbnzKpQ/BT3Mo899nGv0Bn6ifMjACnc7JDINjAseFNGqBnX
tFMHZsTrFiucawFYOpt7ZRVJX9/IKqD9q4eaHpHw7AC7Zyp9/WQy49OQSX/7UyZh
WtbDoJuCMUHMNXmfep+NYQHB2im3QdNsaXs+HLwJ61ACcxAf7KGI2/9gyaOs6ODR
zcQoPljKVMZaojPzHwoUJajpOQnsNHKUUZPJ9Rzn3jb2if5ZWmQ3CHT/23sZfiYr
vLIf9dqHacuG31D6QD5+QdU9gv2pZOZJOYxyKv1HNLDdxkDfeVxhrM6zAJQIs4Pb
l5ydKcbo4OvuRPJCED9wFWhuGNw3GrXGoMPwYBUnYORUfG0ZuxkQ3JX7sMeO37pz
ZAejLZAFxQSV+Bp9fD5P8hkwnNLDzyrnCCUv0UTYtphTzCrOtPV+TNbYd9sGiZFX
7YgdF1ww1qXcz1omKpQglH9T78z6nqfMrt299YFq/FvLq2v1ndM4lPBf6hHIaVYB
hpOgYfPK5Demeram6iuZhcGS24wONPDVPujToVto4qxflgaC5IQA2ERJ5pTrRj0Z
tBdzxvjrkHmCRitkgio6Mxy5H7c8Rx+ScOGmPb4rGF8D7oR2ZU8Hv3DqvITe2khn
QjHcIcdQhVOghpSV9oNhBVPHMsk+HpRW840VEpYUjXDWV/IIcLp8WJZd7V2+rK3S
QH14G8msdIE04Q9kFMRvEwHGUG1gml1ImthTBlO12Om9G/VnqdNmwnXXE2Ta91EY
4L6KYHmwIDkNa3MLV48wsdVJxan8/oh0phkJ1StvRZmwHJGW5z0RNYyjaVefGS63
RqIlHLm4l8XKiK5y/mgjetogBEPkcWje7tvhFztVk6qkHVADohskBzqKi5D1jQwr
QNjPkGQG3EINqFTSKdey9sGiurXk1tWNLGE4W766ywVKKe2O/Meu6f1poINQCoOy
pBY41HfNSQln/ZdRy90Gcm1FBSpe29AztxLTSZZJU3SGgJuYeQ/A8Aqr7oSuTHY8
KtMXKHqU6YkwwL0DYwfG0M5BkV70gODa+q3H6d11Wchqss8VaCDAgustHSdiReHw
IaAMQmbSOOAkSa5laLWeuR44+4S6GN98OlJcwiH/QCeQcr+jML/+/1dDoP/SPoUb
4NWsCPzIcGP/a+MjNZDUojxtiMLw7rAJ+jWJW2eUAHkXTT9NN4TQIyfOggaaierF
3djKD3L7Wc3lR8FPopepsQTfzldMERv0Fjfu5yQyv3GaDBnX5ULgORU8TReb7gc8
qXqs18rI6ELuexfb1Bsv25r9vDVcU5GeFlSDal3dCMP1NnFRsHRGUR+bbjwYbiYU
uEwLiGRaex9kPzfaIWdrROvKeOReAZzCTyRAsHw6zk6Xn9ds9YDR2gTNjvZzIshG
uw9ssgEQbiAGu1dLWuL6wJ3LDgQe2xibwZizfcrMYYsIH3Nu6wvy0w7TaJJTcbMj
zHe8A5Ai5mJ/YodnuAjTW86M992DB4aXW8DZTyqIGfjrEIciVXf+m35ADOMO4l73
KjtC4bG7C/GFJ3E8WZUqY8Eseg1n/1a9oznIrFkfBSv+dI6e80yTow9Foir+ATTn
ChWKxbyAyamGbiXIF/0SckfC/1jB3f62tnD5NHtkwCrgMxHx7y45fL8ielTAvRGJ
28XdS82gJF0xO0CRUp3eW5xfLGEA+TUjhvAzwgBj04/nRMEtpRWt0D53r8neUSgX
kPr3N/CT961Orlg22IQi4DzomSuSaGHkj4JYwTzt5NR2gwM3/e+ifF5KoMslYDcp
2f0Y8orAwNf4YSRUoC61BzCTVJ3l3tNSubFIvF5VQzb1KJstpR80Rsp4iRPlWqQz
1QID7SAraQRCByaAL059BLs5csWvX8iFkpKjWD0wDcoKJ4PqGxwVbV7HDL1rn0c4
FzpQjqrldrGSMvn+QizMhnJmyUTy9ld7O3NhZ4bEMBIcPsWMC+GlJ+zcwzULPRP8
3uL7CRdgc44SRO5LtDvi9RklJPD0utYPOV9yandvV5rdf+4DR/ZTBIXsXzEURXXe
Up2ln13KdeCRRMiHs2yin4dzRyORlmORrdRardSmP3hs9Fhk+EpSKkbTbozTCKRI
EvHkZVsUlTpTei5V4nqux10UcvEKL4yMgy5Sm6/WSR3lt8na1y3AMRYfaC/aa8Oz
vMLQkFH8LZlW98Mq5Nne7y95FUqhvbrRzs2m3OnmWPs3h1VKUTfUmHknYiGU2pw+
PL+b5+KgoNDaNiHuEpwOJumCliEC0M8BH2NOQVRdlZwW/duIrND/m30PCPwds2Ns
lnEHFEhbuWNAmrDjQabtaR/pzEL4U0RNwWhYsVfggvCVzWEjGBxRTBBcux7RKR8Y
/TNx8BeqdFfug8Bvta4RK4RqF/IVCxpTQfeTtLemEzYLLR/xVLHT3vvlxJiXLWGZ
NuuRFppsP1FAfha3jEkORkip/ZEEyItXl/X9PxTmghzw4XFCKop8UBDf/O8FMdVi
jA0jx2gIfqqa15nnjWBTB1yhlDCfE8c7RVwy7W3h833PWpu5J8dEpbc7MHOpppuP
lgtAQBQMv8zOOfFrjVmed3GU3HPgVqKM1sKfV88h3dLM5eQMJmJJasNfn8xtSdme
nXwZQTYZH2lHRNoGymKSs7y0OhvukgeDu/EwFSdJXg+SQ70vPw3l6tTNxhf+sq+i
c1FyS9HPbpcCpxCc4eLF+D2GkVjpX41LGi7LVmTp3lwk5C9+QY3HWw6wxW0akkuU
OmRf9gSYN0e82j8vwt1fhlmMScJOI6+Q7R/L2zqquCL5GdngqZVnfqzXbUSTphTR
86nwkNEsi6WHC5NMbIgv0GGdYOEkxxZuwsJyu3wiEQ6D/xw+45h/KQ6GCvCWNPbr
8h/y23riiDO/L4hqb5ugBrKGv58QonVmyI2mvWUhDqh4ZMbTGe4YTQFmfNPIsHPp
Rd/YsIiQbgRG+dRzsExfZbwconYpvqlj/IWBdaRXSb0+74u6/F4woqbXISAA0ZkD
8p9frvGIgTgeyKqG5nXyeHZoiVuUe/DekfDgAzSgjAudXUMe+vJuYL7uEifh7K0J
yP0+OYbrThF4kgUl5joAhjghywb4zMrEpKABERej+7eOnLwN0TGpbh80jOJjpliy
qYjyRkSQHn5LMPuhUDIhAdhUTk0DgLCQUIP3O9aUPLxVO0l2GYNYQgjp3kcS1u2n
XwRBL/YeJDko4HB/EWuCa0DdRApXcnzZG/22M5xhwcygySeFkzIxHAbh2oxS/tky
rft8Hp+IdyCAoHAD3/IDFQiWwDvuVot1gV2xKW6h+83Kv46lmhTL8hnFaEY9zPlI
4hZH/n7Jp2UJCfm9yvBuPOxI8f40HJ9hM1O+vTjcE8V3Rm9dReJ5U3HQRc6EO6M1
Tta/dLWytoSHtFT5TAwAV+MgJVYohzAU+iTRMrhkduUZ1uJa11tH7442K3W2Mw0/
M24Hk0XKCfyV69ufNZ/1CHpn2WzJ8mwvhdJjT9Ab0QuPbEm6zroJLHvNO4eOek/2
l8cVUsBvl46jVIh886PQeDZ3M5QjwRfs2DGybnSKq/PO9uUTK6IckNi63vqy/SSy
CvuWTmtHrVhfIgokZF27eEajOLqotrU7RZlGKZoO3WD13EyrJf8+Epp6DBcJX6TB
i2tvct4iHDC240JcEwvtut9RRhPQIaYJTYc+pCqBEQgz3o7ds+dN2FZOBBjxd7Ew
8tydHVlafuHPH6etYa6KsA4mfjcBxx4HhsvCF24lMuGTvHJiS3VlxUAvH3GvzNGc
eM8SnjCi4dStfrdx+VSzGRmjyq4N0/yPPhE6ADWmjiZF3A4HO6e/TjLOteSoN8/G
vZYY+2JblNZ2eeGVXAe1mQ3YPZtIJo/4qE9CJfDoCR/eLlgV9EhX1vEP7dNC7teH
qFPcadzs5ZYQ6ox4jskDnjNt7UZ3KSCNlt7+3nUkH7RQDWmLm4NLu/g9hG82kJNx
rorv1glQItgvxI4O6x4DwSokREE1UI77OXS3gIwU21MwFlMllt+LV0GCQxbxmT0D
ItxBDyIVKeuE8sejE6+EO/mGk/qk6Z999rBYrbDUNaVDJyKBWmOIeqvyOwtkiMnw
bsrhFtgs5V1IabuwbI7aHM2bOCkiqWdrcG7jS4XDBt3LjkYyA6mPTDiL0PrP3bw/
u4qhHdzdGZqIholBVqI80cyQzqVqXavLPq4znBcgUDBFI1CNIKR2BIwalQJVXZzY
yKaGo+2edwuXDLyxCdCt1+1SX2wHURChOjgleKe1T0Tpdfl8cYJtTxwDriDpDIdL
0XodIrdnOnqikb+gMUdM/b1JWdsP8IQckAtAJcVfr99qYXmn5VbIweq9KxTioyM0
KsxjP6SGzw8PHdUjCGr1kOkq81bBD6k7HQL1/vFmvUWtNPGmFHfpnpooP2Bi4B64
NWPXMSqRFmybU4AfUKT7/oIwkv5lg0fc7QYGU8ZiidgFkLKxqfPgoIRTBS9UBV0r
ZO31HYsTzLIbJqM1PWIpOyezCAJV+dtKCDR2K8sRBxMohVrFrvrqyCK4f2k4WfL4
cvuNN1Ypgb3HIlc4y+4ou3DgaUzUOCvZwkCrd0zYcpqpbz69aN+jTzsDXncxyexe
lfaJfZdWeRcZkmM/9Eh4FxPh0jpba2ZaJeYblYt+noiFbGk6wBswqo4xjr2y0e21
xHBOX+c65Rn/MyC+8zNyRPUydvjoKanVjmgyTuj4fFaSi6h4qtzJokjjir6Xm1U1
QbrktMFzS4sRfRzWb/RphNRpjzvXNoxbXb2iVXHGVz2KYGJki2Wt9jRcVaNaErJ/
NnstbHEkHTAWFAoTN5BfJLqYHNu1VIa5k2mdEI14Gn0JcBe8jFD0VZQ4/PrU70iB
jq360jCNAOTVAjduFDvFx4tY3J79wHivewbDLq/r7jrDwTYrbnP96HfEo4mY7JOj
/G1/S9V2UfggUFzG9v9zWOBK9XuHEmO0QzR3eJrc099FXnJLrbpc4u/TaVYndmre
`pragma protect end_protected
