// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
0Wvqjbcxj7NdFs//tOCIEM6cWhwRJlQtcr9U8gVvuRL3/BUqe1K69k4pw9wRnS+i
GHTxnuW8Ta/C/Dg//9icpmX+flrAu1fFePlNJ050oZkMlP0nLNgQ3X9xd5SqQ3L2
E4t5LmBW5OQ+JYQR+NHM2zjwm1o/LdWMuCLLcpmxHOyKNKLwD5tP+Q==
//pragma protect end_key_block
//pragma protect digest_block
Vun1S1WvnqVFd+JPlwjy3ZYmJeg=
//pragma protect end_digest_block
//pragma protect data_block
N51ctTIVlqaZ486k+mohnhErCi6+K55dkEAQ392IKqDpJj5Sg7Xb6SEytrW1z3yy
ogX2VtYRmZ8g8mYIA/KLBj9SJjSZTINaVeGsDjHkTajV8OjA/geTfKt2GnWM7xuk
Cc6Vsk2/YonQAEO37qx5vACz1qFlOdU2S1DKNl91tx9K2sHypIlaJ92QWj0u2B51
MioAp4UrW5fKpFZtIDNulmKuLUQiLq6vrUeMc2riC3TxRTcUMcmGH6F2VcuUdRlW
6ZupAc8KYPU4WJVFBP/Z0HMd3Sty+UdJm0foJxSDKAUA51VNtGbjVJpkrgDOp/ku
s63len+Y/2FX76yUQk4ApD7dIfHCPnnw8I/Z8MWA8oSzNm3QTJN5FrWFrGmWEYft
nyqAugEqBTp+txz6MkEXyabXyJemyveuGKd3VcwxcMDO/AXwz2Qhr1PJJByvJYgw
B3+Bv6vqF8g/qvmL454KHGe3D8dx79jtyT9bGCrbD9dOkM+RIIbIDlxt31srRfUP
RVZI9Y3bbG7aKv8E4fWXnDljQ00Td+e6E1ALXujFzG3IZIqRnhnfJHzJGnibtgVB
RUDzz3R7wY5pMiSCZ48f1T7bf9Phct1IZxDHd4AWjGITmzB5RH/XrqH/vX8ttLAw
kX1mnbKYu9Hl3dcKQU0Xe98aBo59SLcnCWN9dNQwB5zF08iiwypD/9tdV5PyO2cb
WfjTiCPoPj7IBVQtOdYx8T03lhuzmVWtL+aupCbm6HVmOdG51xHuCuK9YTHqLGNy
cJ4oCdoN3E1zBuGKMVfk5zYRbBDJKrSTJcqq20zrbcFhfexxjIbyTD09XhxyeLs+
wv9IgiGF7UxSZNrFZR7UIrDKi3efMZeulTxdct7uGbQFtiTWLRb2KaonYpdbUme6
tDOUU0ChINyaadjlhbvC4qmb1MicxYVX15UqU92VvQJmkCMmJMtITBsaoHd+1JMv
eRJABdAOMbwdkjsLb/XFv0eqebijikAs3Bk9J5Byk05I5RY5A6XhPo+ysI3nAEZD
iPQ6LqUTrjtBv7+DgviSmvDf8Flzg+BoeSakSqANjogFCoCi1wS5sTHOgAejwjBg
UVC1vo8FS6+NQSQL/twjMvbVXZGc2oD02qpDf1SL3QfSJuUkvV3M727PiCIYI1BH
FA9qERiQNMfL1EMowia52frSi4PZWUcFtXjW2t16AOJVdIZ2ivTcAyGIhD95hGmN
y/xBBpPXsaKqB0Ip/BRnWNkKiBPFelSe6zy01Zohyj9pdasfr7bJLWxvpVG5QKIQ
uvaiRv0i1M6FoggqtaoZYrC3zg3aclum3WCQjkKxj5iJj4AoPe1rD5CJoS3QTcZK
EU9rGC0pStGSXd/d4tOFceRHBVyaQIJQ0B2EXLniLceTHBFFumpdIQXngTo95YeV
2y4CLXENdT/BeKDtfMTNqBR3DPlOTR2spJ42NiGa/fup6rq23CnSNfltzK0N9H24
O2nKngNLR9sTZiXO/PPnd91KffqidS9rAELRyWQkTA6kkfWjV550/6LrC6wVYA29
8daV/g1XW/S981VpzGLrWwjNoNu3zn+7Brvw16e32Sy4YH9o4qQmdiFvA7aH0OHV
PYv6UOjBznW0h3ZFnxVIpy+xjY30DWz0GJNu2iYdTd8W72lWEHT9P1pK+FUa8Fiu
3iEpAFRLd5AtvCsx4hwkNu3hhs1NMKLM5cy47aztj8CwGhPF2CLfc+ZtXroNXKVc
brkxrKXSGZWYdBnG1HLenhYKnfdbZG2IvWBAaEY9vcp5szYyfsqTbgdJ1dGdc43P
zbHf3nDJ0tDNQXQE9G4K+URDI/g1P0VyPq3Aj5FRTk4Eu08TLw6szZdf2IYiV2e8
c2QGl8qmEqWzUAFLkSItDztIBJWJhcV0L8VjpWZVjCpSZ4/KBM342IGnRy63zRZo
lE2kK/Je8Rrtw4QpAF12YST/t+NEbzFOfw6+GTQ9TDtEiNuKOhiO1iCr9AlCWK4a
GTnuGXmRJdFkr9l8KTR5KkqOKWy+O7HrgM644pwq1Pr+l+wN+NhvZjYfTQV/Mnhb
EVYPBIlu7Zt80Yi8mbowpbnjKCmYUfEnsejW1p9YFuxxBg7s+hNhDh5mBeiD0evd
W0b4ROmZyhroVdyo3jCcr2F4V+wKMKxvozqohLr+5TT7qRqneZ7+5+6V0QvEcejL
G9U00bCELW8Q0MF9z+Cyv8kP4T6SdPtNHrrIIxMdPEx+EevEy1tSivp4CFTkrsSe
esqaGB5tRnmyzLznNgkDy9GZ4s90P7qMx79zIu/2kcNrQwvg8v+D6nWjdgCAJI7B
crrvs5VFglL/Z2ZxbatfApdUgmYpnmxwDuT2nQbSo+jeQTuXZvncyBIFHhIioIpQ
xN5EJo7Uf7dw6bxH4UtWzRwAH/yUn6Uy0LP3nMnvE+qdPWmUn7bKTJyZhELJJSem
ZMHW/4XThZVZQLOU6EtaXUr3F5v7sj3gc8btRyo13RgsZY74Utlggwm9LosvZbGG
LND0XdO0yr/amtDqm2abazYqWOHb5fkj3l4YAZxSqmdSv8R1cdMC9duTKBGXt66H
7cIr/K5SbRMr9eo2Ol1LRMx4yHdfAh7uyHSHh5CCz23q7Rl7pU5sxw/mNQlDzFtT
0HCYD5XkoXoDLA9gXVsas7PpXgna0aVFL9MR+IkPfxHqBzZ/qsdyIAeNNxDq/djL
meXgwkRUHSu5Zyr55o3V7IxQHDZltvenZr6/bDaNc59AyvTNYnc9fMdspUF5A1xx
5iP8lh36BeE7lbFomG9bn5xlNZPEQgNS0EgmroxcOkBbjzrkRUTB8pRjN2ttuVYl
LdnodKWflMGQjBWSFYtUEGTTDjCSwAfE3KQkP0NadzL5OCctwRVmBsgFeD6kTYMo
X3EZOjc+iIV0onSCWwos+9N92i0VhV+1AvKv95rNXa1UZJijWoRT0IZBzKFAzH6i
7F0p0H+BH1yOs08eqqhUBmjpXJ59ID1CShguQl5vHJAgho0FqaVpjcs6Lqs7toIV
QAKZ7uux3Y08BcdRoeR5DlT/KwaMxgRTvmdoIBWHus39xZzUZMu/lMNZ+Dmp8yoo
+LuYHZ6ToL9LfglPzYHN/eXYV++PwkOvJ2AS8j4qkxO37LMqpi7PjJQ/qdxHkdDe
vLJ4UHR+9aWEe/9l6GcgnyWqpm4YG9laWtkB3nEdpCNvUfZROX+S025W7pKuSx1Q
taYy0EDb5o7hgHHn69sY4wJI4kOs5FYf0TeG3DiVqLmdBn++qTOwzNNFUwDMHoYw
ZQx6i9XHMyJ4Tv1wGcvvBlvfk+Qn86Dlq++8lUx9rOdoAMWvva/Xh0tKzYGMxqrQ
k3LYJiZb1CUlvXAETYAYzo1ijkZkRSarhsC12oIYw/HoqUZrCZO36K3E3VGreJQh
Vru1ixtS6SBrfR2txvdMfivfA2a8h3t1MYm59ixNc/akRITOcrPVcLOpySQpvdvs
rSr16FcrnHVdKhykWmPLXgfXWyxmrT10h1yCRpTBH0i4xWtY8eJ6Okg5UeMI8D9x
mm17Vxb2WVkbJl8x6d52awYQxAzmK+m/sukgYqVQusH6Z9ZHfs29dAUsOG4ih8P5
RQ2NNGGk5lgLDOtO98qToWdkiwbmPeSrhPSPgsGn9foo7cj75kbylSh/GUySST35
3KX/PmZGLLHYANdx3s2dUW3y6x/OXkrd4w1tk5vnpj0+mC4feN02vZBEE0iZjI0u
OD+4gnMGyrv5xNbNsEwG9qX+asiFxYV0FCOvGp4PL896dXc8wB/0n+/cgNYYzfcM
mF7HbFyeqMgJ7Y8fO5QKvBUKzVEC+PaDXiuRilw9hVFVBZdPxPptXMgyDVGz/pB4
mh8kMI3cHPXTz6XoMNpWK+Yi0RnfbHKVTbsOr8nI/1I4LqkygAv4KyAHO1wqHHzH
BIbe9kpR9UCa35UrgWNTf5s3uyf7Fu9yRc9eUg9nzhocg2KTG5XvawTq22Ah3y9c
aMxe812zTYFygPMs9OoTPnGmu3Jz5D2og7QAYUVAP8mjQ6+v5sBv6GNeAYMvKRrf
dglxfq+zaWHCngm6diHXK4Cy1OODgNucgx3mT4MUaUbxMM0bBoJ4O7t320TkzFqk
coZjUlyH2Ah+Ufftg4Pza63HigX9V+1BFwzz6XrTypgvst9FeSuIMAgALJqHiXLt
5bU4B24k2g/rH2wr5gils3bKAGEICEMj+zPAModu23RBxE2kodc1vSWkqnQfWeS0
o4icxcLeA8z73S9HpboinvoAy0G4oRAYIz5LzFwYvbbbVo0/699gAWrtnxD1PIbo
OJN4SDoa/cQiNi1YxA/JbmkQFe6wWarQS8ff6bLHTdStZ/9lZJfmVdNsmF4k/bWK
NKcQfwpZlSG/PW1gvL0g9Y1qen1wsqTBq1QLk5MtQnhtNOp4trgq+w6kcsYQ/EGx
u/J+xlHnkZR0bGc3GNXA/g5Q/GtGc544scJKh0QssRhcmkweRefYxrGmPfZQ1ZoU
epFXwixVO/0vomLWJ8QINm6DnGJdkSy0ktPRtr26ljhK0knb1fEopiKFwayjEyif
Cen639FI6fGDyA7DpXR+TLguihle0SbUIH7uafPi8WR5s47dQuiwbuky8hTUEhOZ
6idgfDQ3YpOZtp+pL/eObMPn9oryi/DlPcxirjLRDEXzhOIbqZR6uwbAkoo5SM63
miFjHiTBsqEnu6Fuh4q1gkK0b1ox/l06Qp4fxLAXrwL79PbzJ/zMj5qvDrQETcAR
4gyoQkGJqE7FRfUkJzW+jpjKTzt3MxQjLXRGNsxcJzku1R9pw2a6UQTYYQHsFc4E
i6CpuSYVsMR8B+nSOs5iemrgMxcM/iwEXBzqujqza3FPgaEXefWbNGfxNGeZRDPL
YVo067kIKMsdAW3QBibH20K/m7JGoaPpxru/DlNeP6Zevy2O7F6fb/2yqYM3PwyU
dv24kSJ3/sb3MCeQ9N9b0+E/q3EaykAN4bO/OluNr/D7md6nEOI8RDxECW39cm+K
T6XdC9YZKFUMtnUSpHkIiWHYJfBdXZx0ziq3AvHL8sbb+LPqVRbvh0TgXCmNk0Pj
kT1CUv5xIrTJ/ZNK0AozB3NN8mLOkZqfLMJjygXMJ6z/z0U9mr/PuvWnAFj6bEcO
R54Zabz1tFUeof1Oo9IfxAsMoxSCIOdmd7RmTBlhhLkQwvaDrihDCrZB5knLJ7TB
hkeSZxqtbv1eb2tiMLON9PbZPuylP2rSBvC/PbwfbYruYimru4yLPSM25r0rwSu5
RRznC3lJaWMaM7y0zjY0xRo/UzFl9B9YNOqR+loosXM6aTPkZVxWt7thvHJGh16b
xDF5JcL/FZ8ySGWkkTzWJCYP/z0dYBEw8lxjkbCSwDniOjnmfvr5+7lnNggoplmz
oPmH98cQXJ+7byRrrNpppQZ37Rb0PEixN6sCMBoHhPhi1bcffJXoZxFerScsLtkx
REHSxfODvgtYwpZOjnixeucBv3Kxqy4zXyfmethwO+NV52aL8npd4b1rYAmnTJwB
BNMu+VzdMK1/d8XWW4io3N71u7BZMwVJZX51DXBArTIexEurPd5lh4B8R/8S2B1M
cn0ayqm3bo+jO9SPEMLgoyfQMjN6WxKsLZnmWM6L1pnpAQUEvMtCZ481OTN0RetT
aIUzxXKx9s15qgKF9BdWJzDJmspM2HQcAaqhHoModhmrRPD+y1MC4Ed4w07Efre9
K7qhHah81OVv96rc6wzX3u4v0d9MLHO/pkGUNHgy7OL8faGwZfu5NmyD+vXLpT8p
+I3iH/F85GI2ntSJGUiy6NmpPXgl8VnMKhAsjoXmlD7bZS+mBIQOsbo9LAflE6V4
rpRUqHQqQLLpIrAnSsh/g5Vdzbrs+iJa4YIrdu/cU4yb2rpV32IJVA7lzyI3oucu
jMVZKSmOfq60FRtTRz+HKbicSZCfZxAO27lgalQm+ArIfghsObrGHSUwrSMS9m53
47Uy1z5XMIDyD3axlDqn6ONzgNN8hTFnWVtFg5hCZ6BwUwoY6MPFnh93knKoVLrj
QWfrpkXS8/7paJ69okIj6Z3nGz+jxT3R/Vxw4RaYrflvQVCh9GI/KM+MksWwDxIR
h5IU+K7vSL2ZGRQKszFbqaWhl5b0oefn5Nn2lTfAnLQpgjftvl2TnSFa9r1MXMKn
9h9luo4K2d12NRf4GKK1teE0zBh78E/+CJ+76gKtNl+ouKma3zrZDkT68McoWWH3
8VeJTx1/wMYzAtl/tr6Zmrn0jq3+fiQ64WJk2FKCduxy4IzHoRMDyUNwuS+M2wZS
lfZGHrYJlDSFu2yFuEc6fKjBjy90e9+AJ5ajS7PqDpmKtkgAq/oWl27VW67kbV9x
0Ifoi8uGrrQbIRC4r15xwnVtSdu5G8T/Wt4Vs3lneYbwMkgJ0On4NRU5n7nQnfWr
jSdMMS6omHh5KmVAEdoqLznHVPBTiBCfVUXGy8eg3Fn2BbRn6ph52V1zGD5DSIEP
ORwCWjOzlvMed1NvgPZ+16rq/5Za6QZHqefT1CkNF5hxdKzGi0ORysyEYCr02Yx4
Zo3vHbzr1sl4qox0F4qcfUnij/Xux/aUMh/2RV1IDhxCzotZ+WPS++enSMgZkRam
wJhWaqz5IQxDokFyZKD3oEejbz/R5SAnRm0whVyay0lgSEAiFjfniCVJ536kwPr1
fpxasDOd+HGYfPVnDBXnpuYuuhX2XVxTYeZLFw0bE1/6l+8UyThZ71lSaPBGNsRq
U9ITVPrwNb6iDDhtcuCAbgjKU1goL4ao4/lxDn3ZDm+tv7KABApi8fEgBBKHakub
csn3aTIrKWUc6lg/JIeTs1nDYtI8ZNwOaEnjdX1pTVFsB7gfOs0v35SvhKFwTrjf
QsL7R0x6qWzFOlD5/YbriebsjlWSy7xoCkozSGISrTjEmj6PzzVj2ODmjhPme9Gp
Nxz112tLHC7QN168qO5n60+WMq7LCnSd29nO7Eggku0ZP6uWRwe629SEBBwIuLZv
IGKLavsNoSKSlOHmgI9R4knDt5oJA9lOC/ScyK5UG6OqlzjzHvKpkk4luQg3bQlO
e7SL2pmqpNMAcvN7NZffp+gx1vX8hF2WJ0U7OtKft9nKTAQB43dqhRUFEvmtkd92
WFhYGOA9cd/a8ngEp3LguqIEqOJ6HIxw48krK3PnTLQPB9qjnrAbVooIXKmudzNS
ICgdvXHMoQV/02YqBgOG7QQXoSRV7w5PdboLYAfPAUSumM/WLOg2m3bM9sXDXeBf
bTJHxhfJLsM+VJN1wqLzr+njjtIfAb7PuiPvabI52GDWajwAb2Y6Sh4FNHbwvWY2
/0awRKpSbvgyAEqN1Ng+oi67TYywTu8R8ei2sIisQ8OA0JmuUtyB7gqI70Dm8JV7
6rXcU3kD/4+nmfbT+O76VHpU2x2WQxRh6IjF+jYjS7fbbJmSO3v6bKtq5M9cauuR
+k+MJYR4bwMZasfo1FrcedIFFXka+zERrLmPtC98s629NhbOu06lZiRh+lYlP39C
zt/t9/Sw1tJeFTM68a1ZSlaElMNqJISH7Asg5LAHAg04PeYYOfDD8YWGLaQerf+s
HEwe7Fbz01JaPLfmpVWgZe9tw2DFfzrSkC8RhwGemyIuc+QICCXK0GlpoUvcknEJ
Lqj23tQY6uTmzh9fk41yLcHdkHS24H3RGJ446SSN9D4WFtaXpFDR7B10g14uoI/E
O756WGRQIJs5I/nyFCp09z5RIE7iCz+yaCEnHEQOJHa17Ftgz+Mf0KEU2uc+KKZW
T8zK3FNeff6d/ifdxvHJloHJlKGeIvsH0SVH008BDzdZHZwYMO549fJJ+yJxYuR8
LcXqHhe9pDH0fjqotctlUYr0PuGCVMvirGAJwb6MCjEaSyG4j8zeOdiuPpSo1t7J
wx6RuUMrrZesmUns+ghDw3lCl2Vyk5+IHEZVjC0uABgA/ZvxgEL2BGJQPJWpvIwa
uC1be5I/tQHxCq4sdIA8M6tIFLlfXeE8PxNpQp9w0p652m9rLCfZDliKVQsRoXBf
4tK4fwEMyXdp9cX38uaPUy1WXEnDIn3/w33Pgg00sshQ+jMAIsHKGGj8dXttOLNQ
HUBVbgf2cbDJd00WQrlozEotIoSO8Z8sKVGLOpt9lk9L2Q/rhcV+lxNDnZDV3Dq6
68iZ3qZSNVeuVD/idyGEBvSHeTrlI/jMtjjuyiNkETGa6FPlW2ozm3vYhFqFqGBn
UnsRt6MejM0KXUccIPfajf/romtws7FsJT//ojS+n6U3wcEmVH8V7rjArWIts2Jd
FgFM4y34dEskr7/t4M2N9XiJPtwv9Z/rDyvmcHc3TL/GHamn5jY931zNvn9rfpBH
evZw8skfTmMT94aW2dUrNMlpPvjUops8riSn/4wXaNCjWXgxEsAQauU7FgFOdd85
SEmcktNBR0sE1oB0fa1l/99rtTDiTrgNgmaJYohQqW0sGOiAX/P/mY1evo8bmj7J
oem3dE11ziPJF1SZfDhXmjrFuYmDlUHBRxbYPmtIzRWXGKfBdmwFWWJtjaAYUSlU
1dV+xwCmL4BpTSQObdZABFCQAnnkyice/2k/Pk5wqKqzDX8U94k7bw3v1X989X+/
xldM9su04jS3Cc2RGtSXYdvWFTHc2goMaSwVqwhgKRRTb7BPpbBxLmcpFns6Es+E
kC/r/r3v4U1s9FlJ26jtJmeimWyWqOJZ3HuWyvFK3S7y1b4+5/dGzzKHod6nTMiE
NBIgIjcmAJ4eQOYCGEQNjJJicxh2n9Mrsk7QNC34PYgrSXTl0Lx7+EwzsG4P3pSk
51OW3Bxk8H04gbUNKKEBjcOaDjUT/goNtyV6VACpVzx0jujoHDKgt5QM3VRQqzsJ
NzyBadguRu0tlLyHev7EmIREo9vwJV2OGZ5uIbCCBQvsetn5V96c01B3Ya3gYw1l
2gGsYcmyZCiqLv5Rq+ZbsdH6KE03m1kjyv88ke0uCP7z4itd3YUVqZctbZe9Rl9N
FDtl+OLCz1pQBBtCcfU7OGfwUPtdI3w5oaSOO4kyOE3O4NMGayOtzSZGWO2gOg5C
KDc6uj4wpW4WDof1gElwU9d6gZkwTMykV0H2opVJ1GYV9aLwSOW0gCUnXVecc9hh
WpFbiWKmfrHF9z4y4Ohihjwq4Th6y74yDSlhFZYdfmNa5pMIVeO0chDuWJYrojtC
swYa9wc1LidcUrAr+F3cMv3ZIcUh5RNuDgbQ6V2+flSamOnz0S/n1DQABbrLUm3X
E+UKC1ZfuDeFMstM6felUbvNTVBhp6Q82KE0/64lokEmnMiA2H7wJDiq3VocH4n8
kyfidLBLo1fcq1EiCZScGD4CmjAiT+6htxb752XyTnn3V1a4keX9qa9bTLHpltOJ
uj3cxbH9rGQ9tZYzaFw91vGdsPqIbv/xfc6EEnAxW4epYNnKDT+MVtHX8bOqzO/O
ltFXnlyhWpBB95wiZkibcU/sUPcROWO64jqaDcFhionMtM8JpKMo5lengt9lcJrs
GescTCVXTx8XjVTq7eFLB/qqvhM5GaaXBhgerkK1wGIe77Yur9ENCSQ/xqz7zST1
veW797KLlxprM4Hou2mSqciRD5Evl1mOJiA0CXjsUWRH9SeTkU4Q9EBAaoGURIPB
fb5gVdAdKpbe6qvkde1KEINf9O0ehrZ5FL3D0E8zgTpt0rdGuATuqtptv84BU4iH
/Vn767AXKjVJcCP/hQvs92htbcxXuY4Vz6dNo0O5HmFgLi1buKbTAQPhWRAZBdCb
WoeGSxJKZymu1yKctm3fgigSmUMaapBokDRoEZvDl9CIau9KJ96zV8HtJzQx/CH2
tlWaYa8Hzr5rOOBlvwo6Hq2/cPkSPAH+ifPNVPVTXl5SuHn4KD7KvOhcezLQ2Y8G
CEM4KgL7adr0DlkaroZHTK0tDMXNe8XRkYlmFKXqX1iZ5iOeHkzwoCv8+qpWVO+M
fdGi57pmwg4qBSM6akFAJ4ElfAreypJIVHdMw/+8yAOWMleDtZY3f+oVq0lK2/Ji
5/HIGeR88re4CJVUeD6Wurg9ZywT0XvXbJBq0/PmmLdZdiTTW+LOCNjhhdKxL7z1
bkhYJpkxZVsL8fcMdA+g68xuFPMxzaXUYT0XVrukc1IBoIIc13PUZAQH9isNLdLk
X+OzlYdUjvQOUI2Gcr3kIzJE9eOmNvflzQgDnGDanyATCHjeR32YsDAq8JCwvZDt
7mSPoZglMr7TrOM5kd3NC+F+NwX21Af3iJEKHp6CQJk2Jl2cFV7gceB5R3+7rQST
sxDfkrzx37C6hFJhJ3lf0A8KmA77S4qP2hdElpG6M18B+tMvz9J49YOMDOW16HIe
m24RCzeV/7hi3rQu8BE2uXdtQ7mMD8BIw7SZZXF8EDCpv3fTV5f7BIOU0ebbWo23
E4Gy5KpPBmuiFAWExYToLvswtruq7UM1+pIphOxg6qw0ODGY1g/SFeT57ReyMx/y
o2w0Rx8oGoA93S6mRi76grc3b8hOyhP2NP5RWICJjs24ll9laMEmfEvWiwpyELsq
hDpSCB9a42mgxJCJSjSfJsKzy9Tcq8wnNWF+VauOP3U/ZnYyjIc0aYAZgiAZWrmS
R2cpfXcdkt9tMC3X0uAbCzIGKN7PiAMbmPcfzT1CIN6jMH1quia4MSDck34o8wY+
9i6FxwlJ3Ft/cSWVb/TZBxSWQiiZC5XnbleYfSoezQZNGTgiB4TR4+Srb8BfsRzT
7i3YIrt0V6Xs7pCKDTWws7LPkDcRSdvnfpmc8+RZYO58HtUq0ocTlTfIOhlRGZec
xl7gOyCqqeaGuYSD/sfXE3gHPoQhquT3vXGmB/E4t24puqcwcHmuIkNl8ES+/kpq
Lt0EsV/Xo916u75svIGVbezC6IFDA4lfEwzs1oXA8x9NPMekzYZU3s2YpWapEMw9
Kxr2QYjYd09MnGeCbm02nWZEgNUW+wNFONCnO+7tURpr2780TcpIk1V1Od1y2CuK
wwtkZXKv3TRastQrax/kJG/jxVoDO1Co0UiV9uzBZPtl5B1yBPOPbXElQV+zX3gU
RGTS/Fc6ImPjF4QrXwlY+59a9PKSf6X5c8QyYcNgivKypTAelLsVLYY1yyDCWq04
L5sSHtx0UIfVKeq0kXiSBguldczLbA+NjCuDyn35TYbWkG0JPinfk+/E90lf2fCE
MMQE23f3nZvjPtltjQY4SiP9BNJ99IYNMHr5N18dOq/KxVyVVpezSAlinBEoZQaf
sBq/YJ3y9gP+mmc60y2fdjm4eTroDugPnPPi6mWXYkCSpkDsHrM1ooE0Y5h6tJ5d
GSMMPbsbm+EwnuTSkUWZwNEIPFdDOhHGwEH1FIKxSEB/b4GzVu+ykoixmQYHr26Z
s+pf4GS8/1P7sCZKTTvBJ/Oo0uW09qtlldjC+mOxExfEJZ5bt2W4PDASVCI7QMYf
NkgYChZUWXqmNh8oI8W+DU0PBpDr66IhXwpwjFBAMVwfEhp1FXbSecRQeix2wMij
xroIhmSDHeLgXsb4Q69ynV2sQd6s0336bulsTSVQvmaqtPHsf05+XKCNwftRvQso
l9a2JRp+skpGj2RZ5ChYm/PkcW5M1X9dCw9T7i3I0/nJOS3fB8ihl+k/p00stcr+
iB3LTqwGlfROE8WYYJ4a0+KnO8y1VI9B8mkZIpOJh8fmL5gv2EsInpjHV3y0l5Ml
XR0L6tjYO8cBv2e6fwHDZE9GJJRBM8A544+DfNl46XQu/l3uodQhAGF35Z8QmCQM
+1cZYzeIC6/nr0AGt/PjHo9rYiGKaBG+tEkkXXRZheXSSV9YkjW3xygf5wm6YLu+
P0Ih85ChRF5McGzLMNI9YWiUbueSDlL+8nPX0kYKlp0JfBb2q7qDpZ/A3wGEW2c4
nxVEc7DzSZF2whtrGVbNHCV/SlQ6auKz56aP6bi/O7dzpbq8+YKnVQthADXZ/+u4
C8ts+3OruiwCRlOa5C1vHBgQ2wqi61/CGjj876FI2arBIFTfrwRG3URKznaqDv5q
oxtpIyoomgWUOCijWwcf5TxZ8yHYShXTrMiWxYKUYRXaKrbRM6wpUk+GoaZKgLGj
szGizgBQt+z850OM7xDK9sOWEmuowNvfqIQbaDZaEKjDd3PLs83vGgs4ySgYBVRC
giLGzLXOJLF9Nxvzmrm6+agwE9Zgckfgg0pTrE3VZ2PcpqoUv41nIIndq27Cogmx
Hg0NXDvKuzDKQRInknyEH7Py8mXXllAFrLTlcVwHYSKQbo7wH1HR7xssulqKZiFJ
v14w5V9eSbMB3zkGwc4DGgTGr4rzKZ67uAdTQk5knOoDTmrFbah+cOGztCjSO9pz
YmZIBB+hBcbFaAOixO7dwgRNCSzwP9VxvUXZ8WtvzA/xvIm5d6C2W9bKR1B+jAT7
+tnXICU3Ip1m3uzbU9BoZbzkYbbgkJ5DV+Ho7uTL+k9jlI2y/X3Cz9unJj0/60Ed
IwfcBolfoUa2UT2cDKa8gefllvkcdbMiUxnYKwJr9f+goPvbUZI//GECL4iSsyXJ
waRNipau8SUE1sBHZyTpT51yv+vX5lgyX6oLYek76MR9cdsxs0v43TV9861o+xUu
CtXzUdxlVk0uxcXUG+ygayYFrMI2nbn00tB7ys60y0pPcimlNBbxmJe3DHh6sNfn
4gDBGNZw26F9w1aRDlD//OCxSJi4gl1k7NvR2Dd7LH2Zfb1W3FxTYOvxpQc6t8kp
92DZnyKxswp3SM0GdTVQ2gbxx+83NQrKTULF6+/mjaX1lBNjQwt83NRaBDWphhwF
toA+iCa1W0aEqbwWIXq6c946jyw/WvnSvSeXQ+tJxbTKDM/nHTxAhtW1IETLzk42
QoI0HHNJ07Sq1WwVl3PumFnRKp99QLM+ICrisTsH30FT8fLPl2Afos9A9KIP4eab
afW0WCGUWZZFdHdwHYyfL8Rr9HZaO+H/CvsxvVeAc/iakez0JCCn4wzRVDbhHssY
Vp9lzHBBHsdZqJP+8f+LCxlhPY1tfObj2jIGNABc2ybbrSt7xaq+TW6f3zMRrhnv
fXHTXM01T0FNStwuNwUtmHc2oyoFrcHwwJNDAX0ubvuqBuOPiGPjeNRZVdGgBDf5
G5RRum94YUDbWKQslH0VR9adOPYdKYZhDFHYWvywZSvwEZZCRBIxjWUCPPDbmdvB
sdK1US1s+gQpfGRk2xohRkge5oYpEKlET9s/CJ/IKzj6btZ3oeMWbTDkSq5+Z++D
h/Itl6crPH/4P3NsECXJbmUrUN8nskV9V7g8bKTV5EGx0zVaXqqB9zkFYQgmTVb7
SbcXGE3eyBRRvDXXUnBlAnBEmXsXL/zPP7JafBfGhl53BpJ4hRZa17iVqWAcs6WQ
tS+i0BnsGBOQn6wBvz6QVF04ioeEJIXpBYhi37BaCnp3Zd8XGOQ8fCOO8L0qmLNG
OOEVq2eho/Lilrx9l6FA22lR9s/SNbsYhknYwF3fMu/Qt/A1XnxMqoadeoUYAUEw
l0ri11oTQv9U4aS1XVGwkbWzg/84X9es3kX/aVyFgxbhIEkTiemZIEuttVZNOWZs
RLFTgu6+/IuwJsEfMXLsWKUMKHVL3WnV+AaMiM4HWPlsJeBL0abGJnXA8+YUzPP9
REQ+gz5ndOu8cWbcWGIL4VL/BxbKBzjqHEdRwfVUhetzn+aSLjyxJETFKZrnHWxx
VhvK97pZfibT0etETDhdi0szOqZXy4QE8hQc7K0/LrsfQO8UJX7eto3/KBnCB5BH
4tVZCn9OYhMyGi75kbNOwnQy0fhlxkCAf7C6NkjW+XMzTdsJ5ko8fWDhdWRiiIyC
eTai+eMSnAsy6Gf8RYnJmqMAlQE+YIsV+Ymjh5JjUNHEW0Xww/GCjAobUUu8GkRN
bdXDs8nVEji/gpVZH14mLuJTGmRKYghM5718MEfy9uau1lwTaM4xGP0yKYN93afO
k/T4bu7UfFe/Ou7DNCeFm4A2PWjZ2mJAvkNlAEN5TSfL9PqXT05zPdlIKdWm8khL
F042AeT6163gS/UrICsuEDPgZXNZqYCD4N3gUZPMqqKOrzxMUp0hYTaYwm/T3+si
qk4iEVt3SkDdPeOeYhsf+WFcnduDfWFaUsLlOikFWEzWKouzknoHNBFTYsP+0Lup
I4WAxM79Y8qistjBXN/vwfhGVmlm1lvSmRnXgU+zPXfQn1osovbTqenjIGRuzeK4
derPStVwYkahtm+fTTHGE8PO9WVfYmcFt3Fktw9s+G1j7CpRsegfdWgcABBNI+bA
U9kIM3+ENiP+dCpgqJwcXIhyGXu7TAAN/CDhynONv8pgJbgBd4gtHu40ZXj4yNtE
ygkv+ijB5MIJpu2VUwidmI1x9IJqO2TQIAu2qBdU9giOV8VPmiMglXEx+jumwM8n
F5MK3nzGQUwyzzOMjOXiay+n1vF5o0OeZ6/dMNkoTbeRB4/yz7TYY85ue3Lp4DTQ
4Mb7y7of1zyKbi1LyZ/PT53LODmfvVprzq4Ca1eruLwsq1BZuy35cp6RkqcST3o5
KYCwZMUnYnz0BrMILX/HJTu31zU1WO1OuYuoRg25j5QJSPddLJsPRpwdrW8vrkvq
5ByJg48jbCX791CANCaocsQJUWj+8aXG1SJVW2j++adRdEgSmxaealNLI1VhoUpe
+DT7VAebJyJeNBA6ZBRTYQJGSJjKzDHYYo4mf24p9nIjmx0rD+45a/ZZEee4+s3f
KpGM8RcF0trbQ53WpF25QQO3h4sxtyYyjprgAVna8sA2iZB85fwe+5cVdo6OnfXJ
zo+POFQ0PB9kRZoTqbRpRTlZ938KE76Tx9xWr9KxCGeNwMGfVC3Gx99KiMI8WFv3
JDdMBbPWymENq0pzmkZlOaOx1jSrUtGZ0iwnsvjYH7r27DGxt3sSOSH7V3/CSBTI
JvwvmAotZXM/7VFXCIPMmB1FiXkJ7YAAc3kbH0u4jeBsExqwGNZwHLVxGMRg+ZsH
gNStqt51ICuHPXNrBozB2bPBQwiVSLwo9XqLqVzm7DILO53fH/tAgO8vAHhKIQ5O
h5QdRCpsaNiCt6sN5RI3Ku69M4FwnoJr0GDZzvegeNxKOzBQ9meWGpOatSXVzbJ7
WPh2QGbDx/WIYj7KDrFsmsyJUANPiVjpg2U0E8SgB5u0+icAVh9/Eh8exdv8LORU
ZVVaAhbRrUMNlIvSvoB1AxdoqrW5dvXf79t2Cuwh7uIr/+jSbi/qIrtPR1l6+mkZ
9iu+SYAEt5pGcvv4wcFa4PbYKGylJyqaBF2aqKJX2L9C2vhYOrtTpRq9IdvhJSSg
G+rjocpTRIsviEPkBseFYHcnXS3DWuYiAnuYAI+l0mRdodFMcSNpIlRxPsycrkvR
lmEUcEozkgdPfEBkz0G5dVG8VrQ5JcF/kAiaSt671FJvgncUDAXCLnilj3/AzS5/
UnoCyewpJq3IypJt4rkfSW1yUwrq/J1AFEGyJ9857nm0wHRPC6TkBipP9XRMDbJr
OihvOEckZse5C6TB6bLY1nR2V0g0c/opr7utX8Zla/XWjUNNi7lqIunnHSoZYBTq
5ZklBG+ZGzt21kDpge5EKVldnnlQQRZd6X/Br1V4yTQJX7KsN8lBKnUDAH5Kq71o
+08ki3WLnD/sxK+ZjS/WvvI1QxsnjQrL6NWvet4bkOd+Wvne65tD/S42pGMUQg+8
ftOQbvwt1A00COY8ryY4GJh/WMbDTA8/d/CGzRYcnj38DHbCNw0cRK55MiX7IhYN
Ls/YYOKYMP9N1TR/aeLndKT+xc1zMOcb29mqc37luScpNhnMW16ILf2/NZKc4P28
W1qMheM4krdC2QDMBWrDskCPpVa4hhfYcyaolWe/94JrsD1AyfttS2AiVFagh4SB
KoIn6K329Zv2pgFDpxzZnlGR+sJdbUHgik9mEG7+liw2uLwMr0wjN5TiT8vyPKBk
P/kmMOA6cy85F7WWLMQxTB+VsfCgUBgfJAcdSwfr5rgn/DeaFXymQPhIJmvqUDyu
Lle+o+KHJICiXi1CH6hb1omNZ72Za0eCouorh1x/eOlvDx9LyqmEC2xItt73/p+d
NZacPpD+2rv+DWN0VetB2FeaISlIH8YFpeUDVLMszWg+zXt8w3hRTdcIn2b5BgKI
hrS2xKRht8fQWL7FEDx1SpvfnHzKvq1pGBUfVQFueloVZgf94QgeYenIZ9JOBzVz
6yWjpT1OpsFvlfXdRgdp2DcoOyf5V45k5g1aSHxmTh+9f+rGv/CKWECOOLCfkGLO
Kh0LKPIFiY8Z3sTuYFx1cikZcodPVhBAZ0Wl7/2qB/DIF/7VSUhmxd42BAxcRANi
eGFhHpMqMrD+XJ+Uy3V0AE7HPkwyEBe2+oIxqPM7Yz2FhdTln6v2DUNcvY5S4w/o
ca4fh5FlgTd6sl1fb9dwiSRml5fwc31sO/d6D0F2D+YkIIlWdj/HIXOO2+UspxBF
qgIPgcPkdjt875kk1GmtB8W+em3gvCTcYN3glbQf9Pd/oHaNA9prhJKLG3PE0BuN
LJSfJmjk6lWrN5kEf5hD1RW8g83OdoZE8me6C1qpZjrBMQ7hj+fcSMR1PpHQFDs2
ZWuCaD3gYhNAl/Mcm/UZ0/H4NfZ9uA6xLOkQAnCgjXccAMu0heMG15JZXWOsmmKD
n0AVeWBaZKDk5Vg84ujzdDCDizf9a2ze3jH1pXk8DuCYTOkerGU4XJBmspVPS1Hg
ElgpLxrAu6InDlt5+fTCTHgxnmInJKp/eDBjgX+i29Xgyj0X/SoRdztd5wuMsbd5
ongfnOaC0xePZ9NwJis4MvZxVLwqBARvJTxL9gSksJ/3/LQwGT0ihEU520CPkBwD
dZtEzpvEDKhhfcEbHJCqkUhNRIydWVk77BxU+wT0qQmZtUMBc3XqdTL+MTBMJ01d
adYuUIIFALncG6UjAa+sTR6G2rQvUMjTRGbqUGupe067gDrpvqdcjOwVTzcCEyne
gDo+liWARMv3V7UWEwQxKEWbwiKffjfqW42cUF3eE4EmT1LpMgAathoSd2a+jSGf
d4nkk7mSZshRAoh37XyyhgvwavP7pIXBlvBH2wnoiFDUMOhbMe1NSp7SLM8jJ+/T
yaJ3dMgxAnUBAA8OED30/MLt35N+oNyIwC4llca5VenGIxVd2szvwW/wwqo/wP8L
Ql7QN5gITK5IfnWxstrf29+gsARUnH3SkLrqcGQBQZtHL6mTf5wzQM6lpU/1vcbQ
IfhdKTVTMcGzEyCLsqjNOxsm3PdNbXRJmVUCuab9VKwU7Wv7PoOj+cvLFXOOV/G7
jd6Pt/4iMBPcMhqhhGBlUcnj9kINcvHn58zmpd19x84SeYnHrGPXwluFVE273Zw9
ZpUerekHIH+h/gK37fjeYFrxIPB0BT07PucLBJPOstVuG8T32WDqu9uy5oMypDru
6uhyOWg348MjAamSXvlwJqhAoengtz6fiTy3bpVYs98q832DB+KvREoxShkH+Wrd
Hw+NOHgbtAPTHCYubtGa4QMGI0B0fyIbYuU8SLsSPkGjLPnBu+Z19yU9/d+QN1xg
R2ZC1Y2UD8opUNNnUHWBC9l2etbEz6RaALgKJlWiCO/dGeKdHMD9RfshJr2akrU3
Oz4YHn/oi/aLxkaUYxsZGJpz/wEns2iiHJa76VOQy/xdT4qUQQ1gVbAZxymmTshk
niYHOD0Xdg3mYjqxGXAJ+nYspaQN+LUTRShxXjQkPayDjfc9x4lTsHgU9zw3shg+
CQKpI4jz+SrrjWBewt7WiHBsN4KzA192PgOPrhwIE5fMm+RhgQb2e5jBcv5nqdc2
oFN9FDcGe0oUJnvuDF7gS9oy566qtbmn8R/2+91eV80p6bg/czWyDDMQWojvRut1
TyP0J2UpZVTcao7SbjzuJ4nEzLH/3AywUpfBDNkLATAq4XsfL67hfjJc5s9X3qMQ
YhvDf7SHO++69eX5cJ6aL+PeY4uGo/wMbexSY0/Yf+tdsphMP+a27FsbBF1fTIJa
1HgyMevj05IoChiagikQBYQQHCrwqljsqjY+6fj1VUty5crWxNy1nF6gd0w7l5Ux
j6uhZSks67HW6lQOS+3a+t2hBquUJc6OBH5CacUf3d7+RGw1HMSta901Cv3sMBD7
Dy/1Gf6sANh95oO28PYZMXRvZmdAn29TlkzgP1kI0OepPs/Hdxb2MEpO+NZ+51iv
C5vH54VM+bSZ45VycQgsaSw3FasIs1+FUlyk0U5IOM8bJtVbM0DWmq6HdzK801cW
emhPOVRL4C97zSVVq25Nf2HghTUJapepIIjjZ1hHqXKJibL1IICBBVhMec4w4bgZ
Njf1QE2pQDeabTGmPii7UlRfVX9dspVGFPcUKnBOccg3ksJ2rUebR1MnG8R8xn7+
2HSNaDT0vGSeJYjl+RUiT1rhF37Q3jGZic/jfLp/CUyS4BoLFvdYXPH0ygpuT9Yj
Hmjlh+DqLJEpDhrTQlcN0NIaRvFLJzTalZ4z8RSG5xhbWEbYZwEQVhHTf5TktXSd
uLnE8iQW0kg6KqsErhbHmbkUByQN/hiZdopxKyPj+mDPKkCi6q0y+Iuv//AML3jF
pViqfMAnpXWitA6SFbg/L+9k5+RhqMCIkGmJrO6+cob2CbpiFmGzMeG+EpQ1J0El
A/Dml0WCEfEucER0y0nNncbUyDaIpSYPibeilIeNHV23uLTfidRgrWaC19pSeegY
A1ZXTuDp313FLBVJuvVXQGkxT/u4vel5SO+0JrgtPlT9n0dZVshz0gN7qUA29ATW
PLozJBzu4Au4lrLZWZeHGUD4kv3lnQs2B6qrVQmjhdJ6lYALF7IYUL+qTHR57qU3
J8Jr2g5ga0ERBexQ8aotPt32AluFSx9kAl0/MsT85Cwm/xCBzHsopB2V7aZxE7vy
CGvU8yARP+RM88l37vlDOQoPV0TFuv6lqXMT/LLh6PvJyH1gTNGOVb+jb59Uw1Zj
omO6vdWt1z2WAHE9IoMxO3HdHEmtK9Fby5Pe3dc8VWrNAjsDWavviRLRuN5vOaRy
oVVALp5qcxLqd7iC6D46bqIqaWJR2VyeSx+AKi/tj2XgvNmFRGNr7kkOIo1bp9v+
fGgJBvMx+Ri8ZOfrwpLoBfbXdxfuAC/SOgD9vgvWgWULS8mVdQWEaFf1oS6mz5Kb
RvkdNrm2/gnVUN2uc7UYpsPqe89XEsvm9am0qU6CSOCW77LIanTOjY3ufFyKLkOJ
UAAq4R00+48MLj+/5y8CKpCsAQ4Juicxm34pXJcfc/ztJSBCl6Kpg/X/KBXVHwd6
oQePWlhdKOQ60DPNPqZK8ExvQbm+H46oU3Wgw4f4PDFEF15hY/B3ONHQeiLBGgeS
zUZGHlX4+G3vTjLE7PJ/pL5NQ1N1lbuS8sYxYUTOAJlyJswCKcntGIaBbml1cAgx
VVmuH6sHtO8QDiQPl+WhXYwVaXMdbuKq3Ak60glosP8pcB3CLZWiYT8fVZPbcucq
9Q7EFhL1sXB0SHAC9tx4zCO1hvzITqAZnewrRmreN7K3tDiDx0gtYDxPBomtvgv0
rE1qTYS0G/M1ZI1RZisfY+Ero5Nu/0i+bv4cVV96R6j4gbpIDNsbqNkVsTXjiCaH
oNTwgWu1mh0nshtNzrQSc77TeDrwpNBZoJeJXNX70c5NU3Tie9IeMAKfPZCh+K4d
NgCna9MhtIssStU+dOnY3VhwrUV7FQPROfyQoldfssdj1nrOVICAOtWEiAiBdwnd
nrr2+s30cJPNXec8LfWXddesX80eSKhhdSJqVeG+V1bTy1/pe/nIm58ZMKX7t5GE
oxVk6UB9cZoZN54eSx1J1Z0AApL2Wi+wSogOO4+XLFqvAITcDhDZZ0jZ2KdNBuLK

//pragma protect end_data_block
//pragma protect digest_block
+v8JIUQchCJbDaIBs0956Zn14gk=
//pragma protect end_digest_block
//pragma protect end_protected
