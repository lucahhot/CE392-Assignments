// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
L9evczmChCH1hiJTW3uQwYR2SJ3yC6sqk5RbLOWgFxYuUjS7+P4cEDYdxFLVWRM6
5XqhV6M49X1DJBAE/j5TFdPI5GiGyu43C9YK3DxXfd1BK1/t3Aqv4QjCtHje7WFd
+zTKovgTTGFyftL+MVch9WLkhZldICVrf2Ch4cPumlc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 15408 )
`pragma protect data_block
D9jYMKAOHVBNLbdfy2H36YCh8q7WDOcalcY9VoEnqWLIuYv5bC4/utF0oUhI7w6D
caqUSGLV5qEQI8Bl15BFSpZWj16GazWY6wKpoB2lEPF1D/N/jTcPk/aAUv8D2OM1
wDuUWGeJhrywCNh7f6/iH/Lh04eh9uOamHFbFdvN5Z9ThRfhrqdr+WlQhlUC4kDE
9wkRN8zQwXs9e0Ns6l5KZQnn1+sfyyPAx0og6cCvlTf9OxapLBJAaCwgElw5MTXU
UyjCGY1kAU6bOOBArZXxaSJqIf5JDu/rKpfFLFbf/DFWKb24rCBZL5vcvd+m82e9
95XINP3LAQ+uMhcJgc+lgCmj92b2rL+cgkcOy+a2G55HgYnvwh3vnmJYnboaKYGx
oHshqf0a9PINpdyw/0NoObP3b/62/jTYOn+BBNygvDZEpvmILpEIsCSrtrWo1TKo
8d3b/X2VYDp5Eiy+65e062hNCA3MAoEUTJrOEFH+7QuML01PP9ERK/2/kI7dfCJq
eSZh6iX/sLZgG1zGNizRsPWE3YV1MfsvqL8uQ9AnKnaA8QiReG1h+xQ7AvDoWB+/
CESo3FVIhqlEWAZ2eoJsT1nR1jgucetqLGr9MK0WmrhB07wnWkFoHFsXBpWcXOAj
cenSfayPI3jwOUqXkuq+TC8P7KPO5zzYQfE4zyvZLSWQ6r6MYqS8/eDv0q934dke
yN4L6JSdgVcW935SyhHiVWaRRoM5e6NQrJl8FOk6IiYHAlvtes0RYIIgSXbf1Zq2
4tivseaW9pEu19REmW2XZPTFf2zHrMiTA6PCLfAQ1J70L++NAe9LYkVQuF3epL0h
Yh6tejN5MV8rFCngiYCTcmZJ6pwn8bqc5E9Tnwt0g2dqQa3s1Pc6y1bLzpuK4An4
VZQ3hE8ExlPTUKvNW1BLocbspCQo2CkBTGddoaKAiY/b/+1CZ/xCsFwYpF+bx4PF
n9d3ExPOzqqT8LoO2geXsUc7RoWUCIc71F+5LRVnrEnBhZrqrCiT0fMaFhPURYWI
pRArhEyquknAz3LRyluKrECgsqRnGJ8bpoGHeyjOaAg+I2Er+ozT+vfgG7eLf+d4
81yYDy8zD+u+fT/aFZu4bLbDhl6LJmrKvG2A/zmYO2q2G85jNPu0uhkGgqDS6cmt
yTpr9C43rH1wQ4C6VswqWfvN9U2noGIV8A4qDBo3OJr/zMmRA1S4YIqSEeLzfREP
HjSfPUiDpIDM+/cketcflXgxds8OKB+LIlzRgYuID1dPHKaO967THeucspRtVx1v
XMBfWGRgf0sX6y5T5+ryvtOJi3Zv0RhUTbXKW3lm7Hs4WDXOvGDxvK8ypa8J5SN5
h/jD+CZ+eaEhSknlVKbbE1p6a88mcqMUUAQVkhUdPv4/n/WS1iFqVaeR63shkSNM
PEIxWGGpMsAnHON+zayce+xg53Dsr+iHX3qVAi+RXGRUWfwW+P/sjYdcLhZGS9/G
w4/bFdL4/i06Fj8BzsHhvJM2xnLmnEY3GiNoamuru/6YCbPNtkMqjKQfUuTIyrPK
+988UOp7xv7pkWL1hcOMk9yU8K5sCVcFFR8RvMCBQWLWudxF8kC2n1LGlNziBXlr
W5Hx6zPYdkVGceyTap6VwxXy8UXhIELLrldbUZhi8bH/4bH0oRcB27ZPDN6xPjMq
NZ8q2TRpSvTbALOLw8evp6tzm3i+RU0k3t6u1LnsHTU3ndwW9usx6nXRgXCWKy2m
UCY7DfjVZvX+J74wM0UmtqrbqceLufK1WCHXNeDmAqwRQAPw6o7LqpJtgOhPBina
pjwigNx8c15zuoOvkR8I6IQAkZ3x1YwR+qqn945ZwLYLZUDCgLqNVLsY9gmC0jQ7
UonIt1XsqFGdXbul+mZRbUnI0Xnf+dQWDcvDqiLwnvDXd6amqVtknhr6oHZ94FT1
cRtuwOEHhJ9wZBpkP59sEVfLJeyDcT69DJVjd+jtTB1o9LUWXEHtWtthRo+x3GfB
SHbZEYDiwCjhAJfsj/dkH+eT7BdfRklaK6OisiqAl67PYSofLAz5L0+cJgKRXuhT
AyEd0/3fV1mdj7SWEgJLmwxNOi+MuRkXjndMgnaGIBi5R6c4zUcbgMddtAMyEPcp
Yk/P6iXsUvIj/wCfSR7X5U+mq6ZKf2oJvqPBSNpaaFEEfmmCF/dKqsZ48F0TuJk8
lHzTdMc5U1HyJsUm0y8o+vN4M0VsEfU1P8ZD4BcFcQtKRygq7XZl87qbT2dZfnDQ
8ixkUwxz8Qy0X/eMjcISDlupGlM/5YoAM9ZUrs1ih1Fabjg2VwhAImdgnXpsLZsx
BPRPHJ/6HHKVgQzFdYOR1K2YvEsBz9PBibFxgGE6xhIt6051IXhd8D7uDSdcD+M5
eaoEZXYmWLu4RLzkl+EQc5jB4TVpdJ77ksGrvcwDdD5UJ0bThWkCDOG8liAnKUh9
HjbZbFmpMC9RxdW2HIJexJuNJCSUPXA2Emv444YvwqDIUuHBs6Q5vuWU7HkAL5jE
vuFaa0L9IqYvh20vjh0MdQvhTgV4g1gRm8LxUALPb+jN8OASOqU4pnEC2zuo0GZj
PeK+eu0LXhBM2MfuOlZPJfvQ93PMTFWt9G64p7UUdYD+4/VsBewirTQqN+UPT6d2
gWzQHkrB7Iuwgx3BUzr6fjHMLJV/+FNvYdgWM11y2/Mf8JdQL/zZW+/YE8AhWiq4
+uUrj3LgFWuwqC4hQWRw0W+OpwkOCQieBF03sbeZ8U0S8x3xQuCaI9z1tfIf39Wc
TJIubnsGI5V6JRKBnqgDFC6DgZ20+Y/6ngVrp58FIcvFRW8MOA87FKc9WWWkj1wP
QwF3s5soye6GQR8C6uXlZWw45KBsTscgbWKxZq7jnlE7PNj9KIKSarAkfZuJjpGY
11iM0Zz9x2tYlXiOMkM0FMp4E9XTjhNG89L7HsK3jvdH16Q2DJJLdQMthF8PIw6s
DWrqaO7okPpHYhdZX9SIj4Ere/1cgpscKKZo3XcA1qkDDhe+J57LqN7ab803sk2f
N1l3Nm67nTDxVqH5ZfVMVlRMUayWM6SPNMz30J6mIMZjpyI59pqkn5sBnyT6961/
poMjRkXS7CvlzK7LxXMBW/vp9pD9BT1jW0oPu+IbsjGzgXgA7BRQyQ/rxm0DC70h
Y4kAhDrxMyvXJF1VlX/Khm4kvdyxS6bMm3qOTdMdYmmSxLDLBUGzU14LFeNY0I6E
0w+cvftWfWTzdG28lHQE9eDBrTiEQAbfVd0KBr1YJ86Is855wRXzjuOlGIxTDidi
HFsJBBd5+eQbbJcg4fZOLfY3ITlEzdjef2R2WZZ93zwXCmLUKlafkJiv6SB48UiP
itCWpQ5OW3I+H7qjKn1heV2E04gr1qwoHqLS+4Z/M/uQq4Zi2cBfY2+M2PejO6Pk
7CVB7/KQVsDSM3wJGjCRdoHqswMyjZnAODz+0e2X4pVOoJo54G3ChJuSd+sI4eUG
1YfN3pDrOGG7DrTV4WQaNDioZ+h7OBNZc8Ab4ihNBMjgeup4XFzYLxEzwLPOB6xQ
yQyISqPW6Iv1Rcqb/UpK3UTYzovLSUvHj4gco8AWA4/oCB1mVaLMHhuFmbfTk8r0
VxnfSeXghp+siECjmSwSwETLKOja5J5BIK2sBw2QSw69Nhf06Xwo2cQBoPnsC1Tz
SMFf/k8abVpiPm6TSXIKczKYZv+nGY4mPrGQQ9IPelGtFCNN0uT1HEFs0qhAnB/A
ByFZjvhXSMZcPed7M+z3dpX2h5Tz4kKDt1YM83Thg7TvGUTxzYW8yUSBTUgG7Vkq
mvPeJuBPFOQ3e5VlRJeNJ+Bdt9i8f7n1IP8rVOFhZ1va9c9S21Lci3cxnFCpp2RP
Aasv/ZE2uupNhUyOSgKykUJZi0XxH7je7O8IOD+nTLEMzCAFbpJE2j41I9B4jAdQ
ipnKXm+5zmeW17gnQE3hJxo3cHm5xUYRGHUVJyXdI+9VARn5vsEirdpMtNWNXflk
Mviw+ykwHqjojbFxt1Eh7UWGBUsIVG4l4fBZvq/ZjfD2OjAGScXoc7VJpwYx+zI2
VSqAo2p5tLfi3d+pxSGQmzJMb+VsagpElAE3JZhPVaHUmvwR+sn8HkAVlJcalf/2
pkPcMAzf1WNDQniIZdqmesNynzUMQ13JP9y4tijMKAfOwYUmdsE5//ngkfBf+31I
4B4ge0FVHTXknZosb42Rco8DhtEWnGd4Yb9KoXvb8ipuciGvnCAaW2GTw3SG+Y7s
pRuNOqYOxjhYc/0sDkDbsWrulbYMBcX0B7l9XiRbayWV34+fFDO1vEBSZ9dEcV2+
5lyF3C5P7OU6XkxPcGkroBGLU0ZsRl5fa3lmWcfcXFjQOf+sppxpnSHK03UDqjzS
z/cAOgXUwo+tKBHodUB2JyYWRPSzlUmGGkX02rZg5QQmFu+lTxyMHKo090Djbu9g
nkeoR8cHFV7jPs/qN562/vlvTSnElLFedWGLis+jv2Hq+s2/FDHHR0i4RhhK4Y6H
GpIu//kQO3oiHGP52IUp1mrBK9gwLAzBvJfU+h2yGCez0GcYF2k3vPyPuqlQihNF
Wf/LCEwi8hLJPMhz/IOA0nF64W8LDI5SO0yqBZNT0P/5Zx5grSx0MFNapsbzdT+I
TUgJC9lvxclfgdVhTps3EQqaJCqmneBd/mv63pTcbFSPkmBRKvD88hAo9IIwDOih
XlyeMGMH6n0d8WN8LBNpv01G5QyfLFgAhtUAr8NKkM9cjpMP0WYRb2i593sXD/lD
0N80+wQKrfJIIE/6sdOIBOlpYfVMdhw9LILy8P+r26lwbalagOVCiV2nSelN9/Wf
11VyinGRKLktazB7iSf57zGlJxZhklHwKxD0N5ZWMbGuRTd38X0mzbf9GDMMg173
OpIjxmTKtq7qtnNdyGvG+TTMPr1Svsgj0Pzrz98TWFJcjjLGihut20KW6/SnAHXy
NkXCRd3dRVCCF+Mdc95LxM0j/oNtKGHvtqYVleiaxijjBzYdUIV1hNUBtt2seeLD
vQ/BW+qaDSJSoJR9t9vJEmArrXu4WwGO6Tc68mNPeXKC6mn+kdsPJrbVoV3p7+kj
reuxOJYUjF6+1L9WWY10wlj2bZtqmOX/rM/tmysC6auBrgR/jbjMbB1EkyfX+bNR
D1O2mz0KEBUtvmMST8GW6Pahyl+DAgSXvkDk918UIkbcfkiBNaPYeN82NOg6LlGp
k6pud4862Yckp+SgcPryZ2GEMwJrB/wgKNfGgiBv9WVV4isqgiM6EhV6Xs9WOFS+
0kPghTghoQ+4FIX28DxUw5IsUEG5HHDhfx9hKHKopvG8IdaUxbf7dFxljN6KSWxD
26cSkh6t6Hq/KA77KLjrNmCdEe4doMqsYcDI/ityE6hupNbY7ZNOMDlLjjg7n07Z
bh0a2On0MrgVxJNzIQ1bUPOHuKm2sJlHtJtNNy68iNpC1MzIwTV40yNw2XrIE/De
r/6Cjl9lZxIdSIdc4NdaQlrcgeEFhZ5X/iwyQgxSKu58oL+5zfFcDEphT/Eo9nbo
OBqWZrTBfJytEkWzVRbAW4v0+KSZ2itJcOX1rBcS6FLL3fvDqdGxJ3CwHByrPFOy
8cON+GGexg4GRJ8Lax9iq8aYDEtwuQYjWy2M1WbdSa6lq6aGuTnQWn5PcUB/u+mL
RJLBXxIzuTnEOp2Z+Y18BPtl3ntYfgHrNYaQeF3no5MtaYh6WHIIOqc2CLxV4sK4
nxl020pyx2dim0WCmNrU/o5135IvHUpLwBPA5ZjMEsl33z1xr3s6e9/2zZjCCnsf
PSynmEIpKFrZep8PVHADqww9jQ18tYpsZ31CuFP57gPCDavKJDRu/k67vgVlDRGJ
VzVesM/epx/4mXc/HRTheWpTpiAWxM45keSeIU6x8SgROl82Dh74h7p2lZQsQ5yt
YbwgHW+1lAdUukWswB3MwldFFOv1SDiCqq9bNNVp1bY1aaCyOZ1Vs+OI3G27QLaq
dca1hpyJ34/KWHzyklge3oySd1nZK/tNnvU+jpTpRhKpXwbNDgIDlQTruWDF6LeW
o49sabIKInOx+/sMlquAZWMvWZ3cvlrUH219BTUh6G/wiaj0YDKLRl5NR8peTII/
slWPqy98yTiVB+jkeRTEgFD5jGpDp4ZWQXz1orODYfp7FjUxHGahIK/QNK+D5nNH
a9nibKGs2zJqngZ2bgjGdXO+avgF3W0MRiybt7gq36QHFlzJQk+rD9IpoE7k6AzH
A7mMe7HBc7kl2Pc4DTeZFNkj0o2Nn2hrhSKi4V53qEnJiAMmayiZBPwA9mPyfDti
6itWpnZspeAzgM0Rh82c281Kx1SHCFLQgru8XWfoLzZWKHIWwZtVwuQ7cnZUdHGG
Eh5PTbO2mhNZa/oMAhfYKrAgrg3U1u9VRUYkKnmHacW+Q2X2nc9j8RJklfvyyTXW
MCL3iJW0e7xucP2LDgqFcA3y7UocValgrPc9GUcmGZ5kHvzvbNpRZzZmwLtaVySg
BJBPQkJton4+XQz/AeMk1N9RcetALD0oBrS8p9xjSlukWcUtZIquUCpqVjcpRfQo
5snu6+jPASYfNCwc/1jajRhRa2/T8lueyXFI0xfB+0O6w+cFUyIj/Lpr00YKG5eS
EUKYkbsrl/nY0fAnx3kjXvouhStnzJlfl4ts11Fzk7Ss4H1DyVbDbLKkm+NepCuI
JavJ36jlQaYWQkaPDakzn2y8nWKLR6HF9gIxGXmuni2Ya+BHUftht7yZRObyv9i5
E9D+A4irMn2/PnYFcWyOL53UEwKDM2J8fzR7deyCh7+2+113PFPUZd02+VEtDDhm
M2KfJ7k0BkTQ/xKVc0NQYlV6pGOq+wvOPNlExMIgveawJoQwIviFeUvRy0BnvJZQ
k4hTCS/0Qh9o0Ek/ADm5S+VrgFj0jkMpyt5LuTROlRkfXWZyhaCgSESjLmp8EY1R
UrT5Dn4JY9LFIiBg9v2noAJynqLoLsk9FDo6ZKkTcCCPO6m1WSQc5CcsVQdEoHlX
8wRgAqBCKiCMLhySHeIbEYWhWek1Hf9Gg6wixPpne11A6afbpz4c2OYmLE9St5a+
UYOsmfuhlbQbj2vuiJOrCdGvmtUea9R8AmzhRMC2T2B9K57jXfC5ycmrEXVQg9MD
w8dYkuzcb+/LNH0VZh2zJtoWMBkHFxWfLenTdgJtnCCxemFQ8gsiAyMNF4NUJwsT
hjZYGv2t8WQoMHSdh83j/N/zvUW1o4c/ZZ29sLGr3BDswhVwjkk8IP86XxJg0Hxc
w7GeX28R1qJc7ZKJmT0I/Q6uS7PycxSNQEYmSgcUGxHYHCxNoU38b1qUUaoKwcCL
9aL9HEPeW7XWLP+1mkx/lS/5KvrAqC2aHACyfujkxG2GgMAH8y/S3lK2Yua0hOoj
qi0ZZ8COsYKNfgSj4xrdk91qKLIKeGEM/mY/ymIMS3VqbglvPyHnzDbaEB8cAbKT
kP1M3w9D6Bsvhy9fnmQxbwvYsHVkFVUlZR2HqlOIR15wVH6ghyX083Ux1DMqgL81
yViR1dS8gdldpNpsx0e+r4Szn53v0Gb/QvtLNuqSTqnaHkVJbiBZXCs39awMLo7u
FBspmd86u2VjPIFiCbFa6dDmAzb0CmiP8BPqDu9riCXyIPdxNMg/7x5HiM3wp6CO
PSTUHw1aVcLZJiQ6GvbgCHj5x6LRQNjTNg9UcdZaEmJmEJki4PMSEGtdcNmfAted
VJKNmbtJ2bhcTUiACgRcwlhcGUOpXHmzjZudgWRcoG+LIQ+BY5BoK1IEt/pHIgkV
5jfRTInhuvH1hD1qYY7eTI6l+0+m6oNOqxojV9aJG8rJn7tgUXJjAw2gHr3SIeqB
Y12WmLeJ/LExmXl5N5ZnlxlKSKd/natDoK+BAzmK3nHtU4VsQ8gv3MRceCh8LmLm
VeGJKnfB5Y0kgid1hBgFj5fkW/eEGAyfWlEIzXPLWV3iCzep6aIVcRovTQ3MC/pk
gV3n02QP+jxb4dbGp7zRchOim7JT7NvsG45bDKF3j8PsOOEmPqin9iEwCwg4PULi
cZ5BaMa2u3L1UcRC1ZFzrHqCbEDgPJYYGCB/z/BdhYRPQXTJVWAPO2rlLMifAg0O
wc6q0sbaGerjGs0Q8JkrIiazPkt/akU43TUU9WTXllVTMpYUwDXHGRmFRltuq0By
YmLjef+1aYnUchrgQRA6dRKMLD3zbLxgisNNiqLSuTLKVrOcOEsyz9EgMHjQsdVU
RqUmhJQG4l0HNSP9XoS+Teq9gFRZ7PYdIvykGmHee/a4MDXY4UmsCXEAa/6tEBUz
vwSTSbqD3a2W6s7WmEX+TVCdmIkY21wZVqTdkBhkFOi7duSTYWbOh0xlclF+KR9/
3a1e+qHnzAV2SKc1MH7WZpdxW/7ftDanIF7d+fbkFUKtgS9YUQEN5hsKnx9dEv11
nRgVzZW8Akr4zUNw/KWFMUD1ER9MTYOLL4KnC6bZpz7NfRysVGSOoKX1xDNHL1pF
PhXbaQ6WGBhADtt6/Bfuzy6AXQMqIXGvvcV96Rv3px2UH9HXJXVfGx1X/tcQBF6n
e1m+3pFUUc+TkcM7GnDLYos8oUXL5uJxK+wjAyuD/9Wkf2FN2e597sV1xwBSFH8T
BI+ZokxfIvzEv/Zz/gvoStbWisP4XCGRxoES3LqTlLhqquQHFqm9/u5cuiXTUHAF
3/O7oDhukeVVHDgiHD05312Q+g97h2rjWNbxrpCYtuuWWgqyMmdIQqd9MNpVRJIy
gU0Q/UhIsctJx6C6U7eGJ0c6jECGXLGyfsrPvs8GPTEoEmhVN6cPgTMoUR9QTabI
v2w8/Nf4jwMuib+jmZRCW+3XVPLuw4CEHnvUCvjGtmolB85d5S2UbEslWZZY9SRb
7G4xAVp0+EGX0yteZSt5m4fgigcTKiCtMB1CY0ryibUlLBaeLsYPwvTpxU3GZQOE
/L9HhH4D5ddJOJ8NS+CmrgXy2vyj4DPpHrwTuDAaFbPzmxFsDG2SullDuHvSmCUK
bxfmbHZ3CkNG83q+3DvxK/JtJgMBCQNCPK4ngiRVbIFhVd5ArqEul6DxBuB7D4Tt
SbYLm51p/ZfXX6XRJ+Q/IQVMwvO8ueSary6JfumYJyTqkCVQ/JRvXn6DuwsFi2Q0
YTZzPRpRsq589hl4s9SAd6yWQbetYQryRbOKkkZA0AUdfYyFOu0mgGNByPVW3Bn7
3dFXXC6iO3fZUUqfi23meCnRmmzogpiy/eoX7xxJzGsKkNPh98tZP162dk2xfX0+
oorG2m9M5Om3tUSHAyqlmT0THfw7778Ymlp/7jFsH3d5d+QllEg5YB+EvTfjd2xH
ZNDmOxfwC0CgNH6taBL4Uy57eE+ryyWbjqg7/N1LgwRwtUZgb7bFdHf4Y5P7HSBW
48brs3++57sC8X3otKAGuI63NWP05JfSJLRuyOxIOfTpvrI99gN19tfPAxr76nF4
6FDXp8EoKd+hpoiIMt+o/q1jX6Kq1WFkhk7v2+DPWjiqyaA429OJqDXi1G4xT6EM
RMRZJXZYCb8ruVXgAFL0RW/3gPovhQ7ghmnQ0ZOCQoXLeYa3ncl46U57D5wyIghq
jty2Uudpy9upgqKeAOSay5/fVAJjAFc18k1ALTwKCILkyreDpbLBwJ/vsjA6R15c
wfd12zuoBCbgAGpHEea3Tg542k9cubsW/5kImdyhsB80BcYBLQ5jTknKLphaVi4q
1hvAOKRwbDaLEFZJZd72e2vIh+oszLYqNd0P5LqGcRhzeZ/LqrGVrd903cyFO8rQ
d22Ys9GrER6/Qnyx9mqYfO/+79JKp/gmX3fDlf2ZBWgF6PF49r6zv5LnkF5z0xpZ
zlRMejqEnyIBV7eqWhkfVETmgHZis8MJ+S+KA/b2qzMrNaexv/Msmtvf4OravobF
Zg22Pg4d9CJsAaXKQAOM5OALRiSZAdOWUlMb1vfuZ1kfw6QF1wYQAvz00vwD+N94
UAzqPRQccpd3Kt/qCklv9xtMLO7C61qjDnSzzdQTsjgWgkYAuBM9fSl1uLJiJngJ
2GdtuczIcePdNEm3O2aP/N3PO1EWKriU/3BrvP4/T3Wdvx8nyM2nV2CNeUim8JVI
d9Og7Qo2C5uFZgGZxdJDTPyWlpphlJx35RwqQsjvET9Lo660YW9n6PhQo6LVA2OV
IQj5IELaayzdqyByYpDEjpZKLrOv5rlwgSFrvlfLKTlE0WuR/wD6KlSSAxsR8Gm1
krYG+X799Atmv2paUuEsbny08869PDzOK/d3vN6SLGK2pr1UHaZGp54EhFzy7XwC
4FkfUZFZbU2k9u+hBX9Jsqgwm3qmFLnukq/SeHF5gavwoKYUyX1lDDde339kY/Kn
oqqfsh6NsQQmBdw7DWtNnfRWMYRD+qZLlF+cSuFVgMih2+VgF28BflUpPIjYQvym
Tbxz4cFgEcXdJxufh0sEh9VlTdyu8fI6ODf9NNWH5pPb9T23+9ePfdTNTb9/qX0b
cDxYozNYXImf/QzhNPQ1ngomVkqYIp2GxPWr3FqXGTdA2fYtOJwsImim9p0975Ds
ZelEmrL+3OQ85O6L109pChq1VMAn4v5k5gJQJvC0qp/k+A51uGLuRwSdRcLj7WMa
ZspiziyYgg4DEzmYXoJdvWXPAOL+sp5tJpQFeJmpYqgD4UnAE82Df1IFkngGb7vO
snW9SlLadwtARWWBgHaYPdFSdhWbyWLWYDY5/tuHX5KuBwtRvs1QtVtBseTNjwzR
zRasLG44m7bH4zs5EUE7WPmi20ciCjQ3ycvPBVx5cUlzbvNPauKaoT/bACa2/8JM
x1VbHR5dYLWvQC+Sq9S/sBmlHWEW63sa+S+jst1kUp5DOyC/fq1hUH0xNfV4JrbT
ynWDTCvU061CPWxRlnH9BYWK/6fRAoiw/aqBjHiYG6n0CPZkkBBRYpDrT1umh4gb
Tm1bB1LzSq98/AgvZCwNEQ7hcmwhquroFum7WKM+M5pVCIGOAYiu613q7sFVo0yx
CC0K3loRzxE+4k6RTYl6u9I87qMqJfW4CmQA2n4xvmChHL1gqzHGIHY4mpZzs2aZ
l0shMxKrpPdIDD3IOOZeS5jhwch+wx2W+Xa1cB3AzwcfnmUaeyW/mLeC+uO+jDKs
3AFpJdS0gCy//J+XokyM0A14wNqP81moYWSUmJ9MtdaSqT5+d5Q6tUlD5Q0XEVxQ
8h+wdxm5VRrr4Vy/bppnxBt7wq6yPMvU+Z8jyrN6l2BiYPfx+5ct47oWVufKwuMi
rY3S9UtAtjbnktffajTXgfw6uMxuhcrn1O82Ug0y4R3sNUQ+E9TXFHMkRXI7UIZZ
D7bKKgbTzLJ91+qACWebOgLJBeuXNwTVSpz24SW94lWzIsVMkMbqCHN2FhiD8d7O
xH7oWgASnYOek/JuWNZHzw2TULAKRd0oP55ObCXaY11oZzwM644T72HKnzJYsVgC
p39mUVTu3mxzSe7XqDozFL9C9zouFfEtJCI2Z1vRJjO+2ko7P69Zqv+Dwj1Ehs7f
xXG+64dPRIz2U90RePyQmdTADuRhaUnHnAi+mSLyRA8jSGo0eC5hk76gETf+AnxA
icmkDquuSWe+ICRFtgIHOTzIS2tUUoliFddCj+30A53BlS1SdL3WgguB49Z0zkts
+O6JYPr6BHGyIT3QjeHBJGMQVObqweO8Yk+U6817b+w1bwhSRO6Enw/IIKhnjz+b
8pjhjRfl23svNCds8YaL8Wou1nOdquSRljIF4DuJwfg/a71qMjsBnaTwJ2UmCJUq
7wpNGulg+3zXY1B8eJuMrD/ecjIT5BOp9dasXzHn2pRP19oneqcIs8bHTnX7WxQi
s4z/vpmlC3ocPQse6RlUTWwZIG/CN6iuCvvjO9PPssVV+gPPcpMWnByivAGvQhkQ
x6HRIk6OGN6+g+VxmujdDCM+rnAA+isY1nlyv3iBp7MoZA7PH6sh2686zTTK/JVb
EOgCAz4x8lXiUZEar5uTgplnv6yVx/3WnVJKRv1W+FAwP9OenRYkKR1sVRVBSlU3
5LmQl54oryUxj5f+bOn03Xt10XXAALB+amxHa2GVIKuh7GFVAI5IBeiIsq3JCJfv
jGwQh+7HohNVcpI9aHJMH+XEnm84egO7VOfgfPl0beTmwZEsAInBP10DBg0VtuVS
1yEXb6glj7lHS8H/dgI5dWRVSWk36gnGIuOsO1Jq4YxwkOzRTNyIcvMw33Ji3cvx
rxTAOrTEVdJhqN7Zs+YmbLg0b7c8sbZkgF++TDLNYpszaPHzi1+GPRF27PgQ1FgO
k6mpJELY4vKg4P9ZnJAvl5BoV9Ev6Qd87JlAIn2in9ZIziPAqrTRhnlBUfV/oxU9
FMTdDakx0v/ilWNAXXlSXHX7K9e6+Q0lnrCCWn3MttvPTA1hnk0u1dSVWQ1lzNxD
EWDZI6fzGxwERgGF2iPKlBzgoaEL/0k4Ed4SmKnSzpQ7Kv4/d942yougsfGJY8AS
emRjZn58BuLhEbpnwXv9TdOOvWsXSxBNUKffcnXxdxkOAVgUVNmfm3VSwjFNeFDz
ytyp5rHf3UTq2UAIUtyxWJXIC7PfIko8FZIj4dQ3+yRVxf45VfGDGghk2LcMi58m
U4siG99UFnh9l3ERBrK6KRFuCeGqbTNkXgNhzWxZ77P2zNyumcr+/q3CvRAJkkLv
qQTSOdh12JPgvKWXUasWiuyh8DKe9cQI+GJ2Mh13c+cTlAyEY3BnmPk44EfmZtRb
cvujGnHViXbhkdYkngr0Kv1pjibsycrK6yhbInVPFBpTKT4myPYlL04TpgGJnAPc
mfxHZMSgkLX+DE7QitsuZx16HDuUob8F9+hjfKPjDSkL+4dwM8G73z1e1LCjwZya
in0e5oiQKzir6+ddPbO7y+sY2XY9LorL/keYj5Z+rR/axF7+BfOvjTcFhbk/5kBN
17waHCxIvn9OhitfSc7qFUJY5gCot0t1itbwGPUpk3yqU0b6oZusVa9d799XQpHq
jc+cNADBFE5vD0r200fx8/EDQsclQrQPCYxUUdyLXKz/cxLAhbWTiJQOnfpL7j7h
hapJMQBEFQpKb18VRiIKcPYeiqaNNmFzbCaGmwwyu0obyy9V2/soW7aAayt2xPs+
diOA72cynUkR3no6Wp19ldoiX2csMYDj7tSVf8aGcEn7fQ+v08p/MEOS9GfCMiRY
D8PCMShUALzf4wTC94uS+qVGKxtCUsTK+7hdFAYTwQdYewX664Gj1JW6ngxZcoaU
ujJiNp6RPAX/2fZ/Q5Jp9mTRZS0WKwfL/IE+iJ+F48Y3UC2Kg167/5RIrEXpSGPM
Zhbexgau1ioehlZFk6qFtM5J9yyUxvYF2Us/FkBBKN6/kqc9S3U3RwU1yzM1OLMp
Yb75S3hMROZNlq8cnRRGIDfN7buuNEox95R9twlQdqY1rsS/sACsyIVfA1OO6N0G
tAvTU/yV6kOuRAULLKHjFBqVY+uvbxGJKB6Z3YcUz+DIEGo8R4wkS46jK4CIXYs1
eIsE8fPPLzzGL3OctWohjy/Vm1EZWRD4oiSmKmgiEYCBb1GFTwP5xoBKkijoD4Vn
SvaJCFe4vqu2dF0LlXLuWE0zw4K29RdXcfYP8PQ6ybfd4hCG2FSKZzTotvJg580P
AeY6RiG8h8HxX4z/qw32xDftU6ZZZxxtmjr6CFz+x3dbCRr+ybY+vC+bmga+Y3wA
/sJyOOl4X4i4fzCQiWwIFD6wmm+6KH4RZrxHpJrij8XYwN/EHI4vMbOdMxAkDqng
83Ngzb/jIlEvKFsEFOcfDd5R5L7DT/iTpvVDBF0EL2cUr9rbZ8h0kJhU/FQOxiUP
qJ4sDtsfXVfsy1QDmbBlq0/+CrBrwvvE1OiRJ9EaYfKpWNNOiFgXJdkjRBdXj1i1
11txn5aAQy5SCRWsPaXzve+fKwX9JxUX0Kz0xMvnI/e6Glqw1SUUnoHySY6vmMNR
ZEBmAF0IpRb7P/J8rDKNzgEeahVuU1tOGL0vyJM8mVtiWMJDv2hno2zaLq1Z0UxL
9xSzLhmR1NMzuZ+tISxC11fZLAI4l7+vWX5PZVFIrumapwnGipR7S/R19UhqHFBn
b2rjkCbrBeqTkqhnEfWCMuqnuRruxKrfpp8dSWBQOfCY76kjIzxuQgEF9KlBjHlZ
sFi/dVBygfGiJVtL0lRIrkVisPpCLpjauV2Qxzn8d8P3AEbYnT3IhFdVkGm8rHSI
+Y/rKHAJ31rDAvPdDF54ZClGi0Opon1vb8jv9/AfLyRPYG+BQnLJtEf8wvUCYGNY
iHMGeuSvoW8tBXQOjbUOnrOW0BsAOD7Qhuy2K/zJvsruSh/qQE1klHcdqXUJUUM7
pyAfC8s6BlAFT4xewUKkVQs4zqTGCP0wRPy1ITh/gG1E6i2/qoHfXjZzlIL5JnQ6
80ppn3qWEPO06+UYpp14YuQNr7dCaHpqD+e4rhEYXP19YIVCVw1qSSjxPQ3nMYWG
usgBLyc64a4OrE86JQMP58K3tczTztVkkUfUgUneEuLa3fcNu3RmaRb9lhUl6yM5
ffJ4ulT4gJrjDIPgwY7niawmiIIR+L928hg4KbXIobVvw/lr2UH99RVD+ujvlZy0
Q9y9hAmUe7CZp2UWFe81YTNFUM1pq9SyOb3Ufd2tvClvUyaKjqghRDU4zg0Z4996
+nka9rhkAhOI/krEX2avmPRwGZm264Rw7mIo8bTl8153U0dVrnKfdkyhvByGufAy
dKe9ufQSDl9Sv5F5Z9Yjdib/75/xaz0WoxY7J6lszBPrOpj+dFAr9NGRp7xuYH50
n8oykOSSOafcIeBVQtqJ9xGroWe069on7hYW5kYlju5EHI/4jtKliWMf/c1tE31V
Q1ybQsSDIEgdfAkuPLVGdvYG26PQxGYkzPtuDfbmUHf8dWx4vj4lHCuyaGpQPDO6
d55wGDtHe0hTrdGjsIxSUAHsC3BKdvxL+/EZ/nE9eJ5hTvlmozigbNLMjfhY/wao
hHO1xne6RfppWKx090rvt7+w+z6BnWlhjVOK/EgCZtsODuh5mOWjhJQs5YIZ36lg
zRjcFYZTt6xJaHkNJZuQVkWetg87/iH//8KFiib9itARGsY3sO5PZAkNcBjYAA8U
vwrJc1vQwCeVfC8NH3aRqQjGtzyAv8pAQfTUyYY2utmLr5SyukIB1NG9qfDTxxgV
JFPgXwpwZAf6ZG7Dq4iYP/rF6gVFHRJlikHNIhedl2LPM8a7oRdfFZdig7VrG33B
LtWEVcpo6i3Px9w5jKnDWUv0DSetLUR/ZY4yaQ/jw0Xg+peoUQvBkvwGeIh/mteJ
Gr9gK1w1JdkcbElYCtPKsFGg4VUcPr1xCq9fphN/WC2xA6zFJVN725o4u7J0y7LJ
uRzfWIajyzVXqk4ICBhYNBWMXR+TncmW/8vbcQmf9QPwLDnpWTEmib0EeaV+2qKw
DkjKGM/bBKJ7ETIKtk+Ea0vxBqh/S10PX0HRanqIxDjaYpfEdNsKbHpFzE2Cx/rb
J2HTb9PnuzaM97U8OMRA5GkwbKP1CPKzv9HlNpOLo2NMUfdTToB6tbwYOszvw2ZB
toWwKm3SuZs9oEEUATjY39dJmIFG/ZzV08gsOTmNACB1YX9iW1I5zsBYuOljfYRf
QGXICA/oFVxHJuYkvJz5K3Pw8qDz+ALUSTus2xYr38pioZaB/71SprODAvQDLJxJ
j01BDHlkX/JxbZi4Lb09AvQ9yIkXq7Cvx0BBjM+6TdbPOkXIBnSHRn+6QQmxtvz8
APhYBW+MVAjVEKPgI8wa/tRIE+0gU3PJBb3/xZoDNSkgu8UeWh80MQW7A6smProW
AhjYB+t50ItJ3QwEE7E9oBGG2H4x9Ks4El23SfKxUdmg13LSd4Due7QqUDTp7l9x
waEYy/qk6ha+9dw0yq0v2mqbZ/77A2A28u9qbHbhvP74GR19UTkJD0kY6uGlnVPq
4wUi8HJnOw4/w0fEkGp4sjaMyGJBU3g/6DsUwqp8ax/4eQv/9UPGSxBNMO5c8oUy
3JBn9k+OUNCa20CTIQxxRykF0SfNxGSZRHsneHSSjiZQt61aDECpAWhDAe7nl90r
Z6W054mlnmGALQqpNfF1yEbh9WlRwlTQGQNbNP7xPpBR+EbJ9isJvtrespDa4lUH
l993F6zuHtB0K6fleU+3xAdp9R6jdAcoV6rABQBRX/yG3+TGjjWys1FTQssZswxi
rx1hyTf9R4ZIR2P/8UJA09tHQRkvN9AehVjZV9XE9nlXBrZxShlJS8MVkJum16os
ECqIFAQOjyGYz4xZii+wHACh3C28sj8yOuQbGGtyNspcS1wtbhqzQOIaUZ5n3Uae
kagXT0l9/dN+vPUNJB6rPkSARYlhYg3hKuuWAQlYrH7j0UrFmHrBwXm7Hm2KTbfD
ayzTr3ClcZa2BMazgTKB8AVZgpKsYYqrLfpwpOGh0o+j7Bo3v4aVOMgi9GE05UmM
mu1rZ/eBHqg5EUgiNmjBefLcmFY5ViySF2WbqjODLWT+Rai+E8JLgCZWlHOiNKD1
tBSI+MuItC0aajH46xGgbsej4H1x8C+CCGAyeujJbUyxn+mqiQv/HvIEzXSqwpte
iHTD2UeNygQesucemsM7I2imaVzNakIhrg2zi2AMmluhSsvJhEsvKjx4KPzXDeBc
L4CBRJ6Tv1QbPgkEodRF7IsILq+qpOupPhqa4nUzUL8x+9d88HVZYZNHxPKim51H
pPUvzV9azpzV1N5ESaWCUSHkGlv4M/+QDsXjEdxYH0W2VLPxNjmIT7LIAMX6j4g3
ylBsPPKMqNhLimkP4yKZPWwWLOiNeaOVah9O/jqcgYTsmvNH33sYtJ8W4Ufuv8Li
H9uX+4uSnC0wpz12TFzJVi4XXpAvqVx/LxWKCjheBpjk5UOuEK4F/wGbQOH0akD+
iUUY/mlxiN8G8IEkT/hYqbhKI6Ag93ynF2LBBQlFGu7f7JWVn/Gl2uzCRKG3EVbS
abs3lnx7pOgxKzl7ISgBtiSn6wEfv/Oz3hGdCvHr+0C95YAXDCQvpkQFB4EeVhXa
tI23tO+DCwpIc7b0tduPkOVozhLVWI2dNq/n8qihFeL+9pa4VvIYpNvXybzVD4j0
c5TKBfVEq4hYdj+3Hw1x30FvtbuOP51hd5Gra2XVGegHlzXEiRdQ1t1j2vpJuBfX
UbL3UCtqOs7xFz3cO8tsNwk6NSDqHOx3XWtUaFrrXtDXsQpISY4IGy2QW3yMtjbg
TrPxIMVicty+g2899AdNovD1EsWIKFyc80SJp94dnYYAkYaOS5H7Y6BOeKY7+JxD
HBvWErMyiJhKFcYu2pFM6pVf+OmbJmqZQuNH0hLal5Isr2n96uVpolyyxW+mOMao
ZdET7IYx9KeU8mZEbxyXMj5soD7TkSdlsF/X6DQ4X1cy6OHw9B/uyE84pULGQEGx
aKdwsyA/fwik8kickoAsFA3E11muE5EenBPk0+LlAKlSByS0/HzPYbv9ulNNK/jj
3Oyx95MrjGvF2mNcxaRZk83fwHo8gX/zW8OlrwWGO32pU1M/kfq936ydrqh7BzF+
y0x2iyOcw6Aak00KjHOJN4FxzbtOdX/qVeN9rLeSM+FVMHu9wBjah8hVD2BNXzXM
/WMh/8AAp4TY8bU4eyaE6/vGbzNyMqt2QEJaP2KZeiPXul9KGh/uB7MwaWxE9Wz3
pzQc3elU3sBGnUpt093owiEQMp5hrtaWxuX2pRnQIeB1wmO5Qvx8k+gSWlByWqvW
l0dL9Pw1qSlR6TUGcgsp5a+WTVuGegzXLPzqYMe1cEjL+a4sPm3lFSZo0boRXq01
j4nwcM9jyfiaxjC4m5/TTO9XAWm33+WvbxYacPA79vdKfcS5xruRFAfULbdS7mlK
tVC0n7ckISLrP4KKQpPp9LaTiGEnP/kx4An9z9agGcPHBoo8MnEvUfs/mHWoG1/B
pR6a3sE25UYdSFy9sH4dr7Ui+va4JiCS9ajkSPxGixDUSllIQAY/QG/3mociZupl
F5g6xfftSIUUKUZY5V1f+LzlrMLZpqFtf6/YQgOFfOq6TjEsCpvQxPekDIsrGQrS
BtEKtzU7Z60WQ3zMH3QZgq42NhNGcxfe1v+r+7HezBos8lPGYdW1MqB5LYS4OatM
cpSzYH3ZkdwFqzH5zUVgXE2dM/yGhTmmGgaYhXeDCVV1FbTLNMMVihJzFof9s5Ta
PRfrYwkriDv6n6+PVi6Q4VqQdXIYxijw2luZo0FBYmVA3C/zVG5Th8FxS3HePICO
q0+TqGNHj3S2uaEpf/ow9aLv+qpVIiGd6cdmWQuwsxBaGEImPkNlqtehSF6S2ZYE
uVUyldhzsIRaefUJ3NOivXHaBUC+8kXPc7P/c7ZDOYI6WjEes7VHhpwTMtt09IXo
Ex1nMsRGaBFHQirarHKJswrg8n+pDa363bo3a5ZQk+4p02eoQOaZXoQ5rTgSirDn
/ZapBe0gKc/MRAJMXl/Rq4wpW+x00DLUfaycBtdED3sG1l2UT+i7ozSDDbrz97K5
XRXJu3scyRpfTLBNyJKniXYKOuYgBf1H0GUyYZCwmUKDnL4Bwfy4uCdnT19KHMg5
oYPm/c2T1OdWF9CHBtF3SkYSY+T53LZDh0gNnclic2+xonPDv3g4lhvzDWlQkIUM
Tl/N/ML1i0gDzzNtHY/hQ973jzaFY8ombUZOJso5xy0tZ0OkkrDmHxZ9ZIxw9uG8
OmHCpNKCBWvSTdhPwhI26DfTvkDmbdJRLpknso3UpteOetk0FicqAQjE5gdyaef4
OG/+QSQlMRL+3EdhZiRw923754XFcYcN5SgIz8XnLfZaf0STBTQ6rcs7u0wp/C9n
TcEJy9F5QHR7XzjCO+yuXOFHuKuhLPqwOKO4bDuoVsl4iO00lfTtcUsf9pskWOfl
Ojw9BUmkVS64k88neUukk9U1q1jH8KR9Mm8Gu+AiDN7QQriUUgZAGnmiBGIvO8cc
8GNrvUAclNLFLKoo4U7MaSgPhtJzM1KzVC/x0uTe/18v0kHkNeLIGUQ9drR4Dpjo
a6rSFGgJMkF00v9zxe9lcw1EJ4NC/91rxSN1+1hMfXNATVaresmEZLWANCmj/GF2
jwl3DtMYDVIoMgMrR1XmRhRTm+luzhlgjxvpDLRMAnwx/YIiJIzYrRenoVo9BKR2
jRaszd4At0fn8KZAfue0wZgBLhxO/AciqxtKnNHiR+HD4Ge0kunYZMd1KTzggMUv
ZiBft4gC5QliYwwQ65bVrypnuuwkJH7h6QkLIxfNsoIjQ51GXuA8+6UasfCDOsNB
Xu+sUduSwQfkTskXNlzfEKrtAqI8zJCs9Xsi+7+oCaqrIixI8Jbm+Sppt3aHRAZ3
U+HknYlSYrLpNgJeMnfP8LthgoPGDdwxpX0pYAno0OZPR0JWplHx8EV1DiANgFNf
tZuBT3l7DDPscLUvjuHDTJpZDABgp8bx8Sof6ZqSUr2T2FdSgwrAHnpWSXbMrONE
iV78JUzs5zlGa2YFjcQPxughADOCOgXXb18O2nMt5+ItfzovrXvRiOBZamYEE+pq
zZNMn1abSVBwpw/75uOk+aJZ5I3s2rs1sGyaIFm1TQul+22CvxmZpFSI3ZJvIXCl
0WrVQcMXZdeYRY7YhRL9fU5X34y299b+gkhR9pKIc9AohCox4G8PNBo1Epv+X1Aa
MUqSxK0L6/kb4OVAPcA7udaTEQuDGqI3BZze7SsN9Jmr20o5UU2YqGqTUgG/pWM6
IeNIU/frKd0j0bazSR2bE9bRCbpNug1hypqsdoPxuu9PYjdSvc6OWxDuMFeu5qNn
ctuMT14wzk4Bw0l6eVhKGSvdjK6tXSc/K2T4qGYDQquqzEmYjW+KtScUTFwhmZ9x
DYdBw4ZNli66DOhToUUPWXpQimSZwWGvZPN2JC1HRJ+oCDZrCV3dDN9w3HMLZX6K
1ltB6fkzZ51PLo3hD5RsiOcSI1SjlYi1ggRhSTQQr49Fosf1LbG85f3cqc46vvXF
8Nrkyl9f0w0bNFaUuneH/097RFzetR8pAomSdrNkU08w9SJTj4UmrvP8Lw5GQapA
plgPIXjpfd78Zq7MNw00HyUjDXYprk0pYVb5NByGgsUdKmyPSjIRBe775GRDlYbs
O038OOwCJJLEkAAEscIEPNdOtEbstFCqw2TUiR43xD0eQeoSTFhe7zUCYilpcvDw
fwPTyCgCiUENLF4Cn1m5o6yuWNM+128UVK26fOr55URz7nr80ceq5Wy21yi8QEdc
fz3mulWfap3i5xW1zoCZCK/lB8CIvrm55XDtaGevOyHJiiKtS7idgkVyhatra2uz
QkFD5/2xDm3KapNJXUOo0Hr80ca53Rb+8KLeHvcEx/Rhr3YComh7qYSdivYSeTry
5+wG8l1CsVZmCg4JWepDOsc05DL/P7y/S2BAyzbkYIRgbjyK1mjlpaXpDwqyjtrk
XRqu1NtR53BAIJ/zNWpDBrWf55r4rpYVaB+PAPB5LG1cLxItwQ02/EnVzK4tii2L
rsOfAPH/TXi8S61I6J34HToykI3BTtfHR1ZPl1nTnPFhrj3OzZvc+XZnOCeIwkB3
GqCxYQnIyNYC5W9CtemZZ6I5WPBAJujXaVCN/0mpZWn1eoI+RzH2gboIl2d3RpWe

`pragma protect end_protected
