��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�:����R����	���^|o���6�C�_@�<��v�H���g��7�,����Fp��p���@�럀}m��X`i9�[������ ����:a���7���\�g�����q	0�,��ߺ���5��+	�K� ���W�te'�V-������O�lrHJA�#�Ay��[� � ���Ђ+��<Q�D�����N��{ ���q'�JBP��,<4��H3��pϐ���`��-�SAO@�<��:�fѲ��o
����-!^��+��4�!��B�i���r�6�lͿ��	u��홓^^_��[�(�G���S��OW��x�)��=.yf2b`7FZ9�y�� ��T{ev'y��"% 3|L$���Z:9*A�\���\@��Zv?�����I���hRą�I�	m{q�[����~ M4K���KN����0��������I�广G	�*���A��a?v�ȒV������/sُ�j���&sm�&u6��Yk��������g�ّɴ��Z����n��Ǌ��NgҎ�Bӵ�<2�W��Т��M��̣3�s�m���>�ldv(�O�9�Y���I��y}� ��|�T�N9��	�Ko什���g�l�9����V�cܩb���h�\�����%F��S�����$�
��'��g$����&ꎡ�7)�Φ.��Smn�e	�:����+�8�l����yXu#}�|g!Լ,�|�j�*zG�0\�2���HMM/�	��b�6�A��X����7:���R�!$��׼:���$�W�}�1�M�%9_p6����J	ZU�[8n�`�0<:T�k{���<rRڰ�a�Z�B�[�.���<	ͮ�Pε������UQxH������σf�<���+tN!��|�VJ,�:mn���E܆oJB�>P������c�?�9���1�nԕӉ����e<0��A����e�9��i���O��1o�HD�=Y~>����+�$B�*dt�⦭!q{�v�㛽
J��c�a��uQ�ds�yC��)vZ�0�3���6��;�F����5�����9�+�X�X��|^���¥��+*#����	c��$�94Ǎk�|O���I��9i�A��͈(������F�¼>w�����>�|y ޝ��uKy��E�iAYSƴ��#�FD�_��I�yG�MT�,���:ܐ���#����ݞz3,�'���p��)uS8�=�/G��AO�f���nBd\N����g�B.^�c�O:�������
W�SF��AT��E(�`E�٪w4����pf�7�Uc)li2T�3?Q��ܥOW��8�5�C�d[���`�c�O���X�A_j��`� _\��O@���>��%e(f��d+��X%��%R�j[���y�~�$��x�T�v]�9]5-�?�o�>�G��L�۔� Mn(������z����A+%�{��r����+��y���?���3�XT+Z쐋?K6���?�3#���U�ڂ^�}�l����[P��1�
�4�
�)H�!s^��:�2�u"?(�r��΃��u��V=��	M�ۡ�J�2�>�8� �GbBR����
�Sc�(r����� r=CY�u%� ������u���m��T�+>˖z�Ծ.5���}���Z�ZI'��� ���f�5�=s?�ș�[�:�Y�5��E�mr�+e>��	��c�:�y�h����2##�M��YUaxต>O�����x=��ɸ�*�: [ˋ�n:3�W>b�����P"a���u�'ED�>���(J�q��r�P�A�d�;JN4�}d�PV:W�1�D�Ȍ�����mѺrh:��&�t$ v�Q��{������XH� J���?{$N&iE�.Ig�w�2/J/m��X���sM���jk�Z<�鳯Ta�AAb_q6�M�}���� �	e���,4ץ"8?�3r��Y�vLo�7�{����)sV-}r]6�"����]A��:;��'��רgB�0����uxG�{��-]���F,67Qup4J�%���@$�U����f Ò���3��8����k�! {� U>�攼&�lm�D~��6c؃S�'��r�,*\@;�F6�Zf�܆��S��A��%oI�t��0c��jg"#j�Mh�Bf;�&����'��+�ʵn���˳u3������'�A�>yk�K<x�{�����Ѻ:X&��	hq����-�1�!5��)o��K���i�/d��?]�; �L����,w���`?��UԨ�"�%S��aJ������!�j�'I�u=pV�5�����7Ԃ��:��ȴ�|ؽ�˧LM�i��gJ�6;��\���2�(ĵ8��F��ۢ]�����igl<_T�RB���.�3�q����Y\�[G�����94C�k�T�����?�nA`�v���X�|����D���^	���_ ��݈�� ���=���Q��6{��;�(%��OE�Qێ��'?�?��{�ZM�$;�����K9�\e��h
ϣ���P#������q>�ԕ�h����*����jq����N�D�v�&��;n�ƟoԢ]�A�<'+�̉�P����x�p�� �++���XQ�RI��8wbfs�fz����[����\A��>�{o��ں�S�,s����B2C������Ec4K:��⁈�W�.#�V׋�e�:�00�B`���
r8s�)��$Hi���S�U��E~Dt�f^d�!�i��v�'z-�YN4~��蒝��ְ:����[<�˳a�>���h,��OU^8�z���BV��}�&Lx�.2E)pǌy��f�qBfB�ԧa�B.rYvߑ�/1)9"�@Ʃ��:7�Cz8��D{��b�{��U�Jp:�m��7`ub�6#!��3^1	�I�	-D��;X�M/O��Kz�ם�n�0����x�e�	��v��w����͓p
����a��K�~�i�8��{��д񉯋؝��~{�b�d��6A�g-p��#���l�)��:kl��OU՝��<��Q��;���ޤ�O���z�����B�1��Y������u�{w��� C잛���K����>y�{UTe2�	�̘���0w1�8��y��v-2��6S�a�G�^'���Y�|~��B�s*dR<8rEK�7��k���f����c�2���ҷ}����ͮt\���н����������eӏ��z�r6{��SUC�K����1aW=^(�d�o�YU��u�"�]p!�FlT)}N
=��*(��R��	į]$쐑����ZeZM0_@GH&�T�lE,�"&�r�e4I�F�>�p���bN#��"�����<�+Mɜm3-��h_@1xk�\q()���~X$�ّ8���At�	���߫�]LP� 
{����Vwde�_m��6RnU�5�qF��<�e�X�@�1��oKg��0E�� ����.�CsXY������}	2߽4 "���-�0)��% ��>HB�+n|򌸣'wDI��4�2�Fmޢ��캕�Q�W�V���CM:p�}���}7#��^���`y]`�$'%���Foq��ޚ����}�K�m�w��C���Oj���ܶ0��B.rP�� n��?��T��}��_.9��Ul�e~��0ڢ�譧�:(�����uۺ�z���ED��^������5���nPSV+Yɪ�2k0ů�#W�;�h��j�2���*o"w���$�f���b��ؔ���W� �=��$��>9�ۮ�sĩ��m{�����):���U`��.�������2��Q���7�P�Þ���{W"���}�=I��ž�@[`v�/<���UcS�V��(�Ow�<$��(GI/��Tw���fp]Z�t)�;�V!\����ض���{�/G�B�/�����::��uq!m�&y��JI{,�Ĵd�-���f����ݷ!r��[����ǁ�,{Z��������b��~'�!�+���̌.%�m�&��ۜf�ԇ�#�^4жWV�*�!z���4pZ�@3VIaD��A���7M �M�����Ó���T6�7D��vN��lY���Gݠ�ńq��QN�ťd�5l�xr�G�0�DT>1v�������t�P!\� ���0����ج�3K'��9պ�ėܰ�6W���F��Y,�%���_e:h��i�J���̸���Q��c k�W6jK�V��ώ��t`���u;��v�\� S�n�.f�� �_�F�3�Ѫ��H���C�O[���%G����G�J�_/g�#�G&-h��a㖭��N��b��R�S����"T�;�qs;*��
q	=�G+K������
�uϨ��5��,�*��e�3�~'G��)��;Zu�gJ/a�
!}�,���ɋE� 7,)���S� N�C�/�?FC�Y�eռ��k!��,��}�e�vy�yEP+{���ec��>�z=��2�];��]ڎ�n��XTh�%�E`T�X>�<�(*�}q�ڵq_i�sߴƈ�j� �؉>enx��3��K�h?��B�F����}��0Q/Rܔ���;�<��/}�`�j�k����s
��^����CW������A]�C!;�́��n3��E�^ة2�c��~+��29���r�.j��m��Gߧ�e�٬�}p�o�:=�9�̘�_�����p�z9�д^��U?<�w>�]�)���(���3=Ջ�t��i� 5-]�06ÖH,� D]2|9boLi���x����i�'�V0>Ր;a�vs�[l^����v{ƺk�:������6����7J���ǉ3{9�_��d�<B$NJƞBI7��=����k!3�
p`IL%���g��/B�G)c��1�ң$�=��Xv��:�/Y�l���=
Z���捛\��=�B���7O�+1P#�դ1�9E@)a��I���8N�ɢ|�m��N��8��8�ƍY���ƽn�X��񬁍p�oJP z�\�1��������"�Е��FeN�8:����fsW��L�O�|bzZ�s��2��~O`��s����/����(Z4���vϺ��K�ШT�x@G�{���N�F�5�Az,�:iI������h�l/�m�@�2��}��7�5L$y���z��/8�#��B�v2��ڷy	I��U�it����kq䍔	q�'g��|�Su5���5r)Pj� <�ʢ������s��K�<b�ň�q��o~�*,�Z��V�!�W�*Pc�����#x'
f�Q���6�qT����R?� U��T-����;K���2���u��壳��٣�T��O�tP��H����͓�4j�2�Yi7Yl
ba9��K4	��&x]Դ��	�L�m��um���[�?f��d�n/->S���Z�*���"ao�0Tp����5y�LX��_�;(e;d4�W�5WA8��J6��LضP��b\�|�4kM���)��d͉#�V��cy�V��΂�
>��p���"�s�q��f5�ܭ-G&��z�ĝ�����p�$�l�`o�a�Č�0�;g��r�7�S����%2L��+�K��^x伴P�b���c���P�}�X-A0g�Of�/����u�����Q���<�W���d�)�����yY��c��� ����F�A��F�X8�w��m)��/i�eӑn� �kz*����{�%/�+WFHZPV�ױ�IBUN�C�.n���L70E�$D--���m�4�HC;��ڋ v/�9E�\=Bw-������E�����)~A]=�Ҏ�t$����̅XFY�$����L�%�P�_��bI����n�s"%��<��<a�6���%
q>5���	�9 C�V`'��=�&9��ě�381�euRf�WS����L`v?`�s��O;&�q�9q�f��!���ao!%�TW<�j�؂K2p�B]g4�%=��,2M��^bG����^fF����X��:�x����3�x�m �;�x"���M��e�<_9Z��j{/$h���@�4�7�l��vNp1�-���%�a�DzT���ݠ��ڋ�˳�t�j墖j�SO�zeG��4�]�%R�L	?� a}�c��@�Gr�ԣ&����k�ڠ	�I�������9�����6bf�oT_���jT���j��~�	�E��Y*�����@��e����Y�ku\}���=)�@��,��R�#n(�zJ�~ǥ���!j>z*��\$��	D�H��x��k���X-D�A<������ҵt^#e���99'�hW�h�-�{/��Q1=����\���&� Ƿ:��ȉ<eˠqE����=��r����H|n�&s��V��՝�X93��)Ey?'Z1�ʃ�%�^[�����8��}Rߔ�yf���l�ڲ{1Yg����'���J
D�w�KZM�+6�_C ��_�xw�oߞ~M�G��޵���BX��PD�|�h}��_5d�A�<����Pe�4b���g��Q�`�`����j;X���(��Q U�����Ɲ#�g���ae�Se��(UA}��ӗ��fJ?-^DE�;���Ț�ҫ�'���rl,��VE�e��ȿ-�Rjc�ȡ�:l��>�F�4���.M��pmJ�������v)��c��
#��� �Yz�{3���Zml��,�R��MX�`j��	,���:��6�~�0e~���	��h��-���3=��T"����|�z������	�]����孌��C�������99����T�xC�'��Z�\�ޚXN����|D�D��	�ܨ��ȮB7ql�Y~�m��@2oλ1W�5�&j؇��t�!B�D�Oړ�j�5�H��d���Xnc��8�oo��M��Ԡ�E���/~_��TJ魳8���Y�m�ofѫgn:G�}v�
�dMD=�6fy�3������;)�6�I�3�ӯ;KѬX�9f�f�T ���|�6韟$�����r:`⶧T����XI�_1���6�1�~�x�.Ab7�u]GtD+�~���w�2EEJH�W3�co��>A��qs�W��7!<tO�Jwb�87�8*Ã�e|�ې�$�#�5�J��׿HB���-��[�ဆ0��"9�^�����\J���춃���&�ų�#$�$3Ϙ>-�ԥ8͆�;�Sv��R�c�Qj]굆�7�" 4�F&�W��p������8ڞ�E��R%�C�6�{��4 erx;Y�jps��L���}D(gK=�9�eI�w�6 ���}/�N_�|d��.�U��(��~5՟`UeX.� '�����`ጀT���mѿ.�*<;�H��+�$�(>0R"}\�%Z��h_<8��+�^���.L���M;���P��.R9�H����ǵw��Iw��Y&����zei}م=��5p�M�bޅ���t%)n��}�PA�Ԭ�U���ʎ��-/��X=��گNR?��#�������t+����e[E��@��� �g�LA���K�t�C����(�E��,$.��z�p{�g2ϲ	c��;��,>a��:k�PF���r�-��K��,E츑o��g�(P�`�:!��x.: `���:[����\�F;�H�8��Km����}qp``J��o����P��^����G����8��*�Ic��[6"����=���C�8�_�|��9��u=4s�m[���ϫR:�@[��P����v9���5�W�f�����ouk*R!����t�� �����#*�E9W�űe��f�a)	#��\V�!)��y�A�T�t9!V��yZE �k���l��U
�c��ʞg���fΕ��F�9�4�=x�BgI+�`�ˇ]��ܰQ��L�����if+&ϳ�p;����0�*��l[`��o����a�OƼ��4�����c{�@W#W��0�v�z3�����y���'$��G��4ƕ�݈	4���!YF��K��c� gU��z`�]��ϓIՔnj�.�g���xem�V.!N$�}Om������`��j���q��Ay��R�MP��/�ϯ�R��e��HB���eD
�哰��Y��Pn%�EWT�,���cy�H����1��^���Y�f�.݁� �
�R ��&ްQ)��m0-�aib�gR��Z ��a}_�{��L\%�,B������v���bT�Wd����h(YZ5�˔b�)�q 8LH%�"�4�VL)���m��lPQ:��XA��;k�
��tB~�f�m����c�8a��ҥ0Q�K�_�er]SK���J�l���"��9�}g�=��Ӯ+
���2Χ�����RW\�FW���t��{a�2�M�m�"J���(d+b�G0Hȕ �g�ojʣ�=�rʇ�0\X_,�5K�K#�f�9�������V����BNE�ޏ?m4r�ͱ6b[�8^m8�	���>��M(N��%k��	$ 嬿G��G�K�BD�6z��S��:�����G!��&{Ձt���*g��y�H���ieǜ��A�g�F��\��ks����G*�����
C�XI��\���@^�=�q�AE���� �j���]�6\�8�ƒ|Z~��ެXܧ^Y����!�����V���c=)�`��ag�*�tFU�):Or��W���v-�X�r	1�Em"Aܠ <��N��������x�6�����;.Xp|��-���؊L�@Xϲ�X�� ٕ�B����i�UK��m�r�\�Mj��S�by>��|7�*D�ջܕsD.k�2��꟦��^'���K��-��9��	f��人������#�?3x��x��3-�\��=v����	y����_���ڙĭ<�����H�()�.K�k.Z��d0yA��,졝}l�jG��6l�&G�ڵ��l9D��BUn��<��`�)�s�ת�[4����wj�i�Fg�op`iĀ�*6 k��$|��^Li���s�:ɻ�R>���U?�>��p�$@q�b�}�0e�3�=|��b�. }�=Px龐�r���G����c�n�<;Pu�tކ-�[8�sh#�)q��I�+���O"
�JJ��-'MJj�5�rBA�g����h�7�A�?����vFR����G�
Y\���C��J&��3�4׊����ʕ����4�;~;2`�(j��(g��/�)����F�Ճ�3G���JK,�8z�6ׇ�n�c�R��_���u��y����f��O��������VQ����Tj��2;�l"
u������]�
0Y��@W%���՘�9̭,E�( �a	��1 ���1>�A��:�R����i����e蒆� �����\i��������j�%n̍���_5�y�}o�n
D��65��u�����b�hz(�!i�X�v�Z�5��-��bGs���	XJG�ށՂ�<(��#��2�L���J�5h����f5�N�-��^��\҈�n�����B���^��$m}�rzXx��Q�%
e4�(Q�b��(��#�P�ۄz��̂"����al�Hک �:��ۨk�35���/+�S�q{/�X)K��l9�Z��c�JSIYP�oE�Kv�F���~Ff.a�t/��QL�q�Sq��kމoë$�h5����$�2�&��7MR�O>U+��g����`��V }�咟-���0��X4+(Se��6_��&9�i�D��rQ���Г�;�=��6E���u#\@�>�Y$ߎז)�0@�uг�f���v��u�ӟ�Vt�K_���9�Oe�����wm>��wV�j���t0df5�.�ty�2��{�=�����>;��V�T���k��<�[�Y��MĻ���A�x��2�7��J�o���,<i�ڙ!2��ɲh4diе!�A��s�N�����]�\Lz՟9�aP�G�0��h��m݅aT�/+1G�ܤʬHMi�uV���o|ܩ+]+�5Rp*�'�g����@c^��$�Tc4����r[���D�uS:I0�#�#2�=�O\��C��HO�2�1~^�����cgw�m��̮ �p�;��f�xq�9-������u�;0����s�n�#��D��;%t��t�~��RZ����ރ�7x���2QO�|��a4��uR��f�,T^݊C�s�x�39�i��H}��h���wO}��g�7�;\�]J-�V�}��C�<��Zj���V�[�?gw��^řC���ؙif˔�F�u���P�hM_�(��+�݈X�g��	�<1n�
� �3�
��&܉HѪ
��XT[$�G�-vz�L��v9�,��WX0��y��b��K���q�"���:�Y1����!���qe�y�29;���M�=�Ճ�r	
��G w��P\Y:,�(V�h0<��l}g�s}�Z��E��z���MI|c({��|3��!k?<����ⳋ���6�!p|t��(|�}��� څ��`��r��Ժr���\��z��4<%�Z'�@[��9ݐ��%�\9
��/t[wf�$)��*�L�G4t��j=� ��f�ɗ�)��:K�U{ ���(V�B���zs�h�fƏ�Y������ W��ʮ!�g��K�@�4/�U��}�L�]S+��%z�v�����(Egj���ͼ�ճ0�Y`���ˈC��f�0:$ܲ��?�_ј~�֡PAG������d����D�b�K��(�Jws<g���E����c׉:�ჲ1��/��� 7��^���0�!�\wG�I0X��2GXE2��tY����.�B-#�5 ��OE6�B����Y�z��3�`Y�zU�^H�� �؏��t�MJ�l~A=�o��"ᰍ)*�0��}o����z=B4~��]'r��<��w�*��	D�%d.+��ݯ����(�2��g$�h7,@7���-�5��{�c�� �4)���g��&��2~c�4c��d�9n�չl@�T���3���~ӠM�N�+���!h��2���9�/�SFu�s9x
w�u,.��Vo��H�w���P+T,�}u��qiZ��q�O=�N�y~vڞ�dw�g1��9ؘ%�Y�&�T��*�q�^{r6M-Cu�?�S�a�c��7;��!��w2��~�!���&#�,M1���C]�ZD7�g��P�;�n-[�#�]6�?<��dƫv�a�`��8|��mۭ]�d� ^�Acj7��{q2��ڑz=�Ir�z�^��k�1���=~b��0��1'i:���F[xd����]?�ö��?]���3��٠ޭ��ߴ�r� 5p�E_F���\�[D��A�H���+�3��, ɱ�RrϞX�D�MG����� ͎��i�#�sS..�QGeS�V��̺!��%.`�O�Q�#���f��[���i�MR���*�L˹��E\NG<���tl�UI>Ѳ�T��8j)F,���\}�����p	8C��?���>NFo��}s>J���\�d>@�(�U�]�H�n�����	W7�f%��; ���MA�7m����2ҙ�Q{��iӈ�m�+�ʪ����&�Y&X�.�Y�2j�͝�8��c�B��YD�Q�ۥM�pu��6�����RR=j��;h��P��$�lq���a�Cr�;c����2�*�]Z.k,�����ھ�W�A�Z��������k���n>ƊP�����;6P���6u���Kz�β�^$˄�Я׌�j)��I�5�{I���8�1=����d�wh�o�O�9��4����!N7�������=R,v�tM�B��Ǫ`FYGvu`�b_d�e�w/��&��7P����1�������.i� �λ�����)�.��J����r�%�oK�!⯙mh��K ���;�����L�bU!�R�$a����g�Z�ɞ7{�}�L#��Q� O�s*���,D�(�e��\S1�u�(<��ONs��!�J��L�{E�4I���CD�o��ZfNtrɑ���7������'2C�����=F��&���z>��@,��N.�
�D�����Le�!�t�ۋo��a�����I��8�͡ĉ����9S��؍mA��J׳(�5����MMG/q84��)=�]�X{�
����&
:�����t�ͥ�v%�{^6vbI�̋GTܨ�&�&�޻��G)r�јZl�C�2S��"(���R��V�XY j�Rъ��=�J�y,`.��n-M�j@Ȼ��*�		dfԮ�'Ρ��ƾy��\�5e~���9�#a�x���!�*�D�|���΍_�\8��9�bX	�q��PaK�r�,���2u��ݯuY�>9�k#�$�nӚ����z�e�PL�_��~׽�O�*����#�(���5:�:?��o�����N�C����MC�"?�_������҅��V�|\z�<���&��B�ܲ͟e��-�&�옮��u�ڪ9�(|+e.��+�D�AW���v�/'.�����֪��?����R8�[!k>[c���.9zy��@�4���g8pr� "�1#�ǘ١ҏ�KWL�@���$��;\�U>�
de�V�d"���v��#�#f�'�`L��2rK/�����Wn<I������$����渲_^�^y��v�Zrf''��+3Ycqy�����Ѧ��VS�s5r��3&����$U1�V2Zn�!��2�o�*��0���W���K���� ��l��g e� ��p[��a�q���4��p�1?�GTb�7ּᰙV��N�@�i�-��/���������Gw{�9�͕��LhEymx7"����?�7�@eT��K)�gC�ٗ��<�T�"
��b;cT�c��lʈ-�Z=������9�$gG����A�3e�ю	���c�d�|xt�?�eK�^��������h}�F�	�2�� o8R3u�d���{���K�r�E���XD�X��-��щ�rH�`�X�. g����a,� 4Ι"Ĳ۠����3Py:�e8k+q�D-x��b�f��lw�g��掿� �(��a����퐴-��fJ���u�7�����K)�녭i֍�2a*p�����i8j=��o@ҩ��F�r��u�3R��C`����i�
*ڼ(Ra&��+� �Iu���D$��J�b�t�M`��|�D�
G��u�P��w�L1�0Աe���=_K�f�O�<�G��!��R }��m}���t�D�M�cv�ɇZ����:��JpY�Ae���e�4���ٔJf�Q(��A�#��~����ݝĴ�K�� Ce��kYD�ߋ�?G�����_3�u�?�}t	���jJl;ƛ2�=��H�k�p�O�a"��e8�7�9�%�|� �q��f���� ̶��}� e�x��_�&�V�r$����{2��T.�Z6Ɉ�3�X���La*be��ҩ-�JӟIr�ַ��y6�}_>�{~�T��<����#p:Qѿ���2�.�hqa�֥/�Z�@@*G7l�"� �ҩP�����f��5ӪRߋg�iӴ��g�Q�A��*�/�'sƠ�O G9��xڰ�\�y�{���w��F����?���]�����nK?s��U�h���Yy	�V╙��O����6!x���4L�F�i~ֈ[_ $��s �vݲ���� 26Y^��E�*�_uߘA��F��v��I�y�;e�f���i�VR�x�R'�ϥ�tY<���n�>-�1mY��8�dw���~�S��s���S��^ݖ`^�<>}���t��P�!5_@�p��0��9��_e���QW����������/�=�a����3/|g`�c���������/Tp�L�)�@�Yv��7ȧ��1��w@�2#����b%�L��8�kΰ�[����_~T��~N+ͻ��(�5?������A$��)T��+�dS�]�y�F����;�
�A4�s�[��f�5 �'�u	��Ï1M��<�dxٟ��mK�'+6��W�ٶK<���f����$�#<.~)��p��f��X� ���`H��݂�Q���I����V��a@�_a�gI���aj��c�%�O�\<��Y��(f�аqR@�]��-�R��>�T����,���:�N���|L+����-�kI�ON,^� �Z5��
��#��/�%\F�(�k׼�)��R_q<�j�����^)<��G.�dq%s��G�򞖅J�О6da��2\�|�e���)��ߪ��=oF����Q�V ��vWu:�o�!����Wī�K4�A���"�U:PB˻(���2���.�B�i^]B�$!��2\�u�8o7�5���?����昶Y�ûRBg�>T�����X�+7�	�[��Ij��#"Dt��Y���eU���V���	�g竦�.dt�
�J
"´S-OWQ�M�)hс`v��\�Π�:�r���,��?kJDo�mQ$V(��I�[P��ȝf�v�-���ٳ��-iy��0�c��G�ǜ�vH��TxI���#��8�CҐ��S�o��ealo8>B@���iE�S|)au����`?��i+&�1#�ΓK7�aq����3!m��\a+�˸2A�\��nW(�������©	V�Ǜ�z��l��/8�� ��aɒ��*46��s{VÁN�M�#	�x��s �_��6c��Fc��/�[#�=�ѕ�ϔTU��Cmc�J��I�n�;�b��-�b!z\�i�(a��ts�
��^�k��`�7b�7h��G�u*�C�sG;��ˬj��S1F�G+$U���=�'�Ё����_ƾ�Vߘ�F����ܮ�Vi�f�"�z��ɖ.Dx��!��ݳ��>��E�z-U)#����K-E����Oç��og�1�<���~�'$?��j��zg_"��q����g�\�}GT�d`�:<�;qĉ�R����#�x��I�큸 �e$���W|��Y.�Z&r"/���=	�����o��u
.
eIdĳPЧ�MS
t��R���xIZg<N�Ԩ��I�_Zaw��xݶsQ
~2�0���]r"�L��mp��1[��F��
ȼT��۴�����t�P���D�af��o�>V�"+����؞L&O�o��Җ� #�:ǖ���-w m';�t�(ӊ$��Y~i��SgI�"X�p���|L�__{���F1h
�;�(�sB~��g�)]��s���q8G�0Vd9X$-	�CP���K�|6��<���B�>��������g��~}��Y[�C*��_S���PR���0�QZd#��:zȮ]Gj���I�m������l/f��و�&ͪ�M}�BÎĭ .Y�-彜i����L7q� ������ЧW(w8-��ͮ�π!ng�'���1ڰ	�y�!�rHp���o�C�&^ J��삦��H4G�"�����hq�.ܱ�o�0;d
ʁ�Au�>Z�ڲiH��8:����o�l�M����s��=�uм�r��ud�=S�Fp�)x�PXjQ3T�����Ui�F^.����-'��!i�򢢞c2���U�z1|����|����jV������W�X�)3x�k�j�D5�e����&�)�f��ј��:��Zd�~��Z/��f��(�'S}d`LloE��gS�?�C�
:�4+;�a�]Ytd�8�7,�<2.���|�GR [7`ےN��M��&i9��M?�9W�9fF
�c�=B�d\x��i�~!�ɴY��~Կ��hrf���+�뀚,�,��%yȗUL-b��0��#��#�u�k��2<{�1*�Td>C��#D\oB������� ���tv �ў��R@�2�F�]�Zg�:רY��\= �ګ~Q|�����\�YeI�����Z "ǲ*2�#��L��TnF_�O)���L�3ڋ��h�����M�227���Sf�
6N o��v�=v�����0����aw��6 ���6�Z�Eĩ�O�N�@H~�w�	y�:T�&�������A�[����3&��@�b��
ҝ�\�������p�#;;�:�Qn*ڦ���|ϰ$Q7��8w��j
�H涨L�>(��,|q1�!�����j�DQ���r1dDtMY}F�.��� &��_���&�����H�[����-��=�8��G��T'h�lb��p_�W�WH.���W���؞�zY����>�K]<j��7�PD}r�i� .��b/X��!9�fl�����S����ՠ�[�ICU�Q���G��e�Y������X�\��!�
�� V��޴f:ַ��|�6sru�~��gM���/�e��^ĺm>w����7���BYN�a3�L��)���~=vݿg$9裼cNvj#	���/�$`�¶v\�'��� �aP��G7��nd� ����t��
��?J0͵��N���Y} ?c�O� Oˬ���{��~e�hA"Q�K���s�"��7Y�Y�3�;?�
)��>�^��oU�i��,�C��
6��J��Ź�	��N��+��:/�Z��Z��@�V�׌Mn�P��![@�9�;����wq�̻F	z��hI�X>����`n�ƃ��K�I+eE�]e� ~��ix��NWI��Ŝ��'�ߛ���g��)�Dfϝ�V��c\� նl5���cc��;�ɴ8j�QſPp����!�K%�%/H���\R���p��+'>ܒI� �pe6�0w�۱��+ǹ��:��u#,�� ��(�VM 3Ys�� �2��n�#�Go���Y(��Ox!Vj�f��E��ڕ���jW��i���e�BG�b��IC�	^	�}P�gN�K���!�)w崸z��Ć�gx*ꌾ� ҳ�'M����n��g���?����X�Lo-LI �ß�zicG�Գ[��5���/��EQn_�Y��|d$E�]�^�M���d�Z8��YTR�?��ܦ�]�{��^'a�=ȱAJ֭��!�B?�fv���c_�l�T�3��>oUgLJ��ji.weh��M��]�钥s\g�p��,s�|��-����.�n�Y8a�`�.���|1Ƚ��B+v�P�X�Q-O�_��j{N������h>a�I#L���alL��.&d��ۓ��o�\�sO\�Vi~v�n�O�)�D�G��5�=�r����!�fD���2�8�o�� ��e���cr�)_%�G'ȏ����������`��S,�jLb��e��"^J*�/Y��Ff���x1����"�ふ	�ݪɮ�.�t풪���?�3N�Q�H�[�Mݨ��*�C#^,f�q�I[bk lv�Ԫ�J�&����4�t��,��%ȴM�%f�ʳ�M�(��;�I?P�ȡ���>e�l�!SG��P����So,_*��o�%l�N�Z�o�����JZӪ{�� �\,�/ի4��AE��p��_����_����ڲ͋���y~;+|H*��~j��z�rbyL~\(�n�fk_����^Ʃ�*ix���@������H����L ��n����e���i���Z��T����j�������^�������>ڼ���J�d��kE� ��X#;7V�m���F���	�s�^�
S�;S���9�̻%Pk�y����d^t���cM4�[�҆�5��,J��Kʂ�z���:�J��0Yr�Z@Q5���7ߢ�-�-^��@�{hQ�������l�H��x�V�-����<�y�����+����ClQ(���yPH�z!�CH���Z�C^��1.X���=�
'|P��r�=��u��2��q�Dޓ����d<��0�-���0de�&��5t�C��C!� T�q�4D�7*<�R�������UYh%����ah�FV�*�����Aw
���0���{C\���)fO�j�����%Ԍ��_�J�}
|��H8ꯜ�����+c�?dOnú���
N�b6e��k�s���/��Z����L��Ԅ�,�r"������	������}���k����Ai�C�Z����p�oO.��y�K�C�h!��4xYO�T|`��P&'fիw��+=�a��JDH&;�\����;4ōj4�Z���PAl��q�{���=^3�5z�pڅ���e���˖���a�|�f��o�i��a1+���P���S�n�<�:%q�f�˨���M����|�LV��� ���eCp����Z�t�������>HY�X����h�#R�;e�o0�1�,}xl?����(�Q}���*<UCϫ��2O���"�ee]!���PF1a�<�@A�ޟ/���2�����]�k+	B��zHE)�7ʒ �E<�1F��1���y�1�^�1|��X�*0�[t`_2�ʌzJh^u澠�$�q�,�������zR��10�h�v%���#�.�$����J!��ϼeٺ(������U���"#�E$i��DJi�s�y�"�c�<.Sl�����m��f	|��B��]�|w��,��x�p^T��bb�p����\W#V<��d �k�Λ�΁��#�&&�T?��:�����п����#�d���ܴ̾i����^�-0�h�� �TZ50w��O���Wm�((f�U9%�o�t�.c��-=�����\�d�e������ǣHc�["�<�&���bV<�KNR�wT[��eu�
�7SO��z��H�&�g��bO�
)F�p�t^�E:LQɝ|f;�>��/^�7���9^
H�9���T���x`��1c�p�aB�V���agT�.'���5Ф�rW��u�h�b�����G��߹c�=�Ż�5�9f'��!V�U�}�/����I9�%t1�SB�4�'�Y:`e
ۈ��x��	Z?T-���(�&�0�#����)���z�C��Y���~�O6�k�2���MQ���Բy�����Ө���Dp��b�����@�������E��{vcg�$��)=?��� @��	uk�&�w�W����>�c���4� ��n��\�y��'˽�g��=��8��5,���JP��<u�4���YOt�n�^�Jey��0+q�zn���֓T��ucL%qQ�a��V0�7��� �l�h%�c R���C�X�E�ࠬ�,�I�)~40�UC��3R��� =�����������+���zن"=!��Z�o�`�Ң WI&�<�fڃ)]�����<�c���$�������P8P�j��e*�BR��k��Y�'��;ޮɼ"����)���φ�Ý������oy�����m�#�K�Y���r��j�sT"����9/�
Z:"C��7-ϕ%-׮����)��#k��2=���3�7*�,�K*���n�b����=�^�l48���ڕ�R���4�Oդ�#����z9�t2HB����9tX݄C[���ǹ"t��w�<N�}ۓ�6�	j�mG���L�.ǳ_�)4Xܝ�����K�s��$�O��i]���ƖN��xY�^r��U8�7{%��}pe6=���|�"p:,�dj�=нÇ�4)�\� �eqF�+�;iҚ��N�Sl�[r�4`�{�(�^m�����Gb�J��v^d�K!�yY�+0��q1���m����Y���d�Z�p����m��\5B[;B�O���g��<Kb�{T_Y���ݗt�! +�%�=�]�fHkw/>��tP�@�z=2�u���ȩ0�=/	�8��KZ7�!SG��|]Em�!��k��Hm�v"I����s*��X#���]e����V�~��R�D��F7κ5�M7����v�XmK6�MJ������0*�����HA�Ђ�Rs��fh���.9� 'z6�7���l��M��.��#����۠�k6���)��<�lZ5k�#h��n�'���ښ�Cǫh�Q/%#��&���e�}MxY#��2r2���@�� Wjw}}n
z��X�-qvk�<�.��B�gF��ڽ*�B�ԩM�(�O�H�>F4��h:�����yA#f�>'`bk� 
<%Q�$��k�H�;�g{�U(Wm��%�"�C�Ӹr̵����̰r�X�?e������n>.'��c|x����@�� *&v����?�L�(D��e�@�ۜ��H-���XT]��5�"��d�o{F<cþ����,<���H�t�t02���Vo�/b����F��qE�v��v~2��d�,X��<��߾�[v4!b�/ �ޝ�f�#)gލ�%g!��s7~ryL�(���J(���t�Ҧf��T*�(���� �U}�fd���*("�7�Y��,U�n�W�d���:��P���֜��3#
�	�>��$AFDf��>,�<uZ���H���~{�����^%���2��	[h�j�ӃL�Ό:�.��g3Iف�ܑX�RJ�����h��[b����Q��0Ё���/�B���}aL6����r_5�D�-�o]ǳ�/��d�)ġ�X�\O��}����")�{`)_u ��S,���;��Tۂ���z�	�t�X�'�8�l3�e��ST��ٝG�/���a���NDķ�qk"��7S�/��M�b�)��pH�Pg��`,��UF'w���v�~���#�yo�ĸr�A#m��xOt'����,�
�ݎ�o qš������&�����W�{$Q0l׬ ��љmelў	8%����_KPF�t)8�,䇀}�+��� $�N�z�K8�E��@�-�����i|R�������K� V�i�B8bM\	>l�_�t8�X7W�K�gh��W��r���J<��5iZ#L��56j�O�\����;�v��U�^,�2(e�,�&7�n����}�͞Y9Ne�6Uc��d�)D\*����d(i���2+P�S����9���[���^Vh7�x�W3�,7U-�~!Zi�bi�c�.��/]�,���4���mI���'�����9���@9�U����W����i머ѪO:�v�y�\1J�����Ih#���~���yw�����"�����}���47;2eZ�,O��Aeg�J�0%��l�nޔ����'&s�?brI�c9�
s���� ��4(H�a�SG���#�:	̅"�J\�{F��յ���v�/�ˆB�r?,���K�~���cӒN�G�d��-@\�kQB�MÔ%����+(Hٓi){h�0>P�'�k,M��͋q����M�&��h3mde��Y�/�T��(p�js�}�W,]%OM��Q���B$_�T����5��,K#�X��F����H��3�;2/b�:��/ˮT���X��-��b{\oB~��sD��e<)M��q%�<��"��=��R����3�Y��J"�U���5�p����Q�M����*�2J�ZL�W���7,U��Z?�=rB;�(P��Pa�R��\�ĥ��"Ov��Q>�e��WS*�t��O�tR�&�8rÇ��[�����5�i�T����vw��!K�.۠1Cv�2WF���Һ�E����ʝ��W4:*0�
q�3�����c��Y�h���K�WN�>���2G��Nhf|F9�〟�<ոj�tE�.��=o�٣�,+R��Np�S��j/�\|��h�k�=��b�FM2,dJ���K֦�z�X8#���N�EG9�,�;(A#Ή���e�� c&� ��d�V��ܥ��#�����V�
��O�9��-�v�Vꙻ�U�U@xA�q[�IC��u;�U�Y����[�q΁�@FuX�&FήY�{Ѧ�̀y�z^�1L��u?��`v�+��#�-1�	�{�꭪�@�ō�H��f[<A:+�=e8֨4�1D�B�Gғ����'4:��[$"V�`��x4@���Ўa� bR�q3�(d���F�Jp�3�����{=Ф��E�L�D��qH�)�;W�ΰ��V\;w�hȫN���1>KD��g�|լ$�<*��6��Ú���}�3}��5 ����T�D��ҁI��Z���<=s���6�3c`�O��������+���:�t���z�\� [���'��J7Xd���C�[4P��.ʒ��{�zvQ�?\���~�)f�%W,w�sjd>�G+B�jXұ��kp{#��
{��i}Bb,݊�I���g; ��ŧR��~ȵ�mDU�A��b1�e�=��
�b��($��1Y�����ԧ��r ̈́�+k2��3F����6�qxOY�K�R����$>(���^�~zf/WG�>xK�N��Lf���;8����'��]D�nL���l��Xе��쌦[&�<�{Rm��j�1��!��ڴ��2��M-���{(�㘸��u4v�O'�_����ɹDV��,�q��R�a����K,�Y��7=VӜ���]?H���4Tם�t��xN(DW�z�]]��[z����X���3ʨ��g[4��lG�����؊.�T�ԛ��x'�:UG>l5�w�I�쨌[�t���R���Ԉ��Y�g���<��-�н�jv�2�պ�J�����A��YK�����ϯ��CS�A��̍ej&��MT%��'�q�Y��;46��1���e}���P��~�'[�6P�.�ԧ�mL~��φx�0��Eό3@ �?@J��X�nZ��٪�#Մp�hSHE8^+]��S�%{b�� �����D��P,���gמ� )-�fJ�$İ��#���	����
��ʹHK��W�Y&/� ]Ȓ�p�o8�C��|rZRD�Bǥ�n #�ӊ>��d�Ѩ��b������l�,��8�0�h��:C۷��y>\e��m�ʹ{�ii�ј[P�-��/��A�g4����~_��Le:��C�{#�=;����h~�Q�S��\����۠���[���+�_��6P����e���m+�?\7<�U������H���8i]�^� �۪��U�����yK�//������Ar������Q�=uˁ�����;\繕�P�յ9Vn%��91�C�IN{���d�zxal�Ȗ���A�‗�������xs��sZ��7��Z3��K�|\��nZM�0�@�±M@�C�z��+Jz��l��sg5�9_Ε�oŏ��%�1�{Қ�(R�������.�fB�	�|��}"�.�,��U��[�37�����s-��wɚ�K��.���d��OpcJdX3���}�.�#�).��1�"����OB���+��Z�&�E]3\��l��{Z�b�d4#�Pyh��|�V�m���-y 2�v
��fi�>���نwTSk�5����^�L3XVȈ.0��3rǪ\6��?�@]�L��?�v��hK�y|�"|��3���d6�F?��D�����#],�Ǟ��|�-1H��:���l�٬�d��<@���95"��b���f�SMuǸ���uO�����P��1u�Ft���[%A�"u�ެA���/$�YY]g������ ��3q�g@Q�
�-��}��K@��x��B�ҞЪ�L[�w��
X�7v��"��{�R�H��m�pk�c�ʔ#u*���0���J�4�<�#@c�9�g�U���K�|��C��O���r'!	��O�:����Ŵ���[ۄ��C��[!��M�'��d*��(,#E��������sh�$LT��:pq�Z��{�UH
L�k-���)b�8o ���7�5����7A�F����0ahG�������[8����-�r��n@W�!e�l^1�v?������20�: �og�U�W�a�ń��Ezw�`@���?�x����~�E�q�A�a�����������/�8q��5:�ݯϺ�R��!��Nf�Î!�9̖��"d��󨢣q����<��'W�w�6����k��#��K+u�J�`�d�N�9��Rh�Ͽ(po���T��u�s�T=�/���Q������*�@T��&188r,���|��3z�ʩ⮖���Bu(����Bح��Q�M��X��S�u���ݥc����GƮ��!Ny����b:���5s^��}��i��`�#ƙ6�����ϳ�7� \L�.3��{�y�����q�1�]YW�Sr���*��lr8��1<l�@&9�`9��t<Cc�]���>P҅b�,���#|�5D���+�	�29]r���/\�JO���������å�ҒU���$�\ە�惧�4��	|E�N���{OA�F�<����`i9�����ƥej��*�X�r4��J�QfJ��[hA9G�R��68� ��C�4΢��2Z5soG����~� sma�<�}�U#XJ�fvs��ҟ#�HL�c�w$�?^0z	R�mC\PW}圶Wr�q�e���o�E�y�f~��t��W��jӖ"zp�]+�y�{�o�`�alf~�ӄq��®�7e[��>�R�Ǻ�<x�T�LG%wh�sr��m��B1Ì�EK��4S�Q� �d���c��Ns�D��OΈ��a�ˑʉ�y\��2Pw6�����pl��7�>�,��XVX�1���]�z\cxڪ)�ܮ���=`J��l��%x@��Q���G����֋��E�\"�?�50H{���Z%#�j�bUwBq>N�e�՞�ɐO��i�$uS'WD����Qʬ'D[�b뗰�2��M4�;��L�Omb$,ֱ� �6��3��U������w8;#��6g)��Ԍy�$�8?R�N����D��*.~~%�;��vt��F+��C�\���{�����u�f��}<gFij�Z<�e�!;%^㤺2�[��?�[�}aZ���3D��zsʠ�V�� �Hij��]�@a�ڌ3�����'��ԦI�V���H<��*D���ȭo���l�ON'��X 8x~��b��g��� L:.Eq\�ԩ�e�T)�6{4��F�B��]e'o,WN�3p�����k$�h�VS���Jc.�H�3E�uC�C��*���fFę��p�π:i}�NWR�b)Ob���5{S�q������<:���m��h5�.�"H8'��F�L<Lg�Qn�	�d���Bt����O�N_$0�tÆ6e��(��2��-��7��Hi�\��.�uٴ�$b��q�w$!����4�����F�������H� I�h�@K���
��&a���H�,_'���q�./�%����[������K�7��Nķ�Д;��\ر���'��D�N�9-�x,��T���ؖ"�Q�՛���H8��S���Q��ⵙ��� �,R��v҅��p��������x;���e�sF�hQ�����e	��WB����
]+$=�Wg�oz�]�H}
�
!<��8���\��>��d�� ��hnx�y�󸐃*�$�,�6|�vw�6��}fuǧ���ฝ�ߑ��TL�Z��AK�|�,3��i���𯝤Ԥ #>���&�ϩ�Q��mG��% �J��'u����䑯��	��e-���e�S��O��TI�CE'6��]�z)1�s~`tN�ً������߃��<���'.��e�N��0E't �k��]�J���l1�aOip����GƋ��G]��u+L�Q�{&�hH���`Ζ��
�įR�_Yu�����l�-5STk���
쾄#x�&-�;�:��(�d��UQ݇��\�V�R�$�B������ǂ���˩��^E� �[Wc[G�d��,�ƸK,�.e��� ����#�>FF��bT@� �~�<�.��9���G���9�O�ZU<OV9K�9����r��ґN�lǯ�2���?�.��d����L%3�}��,�//�^�
���,��
��~4}BCz��ȿ�n[�o;h�<��za�������7{�G�q�M�����If0S�=%��&IH+�]傡@V,;�*W.���=�1��}Yil��X[�C���i�o��I�[*�O/�L�������KEH�h,�9��"sꩌ�Hw��bBW9T���*�b=����ư� �;�8پ���[(�->��=Y�
oz4WCϠo�}�C�!�[��D�m��Cl���?��K�5�y����6��Հ&+����
��وiE��W�}@T%��36Y��s�����! ?��M@�">��rJ'ݷ*se0������>� �����*±y緝��;�r���NCY���̼���2��Z��� j�)Xu��α6+2�(~T�Zb��m9���{��?�����0�����|,L�X�uV��5Y�����&%�e��Zb���&}���*	r���w�+�V�)^�J��8��S:!p�뤠�&�a��sV
��D��Y$�?�5%V\	�Y�	�F7[ÆC�k1Ͷ��4�O��)yaa0���a�2]��.GB��҇���MH��!=���]�M���{�7>s����k�X���2����p˾��n�s���W�`���T���q��F\���9�Bk�Z���q��W_�. plo�����-�-!�o���^,
�:��Ţ���v���Mr���НhW�O_�f�FZ���ۑ�5l�ɿ�X쩬O,��Ct���ސWa�I9�y�.z-��54�P�ꮛY��l�Jae��d`���b��I.6���c}�D�͜��) ��9mq��" )��Ut7�B��#���?Wa %�b3>�Kzc�Er.��2�/��Ih��1���C���.� ����ׇ
O�,m�$I=���ѝڣ	 ����" �{�E`��=���z�dc�ei�G�q�H f��V+H��z�I�����$�@�����X�+�E����P$����nl	Sv�%��M�ʜ�m�M0�����&dp�K��w��j�,i���F�[�K��D�=�ȑ�OK(g\&�<@=�:Z%�93����������~cNێs8-�r��s4z�3���r
�4 ,���w'�M$O8�J��x�$n���! ��e��Ob%k��z�	����\��K���r�A��jAp�/[	ZE�c�$s�'�a�g�|l<|��r:�֖p�Pę��ddJ�0�F`c/+
���:`U�������J����ZR�����'�ammc��f�#WQ|訊`w�V�j��Ԅ���Nu�M�������1��?���as�帳�*ڛ6pC �_���Zu>�),a�$oRYxi��y�'#ĕ�l�n�C���mֽVM�9wz�NB9��%N4(�QY��L�}m���x��;����+���EˡB�iO���KU�Ю�fގ�݊Ly%=җ���Zq�Vϼ4�����bMV�h�o-��3�	n|��eJ��R0�D��W��9�����i@.�����.�ڈ������|�-'�|E����rMʜ���Q����M48����ii@�}����s��r��7�gӮcv���h8�_�/;��w�Ħ)�v�z,���d�dd���v�6�̪�G�LJ���8E�}ܨ�\#��zPz�h�ܖY#���� ���7L)9����� ;��%�&��E�\��"P��P���0�[Qr��X�a�g	���>�4���Z���&��r�LN����Iu�pE���'�4rHAta�]�yШ��J�tu'�+^�c&�r�u�	����r���[�5���O����nF�����k�&��:�W���O*j �y�1I���$�'E����b��A���ƀد%��}C&f���G�>�d�F�[�����]�p¾�z�N�P�J�UҊ��
��k`�m��"e@Յ,�4{@�L����񖞬¹c+P��lI�y�:5�X�I�Ӗ����.	2輬��~�z��1�z�\"L���w�	�mc+W�!���]���x,ʸֳF�}A*z���x$'�DC�5��1�s�f�
�c=�y]���..�N�W�L��@��,�j.�H�*��y�m��I�N,);��&\����N����?)��L���<�P�+��	��ή]���{�n��v%��2�z:׀�]}f�}��)�� �K��2�ߊ�+�s��7?y���R��f��WE.�XE��X
t�W��S�o�H���E��ap�S���(�	��Dβ�����+��BR�[��h��ɢ��Y1bSuc����-�z��k���6�en9QCTj&�`�d���������Gsc%W��B��M�ْ��@�c�F�Ӎ�b�)�E��&��5r4S�]n���%�;%�@Ū��C���T1�A+NXq/
s:��Sg�֟�oe~Qrv7������$P`�5�s^�pr��^P�5�h*��� ?ՕR�3���� Z)q���z�#D�
C`먚����͆?��f
5�m��PB��,���}�8�"�8�	f����=)�\!V�?hJ�D���
 Vքt1���Q��*�V4��B&E�x�n�`K���ʘ���!��� )d>�%�:f�ʜ8z8��KM^v\��c1�e�0ܸaN�b��ek"0_ThC������AIeaѿ��6�#Hx�v&y�x��	�����I�)6�*�[f'�7̧��p�:^��!�٬픿�95��V\��v���~��lw�Vu������3=��Zq_��(q$Z��q�{o]@-U��@���[�Ӫ33#�=�� ����p�YP�#E���D�V<��Gk#��n�ɗ��}��{����:��n����k/�n�S��Ts?����R��s��9�S�\Q����"H�~��Hf�3;+��S����3{-1�)��|�g��/$��bZ�ֻ���%��p��=0�+���6)���>un"Cs:�Z�K`@���o�hp�� Eĸ��0����.�ԕO�[M5^�=<���=(`۞���RKḽk�VM�k�PT�09`Z���GDm+Z	JS��sm����j[y�a䓱>\�I
�����?����o����1�����p��KH)66yF�B�h��7>F����-X;���7�wP]Ȣ�b�ȉ��h�k$�큉����Ո4l1�b�o�$	�q��7R�>D��k�����\|~<��OL/}y$������s$�M�06����YN���znѺ=֋���ԝ��k<��Y�B���=�x��KK��ݪw�MqB�>�֢a�D��0����@�^=�*Ԣ�UhN�M�QA���D���z�Ь��H���pJt(>j�:�lC��<�qp�V`^1�)��G
�D=��j݀��UA��ʤ{��0"i�a����w��3� @?�VӢ?{����u%�BM�Ѕ�����h7w=���pi��l�bT5o����_�5C[�R"ZD5���Fױ<{�����$0]T����h�n/� Z<�yJ�3˹��5(�~��V}	�צތ�0�0}��O7'm���f��ucÃ@�Cj���Z(��Ʉ������3#�����t|2�f縞0�b 4|4�W��Rm�g�J{���t���"�}� L_���	�q=������:��1������U�fwv�J��AY6={���S��8����$�ٯ�u�"Z�/���ePC@������aWC��WƘy���bźQ�}���(�eH�c�ؘ�޳oC����!g�ї�[y�16W�K����L��͝��|�p�Gf`�x߫��;%B��5K�iV��HN{�~B��Z��9��4
ܙ��?���֊�z��o8K��r�5��yk��
����#���S��U]�hx�S6Zn��#n"5�tk�vO��ȳY�"�]T�����"�I�|�w��v�X�#wb���h����f�����BCq)P;��}��٭3t�7�Pl�U��K����3!��`ս��Db�k=_���!p>5z1����nj�z�������§kzn?���=��bq�:�D1�7�r�@^�HD ��d��s����u�/� j++�Qe�������Ȍ���*W�	D��]�]k�����P���!=o�ӣ̶�u��W�U
f��:��9a3�&݅��#>�8\�I�kt�'���L��pED>�@$�ד�y���$����U�S��dΚX�O��U�!�cz<����*yz�`���wx!<e��Sa�WJ�4�G���m�$���]�D�d�����L��GG<	d��܈�=��ن���.^��ì+�ܥ��L�4F�-��X�����p���-��홪����L�R�"1@�/Ȑ�,g�����!���a�`�/&�W��0K���iM)?��Lj"��ݞ�����~���h�Q�/���ULf�K5��#�E���̦y:���u�Hj��O���݉��F�r���t2����A~���P��w��D0�&#�C ��bqJ@��;����CgeL�ѫ�v4�'f�~��R�rܹB�g3��Y<���A�U;8����:nܵf��q��%v�I�?m�1v|D�f5�{r��t ��ꤼ́�rh�����ILo�}��c鍋-s'�
�/;3�Q[���2�SQ�.{��'�