��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�����^{�a�ȝ똭�(� ��[RҶ%H�
�-�� �m#��q���b�!$�uw����lq��ԠC���/��দ���x��~;nM`���d���n��)sǏ���@�ߟE�B9�z�Z$U[��H'ͮ�$��	p�@�l8@Ȃ���R��l�|���G9���el�Z�X:��Ol!�L�	֞���ܟ�ۇ �P���$T`���B�"������bxx��0�8�Wz��o�c���O�4���K�b��f���A,��Uɂ;d�}(�.��F^��!��-��b��,;��E��V��E��샫�yU�;����(qQ��,v�8��V|}�	�Tz(�G8�)(�{O�u����yæ���'���K�h7P��"��+%�y���%�TG�a&!b�|���kZt�ː��Ɗ�U�����6�ؠ�
" &љ�N2*}~{��������!d�%���O���"��S�e�Lоv^UD�Q2��9���l&��J2�z��� 	���f8d8�	<���<~֭�C�{�i������,[8=�zV`�~b��n���������z���Y�4n��Ң��$�����s��G"l��5��]܃�x.ڏ�T�S��k�~��t��ݕ�v<���&��y��R���9��X��lP+��N�R��"�q`��=�d'p	�6�n�{_�Q��k�|-�q�;��_]t?s ��5��`��R��_�$��(�W�h6-?���2]W5�< �U�>���P���w݈���+��"���Si��z���1���,6�=3,����)r�6]�`x\{T5?_'�����]���I	`�q���yU ͔�1�.�$�1�C�.��)�*�&�7:�|�����Vw:����-
��Ol�����3	�\'f\�pP�n.
�.a}음�'���(���DÞ��`AȴB� YZ����y
Q�l@%��@��k[qQ&���i��Aހ��c�^��r����\��1?�Ȫ>����C'\�3j�>>:�N������fDKBcIȊ����t9��+��s�0͞��|�"?31�Z��*��s�����}�X3���B���^��I��u)�I�`kI��;!���}Ҋ��"TT,��	�l�7��m	n�L��
0�g�"�"��(��n��� �<)	�\�|��	�?p��\�YY�q��Pݻ�Lߎ�N�X����M�.�&�