`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F72Ogi4IG+k99+LOmqotYnqMtxWCqTZnVti39hcGWwKaGqLktd+WTOtisf71bzMm
UF5oLVomRMZZxsxbNaqLXbAbwLolTQrznV84PWTviKTM2muKy17ncPMGyK4ewxMn
T+dE5j4R4l2GE+zO0dKJOLPJfN1P2GxrFQ8R4uShsOQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16368)
Gq4NdKNBvEmfBxniVQQpRIs7DlQaLxQWFm+GRKHdbqzi+lSkTzesjU0bKazTtrgq
Js8qIbGogNbwQIr91XYRVRXXKdKNHZ+ziPtTIP380CsLA23iuuT6LGsqs3+HJ6d4
PIM1q5+2Umqqna+QQ3IWDuJB78DT6PqJc/wCoD/YCHwm0vBkZySAg4JC3Svah1bp
N8/uoi5SiUc91uGuQ0iR9skmjXzj/kY14DE8BrboH2Kg52NloOHmc5jGuFV4U9F+
lnbfyd6klyBD9sB1vV92EWpJ8MgqDxz0xu08UuYT/KqmFo8yClQm8c4no7Ew9OFj
zZq+xNihIyzhgOJK9EKETjfkOPZ66QroupuzF9xTIMYkeqoTzS8J7FJuN5JMVHsa
GDWtjuqc/zdhEPaR9SiUDNxs1ID/IkEvBWLXe0DQtQaddI0fHt1iSh/1rk/uD1C9
wsQOrlhoYD/zImEgZVXiPr6V5uOJsvvo+T6L2BGFqdkFizsRpNOpuCU6P4g+U6kO
P3NW7PfxeMTMKRsuvQfnXMfVsaUAmr4gQdQQUUjnHR+BHzoXM0+hr6SccEOu4cgr
3WRx21jswK4et3fIeDqYwGL8ZbMMh/S0kpAHLOyc3oDG60bEno1I073Hj5jsQpLB
lOjFWQlAwMriE4DuPK9Rr2QEDw2vWlwuW9A4IaQK0rJiurGp5O2cUFnHApTxOepf
h7CeRL2o3nBa347GmQ8jPwlWMROEnTi1jN0wHNaa5Hx3vhisVDE0ahludoow9MtL
kWmvoPgkdc82gCN9LjAbEVNTktP3bngzXzQ1RVCslf+SJLaYezIcXChixD2diuwd
lEdiCn/LXP66Uba3XCoIwhW9xN2jwiptedrhniVwkZQ5Uks5GpUhRid+ROzqNnhr
hxCJmtLMykUPbJIC3PaOojB8XJd1eEhExCvI8j3J3394Cbfbm0M/8RXdi0hnOMBb
xP20/PCDXuY+j9y/fSdLYj0Wur/+d8UmbCCjih2kl56ojI5l2bMv5z9MmMn/S+M0
zOynW33e7XaW8JKBJxa2oagfdG0Y7tlhO4l7UC/qUTXxgHY63ncAezI1oxRTs0a+
RJJI8WttAj8tURFGwo6vhDwjutpi9QPEq0SYF4ZUW+QT71mS/zf4VjSbxbGNodId
fH/mQQcXnT3DpbAmQvK0xw292iRl2eJ054DFniproGonBg1AWFHB72yORHml0l0e
Q+nKnlD6gYYXUsoTrO7qdgIGDQ4vRnSy+VEGrKdFJcHpMsOHrotO3Ts982cZdj35
pcsbduuwVGHA6dr4SVej2lz0/OWBKWVY9jZpz5HlqvMTZlj37SBnV7iHHj7f1wtB
H3Ts2441Zwm2JUmievIMvDHnmzP4YJEgnpW2mDCNxPyNAHp49juvYS0r2vSHzPUj
HqXVHm43yMG6YWqh3ZjEm/JtzKDGka5n14l+PYL8PyLDDeWU3buv+EF+pUNr7Ody
T1iIrp30vn0NCjxC2t8kqoQHtyZjwk3IZk/OXWPJUoriXRXv7jnIqI76HKOC87IH
Yt4xUYlHR/tYW4qAMSJWyYdT2r679hAcwIzCRtPFd7B6USoA2Oii7zMxqcau8dDv
2XzFtEvy0cIBsAbo+rxXP4+UxDrerlghc0GDoq1xgGiNZXYC5T09r/Ij/ILLznOi
LHd24cxv8zI3K/eCE1eToeIWBWhhjyVVLakUQhrwbK9qlvRMmojKls0Aryv01yXu
0HWZ+lSk5tATo3BeFYRWRN7HCcRQg3HZ8cQjrgrKz/j+XyKwZKT/ixA//J6mZwv4
T5NPYxCqFzHSK8N3pTRzZHi8Lp3Rfu9ohCv6qL8DD/X+fEv/GnYrArnIimo7xbQZ
6EkqyZASgJweY63IOil4fSx2m/43NZpHtoT2fxcJJnrGieBHJTDvelk+yxjFKCr3
XNHxevNGvWs4YWes+uj1hET2qK6NGydAjLFrYNRDtkkSlTtHa/rgYR39FVBhJQhq
zskh1t6+4wiKtUT4Fxh9dAB13uXdocSubYP1Ua/BrE3bVQsOsiJ0QWDky1IdfOXy
ry22OyDJUn4xJ5zhkOA6dKy2qEbYVoGIZYJ/58wD3mn3NRFuRGXBiRXEIE1K4Nsk
mO6lUBWh66RfEAS8HmBFqvKXITQWir0rfuu6+Y/FU59nUM7et41WOv+DyEDfBakH
wGRhFnt54D9XKetUoxHJZkK4H5VegpgVIYdWiLo5KlMGa1a85MYnXTcF+xaR2mZi
dNFDWFcREzK3ay5mZEsag8YX2E+FlMijUVmU766OZpstkyhu+cWjrewcL4SpEWnI
dKPsU+MECeWQPdq8WHkeqZWjj0N89hpKjanwlq9/Vz2WiKP7PwjTl6l9fq1hUeYA
ga+olmaFlGAjb9kfX0LjzMvvINYQIhRrxP1t091JPsYUyy9y7ieI/SEIW1YqdZLa
38YjAh8zFcuW3l9qhJlWxzjYBYFfPmJIsioIPyecBolnghcz4li3WcXfe5AqZ8uF
1kG/7J7N4/b0nNtofM4PV+PKsOm/fAUF0aqEdqbSm1EajvsaBByBv4ca+BLx/enS
EMyAV92dxmtxB/Lx5gcK/ue+i+ahemXJoSiO0k52Ta/DqtADXA9qtx2FHn9ZwYXo
6hQ3I7ngSvKa1RYMEE/5qUjJ5O/Qm8qH4DfIb4Dw2ejPBgOK+DYyC+zyV1NtyP/l
Y62jwi2DfcikLonSd40y2wsn1zrJIPkwNflt7TrnYeqwM7AauVY5FZsIMcL2oanj
Wmx9BkwY3G1XBjFannS5hB1Anjeo3eHLD6LMfT9lIMTXjfLxMA9kUYGip89zuEvl
f90tzyL/HKY+akKJtFIgTAXkc0JW1vEmPVdgnTOu6JcF74MRkIg/sDxJFd9SIxNE
0jhXRZzMnp8bgqNlvB6WTn+YC5SPUddFrcEg+vAnz+p6sAezMHVFFPpit8fvJLVU
xiej1HqEp4xIUzBgpdIO7N4mqWg5HG3Yv9YpWF9yh36GYHwG9PFkOI7YnPdl8iyh
vyPGVUpwGLsPoSdV4WUkKHppOkCvkd5scUuPzMD1pXwYB8sjW/gM5C+PkqlqSb5p
tL7/FTE9CaJZH9wLR+tG7K+QI3Vy54PSkUS5Rr/nsffiEYXtCKeO7uV52GZpbWwz
zyYaJXoKBTqSU7yKDloG4YhvspCYKf27Yi4XLvtRVwsMZjnJyjal1rHoPjAvrXD9
GDpVjCiF22EjpOBwDaK+Y0KGOflpRQtujgSvkqgnIUeZfE9M9thVM2Z/KlXfLfQd
/TPvbwp8LsT1siOjCGUrfCPsrpJd6g+z5aIHcock1EK7zuhrnmk0hLzo3QBb94rz
nJMJIuBRziQaT+u4RqwzyBlrfAClSy1Kk0XbVRQsSE1LOrYI/QeDzAjybF+w1Tww
oI5LwBn+vVyU3IgmXfeHnMtnWlnoW0R4xlL8Fckc7VDZ4roy07JUauK4Nf2DoAMu
gqX8S27eyxkekdbpDwg7gkqwCLRfbf/CEq7GmeG6QI2QQFnjdl6h1y6QdiRvk9bw
yfcPP3ygrkhJ2hrjWtNuaPYHva4WF9K2dQXSp4ooF7B6tRo3goFa0E5ThvoZfw0L
QnaCKVB+ajmqeEmBRqxR85dbOjD2XIDVbAJ9P/pHt2ttbgPD2w68MAeEWcLgxI7r
bOfErbxcOKrTtjoKUaoz/DXZ+lEFOk0l8dJd8ML6lLxuD9aaVsbwCfPbXm1O2uWD
ICsm2KSLC+uqtgcHAYnoIOIia8RKJg5KQOCvDkmVa8IYKz45ejSpj59wBd0LEcLY
0Stkq1gFbY1WkFIDjFUYXcZz2fs/cwcxDsmSzlcUjihXd1FiMKopwUYhi5p0bj66
i91Kqz1MruiyOrpG2Z8C7KxrSSHE9VrciYlYYiRR1IRsmkBfXA8TiIKiinG1Uxaf
nXXbLbGY6DdpTfPcqcImgKyxbZpg4xsPveFW4KqftwwntOw6HPbK8OMFOSI6ShCN
YHORUECAZotAZgySUsn6yYGBxea6NR98LDvrTvoyagYkKKLMTd1noRh0hR72kr3x
KngT3csfpEDjnuoIkSCxp+5c0Y89taroHIH6A0TKFZfKnW6Gsv4qeahIL5qVzsrh
3yn+V5qwlECN0xZL2X7tlzULgbNT9E7g1IKelt78Ofzte0JgMqQ4pOOIEq+C3YyM
+f8Kwh46EDohXrf/r3cFDwd2og4tNiHD0EIbOxSQLeVLBk9zQnR+5e+dVd3rWtEF
QcYde4Kaw8RplC8QLccG/Mb/X7KlVX0/FG9gurpFiXUahOXQXEhfvJteTJyRXhjy
NgKGuu4ljSMDUNsUjo2lMvEeX0LnMnjuAMZbZcP7ZHoBnajUWoq1vzKZDZdZf1u6
APkcWxhF8ZbzeTrhKwk5dvyzkePlkyYqV/bAs6+q8C67biNKPeo7cdVRF5ae2u0B
qSwv3kYAJqMohwiNpzRt6vj8V1Ki40qmoj1bk5TfCYVXofVXrBc9R226G70g0iRP
EvrUJD5HZTP4e+t1XA+JSf4OWJCajGe98pabWV6u4OCkfPDb9Vlp0mvk3WT6k9/X
1XI69iSYimZbAKxDlg6ApzV20kiZEplu7HJJFis1LcufSv+iMDQGWa9YT1ksaK32
6vkGPX8bBS9SvF7hW7dTq5Z+O76jCrtT3P1dDImHWWfqFSZ3c8NdEfhxA/NEIzgF
Pyjt5jcM1mFqhlOwjRTkdk6tMGfwSeYpAxudOlKCxCzVQrj6evgnJen6AX8UoHMR
3VcWIIbgbs7qtUs5vXqSI0JpSO8oI04VHY9QqYykRzs1unFF/6UkXEtyCCvIWL7/
4Xzi/FR7lIKlBtCs9n1ZHa7LCwmGsnnmCW4n5xMIgDMrzZiXQ/yxHrYDKtcWwzZS
tSPPm/gg99QGv8WdjPywfsfnfI+vsZFiFXtQsRqVfjAER5+W+lVoZYJonGNSVSV4
C4a9IjkOAW3XdLSka3Kn0zzjaqBSBLeDwedhZ7A8XnBv/bFDviM9AI538XE33Y5T
zdnX3COV1mJ8RvrwZGmSsu8fKtf6/L893nNU6FJTQtyxhvlEv0ZJq+wl21v4XzZO
6JQH35FEWU4wlAcDfwANpzJyO++pVhxA2VGwa1yCRdfsLrAuAdav4JTt5vA0evrJ
ZfSTK1VF8WbAJIxr1w2xeG/wQcMAYpqmHP/UdL8r2Y/NzBaEgeIb0pZZCzDd0dI8
i4DPcWq1DUPVvaHQgitvfRv2tofySVx+aF+ISN+7Ywlb6iur3YMcqFvINEtLnFPb
dvx/FdS8RFc6bSt+FzsfouDqVpS9KYlfBVstX+l6txdsHxqyTpgHXsQl76xm+jrR
9q4LsCIpYwdO+Rxdv3Rx213o1th34cop9a2HouYDJIinWeWr0emzQkFB8QXrP+SS
aMjIsWnfN6tKJ7Tkmsk2teDi3VsgDsT5bUXS7FugoGCtCBkZ/R+SncK6sGHhoMJS
BjJAzkABbSgROXcnjxhrvtr0R+rOGAomvHEud8x7RZ9d8heWidV7c2adVrEPWjlq
XdiDttMncwIGJC+lg1TOZN87ScLCEfLDmMA51xde+ZCw2n7u9nnKOCZ6lVlQR1Az
0DnKyPSwAh42ysQzYFx7/lStRAJAU2B0TL3pL62L5d9+e3sJSdBMasic9upxIUAY
1gwmO22Qf3Wr11bdOK3PEYj9houoEBxYmoH8DFf78Zcf8glykpSL9U3HlrpTn6h9
TPJid5oAq7h1JxbqWZPNy+/JJOyDHT12v6aOdlKSqfxG8wgOu9p6PdCr0Eiw5t5w
3HINrXw5qT3JYj4xovtu9eNgUSgdjulX8xkqyzWmEFfsJIg158vxX5lSnRaBJRc8
/G/drT+dB4orc6Xwu6IoCS1kiEQHX8g1TStFt/k8vWR4rf4Gn5MGPiPuBQQT4KU+
YvwVDCRoMf3AdgN29reI/wCZSLMxJqDoDVDKjRK1I2Pi/PSPENGOYAuqlFleTgzN
UzQr9hotx54ORFfFkQrP6IQNphtj53PHl1anVqjffCacuZUT++lVHQIDMZbfDJSC
6vVm+6NUx2X7QIkc4ojQjCV8iQ1xffqKCEJ1BLlURmx8tac6iU3bRhBzA6GHP8V2
gA6zcYWgHHGxfyZ89Yon7Z5x0h2fiuxG6uEi+l6rngBh19jjZ1jj307kFygcSKNK
Xb7dj8BMlDpHamlaZkCcJn9gYV+iT5hdH4F+NQ62tEQwyYkXk4FitQ1JYTu3LuPZ
CtwKpUqp2GOa/ZMddDq7CkuLZPj6CuXJcK0HiCFS/3RupKHTqqFZwn0J6BGXWPoY
iRkoh2yKL/lLmt4gv7GWPkNiz6Kr6+GGvi54ZHYQbAx8LvKb+WawYGwbX/cUklXq
AEm7k05KSL4ettCuVVL0sWX9rh+HeyHHwBwPLpYWgqT2rtC2oPk2aIIsInvz+noP
qVrMF/u7w66GZ/mnl2k30LoHEcwtAmTP71REFqgV98c7VVQ6OADpdUi4eLl/GND7
KyuLVEg5oEGyyCwvjfptHQcJiztWnmkl7oyr4sLBRUR5zavHA0PlJLocia6YlJwo
l9q3fzKFfXnnpXeO8kUkXP31IzUc3EBNgj21aIhRaHj+KZ+UMR6038ZHGlrel4qR
QuMDNyXECWauGQsH06sLFH8M9M5LfE/eufxoX1XRYg5XyXPw+KVql2vFuRz+v3ld
2dQJMS+kHZuERP4vOSuJ+d7v9614DJryHHWTh7VX9w99KWch9mvyF+QDPybakmB8
KV23HM4ERGmgtzsVOooZAIK72b2YZPAMDr4PfXjihQoGf8t+O75wtLGTUqXer1st
6oGFIRqayrwoo0xAtTTT6vRBbeJNncbLiJ68vMqEIy+1CPegRXcotwgpL7rqMcS9
9ZQt90TjObXu0pIklb26LZh3RHIKEelml/6MYk/Fxn4q28a5tKqbxOrJCAo0VpyV
nxGfgotOHJBnHiAvM2wRsOVlJ9g7uuXYKArOzV4wfV9MtA51W8adePcIk6bll7MW
/txOCcV6kA3MMcyK++7klXx3HduGqfd1eqwvkxJsZlBqO4QIBBwqPf/dbRvTNLnN
cSLM1WxXcSZ1BtU07i+tMdvD7fNI6iPpnFYih22UAfY8+uL62YgudPF2848MmVr8
gupnsPLciIl0u8BQB1XNKAgmVDr40U0V/RwcFF9yvKFUWycDuGqvUt7cZYZ6ne45
X3GH7c6uFTMBEZZE+/BXIXUgZeJqFzZQNO99hrGyijYlNgUSIS/FHIHlsWQ7zbkt
hD2ISKYl20lhA653PBYpAjdoGXTfO89zxWFhJaXTHjviZOTZ6I5xiCKfK/Hb3N3E
IVr09m9golDW/G14ZA0UKGTUsyXFGuZ35i8+VXvoUziHlp7rYxZWrA9V6vOQ4Ohc
VdLRbXjP7kOGiZnXfpWKro2s4A2l2pw5/rCn30Tpo0X66f0Vl2clDk1lNWmvSwod
dNS6dTvIs3ghP2SBR93bJmOtdMZfTjx43JPzDwc1HHsi67e50rjv5HOfwSQ2J259
9yVZbmAE/FwX50xv/6+WJ7ZDLn1hSlQVuedSmBpLdjEld6vJQvJXB6M2YIDh0egD
sqB1Tpb+zWGAtf5cPfV2Q7/EunlSeDwyNrx/H2uC+sVE08iiyOiXG5vTP2hhYEnw
ejgUkMM9iF1bnp3Q4jBdEstQnHLi/awTL7y7ss5J0pELZbEO9UuKmOGh5MhC5Aw4
hJd4NRla7JS2BgKsPsl/oWXMUmt12ADMmupimjDTXKWiAT56s0d6EzOfO5n6svQS
43DE3BbkuhBPdH8um4Rhofao6gi6pe9f8xSrsFY0np3uoAFmFIWvF5GiPefMurqj
Bhjm2F/lHZcAlCoHsEuWvMBrcRqRRNWMI/aOrdvF5WCwg9keiuurujzjSePxq0Eb
il0TXo3TtBzJTLaeZVbqMGqFycHdugUJk2V2FaCy9y3jiwOHsEqkavBrm6tkqqVz
vJHn7m50kaVk6ogXLKcTMnhkXzFfPD+iILyjZ3q25Em4GIJ2Edh0BxRiIz1YUp9w
xi5mLSWxBCz5xWhKLbc4x3JWG0fUA52EIKZPzuv1VYtr0b5NWBhglvMhA5kkn3X/
IxKQxG0WPSmRf+nnBPtYP+sRvfZ5x+qwYK9MTJ+eYTM4gKJBQMKkhRRz8zcSzRQs
Qsk26rTgKhfWkRhEATYdWI8Mdgxs1CspfHCT2Qfhr+Ge1yZxhaYKBvl+fE3YCc3u
nUMnyApjfzWy5kmo91XXDeq2Xnsb/GOcK65ssJvwYdr8nvarlCUWVaNS6DSK+mZ9
tBiHLLaw5YEGbfhoHn/RF1r3VEgDCDj8K46KdON5p3ha8lO5B8jpcaZ22TiK4GKl
Qnhk+XmnFsjIwBcas5qGWaakrLYf1fLbmPOMMOrB4Jyc9pET7kBxkJYTHVnSzUYF
bnQ/TQF9/js6dbagt5Zr0NXE2dtoTkxbFS6yuLomqGYL2GxQ0SAczwRsf414Iurz
Dts9+UNo0oAQX8++mvbzUsPgSqQrgEICyFR8OvAlTpcdTNdKekSiZBpdi4VW8xuv
Dmt2wJaw6KzKTqwVR4mFftnBxupnQSAiWWQQj/GJpWJnAFJ8FvQGF2x/qwi85k95
Wjq7/FTnOfj1/USGQYoaUW+I/9ZHIo2MJSJRJ53mNdpIcz+YmqI50jw5u0r8X6VR
NbmEW5eHs3uaTlq1ZhubVDLiHq6bb0Z8IlZpxtU0pnwCXYprE9svP9npV5EGxF/5
IUCeqVdLwjEn4M3a1WqnxH+E0tD+Ntj/oovtBHh/E5c0Zudosb065jyPjdTJLiwj
JW16v95Izf8uYLb831Tz742nl3ikXq2PHhNEhbCCz2P5Da/VaopHMhwuL3ksvwbR
UMShtvkaZ905apxxiY9zP9DZVyCB/OidEv+Kbf9qvrBjta+/NvN2W2IuWjILVpy0
vuT0Hk/2OII3bpoGM9SldtRS8yTbvgy0QCYAus/vOfXS0t66agtPPmcYrS/dcZRh
7Lms10rE6kXdWuyZF2gWQtGROf1ngl+TioVcAPNXFut3yMSbm032zHS8F0z1uTt9
ARpDpm3Cks38IwJagpzKNeJvT818LA9RXYFBavXdN4TY9Fq9cPczJ1oJ797weTsg
uF396/jyrBFJOOkQS9dhzE4Tt9UyMqN/34RiaatT9+xhn10IVpTY3nFBrVqc+8VS
0iYrSuSCc9CPqPwdfQbAKvTTMGtoUiFolF5ry8t6CQi2IupFCRAHyJiay1ubHWJT
QrxrynOX/dSnla79ycjQ7i1oQgrpDKO88h80p+iCNg21QJ8e9F5lKRCcnyJTy+oc
csCfsAZU6bkh9qSCF+hi6i+ScOwMqbvrGWlZMp5uovn9RC/F5I3yiZHvZKitKSbc
y69+oOIq+SRPKxeNBEw/dSc32lPjT9kKCsiK3nUY+nhP62vHU5XmIkrokoVD54zX
xZynHZ3P8/n7/yzBOldQUQbXd/dpNO9UDgPCMA7zZhxu5Fay5VuIhtW3ISu9KX0A
lmFO50RHRKpAX5jpj5jnjIdqeJSNz8s99/Qdf3R32iwXPBlZnB0ZTmySmsevS5IT
Lzb6wzYlFbmri2JIXbL6L4STREwrl4Z+uQegduZ30Q+wXBVqK+X48u7U/db9GNfH
5TnII8vxeaA/6kAYPBwlbrAb7/SX2bd5shjYxVoWbdN/iOl8OGiADhMwbG+wOcH+
Vx63eM1FoydTxE/oSYrDJ6/A2JPoKGuaEe77dG/qRIcU98Qsw9XMKyrBLmKutBZI
0RZoZiSD1jD7gP27eLRylcmnZ/vp140CeOAmOVcFYmoDDm6zCzJL71yKrP9ov5St
wKtc0YSQlQH9owSF+RM2Dc4UvWfFOENLvurDxkzVpxnn6QOFfkX5oVora5bqpeCv
FKd7hpSiiUjCglXYBXEZjrwm2ZmbMhWtabN4GlwCITkSwe+iSG2pWKpSNKdgwJtV
IerhqxUsnuJBjgEBos3WDoAnZEDL+uYW4vDn4DatZKNAVKQL8n+FMawVdafqhw5Y
W6MwbFGQ648zY9xf2oakOTv7Uwi+X4pnM8XC3Vbnvom65fS8BNGo6orHj81Z1sUI
dKlhY3cURIPETrzqJIJfG32LkkSLQu66hirUC/QMnmjw2tVc3R1Fcdlbf9U1Ah2G
3yVHC7a05sVy3rWgUJEZaEpbe+Sw42dVtuJp90ywuVCVcsY0chRRBM0tAP0maeXx
8/wyRrWAQqqvl3tfV5pvKfdAPPiXYbnmlxNUj6CnXQDUpg1dg7vDIKEcKwJVetNK
AqDzYa0H/RUu/uf+AqUlRqeDxYN0lOOlDrzK/5tJ9tBcWLRcy0MPsP/7/KzK5GFc
7VIsl+k4lV+YeGRs1+PdeP7BtHw1xH1KnYbieRffBb1n2BSx5C+eRC7ylz9JVG0d
I4BrcE6w8Lm7VV+6ZvBDutTs1/5oyo7Yvs69k6fxKuc9zNY9VR8vzdZq+SKI/hJV
HAROeAdOqarqfNMODj55Jdh+tGwdq/z3Ac8Mayo/lBHo6u3EWrfdWVqS2nMnw+it
GUwDBGmJjeWOntq4i5Sk8Mn47r71YnhEcbXfM3atgBshPlMOIKWADDGibOlUOqAD
sD4RmXfWSVqKhcGnoJlTmOr2du5PFq2yr2mgg5zHHiPKaM+E5RkQ+7Xyclw7NVCE
Ovpss7+36iZCwO9fhqbP3AKmwE/G88QnMvmZnT+dQQsdFgW5fYwRODHDbX8RguIj
h1UbTL5HVPayBZQpEJrZH9qADy9567we5+DXaraISZueLhdtNTat7fWwt2RMHRkq
vl2g/M6l5gYyP6+7rmkLq/EPTD6CEap9FkooKuvhk1+HXQINkqjFA+E95QxDej8c
bSzJHIxBq/G9UzlZQqlB1nRGRirrlsYbtl3CEwQPh3d6tZDtnZiUdskIED2gsEPN
Oil6cQTyz2ja/sCs6/5tGhk8gYik+chG/fN9xTGpuBFffS/pFWVvfXPJ1W2iXK6M
M9Dfz8tJLMvQzhij2pkrHMnvr4hQanNeGjlTlEaWLzSwnVH1ZX4XI4JPpzNmsDm+
dIqgtH5e5599O28WDyjW+ZfJlhG6wj5TQs1fJ74LC5BEX82jsXZ0YfYJlwoNSp6x
n0YmfMXNNaAM+jUdCC5zeAXsQIBvG/wugN4/uRdSAwiFkP2FFWU2In4IO1SedaRF
1upaAH7UOoP2q0h0ciZuVZHDkkuYSgJWjDvEDu7Y6jydxap9QH/CO8F5SjIW5Zl7
GDtLdKHz8+jwiwPhVM+xfw0nmD8UarCrhgtsb4hanKCKnwY36Dxh6pB7YDv1HEC1
Cr2DO3jSFCjEG9S3cphthidB0/M5mXAQKHcvOpw7LYw+7juFaAo0W7KN7AhxNUvW
q2MWIy3te/8NJDKLPiMBra8x2dhgeToT/fH/VFfZ59tSg7krfvfIhPpAQs3jbHT6
lu2pKXJ8tNhULBK4IKh6g0X6quWHKCZSTNoDnQlp51rdMKUMDPo9PaL8ATjIkr4S
rwc+wJvG1yoaw6zz+NRGzwqi8EjqYfbA6zesZ1XrCsOhdP0Y9FGGVE+29ixin5Ff
Q4jaiV6L9dJRSF98Xx1hc+5ohlXLVKnrLB4Tx/TV7yOHN8tpkSGCMk5WQqi/GnY4
kO/YjucGhPyeOjYKEDWMa1RMyZCv65bdA+z7/4yN4haaOl1y7MjmmuI+/gXDR4To
HaQKiKBHM73H97lPmbt3TnUR7VkSO/TrB+dQD+WisTTxAG1o8W7SM6xX7z6T1K+d
uEESrWoQzxQonZLt/YUeLSLRSu1omEYw16m1e/wJFFNiXwi04MwzuzrEcN1My0nv
HmuDJQvTXXFFgYHQu8YKcH+Oz8k7PYaGamQOECUAPh9jlAaWtHR0rvHfXt2hVUK/
yAZJzgxYmg5VBtqab5dReBDeLf2vGdrP8gLUe8sYJlwiX9qfVlssDlVugHTV9N46
FvHdmuglzhXocxJzl7W4wZowkI2f4Jcb3/HEi6d6PpW6fGjsAYo3XMxnBgWQXmt3
2MU1kHe32fJqj4eQC+g0lPKe3oXP/NNhrBNf0EBL+XH7+YvnfHUTG9LpKaD8AplD
B8UIM8wJhjy3xw/i57jbcZ7hXGzJVfnXqCjnXJGeZ+t84MZ5VIbu3FBXROlpMJbR
TixqNhxxy8qGkL9+ra7yqwCrQayNWVDHLe+/t+F2BTydBxGRlH0nE8iRi7zqpgUH
Ex3XHxR423MDPm32etXPhOy548SS3EgILSSIbQYS7fas7we+Z4eLylJAyHUW3ldr
cAAqXZjkJcvbUTXTC02sF4Dhxoz6C6Mi/OJRaiAjReNQE3eX4aNrFdXrnAaX0xN/
OsqTyDQfG9xl3mKOoVoAQH3vdZJ9Z9kDhKAsjIVMWnWFZ+Rv4sBHBknv40IQTe14
xXnlXlkG69PgessEjky9TEVeOzF/ALmiTABwx9Z8i0Oqnu6+9+60Z2AeN1BPv/ry
y1ENBjFuy0pKBq7IGkdJHwVZH4HDrMhavZHDj6EJc6/68AWhi099mN60JvoD9DRb
x7VkeyMDX9Y1C96MhereLdXR38sBtCps5/Ot6O7kPUCgXDBvAySwC+ZhBRdRaeEP
A+SVQKGIOZmzXDmeGibR3fDqAZ2oP7QY7HOZcrq0oumlYZh0bAAqdd/r82iP8O4A
9M5K+FXkm5fCQd8+ZmfaXebt90CkDynooskhLY+J41NnMAsI/qACjguTdoAg0/ni
2W4gzXRG8QLPCzxB3Ejjuma4uQXuWfTLilrqhGKBP/j8WUVXnduQwnIMBcr1WYV1
SRbqEw73pUrY9vL960tAsu4Ujd61GvVyEJNHSg6yiLugnRCftlM7Do/BVRKCkTfv
20I5QBDRT5hnBZZU+qPRRUZdSNlFUeTBhk6p+mLTkIveDa7s/LaGSrq15O5KRWoV
dGIL8m4H4OKReWCU6NTFtj8ZHtnV+O2aagY9OLYqoz6xuXba91vR3th3Fht0GqLK
kIQdFdIdK8/QgLlD9uI5vrLJ1+dPJeCLj4JOy/X3FHGq2W5leLIeQxKn0/NH4p1R
idHbom0juup1t664/9q+WJh/E0pU/eTOkW3gjTYqIwhfxU0SUqqKdCyqsP9byg4D
wmF6Ifh/orZKis+n0LWcweGqlUQIjlb5ZfIoH4fG2M+SgGMPxDJ1l10GtGe/SaMJ
FtYAdKP5wcrlTCwiKeLQs6jeBCYkNM7cVuCirZuXrl8uNd7ZsqbSIdPWB6GUMKPl
h5YH7CRIbXlOG4KMX+k7aMkpv4GTEbkT3NXNFJOexfWgYNUqI93RJI9fWL9c9sV9
PvuKUtnVzZk4/+cXkKereHx7FvX6d3KEnsKMf2ac13+QeJHoBQ2rg/L+L4UYYjfI
RT2MKcPe7G5jmDuOi8BH6H9W/3ZNRvnAhaJeWA3l4TQDlJagM0oDkPyFsAf7TfO4
66+HZ6nzm/e2F/vyzz10n8vj5b5bwuRplOG1IHJAQqexSqDN4JiwwMVVSMHZHAO1
rsufv38rqPfTHs021JfBUgGEinqETfAhfLIxS0iXDGPMwTrFpkSxcYaHa0hDErrJ
PJzenhfccDv6qfpn910gVMG3G4FylEdrMXqHKhLQY1xSH66VObm3uRHig37JH72e
dKEZ53H3UBTTZrhSi3A6L26KYfJ/167LMqZLDI5ZTMORT57y5Ua5Tl6vQpi3z7P9
/jLKwLJHfvDQWvz8VeQoPSYfDLNQVsns3eM6TW/NubwQyWUOoJXNxgJtml3juMNd
0QJtf1OkqZlxv8ax9gW5QoHgIRaZdC6XuTlnf6yEM/Dnp2+evEou2aSg/EPlIyhc
4Zz6bLhFeU6FRiOOKJymNCbnnScoAygc/3D4AP6iOBgT/jK4mwjAkz6Q5t66imzy
AEx/KYv4+DCUbwGmRyY+EeSU00+d77VzsLhps3WFXW3ubDJ0uYpd/zVKvwHoE0Tx
PLjq9m7YbIW1i3aGBuNtm8YTSgavPuPWCamj6oN5LmoGIqLBj4TKwHx/X26sZLFq
X1Uadi7nxxGGGy1ICVbToXdumdhf2HErbajhWoce0y4B+EMfv6Vi1vNq6s43W9aP
L8/WmazcHRyDsI/2cuuqGavrdCKosmrdmiEIEctdCV6YTCVgWSlNgzFMerw0xgDT
HFuyakhkqTLK5zWvpz/ROoiksXm6liHH+Hf5tyR/z+MMDpyhPoIaz93RRHyNUqef
DBbfyU+2hGkCtz/AGac9b5dbu3NzQDl+WVGpgQz3K3iWvRGegIXcmIwbXQksHJ8m
RbeizMvFe7mc0+0imVmi8ntK3qX0uDlJ6QtgutJpo1WoAhPJhtEboU8fM44HeLPl
bGjVHki0FG20RcdGqZLxKccgMKsnKJEdmFHH4x3G+ZQCeYhLPyjnn82nwfAOAWQ/
DrYSLxBu640UCrN0uHKQoCfO2+nCgNxEjAX0ahiYa99pDOZ14vr6lae3mZ/koosD
xz3rB4F2+tITQpSytJ8hyO0tb5S++alwL512ySNAHi85inlkFSVsrBGBO62/iUBL
T+W4KBuUgvrTIVV6+ZqfPnUdIHuhcls5auWJJxEhgedBsZxweHhuYHglMLvLwWfC
+4QJwyGlaSaW6aGAqhqK/vgjoihTRBX6d26/0oy5iNYHlvxaQg/SwtLdrMDRpOJH
EmwfVDokfMYwYwp4wL4LEX+8q9qA2d1PXEAJvu71QnZSsw933iOzdypH9RlF//Mu
71aD1Wi+3qruJ4QGVmF7TlifUhuEih6eD0MNj02Khjzez+HIX5TdBlnNzOmRK/ny
VQdvqKt6JDzqh3V61OCNoUAxpOagJFZlf+aHKYx3XAkCX7HaKfcp0Xe4E0pZd0c9
XRpX3V4AWR4SHNfL3V6SNCNeAkhIY/qw1reZf6++mgIRoe6NKejdhbAiZ5WyxkgJ
McwOrQ9J1wQHH8a8cLmQghYdkkKaoThb0RVjUO3us8rdCkOgS9pkzsg7bMexUJ5W
/PwwxTi4169cRePMQcifCmMxLmzjnYiYQ+25HdHMDL3Z80/kDnVWYUYidH4CWo7X
zrphoUSLQ+LOf6DdT2v7W1r972SWVYR5TdLbzqWFjGSahxoR1lXJDx6AFvdsYPl8
qEP+G/d4I4pI7E5OFW/kAvGDcCDLTGgWopnTleT1i/xm8Z8aaXtsNkQog3YFF+cw
VP1qEYRq7uReIbhevHb/+V5Wpe3WFJWTkn7agZmfp1/iB0oBNwa409ape4ptvysY
vLqIEEEmd2ISV7oz0qv+Bavjp8PQLBIJD9sDIqBv8PlWNXuu8QvAS0sOnRj0QJEt
4MDUENmeQaMFN9kPsjhikCRAHvgy6i8rH/Yv0WkWDDmXD5GBW3eAoT/oziJm77Z3
2vAggJmsFIi5C0zAUBqsmk7SCOMVeqcmb9dY5+1NqQV0y+TJ5MPn8fAxIpTSiDiJ
Sil/juFRj1Bja1PRCx8ZzbNFTGCpU5dTHYlriypch+PjGxHDzlGzj/BKTUO03IA5
QqEYsp5lsDeA8V1A1Jmxg98hng/Z50hISnjKv61K8bkilM7Dx9zQhe7j76EjNUca
HRf8UjI4fnuhfmOaZBo0FlF64M6FvqcfZcWvwKSBNxbnO05jH8eF+9JtCiMP3C+S
sD6ay39nEXfQFBq23VaGqNw6lgcrn7bOQbqH1Cyr1iwsmR7UlLhaLAcuhYaavm2Z
vLqJM057CmORbsN2Z5Ucw7u5fCwycw2QIX5q9jhR1Hh9h9xdND+ZmHQPoQiYJeaJ
xRqlUX0bkaKSJsKS0b2kzsxLcJTag0YnHjs2gAa9Su2Xm0ixsEELSb9zMpavvTe8
whWf3a/fS1KphIFCinTYPD8TSP1+mQtMfzx8pBGmlILjcDmeBQJQ4d6eLdvgW/3L
NlCLutMl/VxmUCD9hwVIW0n6pJSf7a6YomE6QlhcLlcCnb66lPczONtatW7+22Hb
afYKBgxSYDaI9q9UwUdXx1UwWyaoIO9vWIMqyOVG9NOdJ7M/c3Lq0xO+wxe+H46V
id8Zgb1NA4OhvBqIe3gODQcHVT+ZtxSBmM62K5xnlNT3CfvxezWxkaS4hyxgI8B8
NpZ/470QEsJS+sox5zrw8o+lU4vOS+CksAxv2ujkReCempGD9uJBuiMoLAbleKqJ
TObbJXKMvtPSF1XUAKiUzcoPi70iwdE+RMEltr3zPotHuLR/r/oVuPzA4sR+7le2
RlUY6NxczF4renc9afRIAXK9SO2ZoEzxgbvbQ7wqQgLz92dRm4peX+LaNLD9zJWZ
1iFsszmCxwys+uoqqZZJXd1SPCe1xXxfz2ZdjAxLM2t8KGq+6J2MtRZ1m/hxdz7s
9jz6ayjG8vxVptopUdQSLo6L08MbFBXGOm4nf75jnLmhod8haErDSxDL0l39HWVo
0r7xJYrUCJoUmGtjnP0P/dMbXcJwLBHrZ2du7xWHY34H7OsiA0J2KljF8lX3ei2q
JlUNrEfQGd2e25kBqhYO8qmKJEDV+sxYi4lbnJdg5+MYU68YnAVwJ0SERM0GKCaI
KyxNuRbILek+IyEr66gOFnvHoer6Mjc/Au3iJ3jru56aaD6NrkHrsgRspltisINN
LXLcRdmALaSkHM7cwSTxqQ4x4ushgD6j8TH3dXIrpdHmpY40y+LoTT49E94u8ou9
a7OI/QQmw+ZwLhTA24LxYNCR/pz+lljI1FOVPTD34sgJ/riaW1KJ+4tfBOlmJPLE
rnZkFP/81UhjU2vMEQi5EDuI8gqgJS7wn+shEUvetZ8wyesivm6WZnFgomMzb/M+
vY+GsUsH6ob3bHujFpuvvjh08EFZt/OuH3PJ8RpGPkgAm3Ousyu9Gt24n3O4NGUU
ZZST7m1pgTmn7MTSA3RVJS0b54kP/0fMuf9efRzjaix7Wzth4GUR466eyGtpEAqB
ZTbQqynSzwXhz96T3Qf1dpJlX9pGCxmKflwlmMVGWMVDeL4thICJj1ceK+26YrlF
03StskALBJE5m2ORP3OHgA8C1tEsNfwQXB+Qiwyl9KkpZu47hTn2uB1oz6ciwxeI
XrRRyG8MFMPZnBPg8AM8v58byzx8HY7s/JAqTXats6o2SjN+YltmJiavM0H32L3b
cL11fZ14YJ9D0kSZLglOTwInXFsdB3pb5n3UiGRoj/i9gAkWCZVj6rkgH0QdsmKP
m+fmgLXtF9O0DsdY3NaEvIm4O+XRvCWQnTyYM5Fp4WzpvIm1XF7kwRyHDl0nuZqj
6zXQJgbqAox4tKv4NJT3Ww5SMJw0sT0GEirK0H1W08QJfZ25n7fHewG7DY4TFgph
cKS/1s2f47LYgqq9Ennc/YfEelSrlfIFNuYWO8oc/F4USnwC2fK7uoe/HAJrjGh+
3wTnxEDfkZeWeja9Zwzh2o9J1EiQnZMJzIs8MZsbED4I5wYn+rbXEydjuo9jYCvX
s5mwxFGq6rYch0NGIQbYOcAVWnhu/SPLjGhY23sPzlHv1cAdypgJcRxlmcj+rGzU
o8H65F1+Tj08d5GTyeEQPeodqBMO8qxipQWttS/be2HYywrDAi3xXvSgP3YUEfwP
xdtMHSYCg1dx1emiKYiSlyeweZIgn1BEu54UxJLkFsrRVidxjSXwbjq4Nc/mQP/d
6w7et8+1zrOpwtT9aSkdM3D6HPMajVsgssUb+qvDKcpjwFPKqKl3a7YGn4WXxSOR
ON9AmXqpuKyplN/eQdD3Vi3+379jWiQVyOFysnKR1MiGNHng+6qNBXcv3FPNHVMX
XScrbEAls8e5vFZE04Kb+MAeXDc+GznZxGkzrg103DNGWrMaPao491AhVZ2iRLps
e27B6BZ+pVxKtuZUj+hi2Ei03f/FodMJ0POVzzFPscxz/A+TAHyIN2kM6Xkhgldb
kDfktfP/WqbcI8KvODuITY1X/gPsu/T5L56163OhWEJHZKHm02tCjE4+AeQ0e6Ux
A/h3VxV9bRgHwTcdTjQyASmF5okFrcIgrEduurdiZudpln3+zHu8zynZ113gwBsP
Bg/eMUTYsh8pj/CUF0kgjp+5yxyQ9XED9O2DkjlbqRDKAsds4hXBM1I7dLwbr85o
IeMTU1QWGGjEsj7sQqfz2MnJrNy5q5XlnbU0h6MDemYd5sYspJUs7bKATF4YGZk3
SRb0o5U4Cx5IoejzFcVEjbzoDvg+4SwB0ZhvZKl0pOqqyK7lss9Xe35wSrEYCGFV
jEZ1SYDlrVJzGdjKgJBxqQeR2tKWUFCfwomZ4WvqMoBAaFa/oSH/1exboOApp2u7
duO0D/vffjMqZ7xhSbJxPVnXmFVefQox1A4IhcGkBGmIacdarhCwgg9cNRUU4bjB
nPIAWj6LwSX98ZEVUm5SkvQCGgbTfu9XUyTv3gbm4OkyOut/1Ye59bJdRg64DdyZ
mSQKMk/9fJRKsxDrMM1cp/OEkItNt4joj5Sc1alr39j/FMslqnxY09zhP8d1gTEv
hwB5/d8Bt+B3z636ZDS5hWaj93ClkRmDXxP2uNMHUNVM+yAm3iNbtkIxHjCToygX
jxzJUoXNHwadwyWxy9E5Imoem/VcnkgaIV3zMzeEGG3SIm+VxVSDwBOMl8skKenW
SIdZQ1/e+oQ0eWDrP9Vt/hkU6RpJKKfd4D4r/uGELGo0TiH/lIo7mQFwjzWJ75F1
H6m62TOWmjWMKQjAPBmsVRsKe/0z+odKZzyGkArbkTFuVbaQnJM4bmJmkYuoY0UR
mkuJHrfDjstPRSAlRxJRYNBmhINdeu3lfvPmSbGsSsvhvcZYP+9qJhoYeMNk47ia
tIdIl3Uxm+I3KJEX43D4xuFdh/WPYf1uNNVy31VrC+UbUvdscAH+drhqcK7eR9Q9
f6Ai3BhpAMk5Uvf+rdwGh04fgxCr+ROrIN77entQxRcuI3G05dwtuTGfzN7QZd+x
wymTB14TBPpJAQfP//6QURhvu5Ph3RXYPRCKfHPkKW4fXqDQys5bp/ELhYZKNbfY
gkVKb/9RnmOil0BJMErrEFekhZ6TiXO1Qj5iLi1w+7rI2ajL3qRXpneTqoux15DD
QI4cN/0J+/ussSktcMB2Wk1UD7gRD4TmfVtCvnQXGWrpin+emucN4WnK0v4Jm3d+
IUKF/8R27tQDdy3zjuYDVZa+xcIQ1yQR9dZ66UaXckk3jv+9Gifprgmujj4wC+Cf
RmlW4b2G4nE7z0uypuw7XZ1BxidvjNnY/TRt6MM7T2nSvMc0gRC64zP80p4nUcwL
F8hJHgxOgluhevumtqpraIM3Ws9SSR3m0ogD+uYLs/X+7NzuvdDMAWISV7yEh3G3
bb+XvR2YimigdB9rVrseuC9O90EktXBhd+o9649E5agyia+raz5V1RButuSAEwrD
GnWO6VVcKqH9GINH1S9yICKEeOXboVSHvBnl3Gmq00MuGo+4xMoAGisV/D7cnKAv
1TY1PvdD9rG1mM/FaOoNawx6eqjk9wDCG/nJm9Z04gcixfB6q8/hO5klSWisNF1z
s3a/ZgyuldKaYN6Yas4bdvzmLpGvcnaJoNeYpEMdCHXrIZGR3nuEYqNthT3TcKdN
jIHF8IQ7H64yn2JPWqP0So5vcSbNFhT/kjYujS6XB847W/lArobcHnU8aZ8TQOFJ
hxdUhAFBIHQwSdslYDS3zzAy3i8cO7WWeCDFsjVjpRoi9NzungwCTWTd+0YYfV4E
w3TacuvmpDdTpYvMcMOILv3RXQTGL7e4M5cgEfNt/qv4ZtdIfxO3nPIPQ/I/ND3j
7GieQvoM4HgU4KM69BoZKOwJF8LQRfQF16tmWJi6GE9pZG1ehR27OPvVVA9EPkYN
GzxDq5iih5ruUSR/ZNYKWj16TF4m8TdhwQMmR5HmhFwDUQIa+/i08CKC1LuK827a
0ndwQLYT4IQGfuoA1yCfJrWNYSvy7PrMGudHqOoAsYSpUezcp5CX7OBwWjywL2Mp
5y/KE4PnneIgBfGFvg7jaYEssD29iwW5MD5eV+lo+Sl6KoFrycwwKQ1ihNkBerXh
a81eHpOANmvfI4zhc0uPy3SN6I5LDP5lZw2FhxJQCX89apKww1bNDqwnuZeMk4V8
DQQsncTrPA5vytVbPGUysowdrXZwrhcGE68AgW3W/yMGSfY1/4Ec6BxAQr9eFxNk
wBgR7HHWMEzhDN6YGXEv5cloHxDOwwjZ51GwkoJiGGKww6SIC2XWUS68ZU68XsWZ
Yp1pcM3YwOf7DygCfZoOmS0MDGvJRhCQYC+GcKTOPEEHeGZWcghJHGie51cc6SVD
iAnywVcTfqYvPPdgheiffEH367pon5AFPcoiW0wkxDu8rSmEGf9mQSSQ8NIivxl5
l49JIprKE3giftq5IQxlRTo+X7AVC9UtOj98+ENP0PYC1GWPKVhkVaziNJvisWnZ
936OdUSIBRq+cVvopYT31AzBCU75IvTqtR0yVaOuJmBHxj/zI5JMpYYlnP2A8SfQ
l9huuVXggARjWVbaX2EEOH0k/82iFue7E8O/bAdMiUJYybeNWvEqnN19e5VCSiJQ
/6OR/aX/OaPXxPJTadFdbBAw4od84Q6KW4a6J+biDbHeR2RTsiCPnFkBPTRTNhnh
/VG8TIQPMXxDoQIHSKVn27ANuyw//y373EQTA7pDY7T8//UumeYPc0KpV5cYRouB
q6T1muSRxktbpl8471Bnj5Jkuan0kviFy6c45ZXxb1mB0vYLP+598YFg7KPhn86r
wpmf3bmP6gddxEAB4ZuW43k0PXHMSfF98TWa3J+pkX32PEuKyzb5kggbr5ntOri+
cGOzvSpMP9m4EYaRDYopk00FunD6BHFsOyu//AOoISC345UzO28Jkyyr6JxkhbnN
FxAr0SC3OtvAaDDqlKNRTbBQKpCKYRm2mxNdSodLBvhwURJ+keXNFzv+PTW8CRWd
8Ov3h9EpaVduCIVg/I1FNJdSeVECLXU/22xZz1LWEJsv4/THg8nMVg3cnIXMPf9x
VvF7eq/OGhhUemD26BFbMMEEIBB9pcnqKaSl0MHvlPtLjkHYbycQ3ppYkl6CdpEI
nyaa8L8XTDKQS2kLIN9qRlSIEK/siOyFt4Fvllyyq3vf4Z68TYaKJgy2PQq7BnTf
oZOtcuPLTjqJxnNsgtkzAo0Fm4/pKaBJTD+Nw8HwJtaWvec3ao+WUEVRDnkAjxVa
Ny7Td2L9K6kppDNRhsOZXe4wWpbkbHWgTJfoVXxCsFTLsdDT4cdnIcsp6SRTSCY6
SyYktSvvr8TFWkRWsueVwbKvT7/cTCaBlTelgLJEQE38IJLSzFTtiiBpyBumyjah
VblB63Fx7w8SG/n4XRBPUhGg3mhSqqAJACHsFdxGWbOhePknPmyxD/tDT3Xddo7K
iHP1gh5piTTy4wzyLui+NvkqPpWbUD1xvIrc6KWI+WL+zVNBh5XgurdhOMNbWlBG
vW8BK8ieKzQwHhRCnNggb2GO1RqhvF9KN3bfWQQbkK0IqTb6EIcrSzhGQMWY1wf8
1Tesc9lGizFd8k5rTdyAcJTrMQThpGDb/+bMsJ5gLGDMzSOdR3kuVLjtVD/lC3wi
uf+CviDHW7MqtMmqcHiPLtVndwDr2IiaUfr+5PPeu1P03htsXE8gWExUzEln70fB
hSa9gopb/3mhz1GPWTBSycW4ZJFttqKC+w1d8HLUCS22/KabwI0WajMq35wdG0W1
q7/Tgg14C1a0uQKJ74z6rGNyM6GBdQySKK0BGcjX5sDqnQI2dulBpAXquw3SMu6N
Wobhg8MBKfvj8eA3tbGxC1ki8OcVfIBx13Nz9igz5TB6mJt9FXCzgFV29X5yvlsf
oSX3hXozTlfK0+6fFrbNvazZWBWRRP//m1DzksSBDdWmkfQ0ypkWrMSYHfUo48Jx
s1xWlreOOWrXPm2g3BvaxL/CzxyrwKfN/OOePm2nXXMTjm4QEyI4scWcPRAt30X+
`pragma protect end_protected
