// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
LFYtvJOL5EihDquwpCd3GY3v29pc4FRuDsFV2Ddtp3rfpWRM19dxNLnSHXXwruMao0e533oze8jE
iM8LwZzlnepU9nITYM8AbWaljzWLkBRaiJxqMru3K9Ro+Tdfj0xMLXfqPCPRxHS8GUogDz9trHmj
OSR0mcfEl2RLYj6boy/lSMVGWW9Mrbla97o6BKB+p2Eew8NQCyVuX1WzRh40AfhCJZm0DjAY6vFy
8qpFWcN2GoGdM18D9l8bcHz6zp8uP6CXOFGsvcTlUAc3h21QZ6xL/TTRy0eRKEmBqJSYGyaZBVof
vdk1n2lfsD0WD3BxKFmkzDACzzO7vKAcmmzkVg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14608)
Kvd5SCU82ox93Z9il7sldIQR/8ayGJRtXTQh/7/p6xb+pMJ15wGKscOpOm7KQJgf+4mVIkyN0mSh
gcuQv4IUS+eG3gHaZeoJ9uUKncu28pAiL/OTvh/eNQF4dxZO/Nf88bdDNWPmXq/wrr4IfgRXUCm6
a2cU3hs/o9CyWdoFnt6Lsrdu9cZozeHWhP+9EJnUDcuLgzabIrirEr7GHyx6n0/7j/SrloI/ki+W
6H0inpODvbJeeBKyP/ySAWuwNd8v6vKgW8pezEiMPa7yoRBk04fcD7Wf2rV1t2fLMFUSN3jLe67w
smHD5u1SumCrtvSQzXDpecqg6bET9Zut71acQpWTX5Q6/k5WWhBWmAy4z1nydEHOdxg9eh8GUIxL
PzBARimNa2e3DfBacbn+t83Rw2vo5W6lWeSeWTgKgP/rbgoRil9z0F0ry6ze6siF5UNpRyT4OB/i
o92bHJQOACwH1xMK2C6UN1c5UPLSy0Ublnwk56OdN/QV5sviHEwRMRtq8H21QN3xI7n7hAm0JQMa
XxPqdNDKIWRueFostCuiq+ftw8y0aFu53Vty2a9Yu+BnsbdrhWUw5wjvyhO4jZ4K7BYg7RITLIC8
6dc7xtmUtuX3ZKbya8NicTJ2JxdPfPzequKxrZJQKEu5/YlZnx3YM5A6M95W/vcv3vOpf0+Ja6Oy
JeyTL1zjaAUXXbxndCw2WLZgC7ry+ECe05E1tt2YmV2qX5GBHV9IdtDaMDe1Jc+3eYmQknECjT7E
TkbGbeX8D/MeqFmiFGeZhXzW27yBewTIWP2YlpHlhYzoP/xDJTfWvmjhbqmeAhhM7VP7+VWxQ+pp
NFUl9Rb21sHR0+Tfqf58rMSGtObVfESJ838gEupP4Mfp03gN2GKCFbiIMZKiSLXpN6B6rE3saiM3
5lF9mIxLWchqybKA90YpkeQOOSu1ypFjMvdiUS/69JJQFai4V7F7whizDCwLLwb+DSyVmzTficN/
aWa2HlwZRhhTYgjOu90c5S5wzUh7SSlqwDUqWL06M98x3F6mA1qE3NpDsWTNoUTBWtm584f2lJsn
s9PzkfSMX0G8WdOYx6o+vZC9i6BuMvxBep8fMAady+BomoQEJPcxAsHYuji6wAa6hr19tye82wYK
Kr0WNTmjjwD1i7GhuzdaeC2vWBkdvk4DlpVFaDM1Z20YL7dvWrd1c+lsNw3JWpWx2pCbpqGyOUgA
DrG3QHUyse7GCcOtfzSCN/MPjNw79uJPisJGcZ7hAWaHVW15iFJj11jL7+8vjD5cbnzM3R6A8FVe
1No7QuJzHVYTyL1XS6vinXPmGk1vAmc/qBvZUOHg9tcXNL+c+OKdOlA02D0bTuBPvJTvwRQ9n2rU
rV9FYO5a+8eX8jMeGSnjgCR8O6U0do/v0+3g/kC2icGpxHn+KO7delk5VoqCMkAnBsD/E+V6e4iA
MvvP6DNf4/WCgOTKAZkWJ2ZwgH7xCdQWN15jtfm/alNkQrgRQ5E/F5GAncmd2QoK7IvqtStbxKl7
FP5qY/yQnRd5Lsyo+zFVuAShNos7xtFV/IRLOXTqv0CD6QbasVb6doeF171DKjTy+vyybSlBOVdY
lkNcNzdVKsJincO5YdYo4lDbeGo58bh6vPKFmBu40xWDaIx3ZINbJa7ZOVYuRXKRjbanOyK56xBJ
k+zrnsdI1Uoqg2BQF2zpmlruGBkKX7iNCbMhT5IN6yKzrgODt+HoZOa0+dbz0jMHOZ10Ea7nh44+
Mg5NC8xAOt6U6uGY2t/cjoAc9HkvBudZkEhyE3rYPCNSfDY2rAft3OKbCIElOLeI4wtuKQXs0Ohb
LmQ/ZFNmuaH3tpDxLO3z8FQJRSTI5A/dLYJNY1GSrwei+YTAjAnKUT4SEDNHBlVjiXUk1XYVRi6J
ThS8tFtwAuTtU9ZFRjETiPHI9iW1wcowA8i4p421hDxQ01aiFYsJ7YROlj0Ay7nSwg88Qcs/Uo49
Mj0JSzh3TsK60Ye5Z9PjUy7Y9oBPquQky4p5D2h9GkgWiF7ONjiy2k74Pg/500/nTKDVexWtQvdo
hmhPyqtz3rsXAw8DYwPzzjtXDptSarKGi3t6k4+ZDemGXhwx9JnJhR2Xg55/IOYmDxCA52GUgDic
Ei1gc9hxFOpf3wpz4/ERd6iOxsvhFW9OaTPGnvxhBkc9T8H1FId1c5z/Ej/WQuNpGjFmaYlG2mQz
ZvWj+cQ2HRrVHWNtCSkyY1eLZwQVSwSvBaXy2KOoIsIhsjRUTTPJSWOCgKb+/Ue6nO2vT44ezACh
Y7/NI82O9jrEhhSHMS508Y/X1H0d8vbZKq5o7yhXmR+xOmzNvE3/DosxUB9TaPVGzIgRhe+MNGw9
S9JTFuukSNPM1qujjBYkB3R/k6clr0atKPszEVWJHKZz4GDPKluORoCrR329yJn9MJeXfoJ4+n/k
zAodfth+he0gL9n8ZrL/yEH+qsDpH8b4cQ1gcNbxf2LW5UZk5ZaoqRxz57qFx0Q1WE74OUc53BnO
KMY7F/Bj/vazdto3Pyt6omSQ2g6Mpi0XFPAT3upqkc7Tnx8TdazdO6kq8YDn9XFw9L/YZtFKRRiZ
KsepC0vPDGkQlzErfKMaFhjfYwnIQbiMY1hK1QQH167ZOP/Wc4RsMIUq+0fgIaFPzjQkh3Rqbpya
m9VKHKY8bJ+YCVxOA1RtmOFyKBDTCF2O7UAohP+F0qtvjXMjiMys47BSMnKg9icED1zuk9mbN+Gc
OTj8FthpSNiVgtUujBYFuGr+6fVpz0hLQCfs0pUhfEBmnpeDfa+msa/nKq3lfoHYw6VljaQo04LI
dCtIzvBxHIYjiu/eQ4aM0Uhgwcxu1QkTCNd0JhdtEJFrQOuWZOIZQesnXbrYbUAjs01myRKNdQN4
nSZJLKH1sZ7RQ6Yw28ItA3HMojYvTVB9r8U/S5hdnUOo46fxMfWbxEF9HmSAQfl7y7V3mgSI6DO8
ROvkWVDjXxnyOva0FnwLsZJRyqRfr5z1UgjQgLGV9G0t6VrnNPSojsg9dxSTAJ/6sTOZFJGzQBHR
169lQ4HE8mk2ozMkx9aPG+IFj8HMlHLQXQroPQspUK+dRCVmyNeedZGPL8SQap9leFNxb9JQW25m
BW5ppR2qn0gBSpTnb6Da/L9HfSAPPbCRlAxbU6p94k0j1Pxk31eb59aT8nOLK8FutNButMytKFKo
f8+Q+8dFpFGSETqlc9I+XntYmbdHinYaLEBfPGWr/0iL88Ct1NkmjKlU+QlCC62NIhVUSSfB6mAb
yOMTULpj++m0p1YHlD1aqPShAWepXtsjhTGSEEziBYaPHQh6NhOwLJFwHt2PjhNRkDcOTVAA4sSD
7N5s8wqFf6+u6P1jHs7Avun1+H0sWigj96sJR0TfcXADxD99odq9dFpnpCOVHC1YgGTelXV63Pyy
C6amFV9tIpDcJEqj3pfnpkNXITRG1NYqXl28vY8CDzMZ9Ar7R4iWqvXcjxR5dGZETLaFTaVBE2ti
roCgi33aN2RJoNwhveYkfSnda7hDUzaKI1xk2i9gGOgZCXB0Ma9rBNzgj9wEq5n8hbhA9Du2DEcP
ZNMWjTq3R6zPxSGkQ0OCJv9whHEg2TjE2dU2i0f5nCgjXPBJGQdmx7QwmeDU7soFBrK8Bs9GGr7k
UBslofUg7ihtgpQO+YLQqvX5RGU4ofbMX4hdHefXOO+2hCNi00CnP2Hyr15NI5M4W8VXLybkSHYY
ER3ze7l1iJFtsWQxk8yBHyRAgY4LyL0fio0h7sffXHh3K3tDShequGQh5rAWeYfiYFjBagS/h0HG
6SjbdTfUF6WcCIe6a9i0kKVH3kXriByFLA89HzCQorybJr2wOHfjNoMQy8PnChBADhbWhLpGlm5x
UpvOcvjPn3pbp+rxmiAr4lBKbI1yrXo1Qt2EhL+acbxdBF73oYXwJEnFnNWMQbVtCE39FzQIPZi5
Bb5w0gM1uVuhpPmmHlVemLUdRokrpC436t3SQ95KJUPL+BxiNTLimLOYTEJzgtJmewVTjpcXXp+M
UsyRefwv9U+nzjYyXytXat9XViXwBsTbzChB2nVLrC9op3hwu0pLu0FN3NQu6L4BazU/pvNiYCFW
1pdqZxxCvDyqHotu5xkECgIEDtdWJtrNCfqUJePmRSMI3AGgdxpLG2XkPyt9Emk4d6Mt638LgNW2
ul6DUf/gZaCW+LggzrDXPF9WtlpJBjR64pviiZ3gM8u4L4/8LDzzQ2oSbyppjX7rnVTuM+x5b7Du
EGOiL4vtJ7Z24foaK0xD/Felm86DbBDLv8LffFnI1Qo47/bJTWwauMWMYqw2HoCvNhCif38A96Ga
qxItkmH9wDAroQQCY5A/49v85sDM6r0vTL9VbN2ZQx7AFSmjwKr43/tbFRxr9P38rZWK20lwbpAS
JXiAoDs6fug8ao/YAKnij3xLpgZKfoSm/Zqo6I/+P6Nk6F5qjdti7BORwMtyw5GQrEePkro5qehJ
vSjd5Wjf0hZRDc87h78/QXSV84z+XFuSmHjuOTz4brywpbs+5Ie4Pnjrv0YKwQxREOAlKQMwEbSj
LMiu5bTWlHoLdwJoYuzeapeOk+QyHny3bYLvWFlKc+6ot3MLSiXMKpPZ+NNogq+vFHUf0WJANP+j
IlfeqTv7UXMYN0iXO+3K5qVlG6k/+nDt3cQRwljm4+6bg2VNQyCcwIoY1m4AR3DNujTtk3LyJL0o
til9+kPyzhu4X+Oe1HFDRZoM6opOa2TvpSeFeY6lwpFezrTplXajcmyhDlsM9Y2mzRBZB1Ulgk0f
n0B1m/LjpM5DkuVgPg4PVjIp1G7b7Kf5gHil+ZGJ+PKrfFCvd2vW6qDO1iDyuFfAjipNIQVmbubx
POGaPw8tNNmKqKt1wJOhykEYabcw4vFbiLaQZf3/sRfgGCg8zxd9hJx2tlfvD1WPwUpUlKs3TjW1
IdTVQW5sx2d4IBfGkwThlT4VDJI/SWljJpdLKLry+5aZ+PVlMAsYnz1yv+fHDs0mdx79k9AXo1mv
QFNSrwTd8SIhfX6ltlA3rOEiYS9iHnpLuatc4E8oNqo6BYYSSL9/ZTRjApbjgEuG8hkAnd5fMYas
fO+G/jjfAvnrsKrV+KlhFJEYlxJha1ANmEaJVSZDdVCapyMpcfJiMrUyf3Mzu9Y1UMSOiJX/jIql
OmZV6WbqL9sixwJQleK0D6FAxDzdwMH6UojIHTJ2wamKTiBGdpFcZOxmaUzLOQs53qRuz1tEoLeE
yaoVCwO8JcuoWmKTvNkzR2bX9bD3bTDTXBhoqe7ZJ1p60nP2/E0CJ17zS96A8wGqyh7gSpAgCIIT
LkhpAw1LlUqzW13btte7HC0HpAM0qIt8GJWDG6TddOQhfZu0hLMgcZeRmfI51zthE2d6sL/EAJ8T
OpECZo37rK7iG+KIkW0juf3lDAy+wTtDzUr2k99Ztt287Xg1I4TQLUZaodwq+2K4t1xwr/tc8XyD
Wo+SGaMCUJZrm72DEO9VuodQuouXf9M2A4IBFdfYRIQC2V7us2Wj09K8CaA+FFT9IsOhcuZ6sX+E
LerCGiboFzwKMEIjDuagSzV1boVCLVwqd6DBBSXY9F4q8NZeTH+OAbVD9QshmptSUGKjLNBC0smX
SD3Wqcp3nbvZ7Mvi3aoUvlO7149BRqaGaIxI2V7/HbTGkaedllhdvmAYPwP4SqcYgFcaJ5ycsWn/
kvPTTj02wyWHS38EV8gpQd7e28ROD555CL0kVzmp5jYk18GqE672Ns2g2XLQI5oAipQzFFTberfi
JzsSEYi6YwIMqlQ84kMhLxOX6gt0QByHkw3OQvPtESWLjxNcliiPEIlRVJu9CE63DYs3VGCj32t1
1Hz2wGk8PB9QS2DvNketqlK63ogsAXi+q4DoqCHn3ihSEkwz+QfnmIJXFWDaxep1IzsTq3vBXrB7
Px9x4mmKCv1DInJXkzTavrFPox0OzMYLmdCM4yG7PGx66asVtf7t0CDf7sMSSU1nLow4p1aqZp0V
Q9fwzrdlSUnsIDQ+4ykXLUY1MQbqdhPz9VS/kVA2LLkZW4M8NCe+yO6xRYJiUf0kMlB2d5mZrVdg
wwOLzFltd9bH+0O4CbbiwV/zu2cOvfEvTnPLHnBhMWh93FvENNi0Uyg3iG+FzEEGGuDWu9hr447G
HxJy0F8ezONhb5OITmyr1nQeK1gnHdbWfCRXvDOQ9w2SvB+DaWLEvhzv5bHw8vdKEt1usxhrpOq1
1Cntc2wc+Bw0EYghwHN2m6RJV+5NWTigQlEitESIAbvPzi4rgOg/r+EVyoqQ0ivKcT+fweg+zwI0
d37rnR7sdPdoweEEsuPmmU5BiXwGGUjonxL+obMae7kYpKEycDhtuaSzhaaiWipwXWluP+/wsK9Z
x8Dxb6GD81XJyc4qtlLs/DAB6w/NSxzENS7eI+hkp0bcDoljNLGw5WCqiRBrYy7qZhlIqiOGIh+P
ByvMhn6+SZhpheKLX36HjSmA76XuTPo3VZu/mOtb6QFW7FUxb/Mo4K8chhOyCDG19asg6quDeH/0
yGs1IALM/U6wnK5Vs9+3W++1khdqVBAQoQU+otuI6d3bbptLtRET0+KcJP6v+YaDilZpL53vmCZK
JDN8Im4ajmz2R/0RHM+VOXZ8lojt/Kr61j846+uqbE4Br77/pkfnzX/pqk0aRwdd3tY0mS9z1c1c
GZUzy0ZTUBLXFJ47pu6WymgG62GHvYWkgYiIoxxZ3SYAA1pLZKoq0sKcXhE30MUnPaSNpLX03MgP
sHifBhXz9ilLaxYY5HwV/nzGAtGVXFN7YVmIGB+o41IQmwEHBqEK5D5OJ0NNyMDZTkAGgCLDfLXi
LfHmJIIAAkT02QjFPGh8MMz9Bf9i/XqNYLZjrZlitmRcWK4E95VNpjfGyl2+iWcgPhW5sPTyp+qg
XttcHA/HdtzDums/FNkxT9+mo/c7zObc2nGaFyCfYIvVy0Vmng3qHv+KNioLc9sw/CsTSYMpfQHl
LGT49AGWKL+cTzSdSISN3gZN5g/9DJFqQ/lmb48Tlgf+Etqm7mNSlbTgySqwXGHC9wYrWDyAu+wy
7+FUhQjQlZT8Jky5BS4snZDM7g6rsYlko48Tw9iWwAgwOk9+PYjNjQ0oE7VTfkfbxb3pjvSzXxT/
oGDby3vgQhXYZSky9s778CBUzkmL9+VwrQKveD8ycmjuvH782e49IYVqfWSgb1xXRBBgYnptQShR
KnD7umty4cFNVgNVPOMYFepPXhnkSVcIoP/Puvui5sDe8D4mQNtw3yvZJ2c4XdeBTiYmLzUr7gX/
0OrP9dCQRCr9daoczljlMDnF+7v27eYaCpdIvkYltZVAjofrw6qMh+/PpNIgT7bAf9dG3MlOvq6d
VjtXbo6TqY4Bl0Atc8rxs/G3bGkwAbc8ZKPJkrxyxhUv5WCt7g6WuAcIFJjtIxn//95dYnyRdRMM
Y4+IhXUsN2EgMAqMH9tn86k2nhl8W1eGYIER1jg1o49fAaE5tPI+T2sFH3krzlRVN+krrJhXQINj
cpr9Gn9cHND6Q7gU0aK/9aK5RdtQbaVG9NUoxec2/YhKq4WwuVjtlvqP0ZUcdF6uHmOA5Qf5oJYy
iPZ6UqIweO8ufD0ffgGu3dm3xwEWXisFENK1WDPiaNfXbbrDJmYxjXY7ykXbYi+Xbu0+VfXXqlpe
BeqpH6fOvOgzpW9KKvutjVxOkpqRC5hZH64mDOVlyqHXQPY2ly4n6KupScH1wNMPNDgASmPAmIa8
Gt0PhrXonKbQUGuLIYYM6OUrk3IE1j++X2lqFTJgja5LX1Z8ikhvB/0wHBQ9USSXG2SEGM81lGYj
rgmgCcaTHaPxvqLENFioUZExX05CNsTlyLOu+1WRmAmpmOFiF8xvl5q458lUuTTBNIHXxIW4vojR
kagLoIOSzcHETU2H0kLC+wHa2kTJnsb9WvM6uYlVFQldPfh0lRvcauZFPlgMdDODx3yB5ozOkUqp
XPpYPdmYKP7m/GKLY1grJmTegv4zPflHKsVXyQ8JVAES/w29TmuMzq8LGtJctddv905Wjuqh/wdB
zvnUdQfvcKWA3e6pgfDIJbcTp5MWz8eqKED4WSxZop4wSSQLWdGJq2AcfFVPtBxl7K/0RFZvbjrA
0wt59UzQzMfo+Hl2edRMJdFwSKuovpo2oM4ziXmZ3HJuNewS0GhB918NnyJH3AqH5gJJSiBk0Fh+
yDOAtHRygAStpv677orMPIHCZM1BIEFrzvH8I9SVrCCzojO+2wi1RleMXUEh1qEkup3cjoewzFot
WfFezZXsZ5ZYU3st4lv6rV6Q+6Jpm3c+2QHHOtlpZr1/xBez2kZVd46OSpZ5zGkoQ828bgEv3Ugj
XTIZa3OjuPORkP6hezFkZQpP6h9jjrriwLzloPNyRWXtQfUv4LE05pvLbKDwnKql2G8F0AJfkesV
s22gwbjeSMNRVTGI2MiHpNCAxBgC4PzpnB0/oVxAFUo/wKHk43xhu7mdoFWtMi80So9yAO6F/LGi
sM1dFOX5GuYhKl4wlzwdD7e5CNLI/oGcknsnNb+KfBW+mEB5sAxiIKWVN/16Rx1jjvJxHAkVZ4WU
EMv7hGhT7L5N3otveR12oqoZ6c6P37Ccuw8YWrm64HWkiJ6MXW8ItzaNfbZxqtTVGL3bKUDahYr7
WGi+iV/Al0gxlDknFAhH2hwvFQrZbpk4AIblFgBfQUf3LCZaTiVqgmtFrGb/rSRp9sm+8fTZMX34
e+U8oe3Cd3PYN7PjXoZfAyh+To/VWjElgm//w8yNT1N6oUCbYTTpOGfrC5c0jK0AJIwBf4wEbjyB
FDz7cexNrdcXyaMqhoWywarKa8vfG1nD6WeeGVzAc65+eoS4B2lk4cSqMEnAdcLFYtW/MstqWxTk
61CIykL+QX2mUcIyCyVs2ylvNCabEVGYlebyTgbOjzRZWeGgywzjAxIKUPo2+UCERQJ1nWATM0wH
x3vFhKjlKoxF2Po4Dvml7/Gu+Hmo1/T0gBFGqA68sQmK3DVIfbVrTAlMRE3MTgm6efVqAO4k7q0b
em4Sv6KFcTbZG53RJ4l4OYidS1TxCc3La36NlDG/H9ks8dH/zI2vDHSXsF+2FoEQFq/aXxfVuGCT
bdws0HebdXzQ3B9PTLP4TUbreRjy3KJyqqgLzskL0ZuaE2QyDnbW1gI/6peiZb4Tq2vGF/s51hDM
9ogVIfGzyJMHYQmLrO5PbE2SfrtGlx1NCvMk048WLTN4On1aGD8iORm0rdqpQZ815oG85GY4ISK6
Lw6mGi79Gr+zipnKT98+IcGMeT96e4jGCchb9zkzPMfxiDOUd5Dz9VK9tuKEILIDb4skDPhJ8whH
1m3DEjf87N5fDjhSCzdIbPoh2gft0GrZWpgLURt6cGkTwkQun5AfD3JhyCm6dziR5hZr1BJBDPwP
CctLohAH6/xjqA1213M3kIcek7QB8ZPtnmpOfOh9s6JksgzDqneGU3jM8Sa36HsDrk2RxJIHT8vU
PmepE27HSuCecPsmAQ2ewgv8/XBKW/0lwZr4iiKdjG7MSMGmkCh1BpN+WnTYrN9i0phCZeK6o6jU
4xKM4qv6dYov+OpKiEZ/eiEPJuBdkLG+KHeV01LsVtgm1MPBa757PmoZv6yX0z1us3jFfp1zSprK
XW2tN4Qhal8UyrAmyDO0O3x99JAxiWGs/hGM3EGpjqNIzySZQToa5UaW6Rz4sBcjS6oEcD0h92GG
PwtZXZA21nRMogM3xh8gpe+4BaGSOoXNjYFYCGiDNQ42LKuTAp++gBEeaWhbfKc3m/eF8aHcy9NL
oHacmVYAmQb/XXVFaMYHNnFIpnSB6Vz00f9y7V39RzQyO+RJglQauap8vOsdEbhHtDS8NmIcsTkD
cQkauQt7DcsyXXHTqthRmI7n1K3V9rF9eyKxXksULZcacPmGVFV0fkmsbadvpVFKO5j634dpoj3A
YnIXMiurRGiuGL/LY03ahdnxRTUPB1j1SzEZw6uc6P/nuXhuMaaw7zKH4SaMgqDYrje+KWQQuEAV
Y3mgwvfDXLkq4MFFE28J4oN8Gt3ljD9UmaZTFdA9WMT0Xvusji+2qkSW/XL02kfkriRT6JoiY2zR
cTXrNtlG1eP6zZaeU4PVqM1kGA/KP3rF0Sc008du+C+tIurA9fcWc8NTPnDUKBgCvXEbb/7O0uJV
+HTiProKc1Zw+4b73PvIurvKs8TYF1w8uYSeJNMv9sfPeRAkzHPXrH+GdUGl1WFHsIqJ9dch0mr/
OMyx8oaOZJQpmz3axQtpCLrt/1RUp9ZUq3zaHirZOmgYUd7OYPsd7Ntx6Cwk+71Opr8z8K8t/ppk
/HbFfWESkRy2XoKCzFJ5KsbY9bB6Og7qkclXen9iCBi7EnzLi2eMWjqGPlK+2MuJW508RCFlbAAC
RXD/xfneWSeQq6iO4zGiMlJt+r8dIu20ZjIVr5zZzhXEGCl1ekQRXk0EWL8p77y2Ab9RdWZNA+3u
jjQAYmCbMZbyNNNLUugzfyJU3mjkNLA53Me71YqUwARH57qp0XwscUv+fg6YuWzqHfT6rCfSMZX8
BznGIf7DQtrYFrIvRTiU46SKNNQrJQ+yQOxYGH+sJbaH90vzx11SmW7kcoESyDZvz4KndJzZxY0a
Vec6KJPhqoqsfkA/XPzwIQc5G6+0ggCgQ+Rx42K3CIgwwoPBCkI2b03lg/M2YXddBDDM2cJlQdkV
nCUqThHIK3QsFs5gpe1jr4vFisVAsyg7AJqU9cBPXxL/Lpg5fw8HgMPIje1k9YQ9LiiETypx9e3n
zLOaMxDEIylQTVGtvsTMud0juCGdWY2cueuLMTu6LWACp8Zq/txdueQmdU6sX7HoAAlYVBeSh1KY
kski1kZwWyNdX0C3t5AXUj11iJaEV7ZCV4mE3OTqksZv5tbkhmZnfsfr1LEPYMBS0TQ/Xl4/8eDI
8gvle+JxYnVx1LpQWYTMNSexQ3GVi9ailNC3L37IjC06pNyyoZ6LYH9evVYU6shIeuCMp9SDyVfm
JrRS/PfESYIUoeXU+5qVC7Z0CZP6q73F4tYlshJwnojj0jGRWKGayVufeBmkDCw/8BCwenIs0rEe
aIaaCf1Fja1PA5WJOlgJKi1oxHBtmmoEfdngeozeONuv9zUTBAKb2XK6ejrtiS9Kvh7oAkv0GCL3
wfPvr7t/PLgYeexOMPFWCUslX0OKbNzZIu+4khVRjawBj0BAEvw5bU/2Jd5nQ5uWYHBnXOwl7zUw
AcIA8D0wTrRmvyNmldzcHGIrrJczdZTwqiRE7OhB06Eu6yz+A9yJMBwdaXf1qksT3qXtnp6xnvTZ
SQ2nQ9Vsv6AWuQ60KjIA43e1QPYBqOIt3XMFCc7Erl4ag9O7SeS8QrzrhHAJN9zKw+UGPpFAkxZ+
qMBzh6RiB8cTkSOuoVmDLf5UGTT2LDWdIVZlHEs+aZRt0UYcGv1/6S/Ob+oY67X8nkWauc6q/q+p
UVFuLzsOOPGWjbX5gb/p1xc3cYGLsQmG3iI091HE63Lesmg6H7/N3ovN0PtbnMCANn85VGOdxazw
4c+Kud38b2pAQp5Uubf21CqjApUuxMyrXq9RgCbeEJbYMneJ1s3RutUIJXRuXLJFMKR/gXsZUO2E
SoHNdhDlm+LzKfIhpEcXPkrQNApr8hqs8/fHWwJAYz+4TJibXFGXGvcZOAZ0eiddqmE0KusVPl2N
tjMqWi9cELKZI64UVByiKCneFto63sKro8PgaX9esQyRWhuZyoh0yA/4Pc45L/0Y5qrVB3E7F1SH
r7H+nZe7h+SCzBNOvuNPKQZI58fF+MKdTAXJgMbtHHauOxGQWWcUA3KdePnPmalfhL852oEKiBgi
erjiGl7iVfilKy2728x/ybHRtX+hxA1AzwgrZL4baMUtvhTpF6NtklN1Ln4f+yMoR2oCjxeq8NBy
ApAN6uKZNa2pGPgqF42DnM45uxW+rCpixtgFNd2Fwuxc/n1zmjBkzl7KZLgIGUlfqalzovDbJMzN
7UOy92xUHMme4gPxMI3pmWqBZRdD5Saos+Dok6vvf6OpCXLCh2rRHtrR+2yVQiJ9RbyGly5z9YAm
1s/vu98Ys9grePeahPhbbUFocckUrPgC2kqIe0/Xk7U+5EYSgcRH/XZbuzT9nbUx9LhvD6O/+MOg
TJUDXAX3ZZ23ixXpFQsbXPodudhapbJ5Xl8wfFernJdIXKVqGgs3eV3DO+/Z21SZ2le5Tw1vg25e
ww5mfZ/6FlblIyv5FmzaxX9wEshucHlP1yqt7NbjWSW3GnBFwtvBZksJbzqYI11ebUz78bMye2dH
lt0JyHgFG9rDJQASNEsKx/kSCvLsvhNDbCxMLGtehfVOVkBNIXaL14LPIKkYu/X8UfGxfgfb9Q3Q
igTAqJLXxEXKRVyd+hsZLUQXYIaNsXol5pw/VPeY4FZn1r0cqVMoUk7Ukti9bY+LsvwKd/S84RS7
GLAi6Cdug2mPp134m0HJQr9pal44UmS+p/N5cQJ2Jw2XprNDNdOhxg0MxPHcsgjVs0EmmtYUbXGu
Fzt5wuA0W70NA8poC6mm7q2dQzvbRZpg6L/A0v6YzWjn3MQ30+FC9VVbRF+UI/uViUve58o/DbTi
6MrYO/TEdkFMwO6Pl63AldDBqgTqJeo7YUzuKgEmjSoCpF12IehNV1c/jI6MdGZ9ZTU+IF4peeNi
1mEXpn2dgRMIJ0YgJPcGIgLTT8krUZL3PXD8b+RXVNbachdy1jSB8GoBS4y0phr03xxJKoFdvVHA
hjvnZlycsZ8e67xlXaOrLMWSGoM2WV3cENp7w3ixek/eqWAFx//iFccjXW9du9TxTQPMAL8rSczl
9/cvFDzPIVre+yoMo2/t0kKx+zovIRsplY4tBOi1rkvJxxGEbPgXu17Fh6bZOiderfNTTkm2XkFZ
j6zVlzq71PJWO2yDKkayrEk1NSr9RsmFAetYVHumnjhML1Xu3lIt+jeeNBhohTkdC8eceG5YGH6Q
yoXlP1ZJsPBT/WndAKNTPtFfqDrCGO9oX2Rzl0dYwM1kKiCI70Z87mdq2WWFoFrUcvXtWIkBcBSD
82u/LqoOrLxokcZS4vIwjAPxLqVxemwfXgJ/gU2xNIlz9DNyoFI6NXgaimzRGW/rL11uTbl/udKx
n3YOczT0RdT+ZT8C5FCKTnM6r9keR8fSfDuuxnDx7jbjn9ARR4Z76ZDW1pw3D6WgBW3jhtc1jnEI
3yBYv8LLhZDAlTi14Ri7bTCo2sk0fxarr4SppIr+znLk6TpCr1DzrjnCXpTnjUX6z6QCSrGvH/47
5ixc80mllxjrThtpRBE5iQteifp6kMaxgTKS4J3Fw3KmPrdOm6JUEswkXpIjcEvi7guZU3OET9o+
zOKi7XyRMOklyZ6db0fNpyAKObtzWBfNzfdFRUPEjVOxUa3Yex59m3eEsOpkXTVlgjc8b9a6o44k
cSAYPtQ82ZTS3CfCWlnls+lf8AWCsFYKgljGr4yyeX/MxDJ5fe311moyuCLWKKNa1nmZNSmPK4yy
EToR/EUsiEHDExTHdZEJfoBxdylEPa51pRh8tjkXytwEhQZYNhWBgQ7jOyzsgT7xzi7FACgPrV6Y
4k44jhCfejevUa0LjVf9X2e7zRLKoZ1rWzIXPVqn5q46m/+M80Sbh5JKcMqTO9TqhC1VrztywARL
WyMLznT7DbmJOLQ96sfiF5TgPuVBNusl772EDNwiUhBaAXZCmMANOHr+269GVh20On5BYk0KL+hX
doAlxD1bADSp7gKvdoA7Anxdj01/fb+ZjHqHJV5R+HQ5H/BJk18+vRAByZiCxCEPKZdxdZhE2l89
yYQ2dcvCgIGTKdkPLSZZadMc1NYee62ioKTcAPf22uGV4mC1TkyhN4zkbLoMqSB11qXBiaWmXkZU
pJbPEbMVOKh0gtWxSq9r18UlK3QjIt6CRQy+i4mg3i/ypbRRCLShhtp0KxcMdmeJu4J1HdPaV7SN
mZW9sJpxBwfKFk6SMuAyUy6SPT9xpnGgNA+v7tH7s9vkPkHDEVWNxoZqusuJk80o3zDRQJBLOkzy
EmjB21Uirbkui56omooV7O1sMqhqT6dgk0mJ2j2ylDiMB4B7jr2z1AVQ7036DopYqeXsLeGNMyZY
QICsDM9Ye9TEOYVfwJzUmv1Z+LVbPZY6PAv//UEBzHnolFXzjwZB6tqCPcgjG8kkBT06qtvxv0eO
PuiJlqo0jhUh1OhxpTXMLPkPjxjmmN7LAATRL7ruXGYLrR87VFTbCYQfC3p9bHfnWfa6drM5yAqB
xaGclZqz+mmoACQA8k4UnAeWK/90l77NNEDcYO1btxZUU9mcA6HTKlWswH3n5ndYOolmCeIOJm/X
aqgI3nMvQkeBHzByMdI1Bb+O2Of/LyDU/BzxIusIyj0r9NzABg6WIMGajkszIniw300bRFY18WaZ
A/F/iguasZdD9Aj+Yl8ehaiZ+GdCmtNfcZ4kaZ8huq6exuHi7OOFmDG2obmrWdSZ1oYCQaO7lq8X
g3ADUkRReJqA1kAnxWcO/Ol/5wnePDhTt5i6DaiOH9qXOuXQSR/N9ejEB2DSLj7A/Hx50IXeYRuH
4/UtQY3sFFG7HyrlI9lZA4q5YFJ7QfgbmX5tHkV8Ag6tYmoqaww2RiOO6VNkDQyJJNb8YR59dbON
gpniOuSVr5zL26w+qk4fkfEvyOyho5pd0s+JrjNAzlmGwM4BzlBqLbt0ximt3OOMRgDxrxwrp2YJ
hWcFgo/3UBvurB+625Xo5eB1XHVw81jUt9F6ks9ujJ2clvA/hWNH1DBTpk7RmTPdcK1lIhoyWizr
klkdsuOHIsGlbSLBUFFSXZcQK9Y+jV0a/DZqWYc97zWdQpRervWxjQdG+zn3/RydIqiVLra7FYJa
APhkILnsRaLSZ8XoYKxzx7wAcpdjaD8AoykVDwYUzBWU02qr4yuQ6CChpdMpBygd1rF+nXnTId29
FnRzRF9ztdAvwKW8tLuoV7h9EVUOaTWK+SLmdfDKXqLU1N4qaOKidGXtNVWtU3AfPwRR49lN2iPB
V/fJkyS/mIDn2MEHDQ+sivOxZW4v/EfyaWxLa8qSLLKZwjx7tlR91tzj8Bu/V+RwAVQVUvLycPu6
wArUQe4hThl7yI4i1bjhWr5bi5V6KC7kiAOekRSzCBzCAcGrIZDI98rzeI0ZcKfx+KnZQ1exTcPz
gNfLZGkzYhKRox/VJjl62ECFYy0zGIKX4z9mcsc93DC+AzLYytnH53LHVu77gaiaA31Y3ttWRnhk
QjlYKi51y61XRvPvJqt7XZAqR2UYGhebakxlsL1/Dpca/hp2sgRQmsEUa8ooxoDl3bomYD7L7iJU
7VNqINDL+vZiueX7tf1/foAQPQb/6DmGuJbNy8JjpAmOnLEMbCARajYlv+NMRce/VZnNXQnnRkFd
h6LsmIdFEfK/xFfl/7CFFaL9uH4nTSKKJM/udJ2mbbv/5GXSokxMI2HKGoB4gIysxnoC0dVW3LRi
wtagjpe5ykSUpVsjtXpimD3AqQSlucKCNAysI6qNiF80Y//hmIQ5T+I9q797kQ6VfDawT4gISIyH
1MKeQWbrapM3AWoLHsPdwyQerk78mAGst/YELfFp8CKHCla8NH5YOtfgOZqU8XSDklScPTNrdENw
PqqaCns2t2fKrgOzM2bc9yOc6lYZNIfJIXHEGJ99c+O7/k1Cf1Z4H9Xyi0S07TcKKL4SrffJO4Aq
rkm+P8mMUqyAfGYbF4mL574wycQYwmtOQYQLBEEysQQmPXOcpK2u6dkaPF3VhISlJr1G4LpMc36C
soRT88JvcYjuxjTddGUvMnM+F8k/kD/OTt5Y+sqcTkj34HwtLFI76N75GdCCe5kpgBePpJVOQYwI
oajxlguRzJHEAWExc2yBh4Y4sJzMTofKCl+C1xKy+ZRYkLUlmdn0Xm9IxPFsfVmPLOpfCsC1Mfrs
mwwBvI6wIgE4kRnZPrFo9xM18XAYRR7S6/8B0g0txzmttTggdoxBYiI9Pyd/2hMHYcXu/hjatgK7
FhFj3Sl7y95iuN9kFVN+bYpHVCeNN8+LULmNokUpMB2eQ+cmw2OgVktZL4bFJ0MB4IMbXNQa8vgh
vz+k7J7BO3I/L4zFf9dq3wII2g0+rPrMuIb6PnQ0uP1vZJPLSWWatM9GS9QCOujY9N44bfAZY+hw
otQBdjgpIbUXZYr+Fc5yVYC/9iDKf5qsA7ctiO0naAA9Z85NkCKrcD/UB8eArpzL1HdRMKoU2ymr
k/oDRgSgc1MkiCGAQDjIPxfCr6IGCcEzFGEzr0OTPPsJKsoGO0BjgcZou/wuM1fxUAKMnLvA3q/E
botxZhjwA142Cz90bInk0tU/VLe16JYax7Sn6Zy5W6KtI/ugMW6sLMVeG4eTrB0BtC27RkSQmkce
F0j4DAyMa88J2xKYvxehAXYSfrPPC3zM25/jur0aqgB3T22oQ6wqrEx9LAhjAQXdqulrd1bi7k0s
oQggd8E83LAyWhkA7/J/eTEzJo8tm6MG8r8qd5jstN8AQdI234qUf8fMDsjAhl27SKnYt+UJlcCx
qECZHwP5Mm+h2hCHLwik1uhXLDFccf7LcjR3RXut71gcARCQEEkEAOq53Zz0GY9/cwX/Bwd6ivyv
PxpWUFvQ0pycfp+QWlI1qiL3KiQEgJWoO2XUqBPi5z4fJN7tvzGCLBGYMY6YIW8FCxW8kFJmU1zP
XYngsi0LGvo7wO6f9q2MxRT4gBxX4HfM9ucq6KzL37OvQWNGVHIDFaluA6lxShQTMjS/25ewpMm8
0uxks62ca2fX1Gtd0wxgndvlsjnSGVeb/VoZJX3oOtfPP9lagN3ZXif+8knKKPj46L7oJ8JPPyc/
i2RMM2Qvir42+3t6OyeddgcajSwTIqLFYQn1UdqNk9mYxia3rfp6C9pQmCJIF0q1gwNUjg/97a7E
UekgYD32g97Di4fzOyvPmK0gylmsCJ0cciVIStF2wkg4DQCzK3efA9+IjosDl/obXwL4ps/HSwYA
mjJorIk9YWZ4MgxxqqBddy9ZgVVDBSe65vsKaW9PPIdGr+fr8G5+IXN3xZrIzBpwpOiGyBOkmTLB
5BtCa9NA7zJYPHTlhaK4pbmkA5ad3Q7xw7pwQknR9Lteuq5ffXy0TLQvEeRWPN1yyMy5svEbpbcc
HyaMx+6xaGQ972R511dYUQ4OofWKlTaozjPMvyG03UCIVOg6kxxkMO3q/wMoiQB+eaMwwx0N3rA6
f6vnWnbEnHSTYk8yIz9V0XKkJpXCSY35/P1WO4qrdnZnHKJbJSv0G8lEtSPYLNFlZHHUpgwuArOw
YpL7vZIZTfAHweIhcuRqKmFuRgXw7BQ5+CF0WXbdSal4wNv9e5Z31yLEiw0u8CZJBvAGduJM3fHb
F/lngf6cx5td2KX03Lje55Aw9lPlB2AzBR/30wnB24lFQyVQ9zvoycVXWY8iZKF78hiBjZnzGW8h
bLzvZftV0wZypr/oUAG3GCtNAGY8dIStNt5Qp4rLFfVdOARdnP1Nw+EXQOZSbA/yaobnlYaZ6RfO
kU0moRZL7P6Et24wEq1AvwrbfQ/8V2mSNInh1t+IhdLF6pkia15OswgIHJKbca6HeWOegBUGb4G4
8L7EbFhytmTKu7BpvvCNLFHsGlQABp94EZTdnhBRSM/yjL7WejSESwXRLVaoiw0rVeMJvNzXHxtl
NP58/+0W46v6ktQENkF75DnqaN16A0ZE4LOPG3r6wZIR5kDiyfKkuFwP57rSqDlBQHeK4gQFYcJk
7PAR04AK5MinXQMOyKGdXv/KQYXtqU13UIkLJIkPoroRwuZW5bRbeJHr5XwT6ID529hw3kFTnZRf
wVW4/gSeTC5TLLK/ot9E2GEWUpC/GpXYZQEOBgnqNv9Z/KTiNq/RTyC7rLiY1RVyyURLRflFyONT
KckRFfV7vgpiD7TjNQ9+jTz7tvWUF1GI9zH+SghweDdL523FVINpjppg5Ol2mlUkF7VHOxUr/M9f
1dhFXT/YkOOyfoXsHOkOmc/qQZGKcKjztRjkmUS5iFscBaTdh8cviNw0kfoAKEEeIDFImVwyxvSX
3Ew5G7w+ApDP4tEyaQ63dbhVxWTbV733ydawubhLrACQdK4TQKWS7JtPLC9w3WxO/LsUXhWseSEs
tZ3hkX+dtDS+GxCql0WxCCYrbIN70NtM6LjiGzngd/h2cKr4MivcMCd1FrcyfIfbtyUjLwEdm6CT
mvrqK8NdyRaXcRbc9IBC0nLpKkMhLhXe1klk33X16CHnOSZjIMz+E0wmxIqIKvmBBTLzRzTSCfdX
s1ERtOhhnqYhLfjkkQ0WAPA0ft8QJFNboaN/7b6TouUZjYH+N4NafalSrzKGFUkwmliGssXQcyfY
PJOhFa2J+RgiGViUqydWVkB0KJdZqv+1iLM/1rlIInJzoyh5/HAHKeyLh6F9HE7z0rRIcKLRuZ2n
JB/wBAS0c862SasV9ppMmBdb+pOPYSSNieg4YAzpr5FVAk9I6zw7WHdYW0Vkho2dYmDTDTRPGK80
2Ie6EtblR/OmPr3mSsH/5vNyn2QqlS9el7CG3cbI+aukInSjK8aza0oEMI23+xTU5JoFYQkfrggq
xPs18MyTdBh0IuDsCflP3gM1AKWBsQgDS+HW+hOiqM9h9FjogFRCsaXEZ6cWCSojVzsLYtuY9sRH
IFu4u4jtd82I+8IGYZz/DxNDHuChmItNPQupEaEN1AlatBm17pP4nOTDfJYiUlPvHD49alqe/Nps
Gvo9FkjQrQdGB6Va9z/yrflQxqnYDwuY7B52pQ3g4l4MqsuPfHz24AWCx6jD0jKnWn61uyjHEEop
lJfBTp3Bi58aBNgvFOhcC+ww0Z6TewcMq6Cxchh4P0SnxBbflVjmuFtibxJlKhijRnsUu0ro8nDB
52LG4JZUtt9V2hxIscsae6fhOl7QNYrhFn4Gwdt1+aB3coSQ9MISSylQ2kKmTDy+PjMPVxbmv4sV
nSa45fGYfTB6iQDeJuTNib1c5FE0vZSQKrYj2BdrgBeWzj11De9+10IyA9NRez3kjNLDPx+9Lqzj
RnbqWm/WioGqqyWm5siSs9iYa7+mwJj/W4lnwdsT51eP+vid7CXaprVRPNoMf55u2qke0DzaXj/A
JxtvQ59uOgSTyJKZDW0UISeosuu0KSTtLbEOnaaCJR5YOk/dyt+s9Zy4rqenQtBoHaX44a5pK9Ed
YGjUFkY/NmRoy1vGMg3FtAvN8Zm33z9jIlafISZp+CKA/5YQjOqX7QRG5GnaUjqNeDQ8f4jIqynL
pPBp3dvaatQr7i5lUti7TntYsb2ULOfF2pArJLpbQm1Po6GOcDkPt5Vc2CR9FQrtzcmQzN7MAlw4
ZZaLFkcq7MeF18IXF/HWIyMab/FFcoxfzZYs+KwFeRs8yGxiyG4roEGyh1shkkmm8Sb4x4+S1LEo
2aOHrg32wCgtF577JnlspA==
`pragma protect end_protected
